library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity robotron_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of robotron_sound is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"76",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",
		X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"0F",X"8E",X"00",
		X"7F",X"CE",X"04",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"00",X"6F",X"02",X"86",X"37",
		X"A7",X"03",X"86",X"3C",X"A7",X"01",X"97",X"05",X"4F",X"97",X"03",X"97",X"00",X"97",X"01",X"97",
		X"02",X"97",X"04",X"0E",X"20",X"FE",X"DF",X"0C",X"CE",X"F0",X"EB",X"DF",X"07",X"86",X"80",X"D6",
		X"15",X"2A",X"09",X"D6",X"06",X"54",X"54",X"54",X"5C",X"5A",X"26",X"FD",X"7A",X"00",X"1A",X"27",
		X"4C",X"7A",X"00",X"1B",X"27",X"4C",X"7A",X"00",X"1C",X"27",X"4C",X"7A",X"00",X"1D",X"26",X"DF",
		X"D6",X"15",X"27",X"DB",X"C4",X"7F",X"D7",X"1D",X"D6",X"06",X"58",X"DB",X"06",X"CB",X"0B",X"D7",
		X"06",X"7A",X"00",X"2D",X"26",X"0E",X"D6",X"21",X"D7",X"2D",X"DE",X"07",X"09",X"8C",X"F0",X"E4",
		X"27",X"4E",X"DF",X"07",X"D6",X"06",X"2B",X"06",X"D4",X"19",X"C4",X"7F",X"20",X"05",X"D4",X"19",
		X"C4",X"7F",X"50",X"36",X"1B",X"16",X"32",X"DE",X"07",X"AD",X"00",X"20",X"A2",X"CE",X"00",X"12",
		X"20",X"08",X"CE",X"00",X"13",X"20",X"03",X"CE",X"00",X"14",X"6D",X"18",X"27",X"12",X"6A",X"18",
		X"26",X"0E",X"E6",X"0C",X"E7",X"18",X"E6",X"00",X"EB",X"10",X"E1",X"14",X"27",X"12",X"E7",X"00",
		X"E6",X"00",X"E7",X"08",X"AB",X"04",X"60",X"04",X"16",X"DE",X"07",X"AD",X"00",X"7E",X"F0",X"4F",
		X"DE",X"0C",X"39",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"54",X"F7",X"04",X"00",X"39",X"CE",
		X"F3",X"D2",X"C6",X"1C",X"BD",X"F9",X"65",X"BD",X"F0",X"46",X"39",X"CE",X"F3",X"EE",X"20",X"F2",
		X"CE",X"F4",X"0A",X"20",X"ED",X"CE",X"F4",X"26",X"20",X"E8",X"CE",X"F4",X"42",X"20",X"E3",X"CE",
		X"F4",X"7A",X"20",X"DE",X"CE",X"F4",X"96",X"20",X"D9",X"CE",X"00",X"60",X"A6",X"00",X"80",X"02",
		X"A7",X"00",X"BD",X"F3",X"30",X"7E",X"F3",X"49",X"CE",X"00",X"01",X"DF",X"12",X"CE",X"03",X"80",
		X"DF",X"14",X"7F",X"04",X"00",X"DE",X"12",X"08",X"DF",X"12",X"09",X"26",X"FD",X"73",X"04",X"00",
		X"DE",X"14",X"09",X"26",X"FD",X"20",X"EB",X"86",X"FF",X"97",X"12",X"CE",X"FE",X"C0",X"DF",X"14",
		X"86",X"20",X"CE",X"FF",X"E0",X"8D",X"05",X"86",X"01",X"CE",X"00",X"44",X"97",X"16",X"DF",X"17",
		X"CE",X"00",X"10",X"8D",X"21",X"96",X"13",X"9B",X"15",X"97",X"13",X"96",X"12",X"99",X"14",X"97",
		X"12",X"09",X"26",X"EF",X"96",X"15",X"9B",X"16",X"97",X"15",X"24",X"03",X"7C",X"00",X"14",X"DE",
		X"14",X"9C",X"17",X"26",X"DB",X"39",X"4F",X"B7",X"04",X"00",X"8B",X"20",X"24",X"F9",X"8D",X"09",
		X"86",X"E0",X"B7",X"04",X"00",X"80",X"20",X"24",X"F9",X"D6",X"12",X"86",X"02",X"4A",X"26",X"FD",
		X"5A",X"26",X"F8",X"39",X"86",X"80",X"97",X"1C",X"86",X"F1",X"97",X"1A",X"86",X"80",X"97",X"10",
		X"86",X"12",X"4A",X"26",X"FD",X"96",X"19",X"9B",X"1C",X"97",X"19",X"44",X"44",X"44",X"8B",X"D8",
		X"97",X"1B",X"DE",X"1A",X"A6",X"00",X"B7",X"04",X"00",X"7A",X"00",X"10",X"26",X"E2",X"7A",X"00",
		X"1C",X"96",X"1C",X"81",X"20",X"26",X"D5",X"39",X"80",X"8C",X"98",X"A5",X"B0",X"BC",X"C6",X"D0",
		X"DA",X"E2",X"EA",X"F0",X"F5",X"FA",X"FD",X"FE",X"FF",X"FE",X"FD",X"FA",X"F5",X"F0",X"EA",X"E2",
		X"DA",X"D0",X"C6",X"BC",X"B0",X"A5",X"98",X"8C",X"80",X"73",X"67",X"5A",X"4F",X"43",X"39",X"2F",
		X"25",X"1D",X"15",X"0F",X"0A",X"05",X"02",X"01",X"00",X"01",X"02",X"05",X"0A",X"0F",X"15",X"1D",
		X"25",X"2F",X"39",X"43",X"4F",X"5A",X"67",X"73",X"7F",X"04",X"02",X"CE",X"F2",X"5F",X"DF",X"14",
		X"DE",X"14",X"A6",X"00",X"27",X"33",X"E6",X"01",X"C4",X"F0",X"D7",X"13",X"E6",X"01",X"08",X"08",
		X"DF",X"14",X"97",X"12",X"C4",X"0F",X"96",X"13",X"B7",X"04",X"00",X"96",X"12",X"CE",X"00",X"05",
		X"09",X"26",X"FD",X"4A",X"26",X"F7",X"7F",X"04",X"00",X"96",X"12",X"CE",X"00",X"05",X"09",X"26",
		X"FD",X"4A",X"26",X"F7",X"5A",X"26",X"DF",X"20",X"C7",X"86",X"80",X"B7",X"04",X"02",X"39",X"01",
		X"FC",X"02",X"FC",X"03",X"F8",X"04",X"F8",X"06",X"F8",X"08",X"F4",X"0C",X"F4",X"10",X"F4",X"20",
		X"F2",X"40",X"F1",X"60",X"F1",X"80",X"F1",X"A0",X"F1",X"C0",X"F1",X"00",X"00",X"7A",X"00",X"2E",
		X"20",X"04",X"C6",X"A0",X"D7",X"2E",X"86",X"04",X"97",X"13",X"86",X"9F",X"D6",X"2E",X"CE",X"01",
		X"C0",X"09",X"27",X"20",X"F7",X"00",X"12",X"B7",X"04",X"00",X"09",X"27",X"17",X"7A",X"00",X"12",
		X"26",X"F8",X"09",X"27",X"0F",X"D7",X"12",X"73",X"04",X"00",X"09",X"27",X"07",X"7A",X"00",X"12",
		X"26",X"F8",X"20",X"DD",X"D0",X"13",X"C1",X"10",X"22",X"D4",X"39",X"C6",X"11",X"D7",X"2E",X"86",
		X"FE",X"97",X"13",X"20",X"C5",X"CE",X"F4",X"B2",X"20",X"26",X"BD",X"F3",X"30",X"BD",X"F3",X"49",
		X"39",X"CE",X"F4",X"B8",X"20",X"F4",X"C6",X"FF",X"D7",X"09",X"CE",X"F4",X"BE",X"8D",X"EB",X"CE",
		X"F4",X"C4",X"8D",X"E6",X"5A",X"26",X"F3",X"39",X"CE",X"F4",X"CA",X"20",X"DD",X"CE",X"F4",X"D6",
		X"8D",X"D8",X"8D",X"30",X"20",X"FA",X"86",X"FF",X"97",X"09",X"CE",X"F4",X"DC",X"20",X"F1",X"86",
		X"FF",X"97",X"09",X"CE",X"F4",X"D0",X"20",X"E8",X"C6",X"30",X"CE",X"F4",X"E2",X"8D",X"21",X"96",
		X"06",X"48",X"9B",X"06",X"8B",X"0B",X"97",X"06",X"44",X"44",X"8B",X"0C",X"97",X"13",X"8D",X"29",
		X"5A",X"26",X"EC",X"39",X"96",X"09",X"80",X"08",X"2A",X"03",X"97",X"09",X"39",X"32",X"32",X"39",
		X"A6",X"00",X"97",X"13",X"A6",X"01",X"97",X"14",X"A6",X"02",X"97",X"15",X"A6",X"03",X"97",X"16",
		X"A6",X"04",X"97",X"17",X"A6",X"05",X"97",X"18",X"39",X"96",X"09",X"37",X"D6",X"17",X"D7",X"19",
		X"D6",X"14",X"D7",X"1A",X"43",X"D6",X"13",X"B7",X"04",X"00",X"5A",X"26",X"FD",X"43",X"D6",X"13",
		X"20",X"00",X"08",X"09",X"08",X"09",X"B7",X"04",X"00",X"5A",X"26",X"FD",X"7A",X"00",X"1A",X"27",
		X"16",X"7A",X"00",X"19",X"26",X"DE",X"43",X"D6",X"17",X"B7",X"04",X"00",X"D7",X"19",X"D6",X"13",
		X"9B",X"18",X"2B",X"1E",X"01",X"20",X"15",X"08",X"09",X"01",X"43",X"D6",X"14",X"B7",X"04",X"00",
		X"D7",X"1A",X"D6",X"13",X"D0",X"15",X"D1",X"16",X"D1",X"16",X"27",X"06",X"D7",X"13",X"C0",X"05",
		X"20",X"B8",X"33",X"39",X"DA",X"FF",X"DA",X"80",X"26",X"01",X"26",X"80",X"07",X"0A",X"07",X"00",
		X"F9",X"F6",X"F9",X"00",X"3A",X"3E",X"50",X"46",X"33",X"2C",X"27",X"20",X"25",X"1C",X"1A",X"17",
		X"14",X"11",X"10",X"33",X"08",X"03",X"02",X"01",X"02",X"03",X"04",X"05",X"06",X"0A",X"1E",X"32",
		X"70",X"00",X"FF",X"FF",X"FF",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"90",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"01",
		X"00",X"00",X"3F",X"3F",X"00",X"00",X"48",X"01",X"00",X"00",X"01",X"08",X"00",X"00",X"81",X"01",
		X"00",X"00",X"01",X"FF",X"00",X"00",X"01",X"08",X"00",X"00",X"01",X"10",X"00",X"00",X"3F",X"3F",
		X"00",X"00",X"01",X"10",X"00",X"00",X"05",X"05",X"00",X"00",X"01",X"01",X"00",X"00",X"31",X"FF",
		X"00",X"00",X"05",X"05",X"00",X"00",X"30",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"04",X"00",X"00",X"04",X"7F",X"00",X"00",X"7F",X"04",X"00",X"00",X"04",X"FF",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",X"0C",X"68",
		X"68",X"00",X"07",X"1F",X"0F",X"00",X"0C",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"01",X"04",X"00",X"00",X"3F",X"7F",
		X"00",X"00",X"01",X"04",X"00",X"00",X"05",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"48",X"00",
		X"00",X"00",X"05",X"FF",X"00",X"00",X"02",X"80",X"00",X"30",X"0A",X"7F",X"00",X"7F",X"02",X"80",
		X"00",X"30",X"C0",X"80",X"00",X"20",X"01",X"10",X"00",X"15",X"C0",X"10",X"00",X"00",X"C0",X"80",
		X"00",X"00",X"FF",X"01",X"02",X"C3",X"FF",X"00",X"01",X"03",X"FF",X"80",X"FF",X"00",X"20",X"03",
		X"FF",X"50",X"FF",X"00",X"50",X"03",X"01",X"20",X"FF",X"00",X"FE",X"04",X"02",X"04",X"FF",X"00",
		X"48",X"03",X"01",X"0C",X"FF",X"00",X"48",X"02",X"01",X"0C",X"FF",X"00",X"E0",X"01",X"02",X"10",
		X"FF",X"00",X"50",X"FF",X"00",X"00",X"60",X"80",X"FF",X"02",X"01",X"06",X"FF",X"00",X"16",X"48",
		X"48",X"48",X"1B",X"CE",X"00",X"12",X"DF",X"0E",X"CE",X"FC",X"08",X"BD",X"FB",X"92",X"C6",X"09",
		X"7E",X"F9",X"65",X"96",X"1A",X"B7",X"04",X"00",X"96",X"12",X"97",X"1B",X"96",X"13",X"97",X"1C",
		X"DE",X"17",X"96",X"1B",X"73",X"04",X"00",X"09",X"27",X"10",X"4A",X"26",X"FA",X"73",X"04",X"00",
		X"96",X"1C",X"09",X"27",X"05",X"4A",X"26",X"FA",X"20",X"E8",X"B6",X"04",X"00",X"2B",X"01",X"43",
		X"8B",X"00",X"B7",X"04",X"00",X"96",X"1B",X"9B",X"14",X"97",X"1B",X"96",X"1C",X"9B",X"15",X"97",
		X"1C",X"91",X"16",X"26",X"CB",X"96",X"19",X"27",X"06",X"9B",X"12",X"97",X"12",X"26",X"B9",X"39",
		X"86",X"FF",X"97",X"19",X"86",X"60",X"C6",X"FF",X"20",X"12",X"86",X"01",X"97",X"19",X"C6",X"03",
		X"20",X"0A",X"86",X"FE",X"97",X"19",X"86",X"C0",X"C6",X"10",X"20",X"00",X"97",X"18",X"86",X"FF",
		X"B7",X"04",X"00",X"D7",X"14",X"D6",X"14",X"96",X"06",X"44",X"44",X"44",X"98",X"06",X"44",X"76",
		X"00",X"05",X"76",X"00",X"06",X"24",X"03",X"73",X"04",X"00",X"96",X"18",X"4A",X"26",X"FD",X"5A",
		X"26",X"E5",X"96",X"18",X"9B",X"19",X"97",X"18",X"26",X"DB",X"39",X"86",X"20",X"97",X"14",X"97",
		X"17",X"86",X"01",X"CE",X"00",X"01",X"C6",X"FF",X"20",X"00",X"97",X"12",X"DF",X"15",X"D7",X"13",
		X"D6",X"14",X"96",X"06",X"44",X"44",X"44",X"98",X"06",X"44",X"76",X"00",X"05",X"76",X"00",X"06",
		X"86",X"00",X"24",X"02",X"96",X"13",X"B7",X"04",X"00",X"DE",X"15",X"09",X"26",X"FD",X"5A",X"26",
		X"E1",X"D6",X"13",X"D0",X"12",X"27",X"09",X"DE",X"15",X"08",X"96",X"17",X"27",X"D0",X"20",X"CC",
		X"39",X"CE",X"F6",X"00",X"DF",X"23",X"BD",X"F7",X"2A",X"CE",X"A5",X"00",X"DF",X"05",X"CE",X"F6",
		X"29",X"BD",X"F6",X"33",X"BD",X"F6",X"CE",X"CE",X"F6",X"2E",X"BD",X"F6",X"33",X"7E",X"F6",X"DB",
		X"90",X"10",X"02",X"14",X"40",X"B4",X"40",X"FF",X"14",X"30",X"D0",X"32",X"02",X"10",X"60",X"EE",
		X"20",X"02",X"08",X"54",X"E9",X"54",X"FF",X"20",X"28",X"C0",X"30",X"02",X"14",X"58",X"AC",X"20",
		X"02",X"08",X"58",X"A6",X"58",X"FF",X"18",X"22",X"00",X"30",X"10",X"FC",X"00",X"01",X"30",X"FC",
		X"01",X"00",X"01",X"A6",X"00",X"97",X"2A",X"A6",X"01",X"97",X"13",X"A6",X"02",X"97",X"12",X"A6",
		X"03",X"97",X"17",X"A6",X"04",X"97",X"2F",X"39",X"8D",X"E9",X"8D",X"30",X"8D",X"58",X"96",X"2E",
		X"91",X"2F",X"26",X"F8",X"59",X"F7",X"04",X"00",X"8D",X"2D",X"8D",X"38",X"8D",X"5C",X"7D",X"00",
		X"13",X"27",X"E4",X"7D",X"00",X"14",X"26",X"E4",X"7D",X"00",X"17",X"27",X"DF",X"2B",X"05",X"7C",
		X"00",X"2F",X"20",X"D8",X"7A",X"00",X"2F",X"7A",X"00",X"2E",X"20",X"D0",X"7F",X"00",X"14",X"96",
		X"2F",X"97",X"2E",X"7F",X"00",X"2D",X"39",X"96",X"06",X"44",X"44",X"44",X"98",X"06",X"97",X"28",
		X"08",X"84",X"07",X"39",X"96",X"28",X"44",X"76",X"00",X"05",X"76",X"00",X"06",X"86",X"00",X"24",
		X"02",X"96",X"13",X"97",X"2D",X"39",X"96",X"2F",X"7A",X"00",X"2E",X"27",X"04",X"08",X"09",X"20",
		X"08",X"97",X"2E",X"D6",X"2D",X"54",X"7C",X"00",X"14",X"39",X"96",X"2A",X"91",X"14",X"27",X"04",
		X"08",X"09",X"20",X"09",X"7F",X"00",X"14",X"96",X"13",X"90",X"12",X"97",X"13",X"39",X"7F",X"00",
		X"21",X"7F",X"00",X"2B",X"86",X"0E",X"97",X"22",X"7F",X"00",X"27",X"8D",X"9F",X"8D",X"A8",X"BD",
		X"F7",X"64",X"8D",X"B0",X"BD",X"F7",X"64",X"8D",X"BD",X"8D",X"79",X"8D",X"CD",X"8D",X"75",X"8D",
		X"0A",X"8D",X"71",X"8D",X"1D",X"8D",X"6D",X"8D",X"52",X"20",X"E2",X"96",X"26",X"7A",X"00",X"22",
		X"27",X"07",X"B6",X"00",X"13",X"26",X"0A",X"20",X"68",X"97",X"22",X"96",X"21",X"9B",X"2B",X"97",
		X"21",X"39",X"96",X"21",X"91",X"29",X"27",X"07",X"08",X"96",X"13",X"26",X"2A",X"20",X"29",X"7F",
		X"00",X"21",X"7F",X"00",X"2B",X"7F",X"00",X"27",X"DE",X"23",X"A6",X"00",X"97",X"20",X"27",X"17",
		X"A6",X"01",X"97",X"25",X"A6",X"02",X"97",X"2C",X"A6",X"03",X"97",X"26",X"A6",X"04",X"97",X"29",
		X"86",X"05",X"BD",X"FB",X"92",X"DF",X"23",X"39",X"32",X"32",X"39",X"96",X"20",X"27",X"06",X"91",
		X"13",X"26",X"04",X"20",X"03",X"08",X"09",X"39",X"7F",X"00",X"20",X"96",X"25",X"97",X"21",X"96",
		X"2C",X"97",X"2B",X"39",X"96",X"27",X"9B",X"21",X"97",X"27",X"2A",X"01",X"43",X"1B",X"B7",X"04",
		X"00",X"39",X"C6",X"01",X"D7",X"00",X"CE",X"F7",X"85",X"20",X"2A",X"CE",X"F7",X"8B",X"20",X"25",
		X"CE",X"F7",X"91",X"20",X"20",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"01",X"00",X"01",X"FF",X"03",X"E8",X"01",X"01",X"01",X"40",X"10",X"00",X"01",X"80",X"01",
		X"40",X"FF",X"CE",X"F7",X"97",X"A6",X"00",X"97",X"19",X"A6",X"01",X"97",X"15",X"A6",X"02",X"E6",
		X"03",X"EE",X"04",X"97",X"18",X"D7",X"12",X"DF",X"16",X"7F",X"00",X"14",X"DE",X"16",X"B6",X"04",
		X"00",X"16",X"54",X"54",X"54",X"D8",X"06",X"54",X"76",X"00",X"05",X"76",X"00",X"06",X"D6",X"12",
		X"7D",X"00",X"19",X"27",X"04",X"D4",X"05",X"DB",X"15",X"D7",X"13",X"D6",X"14",X"91",X"06",X"22",
		X"12",X"09",X"27",X"26",X"B7",X"04",X"00",X"DB",X"14",X"99",X"13",X"25",X"16",X"91",X"06",X"23",
		X"F0",X"20",X"10",X"09",X"27",X"14",X"B7",X"04",X"00",X"D0",X"14",X"92",X"13",X"25",X"04",X"91",
		X"06",X"22",X"F0",X"96",X"06",X"B7",X"04",X"00",X"20",X"B7",X"D6",X"18",X"27",X"B3",X"96",X"12",
		X"D6",X"14",X"44",X"56",X"44",X"56",X"44",X"56",X"43",X"50",X"82",X"FF",X"DB",X"14",X"99",X"12",
		X"D7",X"14",X"97",X"12",X"26",X"96",X"C1",X"07",X"26",X"92",X"39",X"86",X"FC",X"97",X"0E",X"CE",
		X"00",X"64",X"DF",X"0A",X"DB",X"0B",X"96",X"10",X"99",X"0A",X"97",X"10",X"DE",X"0A",X"25",X"04",
		X"20",X"00",X"20",X"03",X"08",X"27",X"11",X"DF",X"0A",X"84",X"0F",X"8B",X"47",X"97",X"0F",X"DE",
		X"0E",X"A6",X"00",X"B7",X"04",X"00",X"20",X"DC",X"39",X"4F",X"B7",X"04",X"00",X"97",X"10",X"4F",
		X"91",X"10",X"26",X"03",X"73",X"04",X"00",X"C6",X"12",X"5A",X"26",X"FD",X"4C",X"2A",X"F1",X"73",
		X"04",X"00",X"7C",X"00",X"10",X"2A",X"E8",X"39",X"CE",X"00",X"12",X"6F",X"00",X"08",X"8C",X"00",
		X"1A",X"26",X"F8",X"86",X"40",X"97",X"12",X"CE",X"00",X"12",X"86",X"80",X"97",X"10",X"5F",X"A6",
		X"01",X"AB",X"00",X"A7",X"01",X"2A",X"02",X"DB",X"10",X"74",X"00",X"10",X"08",X"08",X"8C",X"00",
		X"1A",X"26",X"EC",X"F7",X"04",X"00",X"7C",X"00",X"11",X"26",X"DC",X"CE",X"00",X"12",X"5F",X"A6",
		X"00",X"27",X"0B",X"81",X"37",X"26",X"04",X"C6",X"41",X"E7",X"02",X"6A",X"00",X"5C",X"08",X"08",
		X"8C",X"00",X"1A",X"26",X"EA",X"5D",X"26",X"BF",X"39",X"7A",X"00",X"04",X"39",X"8D",X"03",X"7E",
		X"FB",X"7F",X"7F",X"00",X"04",X"97",X"10",X"CE",X"FC",X"57",X"A6",X"00",X"27",X"2D",X"7A",X"00",
		X"10",X"27",X"06",X"4C",X"BD",X"FB",X"92",X"20",X"F1",X"08",X"DF",X"0E",X"BD",X"FB",X"92",X"DF",
		X"0C",X"DE",X"0E",X"A6",X"00",X"97",X"14",X"A6",X"01",X"EE",X"02",X"DF",X"12",X"8D",X"0E",X"DE",
		X"0E",X"08",X"08",X"08",X"08",X"DF",X"0E",X"9C",X"0C",X"26",X"E8",X"39",X"39",X"CE",X"00",X"15",
		X"80",X"02",X"23",X"15",X"81",X"03",X"27",X"09",X"C6",X"01",X"E7",X"00",X"08",X"80",X"02",X"20",
		X"F1",X"C6",X"91",X"E7",X"00",X"6F",X"01",X"08",X"08",X"C6",X"7E",X"E7",X"00",X"C6",X"F9",X"E7",
		X"01",X"C6",X"37",X"E7",X"02",X"DE",X"12",X"4F",X"F6",X"00",X"11",X"5C",X"D7",X"11",X"D4",X"14",
		X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",
		X"89",X"00",X"54",X"89",X"00",X"1B",X"48",X"48",X"48",X"48",X"48",X"B7",X"04",X"00",X"09",X"27",
		X"03",X"7E",X"00",X"15",X"39",X"36",X"A6",X"00",X"DF",X"0C",X"DE",X"0E",X"A7",X"00",X"08",X"DF",
		X"0E",X"DE",X"0C",X"08",X"5A",X"26",X"EF",X"32",X"39",X"4F",X"97",X"00",X"97",X"01",X"39",X"7F",
		X"00",X"00",X"96",X"01",X"84",X"7F",X"81",X"1D",X"26",X"01",X"4F",X"4C",X"97",X"01",X"39",X"86",
		X"0E",X"BD",X"F9",X"DC",X"96",X"01",X"48",X"48",X"43",X"BD",X"FA",X"94",X"7C",X"00",X"16",X"BD",
		X"FA",X"96",X"20",X"F8",X"86",X"03",X"BD",X"F4",X"EE",X"D6",X"02",X"C1",X"1F",X"26",X"01",X"5F",
		X"5C",X"D7",X"02",X"86",X"20",X"10",X"5F",X"81",X"14",X"23",X"05",X"CB",X"0E",X"4A",X"20",X"F7",
		X"CB",X"05",X"4A",X"26",X"FB",X"D7",X"12",X"BD",X"F5",X"03",X"20",X"FB",X"96",X"03",X"26",X"09",
		X"7C",X"00",X"03",X"86",X"0D",X"8D",X"05",X"20",X"69",X"7E",X"FA",X"89",X"16",X"58",X"1B",X"1B",
		X"1B",X"CE",X"FE",X"45",X"BD",X"FB",X"92",X"A6",X"00",X"16",X"84",X"0F",X"97",X"13",X"54",X"54",
		X"54",X"54",X"D7",X"12",X"A6",X"01",X"16",X"54",X"54",X"54",X"54",X"D7",X"14",X"84",X"0F",X"97",
		X"10",X"DF",X"0A",X"CE",X"FD",X"32",X"7A",X"00",X"10",X"2B",X"08",X"A6",X"00",X"4C",X"BD",X"FB",
		X"92",X"20",X"F3",X"DF",X"17",X"BD",X"FA",X"D0",X"DE",X"0A",X"A6",X"02",X"97",X"19",X"BD",X"FA",
		X"E2",X"DE",X"0A",X"A6",X"03",X"97",X"15",X"A6",X"04",X"97",X"16",X"A6",X"05",X"16",X"A6",X"06",
		X"CE",X"FF",X"02",X"BD",X"FB",X"92",X"17",X"DF",X"1A",X"7F",X"00",X"22",X"BD",X"FB",X"92",X"DF",
		X"1C",X"39",X"96",X"12",X"97",X"21",X"DE",X"1A",X"DF",X"0C",X"DE",X"0C",X"A6",X"00",X"9B",X"22",
		X"97",X"20",X"9C",X"1C",X"27",X"26",X"D6",X"13",X"08",X"DF",X"0C",X"CE",X"00",X"23",X"96",X"20",
		X"4A",X"26",X"FD",X"A6",X"00",X"B7",X"04",X"00",X"08",X"9C",X"1E",X"26",X"F1",X"5A",X"27",X"DA",
		X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"09",X"01",X"01",X"20",X"DF",X"96",X"14",X"8D",X"62",
		X"7A",X"00",X"21",X"26",X"C1",X"96",X"03",X"26",X"46",X"96",X"15",X"27",X"42",X"7A",X"00",X"16",
		X"27",X"3D",X"9B",X"22",X"97",X"22",X"DE",X"1A",X"5F",X"96",X"22",X"7D",X"00",X"15",X"2B",X"06",
		X"AB",X"00",X"25",X"08",X"20",X"0B",X"AB",X"00",X"27",X"02",X"25",X"05",X"5D",X"27",X"08",X"20",
		X"0F",X"5D",X"26",X"03",X"DF",X"1A",X"5C",X"08",X"9C",X"1C",X"26",X"DD",X"5D",X"26",X"01",X"39",
		X"DF",X"1C",X"96",X"14",X"27",X"06",X"8D",X"08",X"96",X"19",X"8D",X"16",X"7E",X"FA",X"42",X"39",
		X"CE",X"00",X"23",X"DF",X"0E",X"DE",X"17",X"E6",X"00",X"08",X"BD",X"F9",X"65",X"DE",X"0E",X"DF",
		X"1E",X"39",X"4D",X"27",X"2B",X"DE",X"17",X"DF",X"0C",X"CE",X"00",X"23",X"97",X"11",X"DF",X"0E",
		X"DE",X"0C",X"D6",X"11",X"D7",X"10",X"E6",X"01",X"54",X"54",X"54",X"54",X"08",X"DF",X"0C",X"DE",
		X"0E",X"A6",X"00",X"10",X"7A",X"00",X"10",X"26",X"FA",X"A7",X"00",X"08",X"9C",X"1E",X"26",X"DE",
		X"39",X"8E",X"00",X"7F",X"B6",X"04",X"02",X"CE",X"F0",X"EB",X"DF",X"07",X"CE",X"00",X"12",X"DF",
		X"0E",X"C6",X"AF",X"D7",X"09",X"0E",X"43",X"84",X"3F",X"D6",X"04",X"27",X"03",X"BD",X"F8",X"CD",
		X"5F",X"81",X"0E",X"27",X"02",X"D7",X"02",X"81",X"12",X"27",X"02",X"D7",X"03",X"4D",X"27",X"3F",
		X"4A",X"81",X"1F",X"2D",X"14",X"81",X"3D",X"2E",X"08",X"81",X"2A",X"22",X"08",X"80",X"10",X"20",
		X"0C",X"80",X"39",X"20",X"24",X"80",X"1C",X"20",X"12",X"81",X"0C",X"22",X"08",X"BD",X"F9",X"DC",
		X"BD",X"FA",X"42",X"20",X"1A",X"81",X"1B",X"22",X"0E",X"80",X"0D",X"48",X"CE",X"FB",X"C4",X"8D",
		X"21",X"EE",X"00",X"AD",X"00",X"20",X"08",X"80",X"1C",X"BD",X"F4",X"EE",X"BD",X"F5",X"03",X"96",
		X"00",X"9A",X"01",X"27",X"FE",X"4F",X"97",X"03",X"96",X"00",X"27",X"03",X"7E",X"F7",X"72",X"7E",
		X"F9",X"8F",X"DF",X"0C",X"9B",X"0D",X"97",X"0D",X"24",X"03",X"7C",X"00",X"0C",X"DE",X"0C",X"39",
		X"0F",X"8E",X"00",X"7F",X"CE",X"FF",X"FF",X"5F",X"E9",X"00",X"09",X"8C",X"F0",X"00",X"26",X"F8",
		X"E1",X"00",X"27",X"01",X"3E",X"BD",X"F7",X"A2",X"86",X"02",X"BD",X"F8",X"D2",X"86",X"01",X"BD",
		X"F8",X"D2",X"20",X"DC",X"F9",X"A4",X"F7",X"72",X"F9",X"7F",X"F5",X"5A",X"F9",X"CC",X"F9",X"79",
		X"F5",X"9B",X"F5",X"62",X"F7",X"7B",X"F7",X"80",X"F8",X"2B",X"F8",X"59",X"F8",X"78",X"F8",X"C9",
		X"F9",X"0C",X"F0",X"FB",X"F1",X"0A",X"F0",X"EF",X"F2",X"F6",X"F2",X"D1",X"F2",X"D6",X"F2",X"E8",
		X"F2",X"FF",X"F3",X"08",X"F2",X"BB",X"F1",X"28",X"F1",X"0F",X"F1",X"14",X"F5",X"50",X"F5",X"E1",
		X"F2",X"18",X"F1",X"47",X"F1",X"A4",X"F7",X"A2",X"40",X"01",X"00",X"10",X"E1",X"00",X"80",X"FF",
		X"FF",X"28",X"01",X"00",X"08",X"81",X"02",X"00",X"FF",X"FF",X"28",X"81",X"00",X"FC",X"01",X"02",
		X"00",X"FC",X"FF",X"FF",X"01",X"00",X"18",X"41",X"04",X"80",X"00",X"FF",X"00",X"FF",X"08",X"FF",
		X"68",X"04",X"80",X"00",X"FF",X"28",X"81",X"00",X"FC",X"01",X"02",X"00",X"FC",X"FF",X"60",X"01",
		X"57",X"08",X"E1",X"02",X"00",X"FE",X"80",X"8C",X"5B",X"B6",X"40",X"BF",X"49",X"A4",X"73",X"73",
		X"A4",X"49",X"BF",X"40",X"B6",X"5B",X"8C",X"1C",X"F8",X"04",X"05",X"55",X"00",X"04",X"05",X"55",
		X"F8",X"04",X"05",X"55",X"00",X"04",X"05",X"55",X"F8",X"04",X"05",X"55",X"00",X"04",X"05",X"55",
		X"F8",X"17",X"3B",X"41",X"B0",X"1F",X"1D",X"04",X"CB",X"00",X"04",X"06",X"66",X"3E",X"1D",X"04",
		X"CB",X"00",X"04",X"1F",X"FE",X"3E",X"3F",X"03",X"97",X"00",X"04",X"06",X"66",X"7C",X"3F",X"03",
		X"97",X"00",X"04",X"1F",X"FE",X"7C",X"1D",X"04",X"CB",X"00",X"04",X"06",X"66",X"F8",X"1D",X"04",
		X"CB",X"00",X"04",X"06",X"66",X"7C",X"3F",X"03",X"97",X"00",X"04",X"06",X"66",X"F8",X"3F",X"03",
		X"97",X"00",X"04",X"2C",X"CA",X"7C",X"3F",X"03",X"97",X"7C",X"1D",X"04",X"CB",X"7C",X"12",X"05",
		X"61",X"7C",X"0D",X"05",X"B3",X"7C",X"12",X"05",X"61",X"7C",X"0D",X"05",X"B3",X"7C",X"04",X"06",
		X"66",X"7C",X"0D",X"05",X"B3",X"7C",X"12",X"05",X"61",X"7C",X"1D",X"04",X"CB",X"3E",X"37",X"03",
		X"CE",X"3E",X"3F",X"03",X"97",X"7C",X"04",X"06",X"66",X"7C",X"0D",X"05",X"B3",X"7C",X"12",X"05",
		X"61",X"7C",X"1D",X"04",X"CB",X"7C",X"23",X"04",X"86",X"7C",X"1D",X"04",X"CB",X"7C",X"12",X"05",
		X"61",X"3E",X"1D",X"04",X"CB",X"00",X"04",X"06",X"66",X"7C",X"1D",X"04",X"CB",X"00",X"04",X"06",
		X"66",X"3E",X"3F",X"03",X"97",X"00",X"04",X"06",X"66",X"7C",X"3F",X"03",X"97",X"00",X"04",X"1F",
		X"FE",X"F8",X"1D",X"2F",X"EE",X"00",X"47",X"3F",X"37",X"30",X"29",X"23",X"1D",X"17",X"12",X"0D",
		X"08",X"04",X"08",X"7F",X"D9",X"FF",X"D9",X"7F",X"24",X"00",X"24",X"08",X"00",X"40",X"80",X"00",
		X"FF",X"00",X"80",X"40",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",X"F5",X"D9",X"B0",X"7F",X"4E",X"24",
		X"09",X"00",X"09",X"24",X"4E",X"10",X"7F",X"C5",X"EC",X"E7",X"BF",X"8D",X"6D",X"6A",X"7F",X"94",
		X"92",X"71",X"40",X"17",X"12",X"39",X"10",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"48",X"8A",X"95",X"A0",X"AB",X"B5",X"BF",X"C8",X"D1",
		X"DA",X"E1",X"E8",X"EE",X"F3",X"F7",X"FB",X"FD",X"FE",X"FF",X"FE",X"FD",X"FB",X"F7",X"F3",X"EE",
		X"E8",X"E1",X"DA",X"D1",X"C8",X"BF",X"B5",X"AB",X"A0",X"95",X"8A",X"7F",X"75",X"6A",X"5F",X"54",
		X"4A",X"40",X"37",X"2E",X"25",X"1E",X"17",X"11",X"0C",X"08",X"04",X"02",X"01",X"00",X"01",X"02",
		X"04",X"08",X"0C",X"11",X"17",X"1E",X"25",X"2E",X"37",X"40",X"4A",X"54",X"5F",X"6A",X"75",X"7F",
		X"10",X"59",X"7B",X"98",X"AC",X"B3",X"AC",X"98",X"7B",X"59",X"37",X"19",X"06",X"00",X"06",X"19",
		X"37",X"08",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"76",X"FF",X"B8",X"D0",X"9D",
		X"E6",X"6A",X"82",X"76",X"EA",X"81",X"86",X"4E",X"9C",X"32",X"63",X"10",X"00",X"F4",X"00",X"E8",
		X"00",X"DC",X"00",X"E2",X"00",X"DC",X"00",X"E8",X"00",X"F4",X"00",X"00",X"48",X"45",X"4B",X"50",
		X"56",X"5B",X"60",X"64",X"69",X"6D",X"71",X"74",X"77",X"7A",X"7C",X"7E",X"7F",X"7F",X"80",X"7F",
		X"7F",X"7E",X"7C",X"7A",X"77",X"74",X"71",X"6D",X"69",X"64",X"60",X"5B",X"56",X"50",X"4B",X"45",
		X"40",X"3B",X"35",X"30",X"2A",X"25",X"20",X"1C",X"17",X"13",X"0F",X"0C",X"09",X"06",X"04",X"02",
		X"01",X"01",X"00",X"01",X"01",X"02",X"04",X"06",X"09",X"0C",X"0F",X"13",X"17",X"1C",X"20",X"25",
		X"2A",X"30",X"35",X"3B",X"40",X"81",X"24",X"00",X"00",X"00",X"16",X"31",X"12",X"05",X"1A",X"FF",
		X"00",X"27",X"6D",X"11",X"05",X"11",X"01",X"0F",X"01",X"47",X"11",X"31",X"00",X"01",X"00",X"0D",
		X"1B",X"F4",X"12",X"00",X"00",X"00",X"14",X"47",X"41",X"45",X"00",X"00",X"00",X"0F",X"5B",X"21",
		X"35",X"11",X"FF",X"00",X"0D",X"1B",X"15",X"00",X"00",X"FD",X"00",X"01",X"69",X"31",X"11",X"00",
		X"01",X"00",X"03",X"6A",X"01",X"15",X"01",X"01",X"01",X"01",X"47",X"F6",X"53",X"03",X"00",X"02",
		X"06",X"94",X"6A",X"10",X"02",X"00",X"02",X"06",X"9A",X"1F",X"12",X"00",X"FF",X"10",X"04",X"69",
		X"31",X"11",X"00",X"FF",X"00",X"0D",X"00",X"12",X"06",X"00",X"FF",X"01",X"09",X"28",X"14",X"17",
		X"00",X"00",X"00",X"0E",X"0D",X"F4",X"11",X"00",X"00",X"00",X"0E",X"0D",X"21",X"30",X"00",X"01",
		X"00",X"0D",X"1B",X"13",X"10",X"00",X"FF",X"00",X"09",X"A4",X"F4",X"18",X"00",X"00",X"00",X"12",
		X"B3",X"82",X"22",X"00",X"00",X"00",X"18",X"C6",X"F2",X"19",X"00",X"00",X"00",X"16",X"DF",X"21",
		X"30",X"00",X"FF",X"00",X"1B",X"0D",X"F1",X"19",X"00",X"00",X"00",X"0E",X"A4",X"31",X"19",X"00",
		X"01",X"00",X"03",X"6A",X"41",X"02",X"D0",X"00",X"00",X"27",X"6D",X"03",X"15",X"11",X"FF",X"00",
		X"0D",X"1B",X"A0",X"98",X"90",X"88",X"80",X"78",X"70",X"68",X"60",X"58",X"50",X"44",X"40",X"01",
		X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"10",X"30",X"60",X"C0",X"E0",X"01",X"01",X"02",
		X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0C",X"80",X"7C",X"78",X"74",X"70",X"74",
		X"78",X"7C",X"80",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"20",X"28",X"30",X"38",
		X"40",X"48",X"50",X"60",X"70",X"80",X"A0",X"B0",X"C0",X"08",X"40",X"08",X"40",X"08",X"40",X"08",
		X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"01",X"02",X"04",
		X"08",X"09",X"0A",X"0B",X"0C",X"0E",X"0F",X"10",X"12",X"14",X"16",X"40",X"10",X"08",X"01",X"01",
		X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"06",X"08",X"0A",X"0C",X"10",X"14",
		X"18",X"20",X"30",X"40",X"50",X"40",X"30",X"20",X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",X"04",
		X"03",X"02",X"02",X"01",X"01",X"01",X"07",X"08",X"09",X"0A",X"0C",X"08",X"17",X"18",X"19",X"1A",
		X"1B",X"1C",X"00",X"00",X"00",X"00",X"08",X"80",X"10",X"78",X"18",X"70",X"20",X"60",X"28",X"58",
		X"30",X"50",X"40",X"48",X"00",X"01",X"08",X"10",X"01",X"08",X"10",X"01",X"08",X"10",X"01",X"08",
		X"10",X"01",X"08",X"10",X"01",X"08",X"10",X"00",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",
		X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",X"10",X"20",X"40",
		X"00",X"01",X"40",X"02",X"42",X"03",X"43",X"04",X"44",X"05",X"45",X"06",X"46",X"07",X"47",X"08",
		X"48",X"09",X"49",X"0A",X"4A",X"0B",X"4B",X"00",X"FB",X"11",X"F0",X"1D",X"FB",X"A0",X"F0",X"1D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
