-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "3FFFFFF8000305FFFFFEFA02FFFFFFFFFFFF0AA0FC7F0BFFFFFFFFA8FE00F000";
    attribute INIT_01 of inst : label is "FFFFFFE8FFFF0FFFBFFF02BF1FFFFFF8FD7CFE805500FC00E3FF02FFFFFFFEFF";
    attribute INIT_02 of inst : label is "00003FFD800000008400F000E17FFFFF3FFFFFFED000FF00FFFFFFFF3FFF0AFF";
    attribute INIT_03 of inst : label is "01FF0FFFA800FF00FFFCA000FFF0FFCF000F003FFFC0FFC0003F15FFC0000000";
    attribute INIT_04 of inst : label is "FCFFF3FFFFFFCFFF0C7460D5FFBFFF3FFFFFFCFFFF3FFFFF0BE003C000000000";
    attribute INIT_05 of inst : label is "01600000000002809999999900000160F7FFFFFFFCFFFEBFFFEFFFCFDBEFFCF3";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "10C407D0FCFFFEFFFCFFFFFFFFCFFFCFFF3FFFE7FFFFDFFF2D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280AC6832558";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "9D00999DFCFFFFDFFFCFFFF6FCCFFFCFFFFCFFF701F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "000057FD000007FD3FFF02AA7FFF02AAFFEDA000FFE0A0000700FF000050FF00";
    attribute INIT_0D of inst : label is "00D000FF050000FF7BFF000A0BFF000AFFFCAA80FFFDAA8000007FD500007FD0";
    attribute INIT_0E of inst : label is "0802000E8020000857FFFEA0FFF4EAFEFFD50ABF1FFFBFAB8020B00008022000";
    attribute INIT_0F of inst : label is "6AA90AEA6AA90AEA02FEAA8001FCAE80BF8002AA3F4002BA6AA9ABA06AA9ABA0";
    attribute INIT_10 of inst : label is "E03900030B99000B99E0E000B9B9020204AC95563A1095563FA02FE00AFC0BF8";
    attribute INIT_11 of inst : label is "0015E2990000007E0FF8FFC0EF7F0A88AFAFA288FDFB22A02FF003FF0000BD00";
    attribute INIT_12 of inst : label is "99998000999900089980999000991999000001FF0FFF00AAFFF0AA000000FF40";
    attribute INIT_13 of inst : label is "9990999899909980019919990999019990199999999980009991999911999999";
    attribute INIT_14 of inst : label is "9009DFFFFE79E7999BFD000202DF199B9009FFFD99BD999BBF7F9BF3F999FFFD";
    attribute INIT_15 of inst : label is "5400668B555511BBCF80FFC002F303FF0079799979999999999F9FBFF7809990";
    attribute INIT_16 of inst : label is "B9999999999B9999FFFD999B999B8000FFFD000A9999FFFD9BFF0002FFFDFFFF";
    attribute INIT_17 of inst : label is "00000000DFFFA000B9990008F7998000DFFFFFFFFF9999999999DFFFDFFFB999";
    attribute INIT_18 of inst : label is "00007FFD00000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "FFFFFF00007F7FFFFD00FFFDFFFFFFFF00000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FBE7CF3FFD00FFFDFF40FDBDC000F400FFFCFFF7007F7BF801FF7FFF0003001F";
    attribute INIT_1B of inst : label is "9F909980119F99FFFF998000009F1FEFFE97F999FA998000FF3FFEBFFBFFF3FF";
    attribute INIT_1C of inst : label is "00005FFF5F80800002F500020000FFF502DF0002F900FFFD2F7F02F3002D0002";
    attribute INIT_1D of inst : label is "000F00020BEF003DC00000001F80F80078008000FE78E780007F7FBFF7808000";
    attribute INIT_1E of inst : label is "99E0E0000B99000BFFFA07FFFFF3E85F01FF7FF83CFFE02FFF5F0BFFFFF0FFC0";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000FFFFFFFF00000000999999999D00999D0000000000000000";
    attribute INIT_20 of inst : label is "0FFF01FF000000AAFFF0FF400000AA0000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0FFA01FE000000AA73F07F400000AA000FFF01FE000000AAFFF07F400000AA00";
    attribute INIT_22 of inst : label is "4F5F00F7020400AAFFF0D0190000AB6A0FFA01EE000800AA73F000428004AA00";
    attribute INIT_23 of inst : label is "DBF019000000091F3F9C01900000D1802BFFD3FF0100BD1EF40180311C00EB1D";
    attribute INIT_24 of inst : label is "00B45557BE03017E7D73FED8C000AA800FFF1BAA0005E22FFFC0AB904000E22C";
    attribute INIT_25 of inst : label is "2FFED38B003D00BDCFC0FF800000DE001FDF007F000FA0BEFFC05F8000705A00";
    attribute INIT_26 of inst : label is "000B000000000000FFFF1F60007F000A03FF2FFF300F000AFFC0FFF8F00CA000";
    attribute INIT_27 of inst : label is "000F02FF01000000FFFFDF60007F002A007E000000000000A7FF7FD501FF0000";
    attribute INIT_28 of inst : label is "7FFA1FFF00052AAAAAA8AFAD5000A80001F8001F000000000BFFFFFF07AF0000";
    attribute INIT_29 of inst : label is "FFFF000000002FFFFFFF00010000FFF8001FFDBF40010000FFC0FF7F40010000";
    attribute INIT_2A of inst : label is "0FFF28F9FFFF00A8FFF8CF900000E800087FFF800FFF3FE8FABCE540FC002FFA";
    attribute INIT_2B of inst : label is "16E917E607EF02A8FFD0FFE0F6D0A0002FFE3FFF1FFF00BDDE34AA00FFC02AFD";
    attribute INIT_2C of inst : label is "00000BF535740000002F5550000000002BC01FFF000000009556FFD000000000";
    attribute INIT_2D of inst : label is "955607FF00000000FC00F00000000000003F000F000000009556FFD000000000";
    attribute INIT_2E of inst : label is "0000F0A000000000002AFFF4000000000000FFFF0000000000000A0A00000000";
    attribute INIT_2F of inst : label is "000000F0000000000000F000000000000000000F000000000000FC0000000000";
    attribute INIT_30 of inst : label is "E7D5FFFF1FFF0000FFC0FFD5FE000000E5D5FFFF1FFF0000FFC0FFD0FE000000";
    attribute INIT_31 of inst : label is "0FFFF7FFD1FF000BFFF0FFDFFF47E000CFD5FFFF47FF000057F3FFFFFFD10000";
    attribute INIT_32 of inst : label is "3FFF01FD0000F800E3FF7FD507FF0000A0027FFF00500000A3FFFFD007FF0000";
    attribute INIT_33 of inst : label is "FFFE00570000A000B3FFFFFF043F001F00000BFFFFF40000B3FFFFFF043F001F";
    attribute INIT_34 of inst : label is "FFC0FFD5FE0080000000000000000000FFC0FFD0FE0080000000000000000000";
    attribute INIT_35 of inst : label is "FFFA07FF00000000A7FFFFFF1FFF002A00AF3FFFFD400000E7FFFFFF1FFF000A";
    attribute INIT_36 of inst : label is "F3FFFFD007FF0000FFC007FFFC170000F3FFFFD002FF0000FFCB07FFFAD00000";
    attribute INIT_37 of inst : label is "3FFF01FD0909F800E3FF77D503EF000000022FFFFF500000A3FFFFD007FF0000";
    attribute INIT_38 of inst : label is "7FFA1FFF00052AAAAAA8AFAD5000A8003FFA1FFF00055FAAAAA8FAF85000A800";
    attribute INIT_39 of inst : label is "0BFF3FFF07FF001FFFE0FFFCFFD0A0002FFFFFFF1FFF097EFFF8FFFFFFF48000";
    attribute INIT_3A of inst : label is "7FFF1FFD00050AAAEAA8A5A45000A8003FEB1FFD0005B02AEBE8A5A45000A800";
    attribute INIT_3B of inst : label is "3DFF3C7C073C0BEAFF003FC03C0080002E7F3E7C067CBFAAFF003FC03C008000";
    attribute INIT_3C of inst : label is "3A8D000000002A880CE90000000008A80300030003AA000000300030AAB00000";
    attribute INIT_3D of inst : label is "3FAA1FFF00052AAAAAA8FAF85000A8003F541FFF005F2AAA0000F5F4FD50AA80";
    attribute INIT_3E of inst : label is "3FCF3D0130002DAAFFC0FFFC3FF080003F473C0030002DAAFFF87FFF07FFA000";
    attribute INIT_3F of inst : label is "3F3F3F3F073F2DAAFFE0FFF0FF40A0003FCF3F071C032DAAFFC0FFF0FFC08000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "3FFF7FFF0000001FFFFFFFF81FF4FFFF1FF4BFFEFF1FE1FFFFFFFFFFFF00FC00";
    attribute INIT_01 of inst : label is "1FFFFFFEF5FFFFFFFFF42FFF017F7FFFFC0CFFF80000FE00F1FFCFFFF540FFFF";
    attribute INIT_02 of inst : label is "00000150C0000000FFA0F800FFA15FFF0FFF7FFF0000FC00FF54FFFF05FF3FFF";
    attribute INIT_03 of inst : label is "00FF03FFFF00D4007FFFFFA0FFFCFFE30003001FFFC0FFC02AFF003FE0000000";
    attribute INIT_04 of inst : label is "FFFFFCFFFFFFFFFF2C060616FFFFFF3FFFFFFCFFFFCFFF7F07D0028000000000";
    attribute INIT_05 of inst : label is "03F0000000000140BBBB9999000003F0F3FFFFFFFF3FE7FBFFF3FFDFFFBFF7DF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "01000BD8FCFFFDFFFCFFFFFFFFCFFFCFFFE7FDF9CFFFFFFF1EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF1AA4C943";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "FAAA99D0FFFDFFBFFFEFFFF3FCFFFFCFFFFEFFFD2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "0000007F0000007F3FFF2FFF3FFFAFFFFFD0FF00FFD5FF000000FF000000FFC0";
    attribute INIT_0D of inst : label is "000000FF000003FF07FF00FF57FF00FFFFFCFFF8FFFCFFFA0000FD000000FD00";
    attribute INIT_0E of inst : label is "0505000150520005007DFFFED500FFFD7D00BFFF00577FFF5050400085055000";
    attribute INIT_0F of inst : label is "30302FFD0C0C2FFD017457FC00005FA01D403FD500000AF50C0C7FF830307FF8";
    attribute INIT_10 of inst : label is "9ED9000DB99900B9999E9E00EFEF989807F41D5C1FD0357405403FC0015003FC";
    attribute INIT_11 of inst : label is "00006F9B0000000501A83000019019370451A6D10640DC642A40000C00005000";
    attribute INIT_12 of inst : label is "999999889999899999989900099901990000001F07FF0BFFFFD0FFE00000F400";
    attribute INIT_13 of inst : label is "9980999099989980019909991999099900019999999998091000999900019999";
    attribute INIT_14 of inst : label is "0001995FFFEFF9F9BD9989BF2DBF003F0001FD1999BC999BBEFF9BCFD999FDD9";
    attribute INIT_15 of inst : label is "0000E6F90000AA00D58070000257000D000707991F99F999999999F9FE78F900";
    attribute INIT_16 of inst : label is "FFB999999BFF9999FD999BFF9BFF9988FD998BFF9999FD99BFFF89BFFD99FFFF";
    attribute INIT_17 of inst : label is "AAAA000099DFFFA8FFB98999FE79F98899DFFFFFFFF9F999999999DF99DFFFB9";
    attribute INIT_18 of inst : label is "AAAA07D000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "FFFFFF00000707FFD000FFD0FFFFFFFF00000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FEFFF7DFD0006FD0FD00FBD04000F000FFFEFFFD000707FF007F07FF0001000F";
    attribute INIT_1B of inst : label is "9BF8B980000199BFFE79F809099901FFF9FE97F9157B9009FCFFEFDBCFFFF7FF";
    attribute INIT_1C of inst : label is "0000005F0058F8002500002F0000F5002DBF002FD000FDD0BEFF0BCF00BC000B";
    attribute INIT_1D of inst : label is "002F0003BD6F00F6F0008000E17AFE001E00E000FFEEF9E0000707F9FE78F800";
    attribute INIT_1E of inst : label is "BBBE9E00BBBB00B95FFFEA17FFD3FFE000051FFF14FFFCFFFD073FFFFF40FFE0";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000FFFFFFFF0000000099999999D00099D00000000000000000";
    attribute INIT_20 of inst : label is "07FF001F00000BFFFFD0F4000000FFE000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "07F7001E00000BDF6FD074000000FDE007F7001E00000BFFFFD074000000FFE0";
    attribute INIT_22 of inst : label is "D42F913D00000BDEFFD2000000007DE407F7001E00010BDF01D0001A0480FDE0";
    attribute INIT_23 of inst : label is "2FC001800000BB390FE009000000B3B8FFFF086F00009B3B403EE0020180FF4B";
    attribute INIT_24 of inst : label is "2BFE0A137D03000BFF4FF5000000FFF83FFF01FF00007FFFFFF0FD000000FFF4";
    attribute INIT_25 of inst : label is "FFDF407F003403FDFF4045F800008980038B003F0003FFFEFF4003C00000EF00";
    attribute INIT_26 of inst : label is "00BF0000000000007FF507AF0000AB3B0FFF3CFF100000BFFFF0FF3C0004FE00";
    attribute INIT_27 of inst : label is "003F03D000000000FFF507AF00002BFF001F000000000080FEFF0F1F001502BF";
    attribute INIT_28 of inst : label is "3FFF01FF0000FFFF5F5EFF500000FFE8007F000000000200F9FF5F6A007F002A";
    attribute INIT_29 of inst : label is "C7F500000000FFFF5FD300000000FFFF0B39D01F0000003FFFF8F4070000FC00";
    attribute INIT_2A of inst : label is "07FFFFFE1FF40BF3FD7C500000003F803F5F7FFF01FF7FFFDCB4A800D000FFD4";
    attribute INIT_2B of inst : label is "3FFF0A7F00152F7F3DB5FE7C50009FE03FFF3FFF017F03F3E540FFC0FD00FF68";
    attribute INIT_2C of inst : label is "02B89556101000002FFD0000000000003FEA017F00000000BFF4FD0000000C0C";
    attribute INIT_2D of inst : label is "1FF7001500003030F400F00000000000001F000F00000000DFF4540000000C0C";
    attribute INIT_2E of inst : label is "00000051000000002FFF550000000000FFAA17FF00000000A800ED0500000000";
    attribute INIT_2F of inst : label is "00000000000000001000A00000000000000F000F00000000FC00500000000000";
    attribute INIT_30 of inst : label is "FEBF3FFF017F2ABFFFF0FD55F400FA00FFBF3FFF017F2ABFFFFAFD5AF400FA00";
    attribute INIT_31 of inst : label is "BFFFF3FF402F083FFFFEFFCFF801FC20FF1FFFFF005F02BFF4FFFFFFF500FE80";
    attribute INIT_32 of inst : label is "1FFF00000000FFA0FEFF0F1F007F00BFFEBF1FFF00000000FEFF4F1A007F00BF";
    attribute INIT_33 of inst : label is "1FFF00000000FF80FBFF0FFF00070AFF00AF3FFFF5000000FBFF4FFF00070AFF";
    attribute INIT_34 of inst : label is "FFF0FD55F400FE000000000000000000FFFAFD5AF400FE000000000000000000";
    attribute INIT_35 of inst : label is "FFFF00050000FA00FEFF3FFF017F2AFF0FFFFFFDD0000000FFFF7FFF017F2ABF";
    attribute INIT_36 of inst : label is "FEFF4C3A127F80BFFFBFAFFFFD02FE00FEFF05FA007FE0BFFFBFA5F7FD00FE00";
    attribute INIT_37 of inst : label is "1FFF00000080FFA0FEFF0C3FB07F00BF02BFFFFFD0000000FEFF4F1A007F00BF";
    attribute INIT_38 of inst : label is "3FFF01FF0000FFFF5F5EFF500000FFE83FFF01FF00000FFFF5F4FF500000FFE8";
    attribute INIT_39 of inst : label is "2FFF1FFF010500AFFFF8FFF45040FA00BFFF7FFF010500AFFFFEFFFD5040FA00";
    attribute INIT_3A of inst : label is "3FFE01FF0000BFD55A58FF5000005FE83FFE01FF00007F7D5A58FF5000007D68";
    attribute INIT_3B of inst : label is "3CF71F3301113FFFDFC0CF004000F8003DB71DB301110FFFDFC0CF004000F800";
    attribute INIT_3C of inst : label is "0000000000003A0C0000000000009CC303000300000002AA003000300000AAA0";
    attribute INIT_3D of inst : label is "3FFF01FF0000DFFFF5F4FF500000FFE83FFF07FF0000DFFFEAA8FAF80000FD54";
    attribute INIT_3E of inst : label is "3F033C0000003FFFFFF0FC341410FE003D01300000003FDFFFFE1FC30141FF80";
    attribute INIT_3F of inst : label is "3F3F1F3C01143FFFFFF03FD01400FF803F4F3D0304013FFFFFF0C3D04100FE00";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "3FFFFFF8000305FFFFFEFA02FF4BFFFFFFDF0AA0FC7F0BFFFFFFFFA8FE00F000";
    attribute INIT_01 of inst : label is "FFFFFFE85FFF0FFFBFFF02BF1FFFFFF8FD7CFE805500DC00E3FF02FFFFFFFEFF";
    attribute INIT_02 of inst : label is "00003FFD800000008400F000E17FFFFF3FFFFFFED000DF00FD52FFFF3FFF0AFF";
    attribute INIT_03 of inst : label is "01FF0FFFA8004B00FFFCA000FFF0FFCF000F003FFFC0FFC0003F15FFC0000000";
    attribute INIT_04 of inst : label is "FCFFF3FFFFFFCFFF0C7460D5FFBFFF3FFFFFFCFFFF3FFFFF0BE003C000000000";
    attribute INIT_05 of inst : label is "01600000000002800000000000000160F7FFFFFFFCFFFEBFFFEFFFCFDBEFFCF3";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "FFFF07D0FCFFFEFFFCFFFFFFFFCFFFCFFF3FFFE7FFFFDFFF2D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280AC6832558";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "00000000FCFFFFDFFFCFFFF6FCCFFFCFFFFCFFF701F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "000002AD000007FD3D0002AA000002AA3FC0A0003FC0A0000000FD000000FD00";
    attribute INIT_0D of inst : label is "0000007F0000007F03FC000A03FC000A007CAA800000AA8000007A8000007FD0";
    attribute INIT_0E of inst : label is "3DF72A84DF7F000800004000000040000000000100000001DF7C12A8FDF72000";
    attribute INIT_0F of inst : label is "EAABD840EAABD840F402001FF80004FF801FF400002FFF10EAAB0127EAAB0127";
    attribute INIT_10 of inst : label is "000000000000000000000000B9B90202AD04D557107AD557003F402FFC00F801";
    attribute INIT_11 of inst : label is "0000F7990000001F0150154044DC01FFF7D7F7DF3711FF40054001540000F400";
    attribute INIT_12 of inst : label is "00005FFF0000FFF5007F000BFD00E0000000001F03FF0000FFC000000000F400";
    attribute INIT_13 of inst : label is "002F0003000F003FF800C000F000FC000BE0000000007FFD002A0000A8000000";
    attribute INIT_14 of inst : label is "0FF05FFFFE78E78002F5FFF7FFDFE0020FF0FFF5002D00022F7F02F3F000FFF4";
    attribute INIT_15 of inst : label is "000066DF0055991129001540006801540000000078008000001F1FBFF7FF800B";
    attribute INIT_16 of inst : label is "A0000000000A0000FFF5000A000A5FFFFFF5FFFF0000FFF502FFFFF7FFF5FFFF";
    attribute INIT_17 of inst : label is "000000005FFFFFFFA000FFF5F780DFFF5FFFFFFFFF80800000005FFF5FFFA000";
    attribute INIT_18 of inst : label is "0000000000007FFD002A0000A800000000005FFF0000FFF5007F000BFD00E000";
    attribute INIT_19 of inst : label is "FFFFFF00007F7FFFFD00FFFDFF808000002F0003000F003FF800C000F000FC00";
    attribute INIT_1A of inst : label is "FBE7CF3FFD00FFFDFF40FDBDC000F400FFFCFFF7007F7BF801FF7FFF0003001F";
    attribute INIT_1B of inst : label is "0F8F803FA80F00FFFFC0FFFDFF5FFFEFFE97E800FB407FFDFF3FFEBFFBFFF3FF";
    attribute INIT_1C of inst : label is "0FF05FFF5F80DFFF02F5FFF70FF0FFF5FFDFE002F900FFFD2F7F02F3002D0002";
    attribute INIT_1D of inst : label is "000F00020BEF003DC00000001F80F80078008000FE78E780007F7FBFF7FF800B";
    attribute INIT_1E of inst : label is "0000000000000000FFFA07FFFFF3E85F01FF7FF83CFFE02FFF5F0BFFF4F0FFC0";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFF000000000000000000000000000000000B99000B99E0E000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "00A7353700000000FC00FFC017C0000000000001000000000000FE0000000000";
    attribute INIT_23 of inst : label is "0BFF1BFF001F03FFFF80FF90D000FF0003FF03F8000000004BC07FC003C00000";
    attribute INIT_24 of inst : label is "003F000100000000E3FF7FFC027602800BFF1B55000503FFFF8057904000FF00";
    attribute INIT_25 of inst : label is "000303FF000000BFFFC050000000FEE400AA0074000000BFFFC600000000FF20";
    attribute INIT_26 of inst : label is "000B000000000000FFFA099F007F02E003FF03FF003F000AFFC0FFC0FC00A000";
    attribute INIT_27 of inst : label is "000F02F500000000FFFA499F007F1B90001E000000000000AFE0176A00BF1B00";
    attribute INIT_28 of inst : label is "3FFF1FFF0005002AFFFCD2D05000A80000780005000000000B80FFD5007F2200";
    attribute INIT_29 of inst : label is "15FF00C010C12FFFFF5403004304FFF802E03DFF0000000000C0FF7C00001750";
    attribute INIT_2A of inst : label is "0FA82838F06F00205E92FAC00000200007EA0F80005F5540854BF540D40005FA";
    attribute INIT_2B of inst : label is "091600190010000000000000010000000C610F55015F0036F5D0AA005000D1D4";
    attribute INIT_2C of inst : label is "00000BF50A0A0000002F5550000000002BC01FFF000000002AA8FFD000000000";
    attribute INIT_2D of inst : label is "2AA807FF00000000FC00F00000000000003F000F00000000AAA8FFD000000000";
    attribute INIT_2E of inst : label is "0000FFFF00000000000000000000000000000000000000000000FFFF00000000";
    attribute INIT_2F of inst : label is "000000FF000000000000F0000000000000000000000000000000030000000000";
    attribute INIT_30 of inst : label is "3FFF3FD61FFF0017E000BF40E14056007FFF155A1FFF0AD5E000BF40E1401FA0";
    attribute INIT_31 of inst : label is "082F3FFF11FF05D4F820FFFCFF4417500F6A382F07FF05D4A9F0F82CFFD01750";
    attribute INIT_32 of inst : label is "0FFF005400003800EBF8166A002F6C0020021FFF00000000EBF8D66F002F6000";
    attribute INIT_33 of inst : label is "3FFE000100002001BFFF5FFF03EF5D1F00000BFF3F500003BFFF5FFF03EFF81F";
    attribute INIT_34 of inst : label is "E000FF40E14000000000000000000000E000FF40E14000000000000000000000";
    attribute INIT_35 of inst : label is "3FFA015F00000002BFFF557F1FFFFA8000AF3FFF34000001FFFFF55B1FFFFA00";
    attribute INIT_36 of inst : label is "3BF816FF002FAE002FC0FFFCFBC417503BF816FF052F09D42FE8FF9CFD002750";
    attribute INIT_37 of inst : label is "00000000000000000800082A04106C0000022FFF35000000EBF8D66F002F6000";
    attribute INIT_38 of inst : label is "3FFF1FFF0005002AFFFCD2D05000A8003FFF1FFF0005002AFFFC87855000A800";
    attribute INIT_39 of inst : label is "0BFF3FFF05070000FFE0FFFCD05000002FFFFFFF1D070000FFF8FFFFD0740000";
    attribute INIT_3A of inst : label is "300018020005002A155C5A5C5000A800301418020005002A141C5A5C5000A800";
    attribute INIT_3B of inst : label is "2600338306C300AA0300C0C0CC00800025803183078302AA0300C0C0CC008000";
    attribute INIT_3C of inst : label is "3A8D000000002A880CE90000000008A80300030003AA000000300030AAB00000";
    attribute INIT_3D of inst : label is "3FFF1FFF0005002AFFFC87855000A8003F541FFF005F002A00004B4AFD50AA80";
    attribute INIT_3E of inst : label is "2FCF3D01300000AAFFC0F41C341080002F473C00300000AAFFF87F410741A000";
    attribute INIT_3F of inst : label is "2FFF3FF407F400AAFFE01FF01F40A0002FCF3F071C0300AAFFC041F041C08000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "3FFF7FFF0000001FFFFFFFF81FB4FFFB1EB4BFFEFF1FE1FFFFFFFFFFFF00FC00";
    attribute INIT_01 of inst : label is "1FFFFFFEF5FFFFFFFFF42FFF017A7FFFCC0CFFF800002E00F1FFCFFFF540FFF4";
    attribute INIT_02 of inst : label is "00000150C0000000FFA0F800FFA15FFF0FFF7FFF0000AC00EA54FFFF05FF3FFF";
    attribute INIT_03 of inst : label is "00FF03FFFF00D4007FFFFFA0FFFCFFE30003001FF6C0FFC02AFF003FE0000000";
    attribute INIT_04 of inst : label is "FFFFFCFFFFFFFFFF2C060616FFFFFF3FFFFFFCFFFFCFFF7F07D0028000000000";
    attribute INIT_05 of inst : label is "03F0000000000140AAAA0000000003F0F3FFFFFFFF3FE7FBFFF3FFDFFFBFF7DF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "1FF4BFFFFCFFFDFFFCFFFFFFFFCFFFCFFFE7FDF9CFFFFFFF1EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF1AA4C943";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "AAAA0000FFFDFFBFFFEFFFF3FCFFFFCFFFFEFFFD2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "0000007F0000007F10022FFD3A022FFDFF007F00FF007F000000D0000000D000";
    attribute INIT_0D of inst : label is "000000070000000700FF00FD00FF00FD80047FF880AC7FF80000FD000000FD00";
    attribute INIT_0E of inst : label is "0555FFFE5FFDBFEA000000000000000000000000000000005550BFFF7FF5ABFE";
    attribute INIT_0F of inst : label is "F0F0EAA80F0FEAA8F8220005FFAB0037882F5000EAFFDC000F0F2AABF0F02AAB";
    attribute INIT_10 of inst : label is "000000000000000000000000EFEF9898F4025F5D801F75F5E00F00AFF00BFA00";
    attribute INIT_11 of inst : label is "0000065F0000000000AE0AE0AB10B3390410B59A04EA6CCEBA000BA000000000";
    attribute INIT_12 of inst : label is "0000001500005400000700BFD000FE000000000000FF00BFFF00FE0000000000";
    attribute INIT_13 of inst : label is "003F000F0003001FFC00F000C000F400BFFE0000000007D0AFFF0000FFFA0000";
    attribute INIT_14 of inst : label is "BFFE02DFFFEEF9E02500542FFDBFFFAFBFFEF78000BC000BBEFF0BCF4000FD40";
    attribute INIT_15 of inst : label is "0000F5900000FFAAFE00CA0000BF00A3000000001E00E000000101F9FE7FFAFF";
    attribute INIT_16 of inst : label is "FFA000000AFF0000F5000AFF0AFF0015F5005EFF0000F5002FFF542FF500FFFF";
    attribute INIT_17 of inst : label is "AAAA0000005FFFB5FFA05400FE78F815005FFFFFFFF8F8000000005F005FFFA0";
    attribute INIT_18 of inst : label is "AAAA0000000007D0AFFF0000FFFA00000000001500005400000700BFD000FE00";
    attribute INIT_19 of inst : label is "FFFFFF00000707FFD000FFD0FFF8F800003F000F0003001FFC00F000C000F400";
    attribute INIT_1A of inst : label is "FEFFF7DFD0006FD0FD00FBD04000F000FFFEFFFD000707FF007F07FF0001000F";
    attribute INIT_1B of inst : label is "03FB381FFFFB003FFE78FFF0D001FFFFF9FE97E8157A0FF0FCFFEFDBCFFFF7FF";
    attribute INIT_1C of inst : label is "BFFE02DF0058F8152500542FBFFEF780FDBFFFAFD000FDD0BEFF0BCF00BC000B";
    attribute INIT_1D of inst : label is "002F0003BD6F00F6F0008000E17AFE001E00E000FFEEF9E0000707F9FE7FFAFF";
    attribute INIT_1E of inst : label is "AAAA0000AAAA00005FFFEA17FFD3FFE000051FFF14FFFCFFFD073FFFAB40FEE0";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFF00000000000000000000000000000000B99900B9999E9E00";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0BFF000700000000FB00FFC0004000000000000100000000FE005F0000000000";
    attribute INIT_23 of inst : label is "2FFF01FF000707FFFFE0FD004000FF4003FD006F0000033ABFC01FC00040A880";
    attribute INIT_24 of inst : label is "001F00000000000AFFFF0530011100F83FD501FA000003FF5FF0BD000000FF00";
    attribute INIT_25 of inst : label is "00AA00740000011FFF4000000000FF8503FF00000000001FFF4000000000FFB5";
    attribute INIT_26 of inst : label is "00140000000000001FDA007A0000AEC403FF00FF027600BFFFC0FF009D80FE00";
    attribute INIT_27 of inst : label is "003F010000000000FFDA007A00002A800005000000000000FFFF04EA00151240";
    attribute INIT_28 of inst : label is "3FFF01FF00000BFFE1E0FF500000FFE8001F000000000000FFFA0995007F2580";
    attribute INIT_29 of inst : label is "000009D800003FFF000027600000FFFC2FE61000000000800BF8000400000300";
    attribute INIT_2A of inst : label is "01FFF5CE1EF40ACEEAA550000000C5000F5D07FF000017FAF750A8000000B520";
    attribute INIT_2B of inst : label is "0000018000000080C24001800000600007BC07EB000000CCF540FF400000A59F";
    attribute INIT_2C of inst : label is "02B82AA8050500002FFD0000000000003FC001550000000002A055000000F0F0";
    attribute INIT_2D of inst : label is "0AA3001500000F0FF400500000000000001F000500000000CAA054000000F0F0";
    attribute INIT_2E of inst : label is "2FF81FD4000000000000000000000000002A002A00000000ABFEBFF500000000";
    attribute INIT_2F of inst : label is "00BF001500000000E000F000000000000000000A000000000200040000000000";
    attribute INIT_30 of inst : label is "3FFF2ABF017F2800FFA0D2C0F40000003FFF3FFF017F3840FFF0D2C0F4000414";
    attribute INIT_31 of inst : label is "2FFF3FFF002F03DFFFF8FFFCF800F7C034EA1FFF005F02EAAB1CFFF4F500AB80";
    attribute INIT_32 of inst : label is "07FF000000003FA1FFFF04EA007F41403EBF05F500000001FFF504E5007F7540";
    attribute INIT_33 of inst : label is "05FF000000003F80FFFF041F00000BFF00AF3FFD10000000FFFF041F00000BFF";
    attribute INIT_34 of inst : label is "FFA0D2C0F40000000000000000000000FFF0D2C0F40000000000000000000000";
    attribute INIT_35 of inst : label is "1FFF000000003A01FFFF3FFF017F28000FFF7FD400000001FFFF2FFF017F6840";
    attribute INIT_36 of inst : label is "3FF507D5007F24405FFC541CFD0001003FF50E15007F20405FFC5E10FD000100";
    attribute INIT_37 of inst : label is "0000000000000001010003C00000414002BF3FF500000001FFF504E5007F7540";
    attribute INIT_38 of inst : label is "3FFF01FF00000BFFE1E0FF500000FFE83FFF01FF00000BFF4B4AFF500000FFE8";
    attribute INIT_39 of inst : label is "2FFF1FFF00F100AAFFF8FFF44F00AA00BFFF7FFF00F100AAFFFEFFFD4F00AA00";
    attribute INIT_3A of inst : label is "300101A00000096AA5AC0A500000A168300101A0000025C2A5AC0A50000083E8";
    attribute INIT_3B of inst : label is "330818CC0155090020C033005000180032481A4C01550C0020C0330050001800";
    attribute INIT_3C of inst : label is "0000000000003A0C0000000000009CC303000300000002AA003000300000AAA0";
    attribute INIT_3D of inst : label is "3FFF01FF00000BFF4B4AFF500000FFE83FFF07FF00000BFFEAA887850000FD54";
    attribute INIT_3E of inst : label is "3F033C0000000BFFFFF0FBE413C0FE003D01300000000BDFFFFE1FBE013CFF80";
    attribute INIT_3F of inst : label is "3FFF1FFB01530BFFFFF0EFD0C400FF803F4F3D0304010BFFFFF0BED03C00FE00";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
