-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D352A0B57FEA2A4977BB00080082410493A17FFFFFFFFFFF95FEA7A3D3F3EAB5";
    attribute INIT_01 of inst : label is "208B53050688596AA08094500A24F28449614EA8FBF8F2612971B05C07AC02D0";
    attribute INIT_02 of inst : label is "FC616582249E4F061E45A982F79FCB31445F3CC419F84F3C5720898048BC4059";
    attribute INIT_03 of inst : label is "89BE341034499CAFCD9900090F7AFFA7DC55555E004169FDC262E38A88145499";
    attribute INIT_04 of inst : label is "51A089270943A937ABA93780076A8522A211668162D64C1728AB834409386F50";
    attribute INIT_05 of inst : label is "F34F2110D2108910285499B883E2D415122286315425C47E8BC50541075D544E";
    attribute INIT_06 of inst : label is "4250545C518B4B32A602B64FB4BA4DFDB349E496C9BD51493C0A4D0060B24174";
    attribute INIT_07 of inst : label is "829D5134F22CF4224403505499A48FD17E8F9C5A14936A1964B02AA294A2545C";
    attribute INIT_08 of inst : label is "830615560605408A9137523A132887118145084A0E87540824D26D52CB94E216";
    attribute INIT_09 of inst : label is "54CA121CA721674943381D902702F8DED8D5884236118946074DE28A00013802";
    attribute INIT_0A of inst : label is "0124C9D65DF6D4EBED1FB80AFE698E58E7389223582058A08422A43896244542";
    attribute INIT_0B of inst : label is "E5EB397467B396ACE5D199110A51D6846A3DD99A0867819214870E9F122A1D48";
    attribute INIT_0C of inst : label is "6B64AA0978053234FBB84E2BE5E79653807D913E85137D246FA143C79E5651EC";
    attribute INIT_0D of inst : label is "0065F7E9E00041882DCCBD13E898CBF13E89886EA5A11A3AD6B1955958B5A7F2";
    attribute INIT_0E of inst : label is "85B540000000000000000000000000019ADD56D23D4A4ED942BA0284EDB65400";
    attribute INIT_0F of inst : label is "F4A295C73B654AE89C589DB05B731885559263340305B27CBA5FD229C587F434";
    attribute INIT_10 of inst : label is "27D74148A8F2CC20C9353154A479EDB68DB55592F44F98D5564BF13E621BA97F";
    attribute INIT_11 of inst : label is "EF7F119E3768C5EE6CFBDFF11A5D76E27AF816A69B46E37D78F97539621AC572";
    attribute INIT_12 of inst : label is "0B1A0B4450962510C48201547BBC4D10C674809C06DA3A2A108350F7389A30C4";
    attribute INIT_13 of inst : label is "484546A0EB0C9838649E65AF8E3672652C5C8E3CB5E45FD06081452A445AAA44";
    attribute INIT_14 of inst : label is "8D091895221247ACC00000277646438F3932923D6677632000000000002B4C15";
    attribute INIT_15 of inst : label is "8BC8E48A2FFFFEAA720B26212262E221589B4358CA17429C88993C46D35C0290";
    attribute INIT_16 of inst : label is "B3CF40838708A302315814F5635D52D15505BA343741AA2A41A13CB261A14808";
    attribute INIT_17 of inst : label is "A88551C7AA800570B00337378DF741A66D0AF7DBC646754A7661364651397DDF";
    attribute INIT_18 of inst : label is "200C5ADA168B448DC8AA48A4CCE8D70C5F2D812B88F7399A39CD38191D296092";
    attribute INIT_19 of inst : label is "2E7BFF822726DCCCE49B8C3429481842035F702F1FA084C58267E88402377B40";
    attribute INIT_1A of inst : label is "5110028440684A221250C068413619260C34CC01030D25967F30100000C02B02";
    attribute INIT_1B of inst : label is "232032823233520204401354A798668B10FC11028CBAFE9D9A4640029ED2FE3D";
    attribute INIT_1C of inst : label is "0A78EF5A24BC6E930D0D10402032C320EC4A2C458A8D5406EC19E94100801669";
    attribute INIT_1D of inst : label is "00000009C4067FDFF640080036401F003654204404AD120482E8110842108421";
    attribute INIT_1E of inst : label is "4A5569651FF80000049249111100FFEA01FFD65575DD9E6EEBAAAAAA8A222080";
    attribute INIT_1F of inst : label is "0003FB37A040007FF7B7000FF1FFE95CAC5A1681AA680632A8755570AA74D6A1";
    attribute INIT_20 of inst : label is "7BF7A77B4826D648F836A54A89FFCB19E08ED558FD7FC8763CABA0288D3AA281";
    attribute INIT_21 of inst : label is "994F3A2F708DAA1734B67BED3EE806D34DB687E6804B6F41D75BEBD43C25B01E";
    attribute INIT_22 of inst : label is "75537D2090000154D0D151EA3B56A3D92E0B48F8B7CFC9E23418CA7F49226965";
    attribute INIT_23 of inst : label is "EF561C5008ADAA2BEE638E1870A4299A9E2222FDDD71749C679F44EAA312E843";
    attribute INIT_24 of inst : label is "C40C0008CF0481103A36F19EA8A0000D0400680043000019241475242E5E934A";
    attribute INIT_25 of inst : label is "0000000000000000000001E4CDA07F3FDCF4FE196E9E0F6E87C0E8012A3517C6";
    attribute INIT_26 of inst : label is "FFFFFFFFC0000000000000000000EEEEEEEEEE00000000000000000000000000";
    attribute INIT_27 of inst : label is "F0000001FE00A0000060FEE0DFE000A001FFFFFFFE00000001FE1E00000001FF";
    attribute INIT_28 of inst : label is "59EBDE006B36000659CBDE8A6F3E0F4332842493F7AF3A140522A55840007D05";
    attribute INIT_29 of inst : label is "39AD000037EFFA7DDFF60BFF7F0FAFA50BAF0887914F05E1B5E3D420003F0002";
    attribute INIT_2A of inst : label is "22882AD50003E63319980000000F0000000162FD75CE01BB1D2966FC7C642000";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFAAAAFFFAAAAAFFFAAAAAFE0F77B708468F01009124598E6A";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000001FFFFFFFFFF";
    attribute INIT_2D of inst : label is "0000000000000008438F8FD481806C1500000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000DD1808";
    attribute INIT_30 of inst : label is "59EBDE006B36000659CBDE8A6F3E0F4332842493F7AF3A140522A55840007D05";
    attribute INIT_31 of inst : label is "39AD000037EFFA7DDFF60BFF7F0FAFA50BAF0887914F05E1B5E3D420003F0002";
    attribute INIT_32 of inst : label is "22882AD50003E63319980000000F0000000162FD75CE01BB1D2966FC7C642000";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFAAAAFFFAAAAAFFFAAAAAFE0F77B708468F01009124598E6A";
    attribute INIT_34 of inst : label is "000000000000000000000000000000000000000000000000000001FFFFFFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000DD1808";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A480EAC280DD640080260124B2C96C90016CC03FFFFFFFFF93FBCD6603636BD3";
    attribute INIT_01 of inst : label is "6400615610D5FA3944364C9B2D5143EAAE9FE14B6439A52B5A83497D793D67CB";
    attribute INIT_02 of inst : label is "4D17E8104A28E0228F0030ABDF299E420C06520CCA6306502F8402F90022A00C";
    attribute INIT_03 of inst : label is "B2405B74058EE5E27ABF8409216C64CDE49FC6B81224A3F348000735662AF04E";
    attribute INIT_04 of inst : label is "862D9050B4EE2C0110AC013DB6644885AC7A8B00201A855B41300868DB9A0050";
    attribute INIT_05 of inst : label is "27164A2D02D7662005F04E00E8001D59845DB2BCF268AA84B405054100A28A46";
    attribute INIT_06 of inst : label is "D59785D26A004788D4B56DA2404D14D84DB68A05D51B2A1C599832ED0607840D";
    attribute INIT_07 of inst : label is "BCF36A71645925D188005DF04E05549680E63A814A0907F80E06E52FFD2C85D2";
    attribute INIT_08 of inst : label is "B7297DE27F4BA7FBC2D03362683C97B8AB2146E1C8F734BB0E012039C02796AC";
    attribute INIT_09 of inst : label is "AA92C6EB2C7E0B90F0D2B6E47AD45F18A8A47BF426FD0DB5EC1FEBF9E9EB8164";
    attribute INIT_0A of inst : label is "676B85ECA40002F651392CA91EB695AAB0855FA763523926B6B542C70F12AA86";
    attribute INIT_0B of inst : label is "0110004E100004400178452A93EFDF7274A04C435AEFA3FDFBE8C83F23F9F52F";
    attribute INIT_0C of inst : label is "9C9AC883DF781CA74802204C592B3B8D08965A0B3DA11653A2CF3894ACED9D00";
    attribute INIT_0D of inst : label is "B2D16D424CB2C2F9743200208BD5200208BD51CDDE3C50AB0847462A6BAF4F86";
    attribute INIT_0E of inst : label is "44C980000000000000000000000000054910BD23F63D222DABD3471E9252B6CC";
    attribute INIT_0F of inst : label is "A25E7A18C8B6EF4D84E3D240E50C617622A90540542E880054BFC5E32E4800E2";
    attribute INIT_10 of inst : label is "4079F3A31100F01522FE0064D0B3F9FBB42622A8008215188AA00208557377A8";
    attribute INIT_11 of inst : label is "22142FAF7A81F03E9A108252FC968284E221388B65689FFFB23B8204CDA10E08";
    attribute INIT_12 of inst : label is "74E3D4AA85CB57AF6A75CCB9484621A294FB3FC49B48C45D293DAA90CC435B72";
    attribute INIT_13 of inst : label is "AD6AB1595634D7658996EE5A41403AAF7296C148EA00F25CCEDB69D8BF234D5B";
    attribute INIT_14 of inst : label is "D64F4A47B407F14A0000002CCD98952880403F8A50CC8C48000000000027A96D";
    attribute INIT_15 of inst : label is "7749CD6F415538D55B5979DEFD290DDFFF7F1F8C4D485BD6D5509EAC2D69BBDA";
    attribute INIT_16 of inst : label is "461B9533BB15566118A0ED258369665E6DAF5DEDCA7A9EACFC7FC9979C3DADBC";
    attribute INIT_17 of inst : label is "6127DE6B54B02F2111622CF3A39DC6F9927B114471B108ADBD9A78897672504C";
    attribute INIT_18 of inst : label is "6440C9495CEF7295C3CF3CCC919B9CC5A0524A48C359E64ECF36A5ED636329E4";
    attribute INIT_19 of inst : label is "0D3BFF3FD0CB26221B2CC186ADBC096D007C9361B850E8CE2B4E14E800046361";
    attribute INIT_1A of inst : label is "DE315720857219C628E40572123098668D1EC45551F17EA8FE54AE4292845E7D";
    attribute INIT_1B of inst : label is "86B2FBB044C14B6521E536826FAA2E1AB444555118CFF39BFD8840098B61A3E0";
    attribute INIT_1C of inst : label is "BD1B208FC9B8A1874345821EE025CA72BC944788F3929C992E583FF7F64B6E20";
    attribute INIT_1D of inst : label is "000000179019F0DFE81FF7E0381F80003802E56092E19EA7AB1C8F7F5BD6DEF7";
    attribute INIT_1E of inst : label is "4927D9BB9FF8000016D249111100800001000100000000000000000000000000";
    attribute INIT_1F of inst : label is "00000C1165E2A3A80A88000440F0000C045705C1775C000E1AB031B418B09B96";
    attribute INIT_20 of inst : label is "2E7FABFE6B29492BAA31158CB50011231AD81F92081FCFAA8970964EDE2396BA";
    attribute INIT_21 of inst : label is "25D1BF1163D31C8D3FE8C4D8502AA138B2092FD080032F000F4273FC807FC440";
    attribute INIT_22 of inst : label is "3FE7B124000000200C5AEA35702094126A4C777DF00C462525C84E101B680214";
    attribute INIT_23 of inst : label is "ED980F601C057A07DE4B905482E2492D83A280DFF56291882FFE2DFB995C6DD9";
    attribute INIT_24 of inst : label is "76F2000B1F49CED9BD12C07FCEC0005E0808B04047000028C02876106C1621A1";
    attribute INIT_25 of inst : label is "00000000000000000000005C11AC8CC01157FE5BC4008BA12FC5132A536FBFCD";
    attribute INIT_26 of inst : label is "00000001C0000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "A0000000000000000020206040000000000000001E0000000000000000000000";
    attribute INIT_28 of inst : label is "947A8F43F0790006945A8F41F4790DDE9DADD38E864C6D7807647235E2A3A8B5";
    attribute INIT_29 of inst : label is "D53B000016860CDF865800031968517F534000E08B5A072FED9BE6F151D40002";
    attribute INIT_2A of inst : label is "B6D171460003F76ABDDD0000000FAAAA0000D5A46CA732B603FAA57B7A46F151";
    attribute INIT_2B of inst : label is "55552AAD55552AAD55552AAD55552AAD55552A000A882F142AFDB95E9092E6AD";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000000AD55552AAD";
    attribute INIT_2D of inst : label is "00000000000000016E1EDC2CE590B15C00000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "00000000000000000000000000000000000000000000000000000000009E0E90";
    attribute INIT_30 of inst : label is "947A8F43F0790006945A8F41F4790DDE9DADD38E864C6D7807647235E2A3A8B5";
    attribute INIT_31 of inst : label is "D53B000016860CDF865800031968517F534000E08B5A072FED9BE6F151D40002";
    attribute INIT_32 of inst : label is "B6D171460003F76ABDDD0000000FAAAA0000D5A46CA732B603FAA57B7A46F151";
    attribute INIT_33 of inst : label is "55552AAD55552AAD55552AAD55552AAD55552A000A882F142AFDB95E9092E6AD";
    attribute INIT_34 of inst : label is "000000000000000000000000000000000000000000000000000000AD55552AAD";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "00000000000000000000000000000000000000000000000000000000009E0E90";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B6D02A0085B16A1BB59A00000002090400207FFFFFFFFFFF81F94D7719690A81";
    attribute INIT_01 of inst : label is "62680570D0025A10402486004930C06B44554158A6F8438230F5085D1E2F01C0";
    attribute INIT_02 of inst : label is "91016801061827128E3402B829D646800743AC87540D43AC070269BD40982018";
    attribute INIT_03 of inst : label is "8C6C1017A40B156051A284000834B00DA09D5408FBF683FA3A1A0004A7855407";
    attribute INIT_04 of inst : label is "81204C382523E90221E9020484400021A05186007A0395C3444868000B1A2EAA";
    attribute INIT_05 of inst : label is "C10C3994C294A7800854070328DA05400709A2F85028EBFA86C41D0101659386";
    attribute INIT_06 of inst : label is "1314F514506867A0A700FFEDBFF6E925B6C9759710820A00300A04081A813D10";
    attribute INIT_07 of inst : label is "A7945010C330C521E002D05407057F50D8202A82D281C01D0250A9AB7BA8F514";
    attribute INIT_08 of inst : label is "550C050244382FF903065AFA030801BD3A8BD6F1C4F5140AC810384AE83CA098";
    attribute INIT_09 of inst : label is "A05AA4A1AA4A87E4F14551FAE8E8520823A3A1534850D142881FE1DF51720047";
    attribute INIT_0A of inst : label is "664D4DB7B0D466DBD90DB8B6D9DB36BA71105A0304121AA2A42092824F00382F";
    attribute INIT_0B of inst : label is "23F148EA22148FC523E88D0498B009823690BD0A023FB2401006803F297F446F";
    attribute INIT_0C of inst : label is "5EC2E80BF7557691297204666DBDAEE48C9FE66FBF66DF5D9BEB8CF6F7B7F485";
    attribute INIT_0D of inst : label is "A2CFB77F68A2C7817B599FB37BFF99FB373FFDB77B824C9BBDF6B3B3733BCFE4";
    attribute INIT_0E of inst : label is "616EC00000000000000000000000000039B8F591DBA8DAAAD21A05DFDB2C1448";
    attribute INIT_0F of inst : label is "CE6051AD6AAB08689CB3FB71F2CE7B837B36D67E5E2B666FB7C3FE18AF4DDED2";
    attribute INIT_10 of inst : label is "665973DDDDA8D83799EF3074ECDFFF7E1B83FB367ECDFF8FECD9FB37FF6DDEF3";
    attribute INIT_11 of inst : label is "BBD770F36C85613E8ABEF77716A96C86D3E1B4FDB7ADCBFFDFBBC3336A31CF37";
    attribute INIT_12 of inst : label is "7A120A50052497F092DE1DAD2936050A52245004C38466617FB6C2526C0A1B7E";
    attribute INIT_13 of inst : label is "08413C9B8A690A14CC02AF7145086AE97BD5C500F4C2B069F081400A69520156";
    attribute INIT_14 of inst : label is "868ED684207CA37440000002FFCCD4A4A8A3E51BA22FA66800000000001B4E05";
    attribute INIT_15 of inst : label is "D0950B68C4A7AD8152124891A75AA4915A3762EAA8D552148051E486C1F8C210";
    attribute INIT_16 of inst : label is "2241052BAC524B25A8D5A9052369449541484CA8AA51830F0821F12400214834";
    attribute INIT_17 of inst : label is "B145140330A058FAB22324BBA5DC263504135550110841297512B500543935FA";
    attribute INIT_18 of inst : label is "FFC0524A40E0708156AA2AC4808F58046011462C809064AAC224A9694145086A";
    attribute INIT_19 of inst : label is "4DF2AA2A127DB6864DF6C11429A80849011CAB40881C6087BB02066001484E21";
    attribute INIT_1A of inst : label is "A50637605AF610A0D6EC5AF61190C873E715C02370C168A0DF54B0F69A64CB21";
    attribute INIT_1B of inst : label is "E07A97A03BB00009002100142FBA040D741023704E03F0854B2200008260004C";
    attribute INIT_1C of inst : label is "190A209551B86387D3C40002A055C5D15C2645D8B980CC0F43B8046120004E28";
    attribute INIT_1D of inst : label is "000000002A19803FE05FFFE3C05F9F03C044210084C80DA1286C018843188C63";
    attribute INIT_1E of inst : label is "880639CB0AA806061B6492222201000A02001700000000000000000000000000";
    attribute INIT_1F of inst : label is "00001D9BA7B6F68F9CFF0005D0066828144E1384EF38013560A2C0A160A11C73";
    attribute INIT_20 of inst : label is "3EFFAAFE0A0B6D4AAB11A442A142D23AFA8C5D68733FB82AA452047FDE3B8438";
    attribute INIT_21 of inst : label is "0C8209051241A3A20660C1E25A83E84545542FE480020240D91053D4A875C650";
    attribute INIT_22 of inst : label is "0AA7E80000000074DC91AD255A44A05B4A6C0CFF5068C1C12511461E124E2A55";
    attribute INIT_23 of inst : label is "834D34400C14E258E843C93C49FC908B9AD5DF0888A0810C2B410DF0285A2D29";
    attribute INIT_24 of inst : label is "A20E000A0F50D1DA5A24C9AFF18000040008604003000008357E37656184CAB2";
    attribute INIT_25 of inst : label is "00000000000000000000004C737DFDCFD747FC5BCA9F8BAEAFC57A341A2597CF";
    attribute INIT_26 of inst : label is "000000003FFFFFFFFFFFFFFFFFFF555555555400000000000000000000000000";
    attribute INIT_27 of inst : label is "A00000000001FFFFFE7EE0E0DE1FFFFFFFFFFFFFE1FFFFFFE01E1FFFFFFFFE00";
    attribute INIT_28 of inst : label is "E8DE85CE95490009E8FE854C9149017E1FBFD144BC077D5C0246B317B6F68D64";
    attribute INIT_29 of inst : label is "41B50000030B40DB930A010F9F4720AB7A4F05A10A92003F690247DB7B470009";
    attribute INIT_2A of inst : label is "A8897BF300002AD56221F0000000444400001D0556C6362B015EB2757457DB7B";
    attribute INIT_2B of inst : label is "77772AAD55552AAF77772AAD55552AAF77772A031CFF10932648D1906CFAFFE8";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000000AD55552AAF";
    attribute INIT_2D of inst : label is "00000000000000004AAE4408790E3D9800000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000030C88";
    attribute INIT_30 of inst : label is "E8DE85CE95490009E8FE854C9149017E1FBFD144BC077D5C0246B317B6F68D64";
    attribute INIT_31 of inst : label is "41B50000030B40DB930A010F9F4720AB7A4F05A10A92003F690247DB7B470009";
    attribute INIT_32 of inst : label is "A8897BF300002AD56221F0000000444400001D0556C6362B015EB2757457DB7B";
    attribute INIT_33 of inst : label is "77772AAD55552AAF77772AAD55552AAF77772A031CFF10932648D1906CFAFFE8";
    attribute INIT_34 of inst : label is "000000000000000000000000000000000000000000000000000000AD55552AAF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000030C88";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "924488E0854024AF76D20022820820D4410C543FFFFFFFFF81FE64D6D87889E1";
    attribute INIT_01 of inst : label is "28225067448048026804948001A280505444505B0FFA0A021094015E252C200A";
    attribute INIT_02 of inst : label is "404920A0545101400211283320FA62041511F6D5084C11F4410825A410512050";
    attribute INIT_03 of inst : label is "B0FE105308C95960C19280000331314490F5B8CEE9D241EE30A8A82601255529";
    attribute INIT_04 of inst : label is "014668A0042A6D0120ED01029F260441451D14016895419D0102A24020081C01";
    attribute INIT_05 of inst : label is "8828AD5686D201202855291B2088911D0241014040205000BFC409018430C282";
    attribute INIT_06 of inst : label is "1A1249E21AA2EA009C2EB6DB6DB65B6697EDBEFA0811A820A12A12080C281042";
    attribute INIT_07 of inst : label is "92231A828BA2848848031855291A0017FC045A0852A4420C50742125482649E3";
    attribute INIT_08 of inst : label is "5F2295750A75221CA54F5ABEDD8E1C9E11EA0263A96E3DC9F454880A629118D0";
    attribute INIT_09 of inst : label is "28407241272CB76540C55D9AB06973CE3B51A87EF81D9866E60DF182713D5047";
    attribute INIT_0A of inst : label is "CEB757B239F06BD9DB649C926ACBC234C11A53853498296C9DA63508D400546A";
    attribute INIT_0B of inst : label is "62C318B823318B0C62A08F708A139894A73DD00A63279B0310B6241F132A6890";
    attribute INIT_0C of inst : label is "46C22A217757F73473FC07332CACCC69F74DBB2696724D08C9A1FE52B332F9CC";
    attribute INIT_0D of inst : label is "AA66DBA9AAA27315198C89113709C89113F09872738A9D3EC721919157D8E7C3";
    attribute INIT_0E of inst : label is "D16C400000000000000000000000000496CF6B9D098E4CC6CECA59B86F2764AC";
    attribute INIT_0F of inst : label is "95A51CC6331B3B294A3F0DF6B2631491191262B747233234AE55924C83066430";
    attribute INIT_10 of inst : label is "234D22CC88A25C59CD3311D2A64C062E49D119122444C9C664489113271C9CE5";
    attribute INIT_11 of inst : label is "CB6692304C6A804085CA592922EDB6C6D0D1A07EFA9E4E04CCB8F11923188B12";
    attribute INIT_12 of inst : label is "B254E808028016120262520E73B80538C724D6806D8022296190DCE7300AF84D";
    attribute INIT_13 of inst : label is "69CC0E13626F9B90460265014D4A62652857C54012B5702AD7955E0962027148";
    attribute INIT_14 of inst : label is "9916042DA74283244000009212C4418E383A1419232122200000000000873A55";
    attribute INIT_15 of inst : label is "9890A443136C8B695A48AA95AC1036944053AE2439814ED69A6C42D524C8DEF2";
    attribute INIT_16 of inst : label is "239B39A8314862B4645D4C0CC3AB32120C3526A2A09D0B166825288A20652947";
    attribute INIT_17 of inst : label is "412DB300B090820B2566360810503644821D451118084E2549D685E1984FA796";
    attribute INIT_18 of inst : label is "BBC448C101E7129D00B30FC718812A836A1168B6054C60AA6204EF2D3103CC23";
    attribute INIT_19 of inst : label is "48FBFF0E77AD9806F7B30414A54C1A01021E68A24095634D511024600212F180";
    attribute INIT_1A of inst : label is "CDA3A6828CA815B464D00CA8198144B0601D615240C1693C5E308228CCDF6A34";
    attribute INIT_1B of inst : label is "766AE6383FE580010129A950011034DB58595A400DC2F88549020028D590206A";
    attribute INIT_1C of inst : label is "0A61E1413886404A020504122058CD0342A514B294D4A0D6F32C8C6900020922";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000010A9401145401003D6AB5ED6BD8421";
    attribute INIT_1E of inst : label is "D77802001FF806061FF6DB333301FFE003FFC000000000000000000000000000";
    attribute INIT_1F of inst : label is "0002054B833535084CEC0008D10321A0D00601806718050080E100E080E19FF7";
    attribute INIT_20 of inst : label is "2B67E4794124AD7352B1B9A91942DBB183B871A6413FCA82991A847B8C919210";
    attribute INIT_21 of inst : label is "00A3844E6711B0AD83144BD24CE02924D34D042F00442540AADF03D8C966A16A";
    attribute INIT_22 of inst : label is "233300000000019EB722A104327131C9555A4CFD3050B37589DC258B88029A19";
    attribute INIT_23 of inst : label is "8B290C4008D06620C8B3051428E002088808A2228210940A333E0428863D9CBD";
    attribute INIT_24 of inst : label is "AA5A0019AF1A9B7B53FD680FFD800004000020000100001802201402680E4080";
    attribute INIT_25 of inst : label is "0000000000000000000001203E5F1CE25390BF3133D3E90DEBD11AB6147557A1";
    attribute INIT_26 of inst : label is "000000003FFFFFFFFFFFFFFFFFFF111111111000000000000000000000000000";
    attribute INIT_27 of inst : label is "40000001FFFF55FE1FDFDF9FA01FFF55FFFFFFFFFFFFFFFFE1FFFFFFFFFFFE00";
    attribute INIT_28 of inst : label is "4894306A40A9000048B430EA44A9108741485AEA02E124FC06A7178335350AEC";
    attribute INIT_29 of inst : label is "8477000033531448630009089020A09299280D0A25E802024EB1719A9A840005";
    attribute INIT_2A of inst : label is "449D1899000008442223FFFFFFFFFAFA00010E335BA269CE16903A5697219A9A";
    attribute INIT_2B of inst : label is "82828000888880002828000222220002828280094CEC22A74F4AD88726489ED1";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000222220002";
    attribute INIT_2D of inst : label is "000000000000000A034F204D61902ACA00000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000230910";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "2490381AA55504A6C36A032CBA936DD8518E957FFFFFFFFF8AF96C444D6D71EA";
    attribute INIT_01 of inst : label is "804813E09021701342125A2DA545101141405041203D146B5AA2452061B06419";
    attribute INIT_02 of inst : label is "690DC00908A28A02082409F0080011811A40011AD40340000C004AAB4059A048";
    attribute INIT_03 of inst : label is "1200D92480B10F2E44B673C001800F4C089190A31224C30E9A12001406876830";
    attribute INIT_04 of inst : label is "0385514594A4CE05004E0516910C4885061A288112074F82042A5811B9101644";
    attribute INIT_05 of inst : label is "14514AA5146206802168302F61D2070045058330724051011000188181A68A84";
    attribute INIT_06 of inst : label is "9462B0C61848BC111B074DA69B49B4984892012497C2241145B48C2812846D01";
    attribute INIT_07 of inst : label is "1507184515451885A00109683028222203F101014B04093108E245442145A086";
    attribute INIT_08 of inst : label is "A4204A224858B5B0021E6B94C24D30082035103595E479B120208129886A34A3";
    attribute INIT_09 of inst : label is "019FC089F40891FF8707E41F403C80212C88807E401B942C02981D0127600156";
    attribute INIT_0A of inst : label is "F6081636B3F2CB1B9A6DB2D6FCC9C6304111534C625463CD18C45E017820A8B4";
    attribute INIT_0B of inst : label is "E40F390022F3903CE4008A629E32A99BE617A08C52A84F40226AC430554126B4";
    attribute INIT_0C of inst : label is "970AFD7C802A86182FA845767DCDACC0B3999E6CB1A6D9669B2C38F736B7D0BC";
    attribute INIT_0D of inst : label is "EFCFFE63FBEF5B119B19BB77ED1D9BB77ED1982675060C15AC60B77731FBEC6A";
    attribute INIT_0E of inst : label is "EB7040000000000000000000000000003C9A5BED598CDA52D47451A8EBCD78FF";
    attribute INIT_0F of inst : label is "0D66198C694B51D13A351D68FCC635973776CEE156AB66EDC26BC65AA90CCC11";
    attribute INIT_10 of inst : label is "EE79AEDFBBD798559A6370B26FD81E0C1B47B776EDDF999CDDDBB77E7609DD43";
    attribute INIT_11 of inst : label is "261CB2B3ECB80080D61983CB37BFFF44C411313FDA9CC400DC04C373E1F1BB7E";
    attribute INIT_12 of inst : label is "BA70D10004085A330BC66E8C2FE8462842A39227DDA26665A5D2C05F908C5C5A";
    attribute INIT_13 of inst : label is "318998D7CDF93054CC13411C49090DC088A2C90A369CB42AD5128892A944458A";
    attribute INIT_14 of inst : label is "12A6D6A8C5B002304000004AB6CCD084198D801382AB6668000000000054760A";
    attribute INIT_15 of inst : label is "D370016300E060C58C5200529D5A14522180282A91D18C63114F3608D082D463";
    attribute INIT_16 of inst : label is "6475B038399144B9A08E0888A02A24A2082044C8EA1A294640360D2000463175";
    attribute INIT_17 of inst : label is "1539A2033111011BC64B28D0169126A59651186451BB5884E08A74A92266D368";
    attribute INIT_18 of inst : label is "0451924AD2E9153640E38D58311948066053706404016664CB32C72E2312CE27";
    attribute INIT_19 of inst : label is "498000846FC49845FA930C18C50C03B50120C200A25A620AA9089760010A1800";
    attribute INIT_1A of inst : label is "E8BB1492EE49079770906C480BD8681A7408A751C8C16838E122B3EED8774CBC";
    attribute INIT_1B of inst : label is "D70AE0B833A5ADB501A5ADCB669833D3004751C9EFFC0F066FF6002D7B91BF62";
    attribute INIT_1C of inst : label is "7DDFE5753982F0810300419A40602E0B8094B686F01280D9A3947FED924B2D08";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000002C510144C6DDB70E6873DEE7BFDFF";
    attribute INIT_1E of inst : label is "0040020B00000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0001352B06DA1A04A8C90002E0022A8543D8F63D8060048B120625051205E004";
    attribute INIT_20 of inst : label is "40C04400210DE021FF1410A4124484A0853001A6101FC022A052956EC1851330";
    attribute INIT_21 of inst : label is "8AB3DC01A7041B8FD900081642720F2CB2CB102600211000E884801AF30611F7";
    attribute INIT_22 of inst : label is "0AB748004000838B04026515002212DC450195041244E8D29098B756D24E0900";
    attribute INIT_23 of inst : label is "2D8423FB11418E45D20AD4F2A79CD9FD018820A0A226DF131434402A2D5F67B7";
    attribute INIT_24 of inst : label is "2A420011708F08590324645F03F003DF9C18FCC0C7000038D100511101960821";
    attribute INIT_25 of inst : label is "0000000000000000000000E4D76B2F549D1A00A035648C71302B56F6D04E7811";
    attribute INIT_26 of inst : label is "FFFFFFFE00000000000000000000666666666600000000000000000000000000";
    attribute INIT_27 of inst : label is "5000000000000001E1BF3F7F7FE000001FFFFFFFFE0000001E000000000001FF";
    attribute INIT_28 of inst : label is "E0EA143601890009E0EA1436018909C81284900090D3403C001EFF46DA1A0160";
    attribute INIT_29 of inst : label is "04B600001800F4C040E000CED24318E5001106C100020621A838736D0D000008";
    attribute INIT_2A of inst : label is "451399F300007F7FBFFF00000000005500003543DB01BB8D07088BE6E6236D0D";
    attribute INIT_2B of inst : label is "A802AAAA0A0A2AA82A802AAA8282AAA802A82A0128C91183046AD9C26DD8B2E1";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000000A828282AAA";
    attribute INIT_2D of inst : label is "0000000000000003B490512A781E150A00000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000471458";
    attribute INIT_30 of inst : label is "E0EA143601890009E0EA1436018909C81284900090D3403C001EFF46DA1A0160";
    attribute INIT_31 of inst : label is "04B600001800F4C040E000CED24318E5001106C100020621A838736D0D000008";
    attribute INIT_32 of inst : label is "451399F300007F7FBFFF00000000005500003543DB01BB8D07088BE6E6236D0D";
    attribute INIT_33 of inst : label is "A802AAAA0A0A2AA82A802AAA8282AAA802A82A0128C91183046AD9C26DD8B2E1";
    attribute INIT_34 of inst : label is "000000000000000000000000000000000000000000000000000000A828282AAA";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000471458";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B6D24C5A9B546640512901A69A4924DC0626FA7FFFFFFFFF8BFE82666BEB618B";
    attribute INIT_01 of inst : label is "A4E92042F24B285145924E6DA541014454014449903D040EF2872D2120112509";
    attribute INIT_02 of inst : label is "012CA1172820802432F49021492490924F4A4B0F5CC54A480965EA25480DA001";
    attribute INIT_03 of inst : label is "9900C93794AD0531245A00000126202039B894A9DBB6980ABA5A44944B933C08";
    attribute INIT_04 of inst : label is "3365104094A607409207489090856A9525CA08003A4801090CA96925B068C144";
    attribute INIT_05 of inst : label is "041042210C424B90033C0808B27A49889F2D4C412B61441090000A8080A68A8B";
    attribute INIT_06 of inst : label is "8402FCF7C969260633242000490000490012490414CAC050409E01293A943529";
    attribute INIT_07 of inst : label is "1752C94104410096E4034B3C08428012023348114B82837D282265C42144ECB6";
    attribute INIT_08 of inst : label is "ED6C4C224868A096103639B44A0C141D34AF0877A5683881F0B05229E9389420";
    attribute INIT_09 of inst : label is "0C68690E8690D244C0181092E301516B2B91992ECA4FB32250C215423DBC2B57";
    attribute INIT_0A of inst : label is "0F1036A62480CB53D6292B948012442C03614905225329471084F23BCC45FDEE";
    attribute INIT_0B of inst : label is "08090200EC9020240803B622920208108404203050806B197668608071123480";
    attribute INIT_0C of inst : label is "808A4A280A0234000820997669A988D044181E6C25A6D8429B0978D6A6269024";
    attribute INIT_0D of inst : label is "AA0925485BEE3217D21112225511112225D116144A4E8549284822222DAD401E";
    attribute INIT_0E of inst : label is "524800000000000000000000000000062C121D0510A4938288C071688208388A";
    attribute INIT_0F of inst : label is "490749084E0A2301D62D104AA08424122224944164B244493480105222488902";
    attribute INIT_10 of inst : label is "4428AE91112A50111202202648900A691202A224488951088891222545851292";
    attribute INIT_11 of inst : label is "2A5483ACEAA20C109D129248219248D494B5252024A884029486822253A13A24";
    attribute INIT_12 of inst : label is "B9365024941052020A40424808008828088696EC150044452110881041105C21";
    attribute INIT_13 of inst : label is "6118A05546AB09408A0073452D0DAA711A67AD0FA351F8AA92371A9A8548550A";
    attribute INIT_14 of inst : label is "12A75E9185500F2080000088368CD0840A0A807904824448000000000088265C";
    attribute INIT_15 of inst : label is "00CA50191FE3E88D185B0CD3B57A64D2611424AEF3D388C6135C2C1D82AAC8C6";
    attribute INIT_16 of inst : label is "6641301811534EB565450830A06426C6DB61846C6B4A07D7249301B0CC8C63A2";
    attribute INIT_17 of inst : label is "3728C626B2120C54078C24647368DE54925B28A22C994AA4C48A54A9AA520800";
    attribute INIT_18 of inst : label is "FFC9DB6B9DEEB634E869044D9199DC5C6453526C4A0892664492852422921866";
    attribute INIT_19 of inst : label is "5012AA045001201A00241020848409B501A08A85A05AE50BBF2816E4012B0021";
    attribute INIT_1A of inst : label is "A0B6AE86D8E86616D5D0DAE86BBA5D366CB5CD6B42C16822217C828C08264EA4";
    attribute INIT_1B of inst : label is "156E56922AB2ADB564A7AD8B511056D558A56B42120D09476F08002DC204D350";
    attribute INIT_1C of inst : label is "810C324A0C02D4522A2C934A6001281A129572AE5552AAD082B934ACBB692869";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000026724D5E8DF97E10E900421000010";
    attribute INIT_1E of inst : label is "2080040040060000200000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "00017F7EA7F6363E9312000700FEE80403C0F03C000000000204040402070008";
    attribute INIT_20 of inst : label is "26886E84695B7129AADA158D955D0844C039E8CD84DFFFFD5EA7B57DC365B6A3";
    attribute INIT_21 of inst : label is "3EC4A8714A1A14B0A42A0C33E32A00E38E389C3F801A678173E6900EF31251F4";
    attribute INIT_22 of inst : label is "B541D4000024234A4D321495132494105C1577043D994EE424B556765B68DA6D";
    attribute INIT_23 of inst : label is "0100004300000600C0020012008000180075D77DFD66F12A5C756E1BB85A2657";
    attribute INIT_24 of inst : label is "6E72000130D95E5BC17FC00C018003C41C1820C0C100000800003000000C0000";
    attribute INIT_25 of inst : label is "00000000000000000000004533FD48C9035481E8A949A0E3601DE6F256C6C83A";
    attribute INIT_26 of inst : label is "FFFFFFFE3FFFFFFFFFFFFFFFFFFF777777777600000000000000000000000000";
    attribute INIT_27 of inst : label is "A0000001FFFFFFFFFE5EDE9E9FFFFFFFE1FFFFFE01FFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_28 of inst : label is "417E606A028D0005417E6068028D1986231858604062659C020793DFF6363F6C";
    attribute INIT_29 of inst : label is "1BF6000012620202420C06B9EEA51CC63473058D34A10243EA146FFB1B1E0001";
    attribute INIT_2A of inst : label is "2F1FD12200011B4DA6E700000000FFAA0001AA7B1BA8AD6D021063A626FFFB1B";
    attribute INIT_2B of inst : label is "FFFD55555FF555557FFFD55557FD555557FFD407131233A1522AC9364A94409B";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000001557FD55557";
    attribute INIT_2D of inst : label is "0000000000000001B6D0D02AFA1E5DFB00000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "00000000000000000000000000000000000000000000000000000000006719D8";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "002921387F45729964B604924924924448D23FFFFFFFFFFF98FF46E2C97994B8";
    attribute INIT_01 of inst : label is "111481090924D10C31492124906180145111050CA27D86210C194C818C419124";
    attribute INIT_02 of inst : label is "069344C48C30C18B6D0A40846592D868B0A324F0AB5AA324769013A2A022001C";
    attribute INIT_03 of inst : label is "C82736804A6F6434F2B2000003111804A6CF6B3700002116452530439048C44B";
    attribute INIT_04 of inst : label is "481198634210511040511046CF732650D0730C0045220426223484924DD58850";
    attribute INIT_05 of inst : label is "86186331812990400CC44B982445242640909A24D9041401C24002A086186044";
    attribute INIT_06 of inst : label is "C62802082494A00D4890B24B2592DB2D92D92592CC900118636232840146028D";
    attribute INIT_07 of inst : label is "4028246186618A601000A4C44B8280384E24304C2088E4928C19109084130208";
    attribute INIT_08 of inst : label is "A7972297271615B1C3938CD12171C629836530A3986782140E511C8494C14631";
    attribute INIT_09 of inst : label is "1AEAC718AC618BCC012002B204031CB5988FC5C26D7098972D8A115E83639C8E";
    attribute INIT_0A of inst : label is "BEEDA736B890C39B188DB0B6D2DB16B2C9DC2E729D0A94104A531044401A0220";
    attribute INIT_0B of inst : label is "20890821B39082242086C8980C9868CA17BCB06D18E86724892E4A10755E8C34";
    attribute INIT_0C of inst : label is "C67020282220B7B7799827336D8DAC4D88D95F2CA9B259D6CB3A7AE636B6DDE4";
    attribute INIT_0D of inst : label is "C6A5B679718283CBD98CC9196159CC9196159966633078B0E625911111B9C42E";
    attribute INIT_0E of inst : label is "4364C00000000000000000000000000398D859B1593A4E2CE50D0D8ACB66C344";
    attribute INIT_0F of inst : label is "243074C638B3943409B15974B66310C11112722CF67B332DE6D6B30B838664BB";
    attribute INIT_10 of inst : label is "33C706C88882DC5DCB3B911A245A0D4D89719113246599C4444C9196665998C9";
    attribute INIT_11 of inst : label is "FBF618B2AC61985035DE7B21935B6EC441F1106DB72ED282DF96F1996C189B92";
    attribute INIT_12 of inst : label is "3481188203C70A98E15328AF79983697F6E8D92499A02230A9D4E6F3306D352D";
    attribute INIT_13 of inst : label is "94A62F017029DC704586FB86B41B2ACFDC0C341839F03A409948A644E0A530A0";
    attribute INIT_14 of inst : label is "4916214A531E1B6F4000006E36C44DEE4838F0DB7AE3622000000000002593A2";
    attribute INIT_15 of inst : label is "0DC18C04301FF2B0B504F30C4885A30C8624B2B9042C252D4C2CC4602D20E529";
    attribute INIT_16 of inst : label is "99CA00C0C70C30300424044A40BA9128209E330306A312069068604F30529482";
    attribute INIT_17 of inst : label is "43C329C2DD440F87F80FB3A87D0F0F8B6D8DCF3DCB66B6331B718B66898B6CB7";
    attribute INIT_18 of inst : label is "00662C6C6072394C6114B8306E6B2B84BB8C1B9783F72D99796C58BA9CCC3178";
    attribute INIT_19 of inst : label is "02E95533332DB83665B704DA52B81490028230733181F0E0418C61F00296E7A0";
    attribute INIT_1A of inst : label is "3690C19243590C520A32415908984C122486A50D08C169A4407EE9425EE23025";
    attribute INIT_1B of inst : label is "719119C8445464909A109B1926CD0AC9803D0D0808590E1CD800402452910618";
    attribute INIT_1C of inst : label is "334AF7D5088E30C12122482100352358D2605C0B81CC0E42C854E21349248714";
    attribute INIT_1D of inst : label is "0000000000000F20000000000000000000191093C856401004B64635AD6B5AC6";
    attribute INIT_1E of inst : label is "2000000040060000200000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0003F52ACA505047E527000F910FEFFBFC3F0FC3FFFFFFFFFDFBFBFBFDFA0000";
    attribute INIT_20 of inst : label is "24A87EC794E04D94A879CA104D724233E14A0F16C97FE222BC50C8EA8B31CA04";
    attribute INIT_21 of inst : label is "48DA88870425C142800449DE8E240338E3CF680000759EC1E7B3D034F01D70FD";
    attribute INIT_22 of inst : label is "ABA2C8004024811A18084A60F499495A04071D843A44D9884A0206DC48070482";
    attribute INIT_23 of inst : label is "FEFFFFBCFFFFFDFFBFF9FFCDFE7FFFF7FF00A82A0038708B386B955CC8AA3513";
    attribute INIT_24 of inst : label is "C7180014C0E4633C3C023FF8FF7FFC3BE3E7DF3F3EFFFFF7FFFFCFFFFFFBFFFF";
    attribute INIT_25 of inst : label is "0000000000000000000001CC49259D32449140F2E34302E1C40F5829813CE01D";
    attribute INIT_26 of inst : label is "0000000000000000000000000000888888888800000000000000000000000000";
    attribute INIT_27 of inst : label is "500000000000000001A12161600000001E000001FE0000000000000000000000";
    attribute INIT_28 of inst : label is "DEEB9CA1CC380006DEEB8CA3CC380F499294838F8F8B296C01FE7F2A505044E1";
    attribute INIT_29 of inst : label is "203D00003111804A69820BFF7E5FCFA5239F0C91C31E01E5A1E3C12828230006";
    attribute INIT_2A of inst : label is "1043D8910001C4A25118FFFFFFFF0000000074D13582271B1D29861C1C212828";
    attribute INIT_2B of inst : label is "AAAAAAAAA0002AA82AAAAAAAA8002AA802AAAA0F65271C1E2D80A089245A5CC4";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000000AA80002AAA";
    attribute INIT_2D of inst : label is "000000000000000C914198C1E1C1020E00000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000CF1288";
    attribute INIT_30 of inst : label is "DEEB9CA1CC380006DEEB8CA3CC380F499294838F8F8B296C01FE7F2A505044E1";
    attribute INIT_31 of inst : label is "203D00003111804A69820BFF7E5FCFA5239F0C91C31E01E5A1E3C12828230006";
    attribute INIT_32 of inst : label is "1043D8910001C4A25118FFFFFFFF0000000074D13582271B1D29861C1C212828";
    attribute INIT_33 of inst : label is "AAAAAAAAA0002AA82AAAAAAAA8002AA802AAAA0F65271C1E2D80A089245A5CC4";
    attribute INIT_34 of inst : label is "000000000000000000000000000000000000000000000000000000AA80002AAA";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000CF1288";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "802020307F04629B6CB000000000000D00E07FFFFFFFFFFF91FE0391C8789091";
    attribute INIT_01 of inst : label is "2010010100001C08200004000061801051540558A67986000035080104010100";
    attribute INIT_02 of inst : label is "0C0070800C30C3020A88008024B6580004816DC4A84A816C4540134080680038";
    attribute INIT_03 of inst : label is "8A6692100C62603296200000033534432E882C1E000000044424200204001C09";
    attribute INIT_04 of inst : label is "2021986100024308004308068A22044060430C00E40204078010800109181A00";
    attribute INIT_05 of inst : label is "8618633180200400181C0958000404040000822010301014864002A0851440C6";
    attribute INIT_06 of inst : label is "C62104144090A6010B01964B65B2DB2DB2596CB24C904018600E02100106820D";
    attribute INIT_07 of inst : label is "08344061866188010001C01C09420290CE2518080180500A0C30208084020414";
    attribute INIT_08 of inst : label is "0246061502141520831142C003208260816001830842003004700A005081A631";
    attribute INIT_09 of inst : label is "086883088820988CC10016226001489C98050504254109020482015301411A8C";
    attribute INIT_0A of inst : label is "B4A5A4129C904209080498A24A491290C5182820140B000008423228CC086C66";
    attribute INIT_0B of inst : label is "208908202B9082242080A8100EB0ED8A533C900C18C82210540C0800E5530C34";
    attribute INIT_0C of inst : label is "C2502A808282333679B8173324C4A459CCCB4F25E8B24BD2C96A3A63129249E4";
    attribute INIT_0D of inst : label is "C6A4932B20828901498CC919214CCC919214C86321201838E621911111108024";
    attribute INIT_0E of inst : label is "4924400000000000000000000000000399C8CC914B224E2E441C048A59265155";
    attribute INIT_0F of inst : label is "646244C638B9107008914B20926311811112622C52293324B255160B0106643B";
    attribute INIT_10 of inst : label is "334502488882CC5CCB09911C244E04448931911324648CC4444C91923218C859";
    attribute INIT_11 of inst : label is "CB6630118460805139CAD9630749260E22838884922660824AC2719928188992";
    attribute INIT_12 of inst : label is "2002180002820AB0415628A679B81614E6D050249C802220ACD644F3302C25AD";
    attribute INIT_13 of inst : label is "10842E01A2308860448C8A023C0B188450043C0891F09900A101840CC0842080";
    attribute INIT_14 of inst : label is "09142108430A0A454000006C124449CE487850522AC1222000000000006C1486";
    attribute INIT_15 of inst : label is "88C08608100002209404A2000084220000A4C0C1002004250834C04420388421";
    attribute INIT_16 of inst : label is "8BCA9087070822300064800840CA11204114122200C300040001204A204210A2";
    attribute INIT_17 of inst : label is "61402140C5000FE7FFF036A865490C99248E4515412294210D508942008924B2";
    attribute INIT_18 of inst : label is "44056A62504A252C0018A014AAA232818A848A9AA155248B692448AA14442148";
    attribute INIT_19 of inst : label is "8CCD55E0332498066493045842A018000202102230814040620C21400212A5A1";
    attribute INIT_1A of inst : label is "1610C500431004C218A04310008040302012440400C1694021C7B14274E22225";
    attribute INIT_1B of inst : label is "619219004454400058000930378C0E00B01C04000209021548004000D0900208";
    attribute INIT_1C of inst : label is "1342F750087420830104000020350350D020640C81041806C848A00000000430";
    attribute INIT_1D of inst : label is "0000000000000F20000000000000000000102002889440100098029084210842";
    attribute INIT_1E of inst : label is "2000000040060000200000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0003F52AE492120FED6F000FB10FE00000000000000000000000000000020000";
    attribute INIT_20 of inst : label is "1588188558A0051800388D088CB2461161040832D97FAA281C0028C883122202";
    attribute INIT_21 of inst : label is "2882804F061483A28224338A1E20011041456BC080560E41CF139C05B110785C";
    attribute INIT_22 of inst : label is "A100E0000100013A30102020AA15854E88070880384AD9A42C0146DC48008245";
    attribute INIT_23 of inst : label is "000000B800000000000400200100001000AA002AAA9430041C4B4192A82A1513";
    attribute INIT_24 of inst : label is "8218001080D0533A70008003FC70000B80005C00020000100000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000001884805BD36C4B180C2A74600E0800C482082309018";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "50000001FFFEAA01E05EDE9E9FE000AA01FFFFFE000000001FFFFE1E00000000";
    attribute INIT_28 of inst : label is "8A801C23402800028A801C21402804431084069A1A09112801B45A3C92120CA1";
    attribute INIT_29 of inst : label is "01340000335344322B4A0BFD6F4F8EA1011F0C00810803E00081464909070006";
    attribute INIT_2A of inst : label is "200148910000800000000000000055550000E1C1105422291108228404464909";
    attribute INIT_2B of inst : label is "00000000000000002AAA8002AAAA8002A800000F6D6F18060F008091244B5848";
    attribute INIT_2C of inst : label is "00000000000000000000000000000000000000000000000000000002AAAA8000";
    attribute INIT_2D of inst : label is "0000000000000008030118414080031200000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000CA1288";
    attribute INIT_30 of inst : label is "8A801C23402800028A801C21402804431084069A1A09112801B45A3C92120CA1";
    attribute INIT_31 of inst : label is "01340000335344322B4A0BFD6F4F8EA1011F0C00810803E00081464909070006";
    attribute INIT_32 of inst : label is "200148910000800000000000000055550000E1C1105422291108228404464909";
    attribute INIT_33 of inst : label is "00000000000000002AAA8002AAAA8002A800000F6D6F18060F008091244B5848";
    attribute INIT_34 of inst : label is "00000000000000000000000000000000000000000000000000000002AAAA8000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000CA1288";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
