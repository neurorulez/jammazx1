-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "000000000000BEBE000000000000000000009000000000063C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF00000000700D0960700D0960B000B000000E000E";
    attribute INIT_03 of inst : label is "0960A00A569503C01694028006900000C3FF27F8FC3F2D78FFC32FD864190960";
    attribute INIT_04 of inst : label is "6009096018240280069000000690000018240280600909600B0001CA0260A1C0";
    attribute INIT_05 of inst : label is "3333333328282828F00F2FF8CEB32558C143255863C90BE07C3D096060090960";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333332D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "01400000478D3491234504212375C4212345042101F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "000090521607DE421607DE44000000000EA4C232FFFF206D61202B5CC3032618";
    attribute INIT_0D of inst : label is "7AD1235D6421141D70860B12D683000000001A80490848134997904425580000";
    attribute INIT_0E of inst : label is "52005800AD8A2D524565BD5900040002C4305700492D524565AD59569A95A65E";
    attribute INIT_0F of inst : label is "24DC4981A7126349C4989D710C1A0015B0008000A920BDB046ECDE8800900025";
    attribute INIT_10 of inst : label is "7DC498967126165C49897712636DC498927126265C4985C712605DC498597126";
    attribute INIT_11 of inst : label is "712E498DA712E498D777A0E774FC498DE7126151C498D87126165C4989071260";
    attribute INIT_12 of inst : label is "3712E498DE712E498D9712E498D0712E498DD712E498D9712E498D2712E498DB";
    attribute INIT_13 of inst : label is "D4712E498D3712E498D9712E498D8712E498D9712E498DC712E498D7712E498D";
    attribute INIT_14 of inst : label is "BAB371EB7AB3716E59891712E798D3712E498D6712E498DF712E498D2712E498";
    attribute INIT_15 of inst : label is "C61B966449E499147922455E79852712E24DC4B850712E049C5885B712E341A4";
    attribute INIT_16 of inst : label is "64514E599D472839A6551C6CE699D4708EE5999079E67554E7991572839E6555";
    attribute INIT_17 of inst : label is "EEC1BB37DCEE22C18B342E5E49669E496F9E79E790B34AF12198223B8A26AB96";
    attribute INIT_18 of inst : label is "3B63829334061D2140D93CD555550000F55F8002FD7FE00B146E1E3400000000";
    attribute INIT_19 of inst : label is "B04EE8E089082421B3C24E59810439E6E59E69B987966D59424F948863420AC1";
    attribute INIT_1A of inst : label is "966151D4E288B06C5279EB2C717DE47175C48A18714D270EC7CB3422C1346082";
    attribute INIT_1B of inst : label is "C1D60E68E411C13492191AC1C7B966251D73C20B8B063E4D1C13492090AC1C7B";
    attribute INIT_1C of inst : label is "E09BC4B07DE72C1F716BCB079E6D1C69209E0ADDBCB1797C2C1C5AD5E598D442";
    attribute INIT_1D of inst : label is "5F94F1EE49850758B050825C26CECDF71AE5981475821B2C18209098252C1B16";
    attribute INIT_1E of inst : label is "B5FC4967C1D41709F4E5F4E534253425DDDDCC7BB5FC493333B7BA59505CE5F9";
    attribute INIT_1F of inst : label is "D525519F0A08224E24A39662D0694BA51E175497086C20AA493892B9013FC07B";
    attribute INIT_20 of inst : label is "302BC1FF060000A5F00C816300905A0012301F960B931DDD303835350F611A1C";
    attribute INIT_21 of inst : label is "3301C3FF060000A540CCFFC300905A0030BFCFD2065500A5FE0C87F355905A00";
    attribute INIT_22 of inst : label is "30A5C381060000A55A0C42C300905A0030AFCFFF060000A5FA0CFFF300905A00";
    attribute INIT_23 of inst : label is "02FF1F0200FD0000FF8080F4FF000000002B1D7F3FD70000F000814BAA100000";
    attribute INIT_24 of inst : label is "02F57F8101F900005F8042FDEF40000003011F7F00F9000040C0FDB4EF000000";
    attribute INIT_25 of inst : label is "00FF00FF0AA00AA0C3C33EBCEC3B1694D0071694728D389334061D2140D93CD5";
    attribute INIT_26 of inst : label is "123020081DD42A282BA92A280F78022031342A2813362AAA30302A2A0FC32028";
    attribute INIT_27 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF1F9728281E9C2A28";
    attribute INIT_28 of inst : label is "0DD1222A1DD408801D1C2A2A0FC328A80CC022281FD62AA80FC30A8200000000";
    attribute INIT_29 of inst : label is "0FC32A283FDF0A823FFF0A820C0C2A2A3CE40AA203032A2830302A2A1FD70A82";
    attribute INIT_2A of inst : label is "3FD70A820FD720000FC32A28303020201D942A280FD30AA20FC3282A0FC30880";
    attribute INIT_2B of inst : label is "10040000670D24D1118D042111BDC421118D042132342AAA1B1E20203A3C0A82";
    attribute INIT_2C of inst : label is "00009052054BDC4A054BDD48000000002D28C03AFFFF13A140A41B9CC00F0698";
    attribute INIT_2D of inst : label is "78D9139D44A1075161C2081EE44B0000000028484A0448136917914016940000";
    attribute INIT_2E of inst : label is "40484840AE861C9655259ED501000002C430444C4B25514967A55956A959979A";
    attribute INIT_2F of inst : label is "37906805849E528DE6109C750E12011180C0800088A4ACF47728EE4820100121";
    attribute INIT_30 of inst : label is "7DC4A95241E617586A0544DE53ADE610907905AA5E41B50710687D449A5141E6";
    attribute INIT_31 of inst : label is "43E66B05849EE690D57FB1A377F06B05C49E5095E610D871059A5E4189071068";
    attribute INIT_32 of inst : label is "04DEE690DC791E89AD173168B85043E66B05C45EE690D8751E898D273168BA53";
    attribute INIT_33 of inst : label is "D4711E898D373168BA5143E66B05841EE690D8751E89BD073168B95343E66B05";
    attribute INIT_34 of inst : label is "A8FB72E768FB53E66A45045EE69CD07D1E899D273168BB5343E66B05049EE690";
    attribute INIT_35 of inst : label is "C61B95687924895448E6571669C5049ED389E63050710D889E50A537306B6124";
    attribute INIT_36 of inst : label is "54915E199D470AB195991F60E699D470BD29A85479E655D4E69D1476A31E5595";
    attribute INIT_37 of inst : label is "FC8989FFFF623089893C1F9A59269E496F9E79E7A0737839229402BB892AA99E";
    attribute INIT_38 of inst : label is "18EFA01B05C20C6572113DD155550000D7D78002DFF7C28317620D7800000000";
    attribute INIT_39 of inst : label is "93C2F8A08A0404A1B0CE5E19810439E6E7966AB5A51E5E95530BA640508E3809";
    attribute INIT_3A of inst : label is "94697154E28893E05279CBAC53F5D4B175C48A1853C5078EF60F04E2C1346082";
    attribute INIT_3B of inst : label is "F1161E28C491C13482593849E63D45A91C77C20B890E1FC90C534824A3601E73";
    attribute INIT_3C of inst : label is "E293E4307DE70F9352E7C90F9F691E6123923B19ACF15BF40F907959E694D442";
    attribute INIT_3D of inst : label is "6D5CF3E66905161C90D09318378AFD373969895064C60B6C0860A25007A4095E";
    attribute INIT_3E of inst : label is "B7F45927F114064DF5E1F5E105E105E1FF55DE33B7F4483721FF9AD95350F6B5";
    attribute INIT_3F of inst : label is "C56563570A08138A24A3946AD261692D0D5B65531B2022A24A34A2790337D233";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "7D7D0000000000006000000000090000000000000000000005540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF000000000690B00E0690B00E70007000000D000D";
    attribute INIT_03 of inst : label is "5005069003C0A96A01402968000009601BF4C3FF1EB4FC3F1FE4FFC306909826";
    attribute INIT_04 of inst : label is "069090060140241800000960000009600140241806909006538000D003850640";
    attribute INIT_05 of inst : label is "33333333141414141FF4F00F1AA4CD731AA4C28307D093C60690BC3E06909006";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333331EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "00000280AFC4412B3100082B3118682B3108282B2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "00001AA4B7118682B31104AC2570000000004043CCCCB9A56EB9AD5B1864C0C3";
    attribute INIT_0D of inst : label is "48AB3310482B004488DA1BB1C1AB015800000000120ACCC0021487AC4A090000";
    attribute INIT_0E of inst : label is "A40009009649209E79E786490000000CEA40233059E09249A48679E59E392492";
    attribute INIT_0F of inst : label is "19C454C671153190454C651101880D5800003000D9309D4582F1230D001A004A";
    attribute INIT_10 of inst : label is "90454C641153198454C251153094454C671153194454C651153090454C261153";
    attribute INIT_11 of inst : label is "113654E23113654E21141051400454C641153190454C261153194454C2511531";
    attribute INIT_12 of inst : label is "3113654E20113654E22113654E21113654E21113654E21113654E20113654E21";
    attribute INIT_13 of inst : label is "20113654E23113654E22113654E22113654E21113654E21113654E20113654E2";
    attribute INIT_14 of inst : label is "CCC49D704CC49D3644E63113654E60113654E20113654E20113654E23113654E";
    attribute INIT_15 of inst : label is "6369953B84644EE11953980644EA01153090454C241157090455C25115319064";
    attribute INIT_16 of inst : label is "3A8C4654EA318E195398C638654E6318DA644EE11953B804654EA018E1953880";
    attribute INIT_17 of inst : label is "1116CC49D71109166C48265E792792696E996D8652C49ADD778DE76ADAF38D95";
    attribute INIT_18 of inst : label is "6B169A048524664A066233190000AAAA4001FAAFD007FEBF582FBF1100000000";
    attribute INIT_19 of inst : label is "C59AC5A6979DA636AB024644E2011913688644DE01913784A771170DA05E6B16";
    attribute INIT_1A of inst : label is "953880642302C5916C6938EEF10C3AF10C38DE7AF11C7B73142C48250D05E79A";
    attribute INIT_1B of inst : label is "16640238B4DBC000237B7B1674D953B8067B16AC6C59CB41BC010637B7B1674D";
    attribute INIT_1C of inst : label is "235442459DB591675D34A4599A51E74D38DE091E4245AD43B1674D16644EA00B";
    attribute INIT_1D of inst : label is "62971D3654E62192C5B8DE61E1731205D3644E6019637BB16E379350C5B16459";
    attribute INIT_1E of inst : label is "55C58DCFD08426783434343474747474444444A655C78D888835D14D10996629";
    attribute INIT_1F of inst : label is "B34B315C4A8D225A75A0D050829D8074BF1031218D2634874969D68D032441A6";
    attribute INIT_20 of inst : label is "C2FF3017005A09004293F00CA5000060151523291514363C1010303010140FC3";
    attribute INIT_21 of inst : label is "CFE0301F005A09920BF3F40CA5008660CBFF3301005A0900FFE340CCA5000060";
    attribute INIT_22 of inst : label is "C342305A005A090081C3A50CA5000060CBFF33FF005A0900FFE3FFCCA5000060";
    attribute INIT_23 of inst : label is "AFD003E1001F002F07FA4BC07400F800BEFF0BA106B6000042807EBCA4000000";
    attribute INIT_24 of inst : label is "0F4207FF001F002A81F0FFD0F400A800EFE003CF001F00920BFBF3C074008600";
    attribute INIT_25 of inst : label is "00FF00FF055005503D7CC3C32968DC372968E00B341CB1048524664A06623319";
    attribute INIT_26 of inst : label is "2FEB300C262C0FC32EE8074333342BBA2B3A07432F692C6C3034303025380F86";
    attribute INIT_27 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF2F6903122D6823E3";
    attribute INIT_28 of inst : label is "262E0F872EEA0CC02E2E0C0C2DF80FD2272D0D852FE90FC3253C2FEB00000000";
    attribute INIT_29 of inst : label is "2F690FC30FC72FF30FD72FC30C0C0C0C0FD23DF8030307433A3A30300FC30FC3";
    attribute INIT_2A of inst : label is "0FC32FFF0FC33A3C0FC30FC33A3A30302D7807432FE93DF82F692FF22FE92EE8";
    attribute INIT_2B of inst : label is "00002008BD8C422700C40A2302D44AA302C40AA32BBB2C4C0F0F30300FD72F7D";
    attribute INIT_2C of inst : label is "0000296884DDA40A80DD272014B4000000005003FF00A9E56EB99E971960F003";
    attribute INIT_2D of inst : label is "6A2300DC4A231100BA12287DE227121400000000024AFC000118A72C4A090000";
    attribute INIT_2E of inst : label is "848008049649239279E7960900000300D88800BC78649249A58279E58E792492";
    attribute INIT_2F of inst : label is "3944754241D520D45704449522041E14000000C0C8749D45B039038D02121202";
    attribute INIT_30 of inst : label is "91415D20105729447442415521D05704449D425D5510D419047491414D221057";
    attribute INIT_31 of inst : label is "0176746200D757860194105141007542411520D457040499425D5510D0190475";
    attribute INIT_32 of inst : label is "00D75786009115D8C0A9116D4C290176746200575786009515D8C089116D4C29";
    attribute INIT_33 of inst : label is "009115D8C0B9116D4C2A0176746200975786009515D8C099116D4C2801767462";
    attribute INIT_34 of inst : label is "FD009C747D008D76752200D75786409115D8C089116D4C280176746200D75786";
    attribute INIT_35 of inst : label is "52AD867795207C29185789427622011520D057040491464D1511D01904759160";
    attribute INIT_36 of inst : label is "2BC85518C8B98E19625CC6385786429CD9687C29185789C057868290E19528C0";
    attribute INIT_37 of inst : label is "0156DE01C45D09165E80179A49E792696E996D867148BB5967CDD6AEF87BAD15";
    attribute INIT_38 of inst : label is "499E89488524568A142A02DD0000AAAA4001EBEBC143EFFB4B638CDD00000000";
    attribute INIT_39 of inst : label is "E616E526A75D85BA888E5508C089085769827712201525CC94BD074D9392499E";
    attribute INIT_3A of inst : label is "86749120008EE4155EA13BE2C3C438F90E30DE7AC3D458FF076049210D05E69E";
    attribute INIT_3B of inst : label is "15680238B6D3C00012BF49DE76D1627C163B27685E91D80D8CC1053BA4FD578D";
    attribute INIT_3C of inst : label is "119C5109AD7591674D7496919859D78D3BD20B1651099C8791E74D1657828283";
    attribute INIT_3D of inst : label is "619B0D7675622096E634DC69D0B70149D16C5C28186768FD4DBB905CE4355691";
    attribute INIT_3E of inst : label is "7545BF07E14016B805F005F055F055F0550065227547AE048931D345225146A9";
    attribute INIT_3F of inst : label is "92CF13D46B09129A64E4D050A31991308CDC00E58D2625C35A25E749012C6126";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "000000000000FFFF00000000000000000000D000000000073C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF00000000000000000140000000000000F000F000000F000F";
    attribute INIT_03 of inst : label is "0260A1C0014000000140000001400000FC032D58C3C327D8C03F25681EB40280";
    attribute INIT_04 of inst : label is "0000000000000000000000000140000007D000001FF402800960A00A0B0001CA";
    attribute INIT_05 of inst : label is "33333333282828283FFC0AA03FFC0AA03FFC0AA01FF402801FF402801FF40280";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333332D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "014000001B48964613114116122591161211411601F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "000090106130101161301018000000000EA4C030EEEE4E85844E9D61C2032608";
    attribute INIT_0D of inst : label is "B34613218116209F20E32660D403000000001A00404584C040485B1824580000";
    attribute INIT_0E of inst : label is "100058002482CD28B20B3C9200000002C0304700928E2092C934824B24C28B20";
    attribute INIT_0F of inst : label is "901580E405603A09580E83560C0A0005B0008000D2345A2B118ACA0E00900025";
    attribute INIT_10 of inst : label is "05580E815603A05580E425603909580E425603A09580E425603909580E425603";
    attribute INIT_11 of inst : label is "52B780C0052B780C02407DA802C580E83560390D580E435603A05580E4156039";
    attribute INIT_12 of inst : label is "152B780C0352B780C0252B780C0152B780C0352B780C0152B780C0252B780C02";
    attribute INIT_13 of inst : label is "0352B780C0052B780C0152B780C0352B780C0252B780C0252B780C0252B780C0";
    attribute INIT_14 of inst : label is "E8AB1637A8AB163790C4352B7A0C03527780C0152B780C0152B780C0252B780C";
    attribute INIT_15 of inst : label is "838DE43305790C815E8B209790CC056C3B0D5B0EC356C3B05582EC056C790148";
    attribute INIT_16 of inst : label is "320DB780C0360CDE0330D837780C4360EB7B0CC35E8320DB7A0C0360CDE8310D";
    attribute INIT_17 of inst : label is "9AACA2B1A02AC2AC8AB117AD869A65B6D8A18218E0AB29963A6E97A7E9F04DE0";
    attribute INIT_18 of inst : label is "8418E1450191403FE405424454150000F41F8002FC3FE00BB11F6D2200000000";
    attribute INIT_19 of inst : label is "2B21063844CE3638D19337B0C015DE83C05780FC15E43E099381288E31A9ACAC";
    attribute INIT_1A of inst : label is "E833056913F22B2AC0821419900511900100E5959029A291AC06B11A021A9A6B";
    attribute INIT_1B of inst : label is "AC68D1373826480403A7AEAC58DE83005693AFEA42B201866481443A7AEAC58D";
    attribute INIT_1C of inst : label is "ACA6F8EB1A2A1AC6963A6AB1E28A058CD0EF44ACA6AB02A1AAC58CAC790C4160";
    attribute INIT_1D of inst : label is "A0E9163790C815A82B00EBB25131AC59637A0C015A83AE2AC839EC27282ACAB3";
    attribute INIT_1E of inst : label is "D6280F0B60BC0E8A1D3E1C3E1C3E1D3EB9A888A4D6290FEEEE1E00CFF03A6A06";
    attribute INIT_1F of inst : label is "7B9330329D8E76A13E14F5BDB00FB53E6D014A410E7439D3DA84F84F464995A4";
    attribute INIT_20 of inst : label is "0FFF3FFF01FF000AF5F0816CFF40A00017350B831F961C9C303830301A340F49";
    attribute INIT_21 of inst : label is "0F013C0001FF000A40F0003CFF40A0000FFF3FD201AA000AFFF087FCAA40A000";
    attribute INIT_22 of inst : label is "0FF53F8101FF000A5FF042FCFF40A0000F00300001FF000A00F0000CFF40A000";
    attribute INIT_23 of inst : label is "3FFF0102000000AFFFFC80400000FA003FFF0001000000AFF5FC01650000FA00";
    attribute INIT_24 of inst : label is "3FF50501000000AF5FFC40500000FA003F010005000000AF40FC50000000FA00";
    attribute INIT_25 of inst : label is "00FF00FF0FF00FF03EBC3D7C3EBC3D7C3EBC3D7C382C34450191403FE4054244";
    attribute INIT_26 of inst : label is "0761300C0C842F692EE82F691B3C033021302F6907632EEE30343A3A0F92252C";
    attribute INIT_27 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0FC329380FC82B69";
    attribute INIT_28 of inst : label is "0C84272F0CC00CC00C0C2E2E0FD22DF80D85272D0FC32FE90F960FC300000000";
    attribute INIT_29 of inst : label is "0FC32F692FCF0FD32FFF0FC30C0C2E2E2DF01FF203032F6930303A3A0FC30FC3";
    attribute INIT_2A of inst : label is "2FC30FD70FC330140FC32F69303030300DD02F690FC31FF20FC32D7A0FC30CC0";
    attribute INIT_2B of inst : label is "000000000F0CD04F011850470138D0470118504723312EEE0F0F30302F7D0FD7";
    attribute INIT_2C of inst : label is "0000814000E1451400E147051414000028288421AAFF3C4CC713CC30914A5289";
    attribute INIT_2D of inst : label is "D0CB013CD047228731B240B8C0031010000008081050E14003414F0C02810000";
    attribute INIT_2E of inst : label is "0400080430C38B34D3CF389300000102D020001CE20E30C3CD20D34F24C3CD3C";
    attribute INIT_2F of inst : label is "9045E12050300A9C0E42C50B0A06141480808040952D0F3F2343DB0F20100020";
    attribute INIT_30 of inst : label is "03503909040E80C5E12050F00B940E42450F2039B00494B042E10B50190A040E";
    attribute INIT_31 of inst : label is "202EE10042320E80440C2AA03019E32050F00A940E42450B20393004949042E1";
    attribute INIT_32 of inst : label is "42720E80440FB08894200BE81901202EE10042B20E804403B08894200BE81903";
    attribute INIT_33 of inst : label is "440BB08894100BE81900202EE10042B20E80440BB08894300BE81902202EE100";
    attribute INIT_34 of inst : label is "BFB7002FFFB7002EE10042F20E88440B308894100BE81900202EE10042F20E80";
    attribute INIT_35 of inst : label is "B21C80E3076039002A0E3086E30052700B9C0E4AC50FA03970069C804AE10751";
    attribute INIT_36 of inst : label is "039CB08894322E030039C8320E80442CCFEA2902280E22860E880428EA300290";
    attribute INIT_37 of inst : label is "FF38B4FCD3E3B33CBC3D733CF34E30F3F831C71CF7F328C30EABB02AB9E12870";
    attribute INIT_38 of inst : label is "C35195D1655556669595555900000000C283C143CBE3C7D3C3C60CF300000000";
    attribute INIT_39 of inst : label is "0DFC172D270343B9B11630A89000A80E9046E32060300A9CA10C3BC373B0FBF4";
    attribute INIT_3A of inst : label is "88E20761202A4FFFF1035244C15070501451B4D0C370E1C8CD87D2C6430FCF3E";
    attribute INIT_3B of inst : label is "CFE180620CF35801343AFBF82E038009700BEFEB743E304725C013632FBFF200";
    attribute INIT_3C of inst : label is "E8F3BBB30F3E3C4FC22F7CBCF3DF7200B3727374B3FB252CBCCCFB340E800421";
    attribute INIT_3D of inst : label is "B6B0402EE30063704CCCEDFB4135CFD003EA1900380FCBFBCB3188B20FB3FC3E";
    attribute INIT_3E of inst : label is "C23C1F1E33E03E0F0F730F730F730F73AAF5B974C23C2E3F8BDE734383F3598B";
    attribute INIT_3F of inst : label is "78DF50B3EB4370BC0CCCF2F0C383C3B30CC0594C1C2C2CC7FC0CCFC3021DB134";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "FFFF000000000000E0000000000B0000000000000000000005540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF00000000000000000000028000000000F000F000000F000F";
    attribute INIT_03 of inst : label is "038506400000028000000280000002801EA4FC031BE4C3C31AB4C03F01402D78";
    attribute INIT_04 of inst : label is "0000000000000000000000000000028000000BE001402FF850050690538000D0";
    attribute INIT_05 of inst : label is "333333331414141405503FFC05503FFC05503FFC01402FF801402FF801402FF8";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333331EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000002802F04514B001451CB001C71CB001451CB2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "00001AA4B001C71CB001C72D2570000000000C03333335C2CC35C4B01064C043";
    attribute INIT_0D of inst : label is "504B031451CB010300DC42B0C2AB0058000000001072D004100DC72C0A090000";
    attribute INIT_0E of inst : label is "A40009001041031C71C708710000000CEA40231061801861460C514514214514";
    attribute INIT_0F of inst : label is "31C3C00C40F003183C00C40F01A00D50000030000F470FB710ADC3CD001A0008";
    attribute INIT_10 of inst : label is "103C00C50F003103C00C50F0031C3C00C50F003103C00C50F003183C00C60F00";
    attribute INIT_11 of inst : label is "0B02C00C40B02C00C500000000F3C00C50F003183C00C60F003103C00C70F003";
    attribute INIT_12 of inst : label is "50B02C00C50B02C00C60B02C00C70B02C00C40B02C00C40B02C00C60B02C00C7";
    attribute INIT_13 of inst : label is "C60B02C00C70B02C00C40B02C00C60B02C00C40B02C00C50B02C00C60B02C00C";
    attribute INIT_14 of inst : label is "0F770301CF770302C00C50B02C00C60B02C00C50B02C00C40B02C00C50B02C00";
    attribute INIT_15 of inst : label is "0370B0011C2C00440B000142C00C70F003143C00C50F003143C00C60F003143D";
    attribute INIT_16 of inst : label is "031402C00C500C0B003140302C00C500DC2C00860B0021002C008400C0B00210";
    attribute INIT_17 of inst : label is "EEDCBF70F2EF01DC0771C3DC71C6185148F3CF3CF477188306018060184530B0";
    attribute INIT_18 of inst : label is "70371C5555155540055554550000A82A4001F82FD007FC3F710CBC1100000000";
    attribute INIT_19 of inst : label is "B71C0DC70C0DC03701D482C000620B003142C00C40B00310030C30CDC0DC73DC";
    attribute INIT_1A of inst : label is "B000140D0000773DC0CF71CAD01C72D01C711C72D01C720EC70771C2C30DC71C";
    attribute INIT_1B of inst : label is "DC0F10003C3B4041047072DC0C0B000140C1DC87C77033C3B4041047073DC0C0";
    attribute INIT_1C of inst : label is "F03B00770F3C1DC3C30BC770F3FDC0C030DC73DCB0770F2E1DC0C3D42C000421";
    attribute INIT_1D of inst : label is "2CF2C302C004703C7700DC3DC31FDC3C302C00460343701DC03720380C1DCF72";
    attribute INIT_1E of inst : label is "4B3207DC10CC0F631E1F1E1F1E1F1E1F111111F44B300733331CD2C7303DC2CF";
    attribute INIT_1F of inst : label is "7353C873500D43D81D8870F0C007C01FBC00F14C0D403501CF607607211321F4";
    attribute INIT_20 of inst : label is "3FFF0FFF000502FF429CFAF05000FF801010373C0111377D1010353505411A96";
    attribute INIT_21 of inst : label is "30000FE0000502D2000C0BF0500087803FFF0F01000502FFFFFC40F05000FF80";
    attribute INIT_22 of inst : label is "3F420FFA000502FF81FCAFF05000FF8034A00C00000502FF0A1C00305000FF80";
    attribute INIT_23 of inst : label is "1FD0000100000BFF07F440000000FFE0417F000000000BFF429F00400000FFE0";
    attribute INIT_24 of inst : label is "FF42000000000BFF81FF00000000FFE017E0000000000BD20BD40000000087E0";
    attribute INIT_25 of inst : label is "00FF00FF0000000015542AA815542AA815542AA815542A555515554005555455";
    attribute INIT_26 of inst : label is "3ABA2008377C0A822BA9020227702AAA3B3E02023B3C28283030202025690A82";
    attribute INIT_27 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF3F3D02023C3C22A2";
    attribute INIT_28 of inst : label is "277B0A823FFE08803F3E08082DE90A82266808803FFC0A8225692AAA00000000";
    attribute INIT_29 of inst : label is "2F690A821FD72AA21FD72A820C0C08081EC628A8030302023A3A20201FD70A82";
    attribute INIT_2A of inst : label is "1FD72AAA0FD72A280FC30A823A3A20203D3C02022FF928A82F692AA22FE92AA8";
    attribute INIT_2B of inst : label is "1004200818CC174200556316034123D6005163163ABE28081B1E20201A962A28";
    attribute INIT_2C of inst : label is "00002878C0948259C094827800A000000500481255AA65839D20B46540218402";
    attribute INIT_2D of inst : label is "1346004D2316011332013428E66B020000000040512394005200C27C1E180000";
    attribute INIT_2E of inst : label is "80C048400400460C20C30C7000000200C898448C21C00830431C100114200004";
    attribute INIT_2F of inst : label is "21D393003424024949C093162420090100400080495A686B2264E30802120301";
    attribute INIT_30 of inst : label is "163424014C49119393003424024D49C0D3120024244C4D01C0931A3434024C49";
    attribute INIT_31 of inst : label is "495B9200242549C090004444312392003464034D49C0D31E0024644C4D31C093";
    attribute INIT_32 of inst : label is "246549C09216244C492192B42403495B9200246549C09216244C492192B42402";
    attribute INIT_33 of inst : label is "921E244C492192B42401495B920024E549C09212244C490192B42402495B9200";
    attribute INIT_34 of inst : label is "482B0559882B055B9340246549C0921E644C491192B42401495B9200242549C0";
    attribute INIT_35 of inst : label is "012DC4911E3504014C490113934035A4014D49C4D3164034644C4D21D4931224";
    attribute INIT_36 of inst : label is "0149244C49101F120034417149C0D004DA3534034C49109149C09004F424014D";
    attribute INIT_37 of inst : label is "ABC888B9A2AA63000039A74D24924D1468638A38C0A3291611488565581474A4";
    attribute INIT_38 of inst : label is "04B25905001541114501510045518AA245518AA2C553CAA303D5CC8400000000";
    attribute INIT_39 of inst : label is "828D2C125F0084726055A45C41334C495193931035640449024D2380A2452788";
    attribute INIT_3A of inst : label is "C0911605105402ACE20226D3834120DC08244D378241029B850A20D682189249";
    attribute INIT_3B of inst : label is "9E0241550BE24100012527885B5200046451BC06C038218EC48144125268E505";
    attribute INIT_3C of inst : label is "87A250630A683942865AC039E2A8A50473C1678884A30A2B3901A50849C45024";
    attribute INIT_3D of inst : label is "38A3855B904006E4008CCA34C25F9E3152B40403404B0680C03347A10A00C83B";
    attribute INIT_3E of inst : label is "4C6A260D63100C2A0F5E0F5A0F5A0F5E004421204C69152E4798B10B42F0E30A";
    attribute INIT_3F of inst : label is "40DF8872074466492F5065F581438756CC85D2811D1010D5C96851CB548325E4";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
