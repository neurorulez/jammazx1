library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity xevious_cpu_gfx_8bits is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(16 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of xevious_cpu_gfx_8bits is
	type rom is array(0 to  69631) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"10",X"32",X"00",X"71",X"C3",X"2E",X"01",X"87",X"D2",X"4F",X"00",X"25",X"C3",X"4F",X"00",
		X"A7",X"F2",X"4F",X"00",X"25",X"C3",X"4F",X"00",X"A7",X"F0",X"ED",X"44",X"C9",X"33",X"33",X"C9",
		X"06",X"03",X"21",X"80",X"81",X"AF",X"18",X"2C",X"EB",X"CD",X"28",X"01",X"29",X"29",X"19",X"C9",
		X"E1",X"DD",X"75",X"00",X"DD",X"74",X"01",X"C9",X"E5",X"D5",X"C5",X"F5",X"32",X"30",X"68",X"21",
		X"20",X"68",X"36",X"00",X"36",X"01",X"CD",X"96",X"00",X"F1",X"C1",X"D1",X"E1",X"FB",X"C9",X"85",
		X"6F",X"D0",X"24",X"C9",X"1A",X"8E",X"27",X"77",X"13",X"23",X"10",X"F8",X"DC",X"09",X"13",X"CD",
		X"11",X"13",X"C3",X"3A",X"13",X"FF",X"D9",X"ED",X"A0",X"EA",X"93",X"00",X"08",X"3E",X"10",X"32",
		X"00",X"71",X"2A",X"04",X"80",X"7E",X"A7",X"28",X"19",X"36",X"00",X"2C",X"2C",X"4E",X"2C",X"46",
		X"2C",X"5E",X"2C",X"56",X"2C",X"D5",X"5E",X"2C",X"56",X"2C",X"22",X"04",X"80",X"EB",X"D1",X"32",
		X"00",X"71",X"08",X"D9",X"ED",X"45",X"21",X"00",X"82",X"11",X"80",X"87",X"01",X"40",X"00",X"ED",
		X"B0",X"21",X"00",X"83",X"11",X"80",X"97",X"01",X"40",X"00",X"ED",X"B0",X"21",X"00",X"81",X"11",
		X"80",X"A7",X"01",X"40",X"00",X"ED",X"B0",X"2A",X"20",X"80",X"7D",X"A4",X"32",X"03",X"80",X"32",
		X"70",X"D0",X"3A",X"AD",X"85",X"A7",X"28",X"12",X"3A",X"18",X"80",X"FE",X"BB",X"28",X"FE",X"CD",
		X"15",X"01",X"CB",X"7D",X"C8",X"3E",X"01",X"32",X"02",X"80",X"3E",X"01",X"32",X"00",X"80",X"21",
		X"18",X"80",X"01",X"03",X"71",X"11",X"00",X"70",X"EB",X"3A",X"00",X"71",X"E6",X"E0",X"78",X"06",
		X"00",X"20",X"05",X"D9",X"32",X"00",X"71",X"C9",X"E5",X"2A",X"06",X"80",X"77",X"2C",X"2C",X"71",
		X"2C",X"70",X"2C",X"73",X"2C",X"72",X"2C",X"D1",X"73",X"2C",X"72",X"2C",X"22",X"06",X"80",X"C9",
		X"11",X"00",X"70",X"18",X"D4",X"11",X"00",X"68",X"06",X"08",X"1A",X"1F",X"CB",X"1D",X"1F",X"CB",
		X"1C",X"13",X"10",X"F6",X"22",X"16",X"80",X"C9",X"21",X"00",X"00",X"C3",X"08",X"00",X"F3",X"ED",
		X"56",X"AF",X"32",X"30",X"68",X"32",X"0A",X"80",X"32",X"10",X"D0",X"32",X"30",X"D0",X"32",X"20",
		X"68",X"32",X"21",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"01",X"20",X"00",X"21",X"00",X"68",
		X"70",X"23",X"0D",X"20",X"FB",X"31",X"00",X"D0",X"06",X"00",X"58",X"FD",X"21",X"3D",X"03",X"DD",
		X"21",X"31",X"03",X"21",X"00",X"00",X"DD",X"56",X"00",X"DD",X"4E",X"01",X"15",X"28",X"2D",X"FD",
		X"35",X"00",X"20",X"0E",X"32",X"30",X"68",X"78",X"86",X"12",X"23",X"13",X"79",X"BA",X"20",X"F4",
		X"18",X"14",X"EB",X"32",X"30",X"68",X"1A",X"80",X"BE",X"20",X"1E",X"23",X"13",X"79",X"BC",X"20",
		X"F2",X"EB",X"FE",X"CF",X"28",X"0A",X"DD",X"23",X"DD",X"23",X"18",X"CA",X"FD",X"23",X"18",X"BF",
		X"78",X"C6",X"11",X"38",X"0D",X"47",X"C3",X"5B",X"01",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"32",X"00",X"85",X"AF",X"32",X"AD",X"85",X"CD",X"67",X"03",X"11",X"3E",X"03",X"32",
		X"30",X"68",X"13",X"1A",X"6F",X"13",X"1A",X"67",X"A7",X"28",X"0D",X"13",X"1A",X"A7",X"28",X"EF",
		X"77",X"13",X"01",X"C0",X"FF",X"09",X"18",X"F4",X"3A",X"00",X"85",X"FE",X"10",X"28",X"08",X"32",
		X"CF",X"C4",X"32",X"30",X"68",X"18",X"FB",X"3E",X"18",X"32",X"CF",X"C4",X"3E",X"14",X"32",X"8F",
		X"C4",X"31",X"80",X"A7",X"AF",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"03",X"77",X"ED",
		X"B0",X"32",X"30",X"68",X"21",X"80",X"87",X"77",X"2C",X"20",X"FC",X"21",X"80",X"97",X"77",X"2C",
		X"20",X"FC",X"21",X"80",X"A7",X"77",X"2C",X"20",X"FC",X"32",X"AD",X"85",X"21",X"00",X"92",X"22",
		X"04",X"80",X"22",X"06",X"80",X"77",X"2C",X"20",X"FC",X"3E",X"01",X"32",X"20",X"68",X"32",X"22",
		X"68",X"32",X"23",X"68",X"21",X"55",X"03",X"01",X"06",X"A1",X"CD",X"10",X"01",X"FB",X"11",X"74",
		X"85",X"21",X"00",X"00",X"0E",X"10",X"06",X"00",X"78",X"86",X"12",X"23",X"47",X"79",X"BC",X"20",
		X"F7",X"13",X"79",X"C6",X"10",X"4F",X"FE",X"50",X"20",X"EC",X"06",X"07",X"21",X"71",X"85",X"7E",
		X"A7",X"20",X"15",X"23",X"05",X"20",X"F8",X"3E",X"18",X"32",X"D1",X"C4",X"3E",X"14",X"32",X"91",
		X"C4",X"3E",X"0F",X"32",X"AC",X"85",X"18",X"06",X"78",X"32",X"D1",X"C4",X"18",X"FE",X"16",X"08",
		X"21",X"00",X"68",X"DD",X"21",X"D5",X"C4",X"FD",X"21",X"95",X"C4",X"01",X"00",X"00",X"7E",X"1F",
		X"3F",X"CB",X"11",X"1F",X"3F",X"CB",X"10",X"DD",X"70",X"00",X"FD",X"71",X"00",X"DD",X"23",X"FD",
		X"23",X"23",X"15",X"20",X"E6",X"3A",X"AC",X"85",X"32",X"D3",X"C4",X"3A",X"18",X"80",X"87",X"38",
		X"26",X"FE",X"FE",X"20",X"07",X"3A",X"19",X"80",X"3C",X"CA",X"7E",X"02",X"3A",X"AC",X"85",X"3C",
		X"FE",X"10",X"20",X"01",X"AF",X"32",X"AC",X"85",X"32",X"D3",X"C4",X"26",X"A0",X"6F",X"3E",X"01",
		X"77",X"CD",X"5B",X"03",X"C3",X"7E",X"02",X"CD",X"67",X"03",X"3E",X"27",X"0E",X"18",X"21",X"C4",
		X"C6",X"06",X"22",X"E5",X"D1",X"12",X"13",X"05",X"20",X"FB",X"06",X"40",X"2B",X"05",X"20",X"FC",
		X"0D",X"20",X"EE",X"21",X"C5",X"B6",X"3E",X"64",X"CD",X"1B",X"03",X"21",X"84",X"B6",X"3E",X"A4",
		X"CD",X"1B",X"03",X"21",X"85",X"B6",X"3E",X"E4",X"CD",X"1B",X"03",X"CD",X"5B",X"03",X"3A",X"18",
		X"80",X"CB",X"7F",X"28",X"F9",X"CD",X"5B",X"03",X"C3",X"88",X"03",X"0E",X"0C",X"E5",X"D1",X"06",
		X"11",X"12",X"13",X"13",X"05",X"20",X"FA",X"06",X"80",X"2B",X"05",X"20",X"FC",X"0D",X"20",X"ED",
		X"C9",X"79",X"80",X"83",X"88",X"91",X"92",X"95",X"97",X"A1",X"A8",X"B1",X"CF",X"01",X"00",X"CF",
		X"C5",X"1B",X"0A",X"16",X"00",X"D1",X"C5",X"1B",X"18",X"16",X"00",X"53",X"C6",X"1C",X"18",X"1E",
		X"17",X"0D",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"E5",X"21",X"00",X"00",X"2D",
		X"20",X"FD",X"25",X"20",X"FA",X"E1",X"C9",X"21",X"80",X"97",X"01",X"98",X"24",X"CD",X"7D",X"03",
		X"21",X"00",X"78",X"0E",X"80",X"CD",X"7D",X"03",X"21",X"00",X"B0",X"0E",X"CF",X"32",X"30",X"68",
		X"78",X"77",X"23",X"7C",X"B9",X"20",X"F6",X"C9",X"21",X"D2",X"03",X"11",X"60",X"85",X"01",X"08",
		X"00",X"ED",X"B0",X"16",X"08",X"21",X"00",X"68",X"7E",X"1F",X"CB",X"19",X"1F",X"CB",X"18",X"23",
		X"15",X"20",X"F5",X"21",X"CA",X"03",X"78",X"E6",X"03",X"CB",X"27",X"85",X"6F",X"7E",X"32",X"63",
		X"85",X"23",X"7E",X"32",X"64",X"85",X"21",X"CA",X"03",X"79",X"1F",X"E6",X"06",X"85",X"6F",X"7E",
		X"32",X"65",X"85",X"23",X"7E",X"32",X"66",X"85",X"18",X"10",X"02",X"03",X"02",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"02",X"02",X"F3",X"3E",X"10",X"32",X"00",X"71",
		X"AF",X"32",X"30",X"68",X"32",X"0A",X"80",X"32",X"10",X"D0",X"32",X"30",X"D0",X"32",X"20",X"68",
		X"32",X"21",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"21",X"00",X"80",X"11",X"01",X"80",X"01",
		X"FF",X"01",X"36",X"00",X"ED",X"B0",X"21",X"00",X"92",X"22",X"04",X"80",X"22",X"06",X"80",X"36",
		X"00",X"2C",X"20",X"FB",X"21",X"5B",X"04",X"11",X"80",X"82",X"01",X"40",X"00",X"ED",X"B0",X"3E",
		X"01",X"32",X"20",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"32",X"AD",X"85",X"21",X"60",X"85",
		X"01",X"08",X"A1",X"CD",X"10",X"01",X"FB",X"2A",X"00",X"80",X"2D",X"20",X"FA",X"24",X"22",X"00",
		X"80",X"DD",X"21",X"80",X"82",X"06",X"20",X"C5",X"CD",X"54",X"04",X"C1",X"DD",X"23",X"DD",X"23",
		X"10",X"F5",X"18",X"E3",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"9B",X"04",X"BB",X"14",X"00",
		X"30",X"D0",X"33",X"B3",X"33",X"E5",X"33",X"08",X"0F",X"9E",X"3B",X"E3",X"3B",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"27",X"17",X"62",X"18",X"CD",X"E1",X"06",X"CD",X"0D",
		X"07",X"CD",X"2A",X"07",X"CD",X"D9",X"10",X"3A",X"17",X"80",X"07",X"2F",X"E6",X"01",X"32",X"20",
		X"80",X"3E",X"01",X"32",X"2A",X"80",X"3E",X"F8",X"32",X"14",X"80",X"21",X"0E",X"0C",X"01",X"02",
		X"61",X"F3",X"CD",X"10",X"01",X"FB",X"AF",X"32",X"23",X"80",X"3A",X"29",X"80",X"A7",X"20",X"1B",
		X"3E",X"02",X"32",X"28",X"80",X"F7",X"3A",X"28",X"80",X"3D",X"21",X"40",X"0C",X"CF",X"5E",X"23",
		X"56",X"EB",X"E9",X"CD",X"81",X"08",X"3A",X"29",X"80",X"A7",X"C8",X"CD",X"F0",X"06",X"AF",X"32",
		X"28",X"80",X"3C",X"32",X"2A",X"80",X"CD",X"0D",X"07",X"CD",X"2A",X"07",X"CD",X"3C",X"08",X"CD",
		X"D5",X"0D",X"CD",X"DC",X"07",X"CD",X"AA",X"08",X"F7",X"CD",X"01",X"08",X"CD",X"23",X"08",X"3A",
		X"1B",X"80",X"A7",X"C8",X"32",X"23",X"80",X"AF",X"32",X"21",X"80",X"32",X"1B",X"80",X"21",X"80",
		X"81",X"77",X"2C",X"77",X"2C",X"77",X"2C",X"EB",X"21",X"0A",X"0C",X"3A",X"17",X"80",X"07",X"07",
		X"07",X"E6",X"03",X"D7",X"7E",X"EB",X"77",X"2C",X"2C",X"2C",X"2C",X"36",X"00",X"2C",X"36",X"00",
		X"2C",X"EB",X"3A",X"17",X"80",X"07",X"07",X"07",X"E6",X"03",X"EE",X"03",X"28",X"02",X"3E",X"01",
		X"21",X"10",X"0C",X"CF",X"4E",X"23",X"7E",X"67",X"69",X"3A",X"17",X"80",X"2F",X"0F",X"0F",X"E6",
		X"07",X"CF",X"EB",X"1A",X"77",X"2C",X"13",X"1A",X"77",X"2C",X"36",X"01",X"2C",X"3A",X"17",X"80",
		X"2F",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"3E",X"00",X"20",X"01",X"3C",X"77",X"3A",X"22",X"80",
		X"A7",X"28",X"10",X"21",X"80",X"81",X"11",X"C0",X"81",X"01",X"40",X"00",X"ED",X"B0",X"3E",X"01",
		X"32",X"01",X"A0",X"21",X"83",X"81",X"35",X"3A",X"87",X"81",X"4F",X"21",X"B3",X"3E",X"D7",X"7E",
		X"32",X"13",X"80",X"21",X"00",X"0D",X"22",X"10",X"80",X"79",X"21",X"00",X"A4",X"CF",X"7E",X"32",
		X"85",X"81",X"23",X"7E",X"32",X"86",X"81",X"AF",X"32",X"2B",X"80",X"32",X"2C",X"80",X"32",X"2D",
		X"80",X"32",X"22",X"84",X"32",X"44",X"80",X"CD",X"0D",X"07",X"CD",X"47",X"07",X"CD",X"D5",X"0D",
		X"CD",X"68",X"0F",X"21",X"62",X"18",X"22",X"BE",X"82",X"21",X"BB",X"14",X"22",X"82",X"82",X"AF",
		X"32",X"2A",X"80",X"3C",X"32",X"01",X"A0",X"3E",X"A0",X"32",X"41",X"80",X"CD",X"7F",X"07",X"F7",
		X"21",X"41",X"80",X"35",X"C0",X"CD",X"B7",X"07",X"F7",X"3A",X"2A",X"80",X"A7",X"C8",X"CD",X"47",
		X"07",X"3E",X"40",X"32",X"41",X"80",X"3A",X"11",X"80",X"D6",X"0E",X"FE",X"36",X"30",X"0B",X"21",
		X"87",X"81",X"34",X"3E",X"10",X"BE",X"20",X"02",X"36",X"06",X"3A",X"16",X"80",X"2F",X"07",X"07",
		X"07",X"E6",X"03",X"21",X"34",X"0C",X"D7",X"4E",X"3A",X"88",X"81",X"91",X"30",X"01",X"AF",X"32",
		X"88",X"81",X"F7",X"21",X"41",X"80",X"35",X"C0",X"21",X"40",X"79",X"11",X"41",X"79",X"01",X"0D",
		X"00",X"36",X"00",X"ED",X"B0",X"3A",X"83",X"81",X"A7",X"20",X"37",X"C3",X"43",X"11",X"3A",X"22",
		X"80",X"A7",X"28",X"1A",X"CD",X"0D",X"07",X"CD",X"47",X"07",X"CD",X"D5",X"0D",X"CD",X"6A",X"08",
		X"3E",X"80",X"32",X"41",X"80",X"F7",X"21",X"41",X"80",X"35",X"C0",X"CD",X"49",X"08",X"3A",X"C3",
		X"81",X"A7",X"28",X"17",X"CD",X"6D",X"07",X"3A",X"21",X"80",X"EE",X"01",X"32",X"21",X"80",X"C3",
		X"93",X"05",X"3A",X"C3",X"81",X"A7",X"20",X"EC",X"C3",X"93",X"05",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"D5",X"0D",X"CD",X"5D",X"08",X"3E",X"80",X"32",X"41",X"80",X"F7",X"21",X"41",X"80",
		X"35",X"C0",X"CD",X"49",X"08",X"3A",X"21",X"80",X"A7",X"CA",X"BB",X"04",X"CD",X"6D",X"07",X"AF",
		X"32",X"21",X"80",X"C3",X"BB",X"04",X"21",X"00",X"78",X"11",X"00",X"10",X"36",X"00",X"23",X"1B",
		X"7B",X"B2",X"20",X"F8",X"21",X"00",X"90",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",
		X"20",X"F8",X"21",X"00",X"A0",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",
		X"C9",X"21",X"00",X"78",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",
		X"21",X"00",X"79",X"11",X"40",X"00",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"74",
		X"79",X"11",X"06",X"00",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B0",
		X"11",X"00",X"08",X"36",X"24",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C0",X"11",X"00",
		X"08",X"36",X"24",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B8",X"11",X"00",X"08",
		X"36",X"03",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C8",X"11",X"00",X"08",X"36",X"00",
		X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B8",X"11",X"00",X"08",X"36",X"00",X"23",
		X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C8",X"3E",X"88",X"06",X"1C",X"77",X"23",X"3C",X"10",
		X"FB",X"21",X"00",X"C8",X"11",X"1C",X"C8",X"01",X"E4",X"07",X"ED",X"B0",X"C9",X"06",X"40",X"21",
		X"80",X"81",X"11",X"C0",X"81",X"4E",X"1A",X"77",X"79",X"12",X"2C",X"1C",X"10",X"F7",X"C9",X"3A",
		X"21",X"80",X"21",X"E5",X"0B",X"CF",X"5E",X"23",X"56",X"21",X"17",X"12",X"06",X"0A",X"0E",X"C0",
		X"CD",X"1F",X"14",X"21",X"19",X"10",X"11",X"DF",X"0B",X"06",X"06",X"0E",X"C0",X"CD",X"1F",X"14",
		X"11",X"FD",X"0B",X"21",X"1B",X"13",X"06",X"0D",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"1B",X"15",
		X"3A",X"83",X"81",X"CD",X"4F",X"14",X"C9",X"21",X"17",X"12",X"06",X"0A",X"3E",X"24",X"0E",X"C0",
		X"CD",X"5D",X"14",X"21",X"19",X"10",X"06",X"06",X"3E",X"24",X"0E",X"C0",X"CD",X"5D",X"14",X"06",
		X"10",X"21",X"1B",X"15",X"3E",X"24",X"0E",X"C0",X"CD",X"5D",X"14",X"C9",X"21",X"1F",X"16",X"11",
		X"CD",X"3E",X"06",X"13",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"21",X"10",X"11",X"E0",X"3E",X"06",
		X"07",X"CD",X"1F",X"14",X"21",X"21",X"10",X"06",X"07",X"0E",X"B0",X"3E",X"1A",X"CD",X"5D",X"14",
		X"C9",X"21",X"23",X"09",X"11",X"D9",X"0B",X"06",X"06",X"0E",X"C0",X"CD",X"1F",X"14",X"25",X"3A",
		X"29",X"80",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"4F",X"14",X"3A",X"29",X"80",X"E6",X"0F",
		X"C3",X"4F",X"14",X"3A",X"29",X"80",X"FE",X"01",X"28",X"01",X"AF",X"21",X"B1",X"0B",X"CF",X"5E",
		X"23",X"56",X"21",X"19",X"15",X"06",X"12",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"17",X"15",X"11",
		X"A0",X"0B",X"06",X"11",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"18",X"11",X"06",X"09",X"0E",X"C0",
		X"3E",X"24",X"CD",X"5D",X"14",X"21",X"1A",X"12",X"06",X"0A",X"C3",X"5D",X"14",X"21",X"18",X"11",
		X"11",X"97",X"0B",X"06",X"09",X"0E",X"C0",X"C3",X"1F",X"14",X"CD",X"5D",X"08",X"3A",X"21",X"80",
		X"21",X"E5",X"0B",X"CF",X"5E",X"23",X"56",X"21",X"1A",X"12",X"06",X"0A",X"0E",X"C0",X"C3",X"1F",
		X"14",X"3A",X"01",X"80",X"4F",X"E6",X"0F",X"C0",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"01",X"28",
		X"0D",X"21",X"1C",X"12",X"11",X"8C",X"0B",X"06",X"0B",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"1C",
		X"12",X"06",X"0B",X"0E",X"C0",X"3E",X"24",X"C3",X"5D",X"14",X"21",X"04",X"00",X"22",X"0C",X"80",
		X"0E",X"C8",X"21",X"09",X"15",X"11",X"9F",X"0A",X"06",X"12",X"CD",X"1F",X"14",X"21",X"0A",X"16",
		X"11",X"B1",X"0A",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0B",X"15",X"11",X"C4",X"0A",X"06",X"12",
		X"CD",X"1F",X"14",X"21",X"0C",X"16",X"11",X"D6",X"0A",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0D",
		X"17",X"11",X"E9",X"0A",X"06",X"14",X"CD",X"1F",X"14",X"21",X"0E",X"17",X"11",X"FD",X"0A",X"06",
		X"13",X"CD",X"1F",X"14",X"21",X"0F",X"17",X"11",X"10",X"0B",X"06",X"11",X"CD",X"1F",X"14",X"21",
		X"10",X"15",X"3E",X"F9",X"CD",X"4F",X"14",X"0E",X"B8",X"21",X"09",X"15",X"3E",X"0D",X"06",X"12",
		X"CD",X"5D",X"14",X"21",X"0A",X"16",X"3E",X"0D",X"06",X"13",X"CD",X"5D",X"14",X"21",X"0B",X"15",
		X"3E",X"11",X"06",X"02",X"CD",X"5D",X"14",X"3E",X"15",X"06",X"0F",X"CD",X"5D",X"14",X"3E",X"11",
		X"CD",X"4F",X"14",X"21",X"0C",X"16",X"3E",X"13",X"06",X"02",X"CD",X"5D",X"14",X"3E",X"17",X"06",
		X"10",X"CD",X"5D",X"14",X"3E",X"13",X"CD",X"4F",X"14",X"21",X"0D",X"17",X"3E",X"13",X"06",X"02",
		X"CD",X"5D",X"14",X"3E",X"17",X"06",X"10",X"CD",X"5D",X"14",X"3E",X"0F",X"CD",X"4F",X"14",X"3E",
		X"13",X"CD",X"4F",X"14",X"21",X"0E",X"17",X"3E",X"13",X"CD",X"4F",X"14",X"3E",X"19",X"06",X"11",
		X"CD",X"5D",X"14",X"3E",X"18",X"CD",X"4F",X"14",X"21",X"0F",X"17",X"3E",X"18",X"06",X"02",X"CD",
		X"5D",X"14",X"3E",X"19",X"CD",X"4F",X"14",X"3E",X"18",X"06",X"0E",X"CD",X"5D",X"14",X"21",X"10",
		X"15",X"3E",X"18",X"CD",X"4F",X"14",X"0E",X"C0",X"21",X"0B",X"15",X"11",X"60",X"0A",X"06",X"11",
		X"CD",X"1F",X"14",X"21",X"0C",X"13",X"11",X"71",X"0A",X"06",X"0E",X"CD",X"1F",X"14",X"21",X"0D",
		X"14",X"11",X"7F",X"0A",X"06",X"10",X"CD",X"1F",X"14",X"21",X"0E",X"15",X"11",X"8F",X"0A",X"06",
		X"10",X"CD",X"1F",X"14",X"3E",X"1A",X"0E",X"B0",X"21",X"0B",X"15",X"06",X"11",X"CD",X"5D",X"14",
		X"21",X"0C",X"13",X"06",X"0E",X"CD",X"5D",X"14",X"21",X"0D",X"14",X"06",X"10",X"CD",X"5D",X"14",
		X"21",X"0E",X"15",X"06",X"10",X"C3",X"5D",X"14",X"21",X"0A",X"16",X"11",X"21",X"0B",X"0E",X"C0",
		X"06",X"13",X"CD",X"1F",X"14",X"21",X"0B",X"15",X"11",X"34",X"0B",X"06",X"12",X"CD",X"1F",X"14",
		X"21",X"0C",X"15",X"11",X"46",X"0B",X"06",X"12",X"CD",X"1F",X"14",X"21",X"0D",X"16",X"11",X"58",
		X"0B",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0E",X"17",X"11",X"6B",X"0B",X"06",X"14",X"CD",X"1F",
		X"14",X"21",X"0F",X"17",X"11",X"7F",X"0B",X"06",X"0D",X"CD",X"1F",X"14",X"3E",X"1B",X"21",X"0A",
		X"16",X"0E",X"B0",X"06",X"13",X"CD",X"5D",X"14",X"21",X"0B",X"15",X"06",X"12",X"CD",X"5D",X"14",
		X"21",X"0C",X"15",X"06",X"12",X"CD",X"5D",X"14",X"21",X"0D",X"16",X"06",X"13",X"CD",X"5D",X"14",
		X"21",X"0E",X"17",X"06",X"14",X"CD",X"5D",X"14",X"21",X"0F",X"17",X"06",X"0D",X"C3",X"5D",X"14",
		X"2A",X"51",X"52",X"53",X"52",X"54",X"55",X"56",X"24",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",
		X"52",X"5E",X"5F",X"2A",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"7F",X"88",X"89",X"C0",
		X"C1",X"C2",X"C3",X"C2",X"C4",X"C5",X"C1",X"C6",X"C7",X"C1",X"C8",X"C1",X"C9",X"CA",X"CB",X"CA",
		X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",X"DA",X"DB",
		X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",
		X"EC",X"ED",X"EE",X"EF",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",X"FB",
		X"FC",X"FD",X"FE",X"FF",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BD",X"BD",X"BD",X"BE",X"BB",X"BB",X"BB",X"BB",X"BF",X"F0",
		X"F1",X"F2",X"BB",X"F3",X"F4",X"F4",X"F4",X"F4",X"F5",X"F6",X"F6",X"F6",X"F7",X"F4",X"F4",X"F4",
		X"F8",X"8A",X"8B",X"8C",X"8D",X"8E",X"8D",X"8F",X"90",X"87",X"91",X"92",X"93",X"94",X"87",X"95",
		X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9C",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"A4",
		X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",
		X"B5",X"B6",X"B7",X"B8",X"A7",X"B9",X"9A",X"BA",X"AB",X"BB",X"AA",X"9A",X"BC",X"BD",X"BE",X"BF",
		X"C0",X"C1",X"C2",X"9A",X"C3",X"AA",X"C4",X"C5",X"C6",X"C7",X"C8",X"AB",X"BB",X"C9",X"CA",X"CA",
		X"CB",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"CB",X"CA",X"CA",X"D3",X"D4",X"D5",X"D6",X"D7",
		X"AA",X"24",X"24",X"24",X"24",X"24",X"24",X"D8",X"D9",X"D9",X"D9",X"DA",X"12",X"17",X"1C",X"0E",
		X"1B",X"1D",X"24",X"0C",X"18",X"12",X"17",X"10",X"0A",X"16",X"0E",X"24",X"18",X"1F",X"0E",X"1B",
		X"19",X"1E",X"1C",X"11",X"24",X"1C",X"1D",X"0A",X"1B",X"1D",X"24",X"0B",X"1E",X"1D",X"1D",X"18",
		X"17",X"C7",X"0B",X"B5",X"0B",X"24",X"18",X"17",X"0E",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",
		X"24",X"18",X"17",X"15",X"22",X"24",X"24",X"18",X"17",X"0E",X"24",X"18",X"1B",X"24",X"1D",X"20",
		X"18",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"1B",
		X"0E",X"0A",X"0D",X"22",X"2C",X"E9",X"0B",X"F3",X"0B",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",
		X"18",X"17",X"0E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"1D",X"20",X"18",X"1C",X"18",X"15",
		X"1F",X"0A",X"15",X"18",X"1E",X"24",X"15",X"0E",X"0F",X"1D",X"05",X"02",X"01",X"03",X"02",X"02",
		X"14",X"0C",X"24",X"0C",X"20",X"00",X"10",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"30",X"00",
		X"20",X"00",X"FF",X"FF",X"20",X"00",X"10",X"00",X"10",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"20",X"00",X"FF",X"FF",X"10",X"18",X"08",X"00",X"1A",X"17",X"18",X"07",X"3A",X"1B",X"1F",X"15",
		X"35",X"0D",X"48",X"0C",X"35",X"0D",X"A2",X"0D",X"CD",X"2A",X"07",X"CD",X"0D",X"07",X"CD",X"DC",
		X"07",X"CD",X"D5",X"0D",X"CD",X"AA",X"08",X"3E",X"40",X"32",X"41",X"80",X"11",X"65",X"0C",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"21",X"41",X"80",X"35",X"28",X"03",X"C3",X"E3",X"04",X"21",X"60",
		X"0D",X"22",X"1E",X"7A",X"21",X"60",X"16",X"22",X"1E",X"7B",X"21",X"30",X"0F",X"22",X"1E",X"7C",
		X"21",X"02",X"80",X"22",X"1E",X"79",X"AF",X"32",X"1E",X"7D",X"11",X"93",X"0C",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"1E",X"7D",X"3C",X"32",X"1E",X"7D",X"FE",X"10",X"28",X"0B",X"0F",X"E6",
		X"07",X"C6",X"30",X"32",X"1E",X"7C",X"C3",X"E3",X"04",X"3E",X"78",X"32",X"1E",X"7D",X"11",X"B7",
		X"0C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"1E",X"7D",X"3C",X"32",X"1E",X"7D",X"28",X"13",
		X"E6",X"07",X"C6",X"38",X"32",X"1E",X"7C",X"2A",X"1E",X"7B",X"3E",X"F0",X"CF",X"22",X"1E",X"7B",
		X"C3",X"E3",X"04",X"3E",X"10",X"32",X"1E",X"7D",X"11",X"E1",X"0C",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"3A",X"1E",X"7D",X"3D",X"32",X"1E",X"7D",X"28",X"0B",X"0F",X"E6",X"07",X"C6",X"30",X"32",
		X"1E",X"7C",X"C3",X"E3",X"04",X"AF",X"32",X"41",X"80",X"32",X"1E",X"79",X"11",X"05",X"0D",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",X"80",X"E6",X"01",X"C2",X"E3",X"04",X"21",X"41",X"80",
		X"35",X"28",X"0E",X"7E",X"E6",X"07",X"21",X"38",X"0C",X"D7",X"7E",X"CD",X"C6",X"09",X"C3",X"E3",
		X"04",X"CD",X"F0",X"06",X"3E",X"03",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"C3",X"E3",X"04",X"AF",X"32",X"21",X"80",X"32",X"87",X"81",X"32",X"88",X"81",X"21",
		X"B3",X"3E",X"D7",X"7E",X"32",X"13",X"80",X"21",X"00",X"0D",X"22",X"10",X"80",X"AF",X"21",X"00",
		X"A4",X"CF",X"7E",X"32",X"85",X"81",X"23",X"7E",X"32",X"86",X"81",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"D5",X"0D",X"CD",X"DC",X"07",X"CD",X"E8",X"09",X"AF",X"32",X"2B",X"80",X"32",X"2C",
		X"80",X"32",X"2D",X"80",X"32",X"22",X"84",X"32",X"2A",X"80",X"11",X"83",X"0D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"2A",X"80",X"A7",X"20",X"03",X"C3",X"E3",X"04",X"CD",X"F0",X"06",X"3A",
		X"28",X"80",X"3C",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",X"72",X"01",X"C3",
		X"E3",X"04",X"CD",X"00",X"10",X"3E",X"40",X"32",X"41",X"80",X"11",X"B3",X"0D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"01",X"80",X"E6",X"07",X"C2",X"E6",X"04",X"21",X"41",X"80",X"35",X"28",
		X"03",X"C3",X"E6",X"04",X"3E",X"01",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"C3",X"E3",X"04",X"CD",X"63",X"14",X"CD",X"27",X"14",X"C3",X"EF",X"12",X"D5",X"E5",
		X"5D",X"54",X"7D",X"CD",X"F2",X"0D",X"EB",X"7C",X"CD",X"F2",X"0D",X"19",X"CD",X"35",X"0E",X"E1",
		X"D1",X"C9",X"67",X"2E",X"00",X"CD",X"FB",X"0D",X"6C",X"67",X"C9",X"C5",X"D5",X"CD",X"12",X"0E",
		X"CB",X"79",X"28",X"06",X"47",X"7C",X"93",X"67",X"78",X"9A",X"CB",X"7A",X"28",X"01",X"91",X"D1",
		X"C1",X"C9",X"EB",X"4F",X"21",X"00",X"00",X"06",X"08",X"29",X"17",X"30",X"03",X"19",X"CE",X"00",
		X"10",X"F7",X"C9",X"C5",X"4F",X"AF",X"06",X"10",X"29",X"17",X"38",X"03",X"B9",X"38",X"02",X"91",
		X"23",X"10",X"F5",X"C1",X"C9",X"C5",X"D5",X"E5",X"06",X"08",X"11",X"40",X"00",X"7D",X"6C",X"62",
		X"A7",X"ED",X"52",X"30",X"01",X"19",X"3F",X"CB",X"12",X"87",X"ED",X"6A",X"87",X"ED",X"6A",X"10",
		X"EF",X"7A",X"E1",X"D1",X"C1",X"C9",X"C6",X"40",X"C5",X"E5",X"4F",X"CB",X"71",X"28",X"02",X"ED",
		X"44",X"E6",X"7F",X"21",X"71",X"0E",X"D7",X"7E",X"CB",X"79",X"28",X"02",X"ED",X"44",X"E1",X"C1",
		X"C9",X"00",X"03",X"06",X"09",X"0C",X"10",X"13",X"16",X"19",X"1C",X"1F",X"22",X"25",X"28",X"2B",
		X"2E",X"31",X"33",X"36",X"39",X"3C",X"3F",X"41",X"44",X"47",X"49",X"4C",X"4E",X"51",X"53",X"55",
		X"58",X"5A",X"5C",X"5E",X"60",X"62",X"64",X"66",X"68",X"6A",X"6B",X"6D",X"6F",X"70",X"71",X"73",
		X"74",X"75",X"76",X"78",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"E5",X"CD",X"C4",X"0E",X"E1",X"CB",X"7D",X"28",X"03",X"2F",X"C6",X"81",X"CB",X"7C",
		X"C8",X"ED",X"44",X"C9",X"7C",X"DF",X"67",X"7D",X"DF",X"6F",X"BC",X"38",X"11",X"2E",X"00",X"CD",
		X"23",X"0E",X"29",X"29",X"29",X"29",X"29",X"7C",X"21",X"E7",X"0E",X"D7",X"7E",X"C9",X"7C",X"65",
		X"CD",X"CD",X"0E",X"2F",X"C6",X"41",X"C9",X"00",X"01",X"03",X"04",X"05",X"06",X"08",X"09",X"0A",
		X"0B",X"0C",X"0D",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"19",X"1A",
		X"1B",X"1C",X"1D",X"1D",X"1E",X"1F",X"1F",X"20",X"CD",X"12",X"0F",X"CD",X"25",X"0F",X"CD",X"38",
		X"0F",X"C9",X"3A",X"85",X"80",X"A7",X"C8",X"21",X"80",X"80",X"01",X"07",X"68",X"CD",X"10",X"01",
		X"AF",X"32",X"85",X"80",X"C9",X"3A",X"95",X"80",X"A7",X"C8",X"21",X"90",X"80",X"01",X"07",X"68",
		X"CD",X"10",X"01",X"AF",X"32",X"95",X"80",X"C9",X"3A",X"A6",X"80",X"A7",X"C8",X"21",X"A0",X"80",
		X"01",X"08",X"68",X"CD",X"10",X"01",X"AF",X"32",X"A6",X"80",X"C9",X"E5",X"2A",X"08",X"80",X"7D",
		X"87",X"87",X"85",X"3C",X"6F",X"7C",X"E6",X"84",X"28",X"04",X"EE",X"84",X"20",X"01",X"37",X"7C",
		X"8F",X"67",X"85",X"22",X"08",X"80",X"E1",X"C9",X"3A",X"83",X"81",X"A7",X"C8",X"47",X"C5",X"3E",
		X"25",X"21",X"23",X"1B",X"E5",X"0E",X"C0",X"CD",X"5D",X"14",X"E1",X"C1",X"0E",X"B0",X"3E",X"2A",
		X"C3",X"5D",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"CD",X"0D",X"07",X"CD",X"2A",X"07",X"CD",X"AA",X"08",X"18",X"06",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"27",X"14",X"CD",X"EF",X"12",X"CD",X"63",X"14",X"21",X"15",X"16",X"11",X"B8",X"10",
		X"0E",X"C0",X"06",X"12",X"CD",X"1F",X"14",X"21",X"18",X"19",X"11",X"CA",X"10",X"06",X"03",X"CD",
		X"1F",X"14",X"26",X"14",X"11",X"12",X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"13",X"85",X"06",
		X"0A",X"CD",X"1F",X"14",X"21",X"1A",X"19",X"11",X"CD",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",
		X"14",X"11",X"22",X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"23",X"85",X"06",X"0A",X"CD",X"1F",
		X"14",X"21",X"1C",X"19",X"11",X"D0",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"32",
		X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"33",X"85",X"06",X"0A",X"CD",X"1F",X"14",X"21",X"1E",
		X"19",X"11",X"D3",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"42",X"85",X"CD",X"47",
		X"14",X"26",X"0B",X"11",X"43",X"85",X"06",X"0A",X"CD",X"1F",X"14",X"21",X"20",X"19",X"11",X"D6",
		X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"52",X"85",X"CD",X"47",X"14",X"26",X"0B",
		X"11",X"53",X"85",X"06",X"0A",X"C3",X"1F",X"14",X"0B",X"3A",X"48",X"49",X"24",X"0F",X"3E",X"4B",
		X"3A",X"24",X"20",X"0A",X"1B",X"1B",X"12",X"18",X"1B",X"1C",X"01",X"48",X"49",X"02",X"43",X"39",
		X"03",X"47",X"39",X"04",X"49",X"3D",X"05",X"49",X"3D",X"21",X"F3",X"10",X"11",X"10",X"85",X"01",
		X"50",X"00",X"ED",X"B0",X"21",X"F0",X"10",X"11",X"24",X"80",X"01",X"03",X"00",X"ED",X"B0",X"C9",
		X"00",X"40",X"00",X"00",X"40",X"00",X"16",X"50",X"17",X"36",X"40",X"36",X"42",X"4A",X"47",X"36",
		X"00",X"00",X"00",X"00",X"35",X"00",X"0E",X"3E",X"47",X"47",X"4E",X"24",X"16",X"44",X"4A",X"50",
		X"00",X"00",X"00",X"00",X"30",X"00",X"0E",X"4B",X"3A",X"4F",X"44",X"44",X"24",X"0E",X"43",X"39",
		X"00",X"00",X"00",X"00",X"25",X"00",X"1C",X"50",X"18",X"40",X"36",X"42",X"44",X"49",X"44",X"24",
		X"00",X"00",X"00",X"00",X"20",X"00",X"1C",X"50",X"14",X"44",X"3F",X"3E",X"42",X"36",X"24",X"24",
		X"00",X"00",X"00",X"21",X"80",X"81",X"11",X"00",X"85",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"11",
		X"04",X"85",X"36",X"24",X"01",X"09",X"00",X"ED",X"B0",X"06",X"05",X"21",X"00",X"85",X"78",X"87",
		X"87",X"87",X"87",X"4F",X"C6",X"02",X"D7",X"11",X"02",X"85",X"1A",X"BE",X"38",X"23",X"20",X"0E",
		X"2D",X"1D",X"1A",X"BE",X"38",X"1B",X"20",X"06",X"2D",X"1D",X"1A",X"BE",X"38",X"13",X"21",X"00",
		X"85",X"79",X"D7",X"54",X"7D",X"C6",X"10",X"5F",X"C5",X"01",X"10",X"00",X"ED",X"B0",X"C1",X"10",
		X"CA",X"78",X"32",X"46",X"80",X"FE",X"05",X"CA",X"4E",X"06",X"21",X"10",X"85",X"07",X"07",X"07",
		X"07",X"D7",X"EB",X"21",X"00",X"85",X"01",X"10",X"00",X"ED",X"B0",X"CD",X"0B",X"10",X"CD",X"A1",
		X"12",X"26",X"19",X"3A",X"46",X"80",X"87",X"C6",X"18",X"6F",X"06",X"18",X"0E",X"B0",X"3E",X"1B",
		X"CD",X"5D",X"14",X"5D",X"16",X"0B",X"21",X"13",X"85",X"3A",X"46",X"80",X"87",X"87",X"87",X"87",
		X"85",X"6F",X"3E",X"0A",X"32",X"4D",X"80",X"3E",X"80",X"32",X"41",X"80",X"ED",X"53",X"50",X"80",
		X"22",X"52",X"80",X"F7",X"3A",X"00",X"A0",X"A7",X"20",X"78",X"3A",X"46",X"80",X"A7",X"28",X"02",
		X"3E",X"01",X"21",X"02",X"A0",X"D7",X"36",X"01",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",
		X"04",X"3A",X"21",X"80",X"D7",X"CB",X"66",X"28",X"41",X"CD",X"7F",X"12",X"2A",X"50",X"80",X"0E",
		X"C0",X"CD",X"4F",X"14",X"3A",X"01",X"80",X"4F",X"E6",X"07",X"C0",X"79",X"E6",X"1F",X"20",X"06",
		X"21",X"41",X"80",X"35",X"28",X"3C",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",X"04",X"3A",
		X"21",X"80",X"D7",X"7E",X"E6",X"0F",X"FE",X"02",X"28",X"38",X"FE",X"06",X"C0",X"2A",X"52",X"80",
		X"7E",X"3D",X"FE",X"09",X"20",X"02",X"3E",X"24",X"77",X"C9",X"CD",X"7F",X"12",X"77",X"23",X"22",
		X"52",X"80",X"2A",X"50",X"80",X"0E",X"C0",X"CD",X"4F",X"14",X"22",X"50",X"80",X"21",X"4D",X"80",
		X"35",X"C0",X"AF",X"32",X"02",X"A0",X"32",X"03",X"A0",X"32",X"16",X"A0",X"32",X"17",X"A0",X"C3",
		X"4E",X"06",X"2A",X"52",X"80",X"7E",X"3C",X"FE",X"25",X"20",X"02",X"3E",X"0A",X"77",X"C9",X"3A",
		X"20",X"80",X"A7",X"3A",X"16",X"80",X"28",X"0D",X"3A",X"21",X"80",X"A7",X"3A",X"16",X"80",X"28",
		X"04",X"0F",X"0F",X"0F",X"0F",X"0F",X"3E",X"00",X"38",X"02",X"3E",X"2C",X"2A",X"52",X"80",X"86",
		X"C9",X"21",X"09",X"15",X"11",X"CD",X"12",X"0E",X"C0",X"06",X"10",X"CD",X"1F",X"14",X"21",X"0C",
		X"16",X"11",X"DD",X"12",X"06",X"12",X"CD",X"1F",X"14",X"0E",X"B0",X"21",X"09",X"15",X"3E",X"1A",
		X"06",X"10",X"CD",X"5D",X"14",X"21",X"0C",X"16",X"06",X"12",X"C3",X"5D",X"14",X"0C",X"18",X"17",
		X"10",X"1B",X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"2C",X"0E",X"17",X"1D",
		X"0E",X"1B",X"24",X"22",X"18",X"1E",X"1B",X"24",X"12",X"17",X"12",X"1D",X"12",X"0A",X"15",X"21",
		X"00",X"12",X"11",X"C3",X"3E",X"06",X"0A",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"00",X"12",X"06",
		X"0A",X"3E",X"1F",X"0E",X"B0",X"CD",X"5D",X"14",X"C9",X"01",X"99",X"03",X"2B",X"71",X"10",X"FC",
		X"C9",X"11",X"82",X"81",X"CD",X"1A",X"13",X"11",X"C2",X"81",X"21",X"26",X"80",X"06",X"03",X"1A",
		X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"1A",X"77",X"1B",X"2B",X"10",X"FA",X"3A",
		X"21",X"80",X"3C",X"32",X"27",X"80",X"CD",X"63",X"14",X"C9",X"CD",X"27",X"14",X"CD",X"A9",X"13",
		X"3A",X"8C",X"81",X"A7",X"C0",X"ED",X"5B",X"89",X"81",X"2A",X"81",X"81",X"A7",X"ED",X"52",X"19",
		X"D8",X"3A",X"17",X"80",X"07",X"07",X"07",X"E6",X"03",X"28",X"02",X"3E",X"01",X"21",X"FB",X"13",
		X"CF",X"5E",X"23",X"56",X"EB",X"3A",X"17",X"80",X"2F",X"0F",X"0F",X"E6",X"07",X"CF",X"5E",X"23",
		X"56",X"2A",X"89",X"81",X"A7",X"ED",X"52",X"19",X"38",X"29",X"3A",X"17",X"80",X"2F",X"0F",X"0F",
		X"E6",X"07",X"FE",X"06",X"20",X"05",X"3E",X"01",X"32",X"8C",X"81",X"7D",X"83",X"27",X"6F",X"7C",
		X"8A",X"27",X"67",X"22",X"89",X"81",X"3A",X"83",X"81",X"3C",X"32",X"83",X"81",X"32",X"04",X"A0",
		X"C3",X"68",X"0F",X"ED",X"53",X"89",X"81",X"18",X"ED",X"21",X"81",X"81",X"7E",X"E6",X"F0",X"C8",
		X"0F",X"0F",X"0F",X"0F",X"4F",X"7E",X"E6",X"0F",X"C8",X"A1",X"C8",X"4F",X"2D",X"7E",X"E6",X"F0",
		X"C8",X"0F",X"0F",X"0F",X"0F",X"A1",X"C8",X"4F",X"7E",X"E6",X"0F",X"C8",X"A1",X"C8",X"3A",X"7E",
		X"79",X"FE",X"02",X"C0",X"21",X"CD",X"3E",X"11",X"E8",X"13",X"06",X"13",X"1A",X"07",X"2F",X"BE",
		X"C2",X"00",X"00",X"13",X"23",X"10",X"F5",X"C9",X"69",X"E8",X"EB",X"ED",X"7F",X"7B",X"FB",X"FE",
		X"ED",X"74",X"FA",X"F4",X"F9",X"F3",X"ED",X"75",X"71",X"79",X"D7",X"FF",X"13",X"0F",X"14",X"70",
		X"00",X"50",X"00",X"50",X"00",X"60",X"00",X"80",X"00",X"00",X"01",X"80",X"00",X"FF",X"FF",X"60",
		X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"70",X"00",X"80",X"00",X"60",X"00",X"FF",X"FF",X"1A",
		X"CD",X"4F",X"14",X"13",X"10",X"F9",X"C9",X"0E",X"C0",X"21",X"01",X"1B",X"11",X"01",X"08",X"3A",
		X"21",X"80",X"A7",X"28",X"01",X"EB",X"D5",X"11",X"82",X"81",X"CD",X"47",X"14",X"E1",X"3A",X"22",
		X"80",X"A7",X"28",X"15",X"11",X"C2",X"81",X"06",X"03",X"3E",X"05",X"CD",X"6D",X"14",X"AF",X"E5",
		X"F5",X"CD",X"9B",X"14",X"F1",X"77",X"E1",X"25",X"C9",X"3E",X"24",X"06",X"07",X"CD",X"4F",X"14",
		X"10",X"FB",X"C9",X"0E",X"C0",X"21",X"01",X"11",X"11",X"26",X"80",X"18",X"DA",X"C5",X"47",X"1A",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"07",X"05",X"3E",X"24",X"F2",X"81",X"14",X"AF",X"06",
		X"00",X"CD",X"4F",X"14",X"1A",X"E6",X"0F",X"20",X"07",X"05",X"3E",X"24",X"F2",X"92",X"14",X"AF",
		X"06",X"00",X"CD",X"4F",X"14",X"78",X"C1",X"1B",X"10",X"D3",X"C9",X"3A",X"03",X"80",X"25",X"A7",
		X"3E",X"04",X"28",X"03",X"25",X"3E",X"18",X"85",X"E6",X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",
		X"67",X"E6",X"C0",X"B5",X"6F",X"7C",X"E6",X"07",X"81",X"67",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",
		X"C0",X"21",X"02",X"00",X"22",X"46",X"79",X"21",X"02",X"80",X"22",X"44",X"79",X"21",X"14",X"20",
		X"22",X"44",X"7C",X"21",X"50",X"01",X"22",X"46",X"7C",X"21",X"00",X"25",X"22",X"46",X"7A",X"21",
		X"00",X"0F",X"22",X"46",X"7B",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"CF",X"3A",X"28",X"80",X"A7",
		X"20",X"05",X"3E",X"01",X"32",X"0E",X"A0",X"CD",X"FE",X"15",X"CD",X"C1",X"15",X"CD",X"B8",X"16",
		X"CD",X"45",X"16",X"D0",X"AF",X"32",X"0E",X"A0",X"32",X"22",X"A0",X"3A",X"28",X"80",X"A7",X"20",
		X"0B",X"21",X"BA",X"15",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"44",
		X"80",X"21",X"00",X"00",X"22",X"46",X"7D",X"21",X"C0",X"30",X"22",X"46",X"7C",X"F7",X"3A",X"2A",
		X"80",X"A7",X"20",X"87",X"3A",X"46",X"7D",X"3C",X"E6",X"07",X"32",X"46",X"7D",X"20",X"1F",X"3A",
		X"47",X"7D",X"3C",X"32",X"47",X"7D",X"FE",X"07",X"28",X"2A",X"FE",X"02",X"CC",X"A1",X"15",X"FE",
		X"04",X"CC",X"B1",X"15",X"FE",X"06",X"CC",X"A1",X"15",X"C6",X"30",X"32",X"47",X"7C",X"21",X"93",
		X"15",X"3A",X"47",X"7D",X"CF",X"3A",X"01",X"80",X"E6",X"0C",X"86",X"32",X"47",X"79",X"23",X"7E",
		X"32",X"46",X"7C",X"C9",X"3E",X"20",X"32",X"46",X"7D",X"AF",X"32",X"46",X"79",X"F7",X"21",X"46",
		X"7D",X"35",X"C0",X"21",X"8B",X"81",X"34",X"21",X"2A",X"80",X"36",X"01",X"AF",X"32",X"44",X"80",
		X"C3",X"BB",X"14",X"00",X"C0",X"00",X"C1",X"03",X"C4",X"03",X"C8",X"00",X"C2",X"00",X"C3",X"03",
		X"CC",X"21",X"47",X"7B",X"34",X"21",X"47",X"7A",X"35",X"F5",X"3E",X"2E",X"32",X"47",X"7C",X"F1",
		X"C9",X"21",X"47",X"7B",X"35",X"21",X"47",X"7A",X"34",X"C9",X"30",X"40",X"00",X"02",X"DF",X"10",
		X"10",X"2A",X"46",X"7A",X"3A",X"C6",X"7A",X"CF",X"11",X"00",X"12",X"A7",X"ED",X"52",X"19",X"30",
		X"01",X"EB",X"11",X"00",X"26",X"A7",X"ED",X"52",X"19",X"38",X"01",X"EB",X"22",X"46",X"7A",X"2A",
		X"46",X"7B",X"3A",X"C6",X"7B",X"CF",X"11",X"00",X"02",X"A7",X"ED",X"52",X"19",X"30",X"01",X"EB",
		X"11",X"00",X"1C",X"A7",X"ED",X"52",X"19",X"38",X"01",X"EB",X"22",X"46",X"7B",X"C9",X"3A",X"28",
		X"80",X"A7",X"20",X"1E",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",X"04",X"3A",X"21",X"80",
		X"D7",X"7E",X"E6",X"0F",X"21",X"33",X"16",X"CF",X"7E",X"32",X"C6",X"7A",X"23",X"7E",X"32",X"C6",
		X"7B",X"C9",X"3A",X"01",X"80",X"E6",X"0F",X"C0",X"CD",X"4B",X"0F",X"E6",X"0F",X"FE",X"09",X"30",
		X"F7",X"18",X"E1",X"F0",X"00",X"F0",X"F0",X"00",X"E8",X"10",X"F0",X"10",X"00",X"10",X"10",X"00",
		X"18",X"F0",X"10",X"00",X"00",X"ED",X"5B",X"46",X"82",X"3A",X"47",X"83",X"1F",X"CB",X"1A",X"FD",
		X"21",X"4E",X"79",X"06",X"19",X"CD",X"70",X"16",X"D8",X"FD",X"2C",X"FD",X"2C",X"10",X"F6",X"FD",
		X"21",X"20",X"79",X"06",X"10",X"CD",X"95",X"16",X"D8",X"FD",X"2C",X"FD",X"2C",X"10",X"F6",X"C9",
		X"3E",X"02",X"FD",X"BE",X"00",X"20",X"1C",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",
		X"96",X"D6",X"08",X"C6",X"10",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"04",
		X"C6",X"08",X"C9",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"F7",X"3E",X"09",X"FD",X"84",
		X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"1C",X"C6",X"28",X"D0",X"2C",X"24",X"7E",X"1F",X"25",
		X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"3A",X"42",X"79",X"FE",X"02",X"28",X"02",X"3E",
		X"01",X"C6",X"1F",X"4F",X"06",X"00",X"3A",X"01",X"80",X"E6",X"04",X"28",X"1B",X"ED",X"5B",X"44",
		X"82",X"3A",X"45",X"83",X"1F",X"CB",X"1A",X"FD",X"21",X"04",X"79",X"06",X"0E",X"CD",X"04",X"17",
		X"38",X"1C",X"FD",X"2C",X"FD",X"2C",X"10",X"F5",X"79",X"80",X"32",X"45",X"7C",X"3E",X"F4",X"2A",
		X"46",X"7A",X"84",X"67",X"22",X"44",X"7A",X"2A",X"46",X"7B",X"22",X"44",X"7B",X"C9",X"06",X"09",
		X"18",X"E6",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"F7",X"3E",X"09",X"FD",X"84",X"67",
		X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"0A",X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",
		X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"21",X"14",X"01",
		X"22",X"32",X"80",X"AF",X"32",X"30",X"80",X"21",X"A2",X"17",X"22",X"48",X"78",X"21",X"48",X"78",
		X"11",X"4A",X"78",X"01",X"04",X"00",X"ED",X"B0",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"D8",X"3A",
		X"44",X"80",X"A7",X"CC",X"72",X"17",X"DD",X"E5",X"DD",X"21",X"48",X"78",X"06",X"03",X"DD",X"5D",
		X"DD",X"54",X"CD",X"54",X"04",X"DD",X"2C",X"DD",X"2C",X"10",X"F3",X"DD",X"E1",X"AF",X"32",X"30",
		X"80",X"C9",X"3A",X"28",X"80",X"A7",X"20",X"23",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",
		X"04",X"3A",X"21",X"80",X"D7",X"CB",X"6E",X"21",X"33",X"80",X"28",X"03",X"36",X"01",X"C9",X"35",
		X"C0",X"3A",X"32",X"80",X"77",X"3E",X"01",X"32",X"30",X"80",X"C9",X"CD",X"4B",X"0F",X"E6",X"0F",
		X"18",X"E5",X"F7",X"EB",X"4C",X"11",X"30",X"80",X"1A",X"3D",X"C0",X"12",X"24",X"36",X"02",X"CB",
		X"FD",X"36",X"02",X"24",X"36",X"A0",X"3C",X"32",X"0B",X"A0",X"ED",X"5B",X"46",X"7A",X"CB",X"BD",
		X"73",X"2C",X"72",X"ED",X"5B",X"46",X"7B",X"24",X"72",X"2D",X"73",X"61",X"EB",X"F7",X"EB",X"C5",
		X"E5",X"CD",X"28",X"19",X"E1",X"C1",X"3A",X"01",X"80",X"F5",X"F5",X"E6",X"01",X"07",X"07",X"07",
		X"24",X"4C",X"2C",X"C6",X"80",X"77",X"F1",X"0F",X"E6",X"01",X"C6",X"23",X"24",X"24",X"24",X"77",
		X"F1",X"0F",X"0F",X"E6",X"01",X"C6",X"16",X"2D",X"77",X"61",X"7E",X"FE",X"03",X"28",X"0E",X"24",
		X"CD",X"4B",X"18",X"7A",X"FE",X"28",X"D8",X"25",X"2D",X"36",X"00",X"18",X"95",X"24",X"CB",X"FD",
		X"36",X"18",X"CB",X"BD",X"2C",X"24",X"24",X"36",X"23",X"2D",X"24",X"36",X"FF",X"F7",X"21",X"00",
		X"05",X"7C",X"DD",X"84",X"67",X"7D",X"DD",X"85",X"6F",X"34",X"7E",X"25",X"4C",X"25",X"25",X"25",
		X"FE",X"08",X"28",X"D5",X"F5",X"0F",X"E6",X"03",X"C6",X"18",X"61",X"77",X"F1",X"E6",X"01",X"07",
		X"07",X"07",X"25",X"25",X"25",X"2C",X"C6",X"80",X"77",X"2D",X"24",X"5E",X"2C",X"56",X"2D",X"CB",
		X"FD",X"EB",X"1A",X"CF",X"EB",X"CB",X"BD",X"73",X"2C",X"72",X"C9",X"CD",X"4B",X"0F",X"A7",X"C0",
		X"18",X"2A",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"44",X"80",X"A7",X"C0",X"3A",X"28",X"80",
		X"A7",X"20",X"E8",X"3A",X"20",X"80",X"A7",X"3A",X"16",X"80",X"28",X"0D",X"3A",X"21",X"80",X"A7",
		X"3A",X"16",X"80",X"28",X"04",X"0F",X"0F",X"0F",X"0F",X"0F",X"D8",X"F7",X"3A",X"40",X"79",X"FE",
		X"01",X"C0",X"F7",X"2A",X"46",X"7A",X"22",X"42",X"7A",X"3E",X"F4",X"84",X"67",X"22",X"40",X"7A",
		X"2A",X"46",X"7B",X"22",X"42",X"7B",X"22",X"40",X"7B",X"AF",X"32",X"C2",X"7A",X"32",X"42",X"7D",
		X"32",X"43",X"7D",X"3C",X"32",X"0C",X"A0",X"21",X"02",X"80",X"22",X"42",X"79",X"22",X"40",X"79",
		X"3E",X"1C",X"32",X"42",X"7C",X"21",X"14",X"22",X"22",X"40",X"7C",X"F7",X"21",X"42",X"7D",X"34",
		X"7E",X"E6",X"07",X"20",X"0C",X"2C",X"7E",X"FE",X"02",X"28",X"06",X"3C",X"77",X"25",X"2D",X"34",
		X"24",X"7E",X"0F",X"0F",X"E6",X"03",X"C6",X"25",X"32",X"43",X"7C",X"21",X"C2",X"7A",X"35",X"35",
		X"7E",X"2A",X"42",X"7A",X"CF",X"22",X"42",X"7A",X"2A",X"40",X"7A",X"3A",X"14",X"80",X"ED",X"44",
		X"CF",X"22",X"40",X"7A",X"CD",X"0B",X"19",X"D8",X"C3",X"62",X"18",X"2A",X"40",X"7A",X"ED",X"5B",
		X"42",X"7A",X"A7",X"ED",X"52",X"D8",X"AF",X"32",X"0C",X"A0",X"32",X"20",X"A0",X"CD",X"EE",X"19",
		X"AF",X"32",X"42",X"79",X"32",X"40",X"79",X"C9",X"3E",X"0A",X"DD",X"84",X"57",X"DD",X"5D",X"EB",
		X"5E",X"2C",X"56",X"24",X"7E",X"1F",X"CB",X"1A",X"FD",X"21",X"74",X"79",X"06",X"06",X"CD",X"A6",
		X"19",X"30",X"2F",X"FD",X"36",X"00",X"03",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"CB",X"FF",X"6F",
		X"36",X"00",X"3A",X"28",X"80",X"A7",X"20",X"1A",X"3E",X"03",X"FD",X"84",X"67",X"FD",X"7D",X"CB",
		X"FF",X"6F",X"7E",X"21",X"31",X"3D",X"D7",X"D5",X"C5",X"EB",X"E7",X"C1",X"D1",X"3E",X"01",X"32",
		X"05",X"A0",X"FD",X"2C",X"FD",X"2C",X"10",X"C6",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"CB",X"FF",
		X"6F",X"7E",X"CB",X"BD",X"77",X"FD",X"21",X"20",X"79",X"06",X"10",X"CD",X"CB",X"19",X"38",X"07",
		X"FD",X"2C",X"FD",X"2C",X"10",X"F5",X"C9",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"6F",X"36",X"03",
		X"3E",X"01",X"32",X"0A",X"A0",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"1C",X"3E",X"09",X"FD",
		X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"10",X"C6",X"20",X"D0",X"2C",X"24",X"7E",X"1F",
		X"25",X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",
		X"20",X"F7",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"18",X"C6",X"20",
		X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"ED",X"5B",
		X"40",X"82",X"3A",X"41",X"83",X"1F",X"CB",X"1A",X"FD",X"21",X"00",X"79",X"06",X"10",X"D5",X"CD",
		X"3D",X"1A",X"30",X"28",X"FD",X"36",X"00",X"03",X"3A",X"28",X"80",X"A7",X"20",X"1E",X"3E",X"03",
		X"FD",X"84",X"67",X"FD",X"7D",X"CB",X"FF",X"6F",X"7E",X"21",X"31",X"3D",X"D7",X"EB",X"C5",X"E7",
		X"21",X"36",X"1A",X"11",X"90",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C1",X"D1",X"FD",X"2C",X"FD",
		X"2C",X"10",X"CB",X"C9",X"A7",X"C9",X"40",X"40",X"40",X"01",X"FF",X"20",X"20",X"3E",X"02",X"FD",
		X"BE",X"00",X"20",X"F0",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"0A",
		X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",
		X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"36",X"07",X"2D",X"36",
		X"17",X"CB",X"FD",X"36",X"0F",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",
		X"31",X"EB",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",
		X"2C",X"5D",X"36",X"03",X"2C",X"36",X"02",X"2C",X"36",X"00",X"24",X"36",X"01",X"24",X"16",X"7B",
		X"1A",X"3D",X"77",X"2D",X"1D",X"1A",X"77",X"24",X"36",X"17",X"2C",X"36",X"07",X"2D",X"CB",X"FD",
		X"36",X"1B",X"CB",X"BD",X"2D",X"2D",X"36",X"48",X"2C",X"2C",X"26",X"78",X"11",X"DD",X"1A",X"73",
		X"2C",X"72",X"11",X"CB",X"1A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",X"1C",
		X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",
		X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"16",X"32",X"EB",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",
		X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"2D",X"36",X"1F",X"CB",
		X"FD",X"36",X"15",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"11",X"26",X"7C",
		X"2C",X"3A",X"1C",X"80",X"77",X"EB",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"3A",
		X"88",X"81",X"D6",X"02",X"30",X"01",X"AF",X"32",X"88",X"81",X"C3",X"86",X"31",X"16",X"7E",X"DD",
		X"5D",X"3A",X"A3",X"81",X"12",X"16",X"79",X"18",X"10",X"16",X"7E",X"DD",X"5D",X"3A",X"B0",X"81",
		X"12",X"16",X"79",X"18",X"04",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",
		X"7C",X"2D",X"36",X"2C",X"CB",X"FD",X"36",X"1B",X"CB",X"BD",X"26",X"7E",X"CD",X"4B",X"0F",X"A6",
		X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",
		X"7A",X"2C",X"3A",X"B1",X"81",X"BE",X"38",X"64",X"2D",X"26",X"7D",X"3A",X"01",X"80",X"E6",X"07",
		X"20",X"37",X"35",X"20",X"34",X"11",X"8E",X"1B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",X"7D",X"34",X"7E",X"FE",X"0C",X"20",
		X"06",X"E5",X"CD",X"87",X"32",X"E1",X"7E",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1A",X"EB",
		X"21",X"F9",X"1B",X"D7",X"15",X"7E",X"12",X"14",X"EB",X"2C",X"25",X"3A",X"1C",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"24",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",
		X"77",X"11",X"64",X"1B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"18",X"DD",X"11",X"E5",X"1B",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",
		X"EB",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"2D",X"2E",X"2F",X"2E",X"2D",X"2C",
		X"16",X"7E",X"DD",X"5D",X"3A",X"A0",X"81",X"12",X"16",X"79",X"18",X"10",X"16",X"7E",X"DD",X"5D",
		X"3A",X"B0",X"81",X"12",X"16",X"79",X"18",X"04",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7C",X"2D",X"36",X"27",X"CB",X"FD",X"36",X"30",X"CB",X"BD",X"26",X"7E",X"CD",
		X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"86",X"31",X"26",X"7D",X"16",X"7A",X"5D",X"1C",X"1A",X"4F",X"3A",X"B1",X"81",X"B9",X"D4",X"71",
		X"32",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",
		X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"5D",X"36",X"03",X"2C",X"36",X"02",X"2C",
		X"36",X"00",X"24",X"36",X"01",X"24",X"16",X"7B",X"1A",X"3D",X"77",X"2D",X"1D",X"1A",X"77",X"24",
		X"36",X"27",X"CB",X"FD",X"36",X"36",X"CB",X"BD",X"2D",X"2D",X"36",X"44",X"2C",X"2C",X"26",X"7E",
		X"3A",X"A0",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",X"78",X"11",X"BE",X"1C",
		X"73",X"2C",X"72",X"11",X"AC",X"1C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",
		X"1C",X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"16",X"32",X"26",X"7D",X"CD",X"71",X"32",X"25",X"2C",
		X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"C5",X"16",
		X"78",X"DD",X"5D",X"D5",X"21",X"47",X"1D",X"01",X"0A",X"00",X"ED",X"B0",X"D1",X"14",X"D5",X"6B",
		X"62",X"36",X"02",X"2C",X"36",X"00",X"2C",X"EB",X"01",X"08",X"00",X"ED",X"B0",X"D1",X"D5",X"CB",
		X"FB",X"7B",X"C6",X"08",X"EB",X"E5",X"77",X"2C",X"36",X"7C",X"2C",X"EB",X"E1",X"01",X"06",X"00",
		X"ED",X"B0",X"D1",X"14",X"D5",X"21",X"51",X"1D",X"01",X"0A",X"00",X"ED",X"B0",X"D1",X"14",X"EB",
		X"4E",X"2C",X"46",X"2C",X"3E",X"80",X"81",X"F5",X"77",X"2C",X"70",X"F1",X"30",X"01",X"34",X"34",
		X"2C",X"79",X"D6",X"80",X"F5",X"77",X"2C",X"70",X"F1",X"30",X"01",X"35",X"35",X"2C",X"71",X"2C",
		X"70",X"2C",X"71",X"2C",X"70",X"C1",X"C9",X"9E",X"1D",X"9E",X"1D",X"9E",X"1D",X"9E",X"1D",X"5B",
		X"1D",X"00",X"00",X"80",X"01",X"80",X"01",X"00",X"03",X"80",X"01",X"16",X"7C",X"DD",X"5D",X"EB",
		X"36",X"3A",X"CB",X"FD",X"36",X"36",X"11",X"6F",X"1D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",
		X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"11",X"26",X"7C",X"2C",X"3A",X"1C",X"80",X"77",
		X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"54",X"5D",X"3E",X"03",X"2D",X"2D",
		X"77",X"2D",X"2D",X"77",X"2D",X"2D",X"77",X"2D",X"2D",X"77",X"EB",X"C3",X"86",X"31",X"16",X"7C",
		X"DD",X"5D",X"EB",X"26",X"7C",X"36",X"2C",X"CB",X"FD",X"36",X"1B",X"CB",X"BD",X"26",X"7E",X"3A",
		X"A5",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",
		X"7E",X"FE",X"03",X"28",X"59",X"26",X"7A",X"2C",X"3A",X"B1",X"81",X"BE",X"38",X"70",X"2D",X"26",
		X"7D",X"3A",X"01",X"80",X"E6",X"07",X"20",X"36",X"35",X"20",X"33",X"11",X"E4",X"1D",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"30",X"26",X"7D",
		X"34",X"7E",X"FE",X"0C",X"20",X"06",X"E5",X"CD",X"87",X"32",X"E1",X"7E",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"27",X"EB",X"21",X"5A",X"1E",X"D7",X"15",X"7E",X"12",X"14",X"EB",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"E5",X"CB",
		X"FD",X"5E",X"2C",X"56",X"EB",X"36",X"24",X"E1",X"C3",X"86",X"31",X"24",X"CD",X"4B",X"0F",X"A6",
		X"3C",X"25",X"77",X"11",X"BB",X"1D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"18",X"D0",X"11",X"47",
		X"1E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",
		X"CD",X"EB",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"2D",X"2E",X"2F",X"2E",X"2D",
		X"2C",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"2D",X"26",X"7C",X"36",X"00",
		X"CB",X"FD",X"36",X"36",X"F7",X"16",X"79",X"DD",X"5D",X"1A",X"FE",X"03",X"28",X"07",X"14",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"EB",X"26",X"7D",X"36",X"FF",X"11",X"93",X"1E",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"24",X"FE",X"04",X"20",X"08",X"26",X"79",X"2C",X"36",X"03",X"2D",X"26",X"7D",
		X"25",X"EB",X"21",X"F1",X"1E",X"D7",X"7E",X"EB",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",
		X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"79",X"36",X"02",X"11",X"D5",X"1E",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",
		X"EB",X"1C",X"16",X"7C",X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",
		X"30",X"A8",X"A9",X"AA",X"AB",X"AE",X"B2",X"B6",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"26",
		X"7C",X"36",X"15",X"2C",X"36",X"26",X"2D",X"CB",X"FD",X"36",X"21",X"F7",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"24",X"2C",X"3A",X"47",X"7A",X"BE",X"CB",X"FD",X"3E",X"00",X"38",X"35",X"28",
		X"02",X"3C",X"3C",X"77",X"CB",X"BD",X"24",X"3A",X"47",X"7B",X"BE",X"3E",X"00",X"38",X"29",X"28",
		X"02",X"3C",X"3C",X"2D",X"CB",X"FD",X"86",X"77",X"25",X"2C",X"7E",X"2D",X"86",X"77",X"CB",X"BD",
		X"26",X"79",X"2C",X"3A",X"01",X"80",X"E6",X"0C",X"C6",X"80",X"77",X"2D",X"24",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"3D",X"3D",X"18",X"CB",X"3D",X"3D",X"18",X"D7",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7B",X"CD",X"98",X"33",X"24",X"2D",X"36",X"00",X"CB",
		X"FD",X"36",X"30",X"11",X"7C",X"1F",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"1A",X"FE",X"03",X"28",X"08",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"EB",X"2C",X"36",
		X"80",X"26",X"7C",X"36",X"0E",X"2D",X"36",X"1F",X"F7",X"CD",X"D6",X"1F",X"38",X"0A",X"16",X"7A",
		X"DD",X"5D",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"3A",X"16",X"80",X"CB",X"4F",X"20",X"08",X"11",
		X"70",X"3D",X"C5",X"E7",X"C1",X"18",X"0C",X"3A",X"83",X"81",X"3C",X"32",X"83",X"81",X"C5",X"CD",
		X"68",X"0F",X"C1",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"00",X"26",X"7F",X"36",X"00",X"3E",X"01",
		X"32",X"0D",X"A0",X"C3",X"79",X"30",X"16",X"82",X"DD",X"5D",X"EB",X"ED",X"5B",X"46",X"82",X"3A",
		X"47",X"83",X"1F",X"CB",X"1A",X"7B",X"96",X"D6",X"0A",X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",
		X"25",X"7E",X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"CD",X"A7",X"20",X"F7",X"CD",X"CB",X"20",X"38",X"1A",X"24",X"3A",X"1C",X"80",X"77",X"2D",X"26",
		X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"A7",X"20",X"F7",X"CD",X"CB",X"20",X"38",
		X"71",X"18",X"E6",X"D6",X"02",X"38",X"38",X"11",X"30",X"20",X"DD",X"73",X"00",X"DD",X"72",X"01",
		X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",
		X"E6",X"07",X"EB",X"21",X"9F",X"20",X"D7",X"EB",X"25",X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",
		X"2D",X"25",X"CB",X"FD",X"35",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"11",
		X"68",X"20",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",
		X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"E6",X"07",X"C6",X"08",X"25",X"77",X"2C",X"3A",
		X"1C",X"80",X"77",X"2D",X"25",X"CB",X"FD",X"34",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",
		X"79",X"30",X"E5",X"F5",X"CD",X"87",X"32",X"F1",X"E1",X"D6",X"02",X"38",X"C2",X"18",X"88",X"0F",
		X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"06",X"CB",X"BD",X"36",X"08",X"24",X"36",X"00",X"C9",X"16",X"79",X"DD",X"5D",X"EB",
		X"7E",X"FE",X"03",X"CA",X"E2",X"20",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"02",X"C6",
		X"04",X"C9",X"33",X"33",X"C3",X"1F",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"8B",X"33",X"EB",X"15",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"09",X"CB",X"BD",X"36",X"10",X"24",X"CD",X"4B",X"0F",X"E6",X"3F",X"C6",X"40",X"77",
		X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"35",X"28",
		X"10",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"E5",X"CD",X"87",X"32",X"E1",X"11",X"3F",X"21",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",
		X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"0F",
		X"E6",X"0F",X"FE",X"07",X"28",X"13",X"C6",X"10",X"25",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"26",X"7A",X"EB",X"1A",X"4F",X"3A",
		X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",X"CB",
		X"FB",X"1D",X"21",X"B3",X"3D",X"C6",X"80",X"CD",X"7E",X"33",X"EB",X"CB",X"BD",X"26",X"78",X"11",
		X"95",X"21",X"73",X"2C",X"72",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",
		X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"24",X"36",X"28",X"24",X"CD",
		X"98",X"33",X"18",X"0F",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7B",
		X"CD",X"8B",X"33",X"25",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",X"7C",X"36",X"0F",
		X"CB",X"BD",X"26",X"7E",X"3A",X"A4",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",
		X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"3A",X"01",X"80",
		X"E6",X"07",X"20",X"1A",X"35",X"20",X"17",X"E5",X"CD",X"4B",X"0F",X"24",X"A6",X"3C",X"25",X"77",
		X"26",X"7A",X"2C",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"CD",X"87",X"32",X"E1",X"25",X"3A",
		X"01",X"80",X"E6",X"03",X"C6",X"28",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",
		X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",X"7C",
		X"36",X"0C",X"CB",X"BD",X"26",X"7E",X"3A",X"A4",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",
		X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"3A",
		X"01",X"80",X"E6",X"07",X"20",X"1E",X"35",X"20",X"1B",X"E5",X"CD",X"4B",X"0F",X"24",X"A6",X"3C",
		X"25",X"77",X"26",X"7B",X"CB",X"FD",X"EB",X"CD",X"4B",X"0F",X"21",X"33",X"3E",X"CD",X"7E",X"33",
		X"CD",X"87",X"32",X"E1",X"25",X"3A",X"01",X"80",X"E6",X"03",X"C6",X"28",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"68",X"23",X"F7",
		X"CD",X"8C",X"23",X"38",X"0F",X"24",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"D6",X"06",X"38",X"56",X"11",X"D1",X"22",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",
		X"0F",X"E6",X"07",X"FE",X"06",X"20",X"02",X"AF",X"77",X"EB",X"21",X"5C",X"23",X"D7",X"EB",X"25",
		X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"25",X"CB",X"FD",X"35",X"CB",X"BD",X"25",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"68",X"23",X"F7",X"CD",X"8C",X"23",X"38",X"02",X"18",
		X"A4",X"E5",X"F5",X"CD",X"87",X"32",X"F1",X"E1",X"D6",X"06",X"38",X"02",X"18",X"AA",X"11",X"27",
		X"23",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"E6",X"07",X"FE",X"06",X"20",X"02",X"AF",X"77",X"EB",
		X"21",X"62",X"23",X"D7",X"EB",X"25",X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"25",X"CB",
		X"FD",X"34",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"A5",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"B3",X"3D",X"CD",X"65",X"33",X"EB",
		X"26",X"7C",X"36",X"12",X"CB",X"BD",X"36",X"A0",X"24",X"36",X"00",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"A3",X"23",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"06",
		X"C6",X"0C",X"C9",X"33",X"33",X"C3",X"1F",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"EB",
		X"26",X"7C",X"36",X"1B",X"CB",X"BD",X"36",X"20",X"24",X"CD",X"4B",X"0F",X"E6",X"3F",X"C6",X"30",
		X"77",X"24",X"3A",X"A1",X"81",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"2C",X"36",X"00",X"26",X"7B",X"3A",X"47",X"7B",X"BE",
		X"3E",X"01",X"38",X"02",X"3E",X"FF",X"CB",X"FD",X"77",X"CB",X"BD",X"2D",X"26",X"7D",X"36",X"01",
		X"CD",X"71",X"32",X"11",X"1C",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"34",X"7E",X"0F",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1D",X"C6",X"20",X"2D",X"25",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",X"EB",X"CD",
		X"91",X"30",X"C3",X"79",X"30",X"11",X"5E",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"B3",X"3D",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"27",X"CB",X"BD",X"36",X"01",X"26",X"7E",X"3A",X"A2",X"81",X"77",X"CD",X"4B",X"0F",
		X"A6",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",
		X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"04",X"C6",X"08",X"38",X"16",X"2D",X"26",X"7D",X"CD",
		X"71",X"32",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",
		X"79",X"30",X"D6",X"04",X"3E",X"02",X"38",X"02",X"3E",X"FE",X"CB",X"FD",X"77",X"CB",X"BD",X"26",
		X"7D",X"36",X"FF",X"11",X"FC",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"34",X"7E",X"0F",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1D",X"C6",X"01",X"2D",X"25",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",X"EB",X"CD",
		X"91",X"30",X"C3",X"79",X"30",X"11",X"3E",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"0F",X"25",X"36",X"00",X"25",
		X"36",X"10",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",X"4B",
		X"0F",X"E6",X"FF",X"3C",X"77",X"25",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",X"02",
		X"11",X"99",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",
		X"03",X"CA",X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"36",X"FF",X"26",X"79",X"36",X"03",X"CD",
		X"87",X"32",X"11",X"CB",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"A8",X"27",X"D2",X"9D",
		X"27",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"15",X"25",X"36",X"00",X"25",
		X"36",X"10",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7C",
		X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",X"02",X"11",X"03",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7B",
		X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"38",X"9B",X"25",X"2C",
		X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",
		X"28",X"36",X"12",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",
		X"4B",X"0F",X"E6",X"3F",X"3C",X"77",X"25",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",
		X"02",X"2C",X"24",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"11",X"63",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",
		X"35",X"CA",X"B9",X"25",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"1B",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"26",X"7C",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",
		X"02",X"2C",X"24",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"11",X"B3",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7B",
		X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"DA",X"B9",X"25",X"25",
		X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",
		X"26",X"28",X"36",X"24",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",
		X"CD",X"4B",X"0F",X"E6",X"3F",X"3C",X"77",X"25",X"36",X"12",X"2C",X"26",X"7A",X"EB",X"21",X"F3",
		X"3D",X"CD",X"65",X"33",X"EB",X"CB",X"BD",X"25",X"36",X"02",X"2C",X"36",X"80",X"11",X"16",X"27",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",
		X"31",X"26",X"7D",X"35",X"28",X"6B",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"33",X"F7",X"CD",X"E7",X"27",X"30",
		X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"25",X"36",X"12",X"2C",X"26",X"7A",X"EB",X"21",X"F3",
		X"3D",X"CD",X"65",X"33",X"EB",X"CB",X"BD",X"25",X"36",X"02",X"2C",X"36",X"80",X"11",X"66",X"27",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",
		X"31",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"38",
		X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"36",X"FF",X"26",X"79",X"36",X"03",X"CD",X"D9",X"32",X"C3",X"C2",X"25",X"26",X"7F",X"36",
		X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",
		X"10",X"20",X"09",X"2C",X"26",X"7A",X"35",X"24",X"34",X"2D",X"26",X"7D",X"4F",X"0F",X"0F",X"E6",
		X"07",X"FE",X"05",X"D0",X"EB",X"21",X"DB",X"27",X"CF",X"15",X"7E",X"12",X"23",X"1C",X"16",X"79",
		X"79",X"07",X"07",X"E6",X"0C",X"86",X"12",X"1D",X"14",X"37",X"C9",X"04",X"80",X"05",X"80",X"06",
		X"80",X"07",X"80",X"08",X"83",X"0C",X"83",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",X"08",
		X"20",X"09",X"2C",X"26",X"7A",X"34",X"24",X"35",X"2D",X"26",X"7D",X"4F",X"0F",X"0F",X"E6",X"07",
		X"FE",X"05",X"D0",X"EB",X"21",X"1A",X"28",X"CF",X"15",X"7E",X"12",X"23",X"1C",X"16",X"79",X"79",
		X"07",X"07",X"E6",X"0C",X"86",X"12",X"1D",X"14",X"37",X"C9",X"0C",X"83",X"08",X"83",X"07",X"80",
		X"06",X"80",X"05",X"80",X"04",X"80",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"24",X"CD",
		X"4B",X"0F",X"E6",X"0F",X"C6",X"05",X"77",X"24",X"CD",X"8B",X"33",X"34",X"24",X"36",X"24",X"2D",
		X"24",X"36",X"FF",X"25",X"CB",X"FD",X"3E",X"01",X"32",X"09",X"A0",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"80",X"26",X"7B",X"CD",X"8B",X"33",X"24",X"2D",X"36",X"13",X"CB",
		X"FD",X"36",X"30",X"26",X"7A",X"36",X"30",X"24",X"36",X"00",X"CB",X"BD",X"26",X"7D",X"CD",X"4B",
		X"0F",X"E6",X"1F",X"C6",X"20",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"E5",X"CD",X"0A",X"33",X"3E",X"01",X"32",X"06",X"A0",
		X"C5",X"21",X"B9",X"28",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C1",X"E1",X"26",X"7F",
		X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"30",X"80",X"80",X"01",X"FF",X"10",X"10",
		X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"EB",X"21",X"D9",X"28",X"3A",X"01",X"80",X"0F",X"E6",
		X"03",X"D7",X"7E",X"12",X"16",X"7A",X"C3",X"FC",X"30",X"32",X"33",X"30",X"31",X"16",X"79",X"DD",
		X"5D",X"EB",X"36",X"03",X"2C",X"36",X"00",X"26",X"7B",X"36",X"1E",X"F7",X"16",X"7A",X"DD",X"5D",
		X"1C",X"1A",X"4F",X"3A",X"47",X"7A",X"D6",X"02",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",
		X"D6",X"02",X"91",X"67",X"CD",X"B2",X"0E",X"CB",X"FB",X"1D",X"21",X"73",X"3D",X"CD",X"7E",X"33",
		X"CB",X"BB",X"1C",X"EB",X"3A",X"47",X"7A",X"D6",X"02",X"BE",X"20",X"A4",X"24",X"3A",X"47",X"7B",
		X"D6",X"02",X"BE",X"20",X"9B",X"11",X"2E",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",
		X"80",X"A7",X"20",X"06",X"3A",X"2E",X"80",X"A7",X"20",X"16",X"CD",X"F7",X"29",X"14",X"21",X"D9",
		X"28",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"C9",
		X"11",X"59",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"F7",X"29",X"3A",X"01",X"80",X"0F",
		X"0F",X"E6",X"07",X"FE",X"07",X"28",X"14",X"21",X"74",X"29",X"D7",X"14",X"7E",X"12",X"1C",X"3A",
		X"1C",X"80",X"12",X"C9",X"32",X"32",X"32",X"32",X"34",X"35",X"36",X"16",X"7D",X"EB",X"36",X"E0",
		X"11",X"89",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"28",
		X"20",X"EB",X"2A",X"46",X"7B",X"1A",X"D5",X"EF",X"D1",X"16",X"7B",X"EB",X"73",X"2C",X"72",X"ED",
		X"5B",X"46",X"7A",X"25",X"15",X"15",X"72",X"2D",X"73",X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",
		X"C9",X"26",X"7A",X"ED",X"5B",X"46",X"7A",X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",
		X"7B",X"72",X"2D",X"73",X"CB",X"FD",X"36",X"00",X"25",X"36",X"A0",X"3E",X"01",X"32",X"08",X"A0",
		X"11",X"D9",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",X"21",X"D9",X"28",
		X"3A",X"01",X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"1D",X"16",
		X"7A",X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"7A",X"DD",X"5D",X"EB",X"ED",X"5B",X"46",X"7A",
		X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",X"7B",X"15",X"15",X"72",X"2D",X"73",X"EB",
		X"C9",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"EB",X"21",X"2A",X"2A",X"3A",X"01",X"80",X"0F",
		X"E6",X"03",X"D7",X"7E",X"12",X"16",X"7A",X"C3",X"FC",X"30",X"32",X"31",X"30",X"33",X"16",X"79",
		X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"36",X"00",X"F7",X"16",X"7A",X"DD",X"5D",X"1C",X"1A",X"4F",
		X"3A",X"47",X"7A",X"D6",X"02",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"C6",X"02",X"91",
		X"67",X"CD",X"B2",X"0E",X"CB",X"FB",X"1D",X"21",X"73",X"3D",X"CD",X"7E",X"33",X"CB",X"BB",X"1C",
		X"EB",X"3A",X"47",X"7A",X"D6",X"02",X"BE",X"20",X"A8",X"24",X"3A",X"47",X"7B",X"C6",X"02",X"BE",
		X"20",X"9F",X"11",X"7B",X"2A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",X"80",X"A7",X"20",
		X"06",X"3A",X"2E",X"80",X"A7",X"20",X"16",X"CD",X"09",X"2B",X"14",X"21",X"2A",X"2A",X"3A",X"01",
		X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"C9",X"11",X"A6",X"2A",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"09",X"2B",X"3A",X"01",X"80",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"14",X"21",X"C1",X"2A",X"D7",X"14",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",
		X"C9",X"32",X"32",X"32",X"32",X"37",X"38",X"39",X"16",X"7D",X"EB",X"36",X"20",X"11",X"D6",X"2A",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"35",X"28",X"20",X"EB",X"2A",
		X"46",X"7B",X"1A",X"D5",X"EF",X"D1",X"16",X"7B",X"EB",X"73",X"2C",X"72",X"ED",X"5B",X"46",X"7A",
		X"15",X"15",X"25",X"72",X"2D",X"73",X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"C9",X"26",X"7F",
		X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"16",X"7A",X"DD",X"5D",X"EB",X"ED",X"5B",
		X"46",X"7A",X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",X"7B",X"14",X"14",X"72",X"2D",
		X"73",X"EB",X"C9",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"82",X"24",X"2D",X"CB",
		X"FD",X"36",X"10",X"CB",X"BD",X"24",X"2C",X"CD",X"8B",X"33",X"34",X"F7",X"16",X"7A",X"DD",X"5D",
		X"EB",X"E5",X"7E",X"2C",X"17",X"7E",X"17",X"E6",X"07",X"EB",X"21",X"5D",X"2B",X"CF",X"7E",X"16",
		X"7C",X"12",X"23",X"7E",X"1D",X"12",X"D1",X"CD",X"D4",X"30",X"C3",X"79",X"30",X"2B",X"20",X"2C",
		X"21",X"2B",X"24",X"2C",X"25",X"2B",X"28",X"2C",X"29",X"2B",X"2C",X"2C",X"2D",X"16",X"7A",X"DD",
		X"5D",X"1C",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"F7",X"16",X"7A",X"DD",X"5D",X"CD",X"91",X"30",
		X"C3",X"79",X"30",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"15",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",
		X"45",X"2E",X"26",X"7C",X"18",X"3F",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"1E",X"F7",X"CD",X"45",
		X"2E",X"CD",X"65",X"2E",X"18",X"2F",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"24",X"CB",X"BD",X"36",
		X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"BB",X"2E",X"38",X"04",X"26",X"7C",X"18",X"18",X"26",X"7A",
		X"CB",X"FD",X"36",X"0E",X"11",X"CD",X"2B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",
		X"CD",X"65",X"2E",X"18",X"00",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"D4",
		X"30",X"C3",X"79",X"30",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"2A",X"CB",X"BD",X"36",X"4C",X"F7",
		X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"04",X"26",X"7C",X"18",X"DA",X"26",X"7A",X"CB",X"FD",
		X"36",X"0E",X"11",X"0B",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",
		X"35",X"28",X"05",X"CD",X"65",X"2E",X"18",X"BD",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"27",
		X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7C",X"18",X"A7",X"0E",X"0E",
		X"CD",X"8C",X"2E",X"36",X"30",X"F7",X"CD",X"45",X"2E",X"CD",X"BB",X"2E",X"38",X"06",X"2D",X"CD",
		X"65",X"2E",X"18",X"91",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"53",X"2C",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"04",X"25",X"C3",X"D5",X"2B",X"26",
		X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"6E",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",
		X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"33",X"CB",X"BD",
		X"36",X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"05",X"26",X"7C",X"C3",X"D6",X"2B",
		X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"9F",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",
		X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",
		X"FD",X"36",X"08",X"11",X"BC",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",
		X"7C",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"36",X"F7",X"CD",X"45",X"2E",X"CD",
		X"BB",X"2E",X"38",X"07",X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",
		X"16",X"11",X"EA",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",
		X"28",X"06",X"CD",X"81",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"07",
		X"2D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",
		X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"39",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"07",
		X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"36",X"2D",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",
		X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"53",X"2D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"CD",X"45",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",
		X"2E",X"36",X"3F",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"05",
		X"26",X"7C",X"C3",X"D6",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"16",X"11",X"84",X"2D",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"81",X"2E",X"C3",
		X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"68",X"2D",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"18",X"C5",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"15",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",
		X"55",X"2E",X"26",X"7C",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"1E",X"F7",X"CD",
		X"55",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"24",X"CB",
		X"BD",X"36",X"4C",X"F7",X"CD",X"55",X"2E",X"CD",X"BB",X"2E",X"38",X"05",X"26",X"7C",X"C3",X"D6",
		X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"F0",X"2D",X"DD",X"73",X"00",X"DD",X"72",X"01",
		X"CD",X"55",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"39",
		X"F7",X"CD",X"55",X"2E",X"CD",X"A0",X"2E",X"38",X"07",X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",
		X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"1F",X"2E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",
		X"55",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",
		X"FD",X"36",X"0E",X"11",X"3C",X"2E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"55",X"2E",X"CD",
		X"65",X"2E",X"C3",X"D5",X"2B",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"01",X"C9",
		X"33",X"33",X"C3",X"86",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"01",X"C9",
		X"33",X"33",X"C3",X"16",X"32",X"26",X"7C",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"C6",X"4C",X"77",
		X"C9",X"26",X"7C",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"ED",X"44",X"E6",X"03",X"C6",X"4C",X"77",
		X"C9",X"26",X"7C",X"3A",X"01",X"80",X"E6",X"03",X"C6",X"4C",X"77",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"2D",X"24",X"CB",X"FD",X"71",X"24",X"36",X"00",X"24",X"C9",
		X"24",X"2C",X"3A",X"41",X"7A",X"96",X"D6",X"02",X"C6",X"04",X"D0",X"24",X"3A",X"41",X"7B",X"96",
		X"D6",X"02",X"C6",X"04",X"D0",X"2D",X"26",X"7D",X"36",X"30",X"C9",X"24",X"2C",X"3A",X"45",X"7A",
		X"96",X"D6",X"02",X"C6",X"04",X"D0",X"24",X"3A",X"45",X"7B",X"96",X"D6",X"02",X"C6",X"04",X"D0",
		X"2D",X"26",X"7D",X"36",X"30",X"C9",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"16",X"79",X"DD",
		X"5D",X"EB",X"2C",X"36",X"00",X"2D",X"26",X"7C",X"36",X"3C",X"CB",X"FD",X"36",X"2A",X"24",X"36",
		X"01",X"CB",X"BD",X"24",X"3A",X"A6",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",
		X"7F",X"36",X"00",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",
		X"7D",X"CB",X"FD",X"35",X"20",X"3E",X"26",X"79",X"5E",X"2C",X"56",X"2D",X"1A",X"26",X"7D",X"77",
		X"13",X"1A",X"13",X"26",X"79",X"73",X"2C",X"72",X"2D",X"26",X"7B",X"EB",X"21",X"B1",X"2F",X"CD",
		X"83",X"33",X"EB",X"26",X"7D",X"CB",X"BD",X"2C",X"35",X"28",X"03",X"2D",X"18",X"18",X"11",X"47",
		X"2F",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"86",X"31",X"18",X"02",X"CB",X"BD",X"26",X"7F",X"7E",X"A7",X"20",X"1A",X"26",X"7A",X"2C",X"3A",
		X"B1",X"81",X"BE",X"38",X"34",X"3A",X"01",X"80",X"E6",X"07",X"20",X"2D",X"2D",X"26",X"7D",X"35",
		X"20",X"27",X"26",X"7F",X"36",X"18",X"35",X"7E",X"FE",X"0C",X"20",X"10",X"E5",X"CD",X"87",X"32",
		X"E1",X"25",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",X"7F",X"7E",X"0F",X"0F",X"E6",X"07",
		X"EB",X"21",X"AB",X"2F",X"D7",X"7E",X"16",X"7C",X"12",X"16",X"7C",X"DD",X"5D",X"1C",X"3A",X"1C",
		X"80",X"12",X"16",X"7A",X"1D",X"CD",X"91",X"30",X"C3",X"79",X"30",X"3C",X"3D",X"3E",X"3F",X"3E",
		X"3D",X"00",X"10",X"02",X"10",X"04",X"10",X"06",X"10",X"08",X"10",X"08",X"0E",X"08",X"0C",X"08",
		X"0A",X"08",X"08",X"08",X"06",X"08",X"04",X"08",X"02",X"08",X"00",X"06",X"00",X"04",X"00",X"02",
		X"00",X"00",X"00",X"FE",X"00",X"FC",X"00",X"FA",X"00",X"F8",X"00",X"F8",X"02",X"F8",X"04",X"F8",
		X"06",X"F8",X"08",X"F8",X"0A",X"F8",X"0C",X"F8",X"0E",X"F8",X"10",X"FA",X"10",X"FC",X"10",X"FE",
		X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",
		X"21",X"00",X"79",X"11",X"01",X"79",X"01",X"FF",X"06",X"36",X"00",X"ED",X"B0",X"21",X"79",X"30",
		X"22",X"00",X"78",X"22",X"4E",X"78",X"21",X"00",X"78",X"11",X"02",X"78",X"01",X"3E",X"00",X"ED",
		X"B0",X"21",X"4E",X"78",X"11",X"50",X"78",X"01",X"32",X"00",X"ED",X"B0",X"21",X"4E",X"7C",X"11",
		X"50",X"7C",X"01",X"24",X"00",X"36",X"1E",X"ED",X"B0",X"21",X"4F",X"79",X"11",X"50",X"79",X"01",
		X"24",X"00",X"36",X"80",X"2D",X"36",X"00",X"ED",X"B0",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"F7",
		X"3A",X"2A",X"80",X"A7",X"20",X"AA",X"DD",X"E5",X"DD",X"21",X"00",X"78",X"06",X"20",X"CD",X"54",
		X"04",X"DD",X"2C",X"DD",X"2C",X"10",X"F7",X"DD",X"21",X"4E",X"78",X"06",X"19",X"CD",X"54",X"04",
		X"DD",X"2C",X"DD",X"2C",X"10",X"F7",X"DD",X"E1",X"C9",X"F7",X"16",X"7F",X"DD",X"5D",X"EB",X"7E",
		X"A7",X"C8",X"3D",X"21",X"83",X"3C",X"CF",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",
		X"C9",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"7C",
		X"1C",X"12",X"14",X"1A",X"67",X"1D",X"1A",X"6F",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",
		X"1C",X"7C",X"12",X"15",X"1A",X"14",X"C6",X"01",X"FE",X"29",X"30",X"06",X"1A",X"FE",X"1F",X"DA",
		X"1D",X"00",X"1D",X"15",X"15",X"EB",X"AF",X"77",X"CB",X"FD",X"77",X"CB",X"BD",X"3E",X"06",X"84",
		X"67",X"36",X"00",X"C9",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"CB",X"FB",X"1A",X"CF",X"CB",X"BB",
		X"7D",X"12",X"1C",X"7C",X"12",X"C3",X"B4",X"30",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"3A",X"14",
		X"80",X"ED",X"44",X"CF",X"7D",X"12",X"1C",X"7C",X"12",X"C3",X"B4",X"30",X"1A",X"6F",X"1C",X"1A",
		X"67",X"1D",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"7C",X"1C",X"12",X"14",X"1A",X"67",
		X"1D",X"1A",X"6F",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"1C",X"7C",X"12",X"C9",X"24",
		X"24",X"24",X"2C",X"36",X"07",X"2D",X"24",X"36",X"FF",X"11",X"32",X"31",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"3E",X"05",X"DD",X"84",X"57",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",X"08",X"20",X"0A",
		X"25",X"25",X"25",X"2C",X"35",X"24",X"34",X"2D",X"24",X"24",X"4F",X"CB",X"3F",X"CB",X"3F",X"FE",
		X"05",X"28",X"26",X"EB",X"21",X"6F",X"31",X"CF",X"15",X"7E",X"12",X"15",X"15",X"15",X"1C",X"23",
		X"79",X"E6",X"03",X"07",X"07",X"86",X"12",X"1D",X"14",X"CD",X"91",X"30",X"C3",X"79",X"30",X"70",
		X"00",X"71",X"00",X"74",X"03",X"78",X"03",X"7C",X"03",X"24",X"24",X"36",X"00",X"3E",X"FA",X"84",
		X"67",X"36",X"00",X"C3",X"79",X"30",X"26",X"7C",X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"11",
		X"98",X"31",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"E6",X"07",X"20",X"2A",X"79",X"0F",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"29",X"FE",X"02",
		X"CC",X"02",X"32",X"FE",X"05",X"CC",X"0C",X"32",X"EB",X"21",X"F4",X"31",X"CF",X"15",X"7E",X"12",
		X"23",X"16",X"79",X"1C",X"7E",X"12",X"1D",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7A",
		X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"25",X"36",X"A6",X"2C",X"36",X"0D",X"F7",X"16",X"7C",
		X"DD",X"5D",X"3A",X"01",X"80",X"0F",X"0F",X"E6",X"01",X"C6",X"A6",X"12",X"16",X"7A",X"CD",X"E8",
		X"30",X"C3",X"79",X"30",X"60",X"00",X"61",X"00",X"64",X"03",X"68",X"03",X"6C",X"03",X"62",X"00",
		X"63",X"00",X"4C",X"26",X"7A",X"2C",X"35",X"24",X"34",X"2D",X"61",X"C9",X"4C",X"26",X"7A",X"2C",
		X"34",X"24",X"35",X"2D",X"61",X"C9",X"26",X"7C",X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"11",
		X"28",X"32",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"E6",X"03",X"20",X"29",X"79",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"29",X"FE",X"02",X"CC",
		X"02",X"32",X"FE",X"05",X"CC",X"0C",X"32",X"EB",X"21",X"F4",X"31",X"CF",X"15",X"7E",X"12",X"23",
		X"16",X"79",X"1C",X"7E",X"12",X"1D",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7A",X"EB",
		X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7F",X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",
		X"30",X"3A",X"01",X"80",X"E6",X"07",X"C0",X"35",X"C0",X"E5",X"CD",X"87",X"32",X"E1",X"24",X"CD",
		X"4B",X"0F",X"A6",X"25",X"3C",X"77",X"C9",X"48",X"21",X"4E",X"79",X"06",X"13",X"7E",X"3D",X"28",
		X"2A",X"2C",X"2C",X"10",X"F8",X"41",X"C9",X"21",X"4E",X"79",X"06",X"13",X"7E",X"3D",X"28",X"24",
		X"2C",X"2C",X"10",X"F8",X"C9",X"36",X"02",X"16",X"7A",X"DD",X"5D",X"24",X"1A",X"77",X"1C",X"2C",
		X"1A",X"77",X"14",X"24",X"1A",X"77",X"1D",X"2D",X"1A",X"77",X"C9",X"CD",X"A5",X"32",X"CB",X"D4",
		X"36",X"06",X"41",X"C9",X"CD",X"A5",X"32",X"EB",X"CB",X"FB",X"21",X"B3",X"3D",X"79",X"CD",X"83",
		X"33",X"EB",X"CB",X"BD",X"26",X"7F",X"36",X"07",X"C9",X"16",X"7A",X"DD",X"5D",X"1C",X"1A",X"4F",
		X"3A",X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",
		X"D6",X"20",X"0F",X"0F",X"0F",X"E6",X"1F",X"4F",X"C5",X"06",X"05",X"C5",X"CD",X"97",X"32",X"C1",
		X"79",X"C6",X"02",X"E6",X"1F",X"4F",X"10",X"F3",X"C1",X"C9",X"C5",X"01",X"00",X"10",X"C5",X"CD",
		X"97",X"32",X"C1",X"79",X"3C",X"3C",X"E6",X"1E",X"4F",X"10",X"F3",X"21",X"76",X"7A",X"11",X"78",
		X"7A",X"01",X"08",X"00",X"ED",X"B0",X"21",X"76",X"7B",X"11",X"78",X"7B",X"01",X"08",X"00",X"ED",
		X"B0",X"21",X"5D",X"33",X"11",X"F8",X"7A",X"06",X"04",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",
		X"21",X"61",X"33",X"11",X"F8",X"7B",X"06",X"04",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",X"3E",
		X"09",X"06",X"04",X"21",X"78",X"7F",X"77",X"2C",X"2C",X"10",X"FB",X"C1",X"C9",X"20",X"00",X"E0",
		X"00",X"00",X"E0",X"00",X"20",X"E5",X"1A",X"4F",X"3A",X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",
		X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",X"C6",X"04",X"E1",X"CB",X"FB",X"1D",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"CF",X"7E",X"12",X"23",X"15",X"7E",X"12",X"C9",X"CD",X"4B",X"0F",X"E6",X"1F",
		X"FE",X"19",X"30",X"F7",X"C6",X"03",X"77",X"C9",X"E5",X"21",X"47",X"7B",X"CD",X"4B",X"0F",X"E6",
		X"1F",X"FE",X"19",X"30",X"F7",X"C6",X"03",X"5F",X"96",X"D6",X"08",X"C6",X"10",X"7B",X"38",X"EC",
		X"E1",X"77",X"C9",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"2B",X"80",X"A7",X"C8",X"47",X"3A",X"2C",
		X"80",X"21",X"03",X"3C",X"D7",X"11",X"74",X"7F",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",X"C9",
		X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"2D",X"80",X"A7",X"C8",X"21",X"20",X"7F",X"47",X"36",X"01",
		X"2C",X"2C",X"10",X"FA",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"22",X"84",X"A7",X"C8",
		X"3E",X"3C",X"32",X"23",X"84",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"E9",X"21",X"23",X"84",X"35",
		X"C0",X"21",X"2D",X"80",X"34",X"21",X"22",X"84",X"35",X"28",X"DA",X"18",X"E3",X"16",X"79",X"DD",
		X"5D",X"EB",X"36",X"02",X"2C",X"36",X"80",X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"73",
		X"3D",X"CD",X"65",X"33",X"EB",X"26",X"7C",X"36",X"00",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",
		X"FE",X"03",X"28",X"1D",X"3A",X"01",X"80",X"0F",X"4F",X"E6",X"03",X"26",X"7C",X"77",X"79",X"0F",
		X"0F",X"E6",X"03",X"C6",X"26",X"2C",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"26",X"7D",X"36",X"FF",X"11",X"5D",X"34",X"26",X"78",X"73",X"2C",X"72",X"16",X"7D",X"DD",
		X"5D",X"EB",X"34",X"7E",X"0F",X"FE",X"04",X"28",X"0D",X"C6",X"04",X"25",X"77",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"26",X"79",X"36",X"00",X"26",X"7F",X"36",X"00",X"C3",X"79",
		X"30",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"34",X"2A",X"1E",X"7A",X"3E",X"10",X"BC",X"28",X"0E",
		X"3E",X"01",X"32",X"07",X"A0",X"3E",X"10",X"CF",X"22",X"1E",X"7A",X"C3",X"47",X"38",X"11",X"A7",
		X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"2F",X"80",X"A7",X"20",X"48",X"3A",X"1C",X"79",
		X"FE",X"03",X"28",X"08",X"3E",X"01",X"32",X"07",X"A0",X"C3",X"47",X"38",X"3E",X"1D",X"32",X"40",
		X"80",X"3E",X"03",X"32",X"1E",X"7D",X"11",X"CF",X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"21",
		X"1E",X"7D",X"35",X"20",X"0E",X"3E",X"06",X"32",X"40",X"80",X"11",X"E3",X"34",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"30",X"BC",X"28",X"30",X"3A",X"14",X"80",X"ED",X"44",
		X"CF",X"22",X"1E",X"7A",X"C9",X"11",X"F5",X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"1C",
		X"79",X"FE",X"03",X"28",X"B7",X"2A",X"1E",X"7A",X"3E",X"F8",X"BC",X"28",X"0E",X"3E",X"F8",X"CF",
		X"22",X"1E",X"7A",X"3E",X"01",X"32",X"07",X"A0",X"C3",X"47",X"38",X"AF",X"32",X"1E",X"79",X"32",
		X"1E",X"7F",X"C3",X"79",X"30",X"3E",X"02",X"32",X"1C",X"79",X"3E",X"10",X"32",X"1C",X"7C",X"3E",
		X"3C",X"32",X"9C",X"7C",X"2A",X"1E",X"7B",X"22",X"1C",X"7B",X"F7",X"3A",X"1C",X"79",X"FE",X"03",
		X"28",X"29",X"3A",X"1E",X"79",X"3D",X"28",X"1A",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"E6",X"0C",
		X"C6",X"80",X"32",X"1D",X"79",X"2A",X"1E",X"7A",X"22",X"1C",X"7A",X"3A",X"40",X"80",X"32",X"1D",
		X"7C",X"C9",X"32",X"1C",X"79",X"32",X"1C",X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",
		X"37",X"11",X"7A",X"35",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"22",X"1C",X"7A",
		X"2A",X"1E",X"7B",X"22",X"1C",X"7B",X"CD",X"F8",X"37",X"3A",X"1C",X"79",X"FE",X"04",X"C0",X"11",
		X"A5",X"35",X"DD",X"73",X"00",X"DD",X"72",X"01",X"21",X"9C",X"7A",X"36",X"D0",X"24",X"36",X"00",
		X"3E",X"08",X"32",X"1D",X"79",X"3A",X"01",X"80",X"0F",X"4F",X"E6",X"03",X"C6",X"B8",X"32",X"1C",
		X"7C",X"79",X"E6",X"07",X"C6",X"15",X"32",X"1D",X"7C",X"11",X"1C",X"7A",X"CD",X"D4",X"30",X"C3",
		X"79",X"30",X"3E",X"02",X"32",X"1A",X"79",X"AF",X"32",X"1B",X"79",X"3C",X"32",X"1A",X"7D",X"3E",
		X"5C",X"32",X"1A",X"7C",X"3E",X"30",X"32",X"9A",X"7C",X"2A",X"1E",X"7B",X"3E",X"02",X"84",X"67",
		X"22",X"1A",X"7B",X"3A",X"A7",X"81",X"32",X"1A",X"7E",X"F7",X"3A",X"1A",X"79",X"FE",X"03",X"28",
		X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",X"1E",
		X"7A",X"3E",X"FE",X"84",X"67",X"22",X"1A",X"7A",X"3A",X"40",X"80",X"32",X"1B",X"7C",X"21",X"1A",
		X"7D",X"CD",X"71",X"32",X"C9",X"32",X"1A",X"79",X"32",X"1A",X"7F",X"C3",X"79",X"30",X"DD",X"5D",
		X"6B",X"CD",X"EE",X"37",X"11",X"2D",X"36",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",
		X"3E",X"FE",X"84",X"67",X"22",X"1A",X"7A",X"2A",X"1E",X"7B",X"3E",X"02",X"84",X"67",X"22",X"1A",
		X"7B",X"CD",X"F8",X"37",X"3A",X"1A",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"3E",X"02",X"32",
		X"18",X"79",X"AF",X"32",X"19",X"79",X"3C",X"32",X"18",X"7D",X"3E",X"5D",X"32",X"18",X"7C",X"3E",
		X"30",X"32",X"98",X"7C",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",X"18",X"7B",X"3A",X"A7",
		X"81",X"32",X"18",X"7E",X"F7",X"3A",X"18",X"79",X"FE",X"03",X"28",X"2D",X"3A",X"1C",X"79",X"FE",
		X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",X"1E",X"7A",X"3E",X"FE",X"84",X"67",
		X"22",X"18",X"7A",X"3A",X"40",X"80",X"32",X"19",X"7C",X"21",X"18",X"7D",X"CD",X"71",X"32",X"C9",
		X"32",X"18",X"79",X"32",X"18",X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",X"37",X"11",
		X"B8",X"36",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"FE",X"84",X"67",X"22",
		X"18",X"7A",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",X"18",X"7B",X"CD",X"F8",X"37",X"3A",
		X"18",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"3E",X"02",X"32",X"16",X"79",X"AF",X"32",X"17",
		X"79",X"3C",X"32",X"16",X"7D",X"3E",X"5E",X"32",X"16",X"7C",X"3E",X"30",X"32",X"96",X"7C",X"2A",
		X"1E",X"7B",X"3E",X"02",X"84",X"67",X"22",X"16",X"7B",X"3A",X"A7",X"81",X"32",X"16",X"7E",X"F7",
		X"3A",X"16",X"79",X"FE",X"03",X"28",X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",
		X"79",X"3D",X"28",X"17",X"2A",X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"16",X"7A",X"3A",X"40",
		X"80",X"32",X"17",X"7C",X"21",X"16",X"7D",X"CD",X"71",X"32",X"C9",X"32",X"16",X"79",X"32",X"16",
		X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",X"37",X"11",X"43",X"37",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"16",X"7A",X"2A",X"1E",X"7B",
		X"3E",X"02",X"84",X"67",X"22",X"16",X"7B",X"CD",X"F8",X"37",X"3A",X"16",X"79",X"FE",X"04",X"C0",
		X"AF",X"18",X"C8",X"3E",X"02",X"32",X"14",X"79",X"AF",X"32",X"15",X"79",X"3C",X"32",X"14",X"7D",
		X"3E",X"5F",X"32",X"14",X"7C",X"3E",X"30",X"32",X"94",X"7C",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",
		X"67",X"22",X"14",X"7B",X"3A",X"A7",X"81",X"32",X"14",X"7E",X"F7",X"3A",X"14",X"79",X"FE",X"03",
		X"28",X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",
		X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"14",X"7A",X"3A",X"40",X"80",X"32",X"15",X"7C",X"21",
		X"14",X"7D",X"CD",X"71",X"32",X"C9",X"32",X"14",X"79",X"32",X"14",X"7F",X"C3",X"79",X"30",X"DD",
		X"5D",X"6B",X"CD",X"EE",X"37",X"11",X"CE",X"37",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",
		X"7A",X"3E",X"02",X"84",X"67",X"22",X"14",X"7A",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",
		X"14",X"7B",X"CD",X"F8",X"37",X"3A",X"14",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"26",X"7C",
		X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"C9",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"0F",X"0F",X"E6",X"07",X"D6",X"05",X"C6",X"03",X"DC",X"3D",X"38",X"79",X"E6",X"03",X"C0",X"79",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"0F",X"EB",X"21",X"2F",X"38",X"CF",X"15",X"7E",X"12",
		X"23",X"1C",X"16",X"79",X"7E",X"12",X"C9",X"25",X"36",X"00",X"26",X"79",X"36",X"04",X"C9",X"60",
		X"00",X"61",X"00",X"64",X"03",X"68",X"03",X"6C",X"03",X"62",X"00",X"63",X"00",X"26",X"7A",X"2C",
		X"35",X"24",X"34",X"2D",X"26",X"7D",X"C9",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"E6",X"07",X"21",
		X"58",X"38",X"D7",X"7E",X"32",X"40",X"80",X"C9",X"02",X"03",X"04",X"05",X"06",X"05",X"04",X"03",
		X"3E",X"03",X"32",X"12",X"79",X"32",X"13",X"79",X"3E",X"58",X"32",X"12",X"7C",X"2A",X"1E",X"7B",
		X"3E",X"05",X"84",X"67",X"22",X"12",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"FB",X"84",X"67",X"22",
		X"12",X"7A",X"3A",X"40",X"80",X"32",X"13",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",
		X"12",X"79",X"32",X"12",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"10",X"79",X"32",X"11",X"79",
		X"3E",X"80",X"32",X"10",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"10",X"7B",X"F7",X"2A",X"1E",X"7A",
		X"3E",X"FB",X"84",X"67",X"22",X"10",X"7A",X"3A",X"40",X"80",X"32",X"11",X"7C",X"3A",X"1E",X"79",
		X"FE",X"01",X"C0",X"AF",X"32",X"10",X"79",X"32",X"10",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",
		X"0E",X"79",X"32",X"0F",X"79",X"3E",X"84",X"32",X"0E",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",X"84",
		X"67",X"22",X"0E",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"FB",X"84",X"67",X"22",X"0E",X"7A",X"3A",
		X"40",X"80",X"32",X"0F",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"0E",X"79",X"32",
		X"0E",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"0C",X"79",X"32",X"0D",X"79",X"3E",X"88",X"32",
		X"0C",X"7C",X"2A",X"1E",X"7B",X"3E",X"05",X"84",X"67",X"22",X"0C",X"7B",X"F7",X"2A",X"1E",X"7A",
		X"25",X"22",X"0C",X"7A",X"3A",X"40",X"80",X"32",X"0D",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",
		X"AF",X"32",X"0C",X"79",X"32",X"0C",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"0A",X"79",X"32",
		X"0B",X"79",X"3E",X"8C",X"32",X"0A",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"0A",X"7B",X"F7",X"2A",
		X"1E",X"7A",X"25",X"22",X"0A",X"7A",X"3A",X"40",X"80",X"32",X"0B",X"7C",X"3A",X"1E",X"79",X"FE",
		X"01",X"C0",X"AF",X"32",X"0A",X"79",X"32",X"0A",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"08",
		X"79",X"32",X"09",X"79",X"3E",X"90",X"32",X"08",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",X"84",X"67",
		X"22",X"08",X"7B",X"F7",X"2A",X"1E",X"7A",X"25",X"22",X"08",X"7A",X"3A",X"40",X"80",X"32",X"09",
		X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"08",X"79",X"32",X"08",X"7F",X"C3",X"79",
		X"30",X"3E",X"03",X"32",X"06",X"79",X"32",X"07",X"79",X"3E",X"94",X"32",X"06",X"7C",X"2A",X"1E",
		X"7B",X"3E",X"05",X"84",X"67",X"22",X"06",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"03",X"84",X"67",
		X"22",X"06",X"7A",X"3A",X"40",X"80",X"32",X"07",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",
		X"32",X"06",X"79",X"32",X"06",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"04",X"79",X"32",X"05",
		X"79",X"3E",X"98",X"32",X"04",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"04",X"7B",X"F7",X"2A",X"1E",
		X"7A",X"3E",X"03",X"84",X"67",X"22",X"04",X"7A",X"3A",X"40",X"80",X"32",X"05",X"7C",X"3A",X"1E",
		X"79",X"FE",X"01",X"C0",X"AF",X"32",X"04",X"79",X"32",X"04",X"7F",X"C3",X"79",X"30",X"3E",X"03",
		X"32",X"02",X"79",X"32",X"03",X"79",X"3E",X"9C",X"32",X"02",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",
		X"84",X"67",X"22",X"02",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"03",X"84",X"67",X"22",X"02",X"7A",
		X"3A",X"40",X"80",X"32",X"03",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"02",X"79",
		X"32",X"02",X"7F",X"C3",X"79",X"30",X"3A",X"28",X"80",X"A7",X"20",X"59",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"2D",X"36",X"00",X"11",X"64",X"3A",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"1A",X"FE",X"03",X"28",X"08",X"16",X"7A",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"16",X"7D",X"3E",X"80",X"12",X"21",X"CD",X"3E",X"11",X"B6",X"3A",
		X"C5",X"06",X"13",X"1A",X"0F",X"BE",X"20",X"29",X"13",X"23",X"10",X"F7",X"CD",X"C9",X"3A",X"11",
		X"99",X"3A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"C1",X"16",X"7D",X"DD",X"5D",X"EB",X"35",X"C0",
		X"C5",X"CD",X"7C",X"3B",X"C1",X"16",X"79",X"DD",X"5D",X"AF",X"12",X"16",X"7F",X"12",X"C3",X"79",
		X"30",X"CD",X"09",X"3B",X"18",X"D9",X"5A",X"5C",X"50",X"48",X"02",X"12",X"10",X"04",X"48",X"2E",
		X"14",X"2C",X"18",X"30",X"48",X"2A",X"3A",X"1A",X"A0",X"21",X"E1",X"3A",X"CD",X"48",X"3B",X"21",
		X"21",X"19",X"06",X"07",X"0E",X"B0",X"3E",X"1A",X"CD",X"5D",X"14",X"21",X"F1",X"3A",X"C3",X"62",
		X"3B",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"DB",X"E7",X"E4",X"ED",X"EF",X"ED",X"E8",X"F5",
		X"EA",X"DB",X"DB",X"DB",X"DB",X"DB",X"BA",X"B8",X"BB",X"C3",X"B8",X"C9",X"BD",X"DB",X"C8",X"B1",
		X"DB",X"F1",X"E0",X"F1",X"DC",X"E7",X"E7",X"DB",X"DB",X"21",X"20",X"3B",X"CD",X"48",X"3B",X"21",
		X"21",X"19",X"06",X"09",X"0E",X"B0",X"3E",X"1B",X"CD",X"5D",X"14",X"21",X"30",X"3B",X"18",X"42",
		X"F2",X"F1",X"F5",X"F2",X"DB",X"F3",X"E7",X"E6",X"DD",X"DB",X"E9",X"F5",X"EB",X"ED",X"E8",X"EF",
		X"C7",X"BB",X"BA",X"B1",X"DB",X"B5",X"BC",X"C6",X"C5",X"B8",X"DB",X"E8",X"F5",X"E9",X"F3",X"E7",
		X"DB",X"BA",X"B8",X"BB",X"C3",X"B8",X"C9",X"BD",X"11",X"80",X"84",X"06",X"10",X"7E",X"2F",X"12",
		X"23",X"13",X"10",X"F9",X"21",X"21",X"19",X"11",X"80",X"84",X"06",X"10",X"0E",X"C0",X"CD",X"1F",
		X"14",X"C9",X"11",X"80",X"84",X"06",X"18",X"7E",X"2F",X"12",X"23",X"13",X"10",X"F9",X"21",X"22",
		X"17",X"11",X"80",X"84",X"06",X"18",X"0E",X"C0",X"CD",X"1F",X"14",X"C9",X"21",X"21",X"19",X"06",
		X"10",X"0E",X"C0",X"3E",X"24",X"CD",X"5D",X"14",X"21",X"21",X"19",X"06",X"10",X"0E",X"B0",X"3E",
		X"24",X"CD",X"5D",X"14",X"21",X"22",X"17",X"06",X"18",X"0E",X"C0",X"C3",X"5D",X"14",X"21",X"00",
		X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",X"21",X"01",X"3C",X"01",X"01",X"64",X"CD",X"10",
		X"01",X"F7",X"21",X"60",X"80",X"01",X"04",X"74",X"CD",X"E5",X"00",X"F7",X"3A",X"63",X"80",X"FE",
		X"05",X"C2",X"00",X"00",X"F7",X"21",X"02",X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",X"21",
		X"60",X"80",X"01",X"04",X"74",X"CD",X"E5",X"00",X"F7",X"3A",X"63",X"80",X"FE",X"95",X"C2",X"00",
		X"00",X"F7",X"C9",X"21",X"9E",X"3B",X"11",X"F6",X"3B",X"06",X"0A",X"1A",X"BE",X"C2",X"00",X"00",
		X"23",X"13",X"10",X"F7",X"F7",X"C9",X"21",X"00",X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",
		X"10",X"80",X"E5",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"56",X"56",X"56",X"56",X"56",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0B",X"0B",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0E",X"0E",X"12",X"12",X"12",X"13",X"13",X"13",X"14",
		X"14",X"14",X"14",X"14",X"14",X"0E",X"0E",X"0E",X"10",X"10",X"10",X"10",X"10",X"10",X"14",X"14",
		X"14",X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"0F",
		X"0F",X"08",X"08",X"08",X"08",X"55",X"55",X"10",X"10",X"08",X"08",X"08",X"08",X"11",X"11",X"14",
		X"14",X"15",X"15",X"15",X"15",X"08",X"08",X"08",X"08",X"0E",X"0E",X"78",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"23",X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"2B",X"79",
		X"2B",X"0D",X"34",X"F8",X"1E",X"00",X"20",X"18",X"20",X"36",X"22",X"C4",X"21",X"B1",X"21",X"E7",
		X"20",X"A8",X"23",X"87",X"24",X"67",X"25",X"D7",X"25",X"2E",X"26",X"84",X"26",X"DF",X"26",X"36",
		X"27",X"4C",X"28",X"45",X"1B",X"18",X"1C",X"00",X"1C",X"0C",X"1C",X"61",X"1E",X"60",X"1A",X"F0",
		X"1A",X"89",X"1A",X"61",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"1B",X"39",
		X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"2B",X"DE",X"1C",X"D6",X"2E",X"00",
		X"00",X"00",X"00",X"DD",X"28",X"2E",X"2A",X"00",X"00",X"00",X"00",X"96",X"2B",X"A6",X"2B",X"E4",
		X"2B",X"2E",X"2C",X"77",X"2C",X"C4",X"2C",X"10",X"2D",X"5C",X"2D",X"A3",X"2D",X"B7",X"2D",X"C8",
		X"2D",X"F9",X"2D",X"60",X"38",X"98",X"38",X"CD",X"38",X"05",X"39",X"3A",X"39",X"6C",X"39",X"A1",
		X"39",X"D9",X"39",X"0E",X"3A",X"25",X"35",X"81",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"35",X"4D",X"36",X"D8",X"36",X"63",X"37",X"46",X"3A",X"5C",X"1F",X"06",X"23",X"AC",X"22",X"00",
		X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"05",X"00",X"00",X"07",X"00",X"00",
		X"10",X"00",X"00",X"15",X"00",X"00",X"20",X"00",X"00",X"25",X"00",X"00",X"30",X"00",X"00",X"40",
		X"00",X"00",X"50",X"00",X"00",X"60",X"00",X"00",X"70",X"00",X"00",X"80",X"00",X"00",X"90",X"00",
		X"00",X"00",X"01",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"50",X"02",X"00",X"00",X"04",X"00",
		X"00",X"10",X"00",X"00",X"40",X"0C",X"3F",X"18",X"3B",X"24",X"35",X"2D",X"2D",X"35",X"24",X"3B",
		X"18",X"3F",X"0C",X"40",X"00",X"3F",X"F4",X"3B",X"E8",X"35",X"DC",X"2D",X"D3",X"24",X"CB",X"18",
		X"C5",X"0C",X"C1",X"00",X"C0",X"F4",X"C1",X"E8",X"C5",X"DC",X"CB",X"D3",X"D3",X"CB",X"DC",X"C5",
		X"E8",X"C1",X"F4",X"C0",X"00",X"C1",X"0C",X"C5",X"18",X"CB",X"24",X"D3",X"2D",X"DC",X"35",X"E8",
		X"3B",X"F4",X"3F",X"00",X"30",X"09",X"2F",X"12",X"2C",X"1B",X"28",X"22",X"22",X"28",X"1B",X"2C",
		X"12",X"2F",X"09",X"30",X"00",X"2F",X"F7",X"2C",X"EE",X"28",X"E5",X"22",X"DE",X"1B",X"D8",X"12",
		X"D4",X"09",X"D1",X"00",X"D0",X"F7",X"D1",X"EE",X"D4",X"E5",X"D8",X"DE",X"DE",X"D8",X"E5",X"D4",
		X"EE",X"D1",X"F7",X"D0",X"00",X"D1",X"09",X"D4",X"12",X"D8",X"1B",X"DE",X"22",X"E5",X"28",X"EE",
		X"2C",X"F7",X"2F",X"00",X"20",X"06",X"1F",X"0C",X"1E",X"11",X"1B",X"17",X"17",X"1B",X"11",X"1E",
		X"0C",X"1F",X"06",X"20",X"00",X"1F",X"FA",X"1E",X"F4",X"1B",X"EF",X"17",X"E9",X"11",X"E5",X"0C",
		X"E2",X"06",X"E1",X"00",X"E0",X"FA",X"E1",X"F4",X"E2",X"EF",X"E5",X"E9",X"E9",X"E5",X"EF",X"E2",
		X"F4",X"E1",X"FA",X"E0",X"00",X"E1",X"06",X"E2",X"0C",X"E5",X"11",X"E9",X"17",X"EF",X"1B",X"F4",
		X"1E",X"FA",X"1F",X"00",X"18",X"05",X"18",X"09",X"16",X"0D",X"14",X"11",X"11",X"14",X"0D",X"16",
		X"09",X"18",X"05",X"18",X"00",X"18",X"FB",X"16",X"F7",X"14",X"F3",X"11",X"EF",X"0D",X"EC",X"09",
		X"EA",X"05",X"E8",X"00",X"E8",X"FB",X"E8",X"F7",X"EA",X"F3",X"EC",X"EF",X"EF",X"EC",X"F3",X"EA",
		X"F7",X"E8",X"FB",X"E8",X"00",X"E8",X"05",X"EA",X"09",X"EC",X"0D",X"EF",X"11",X"F3",X"14",X"F7",
		X"16",X"FB",X"18",X"00",X"10",X"03",X"10",X"06",X"0F",X"09",X"0D",X"0B",X"0B",X"0D",X"09",X"0F",
		X"06",X"10",X"03",X"10",X"00",X"10",X"FD",X"0F",X"FA",X"0D",X"F7",X"0B",X"F5",X"09",X"F3",X"06",
		X"F1",X"03",X"F0",X"00",X"F0",X"FD",X"F0",X"FA",X"F1",X"F7",X"F3",X"F5",X"F5",X"F3",X"F7",X"F1",
		X"FA",X"F0",X"FD",X"F0",X"00",X"F0",X"03",X"F1",X"06",X"F3",X"09",X"F5",X"0B",X"F7",X"0D",X"FA",
		X"0F",X"FD",X"10",X"24",X"00",X"54",X"0E",X"40",X"1A",X"64",X"04",X"2A",X"5C",X"0E",X"04",X"38",
		X"54",X"1A",X"00",X"11",X"12",X"10",X"11",X"24",X"1C",X"0C",X"18",X"1B",X"0E",X"2D",X"2E",X"28",
		X"24",X"01",X"09",X"08",X"02",X"24",X"17",X"0A",X"16",X"0C",X"18",X"24",X"15",X"1D",X"0D",X"50",
		X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"35",
		X"C3",X"65",X"01",X"12",X"42",X"21",X"00",X"00",X"87",X"D2",X"58",X"00",X"25",X"C3",X"58",X"00",
		X"A7",X"F2",X"58",X"00",X"25",X"C3",X"58",X"00",X"A7",X"F0",X"ED",X"44",X"C9",X"33",X"33",X"C9",
		X"EB",X"CD",X"05",X"00",X"29",X"19",X"C9",X"FF",X"EB",X"CD",X"05",X"00",X"29",X"29",X"19",X"C9",
		X"E1",X"DD",X"75",X"00",X"DD",X"74",X"01",X"C9",X"3A",X"03",X"80",X"A7",X"3E",X"03",X"28",X"04",
		X"25",X"25",X"3E",X"19",X"85",X"E6",X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",X"67",X"E6",X"C0",
		X"B5",X"6F",X"7C",X"E6",X"07",X"81",X"67",X"C9",X"85",X"6F",X"D0",X"24",X"C9",X"0E",X"12",X"1B",
		X"1B",X"22",X"24",X"16",X"18",X"1E",X"ED",X"45",X"11",X"17",X"93",X"21",X"16",X"93",X"01",X"13",
		X"00",X"ED",X"B8",X"DD",X"21",X"60",X"01",X"1E",X"00",X"01",X"04",X"05",X"DD",X"7E",X"00",X"DD",
		X"23",X"6F",X"26",X"20",X"7E",X"7B",X"81",X"5F",X"7E",X"12",X"10",X"F0",X"06",X"05",X"21",X"04",
		X"93",X"7E",X"2C",X"B6",X"2C",X"2F",X"A6",X"2C",X"A6",X"2C",X"E6",X"0F",X"20",X"04",X"10",X"F1",
		X"18",X"40",X"05",X"28",X"4F",X"05",X"CB",X"20",X"CB",X"20",X"0F",X"38",X"03",X"04",X"18",X"FA",
		X"3A",X"00",X"93",X"CB",X"3F",X"5F",X"CB",X"11",X"C6",X"01",X"6F",X"26",X"93",X"7E",X"CB",X"41",
		X"28",X"04",X"07",X"07",X"07",X"07",X"E6",X"F0",X"B0",X"CB",X"41",X"28",X"04",X"07",X"07",X"07",
		X"07",X"77",X"3A",X"00",X"93",X"A7",X"20",X"02",X"3E",X"02",X"3D",X"32",X"00",X"93",X"7B",X"A7",
		X"28",X"09",X"2A",X"02",X"93",X"7E",X"32",X"01",X"93",X"18",X"42",X"2A",X"02",X"93",X"3A",X"01",
		X"93",X"77",X"18",X"39",X"4F",X"21",X"00",X"93",X"CB",X"41",X"20",X"2D",X"7E",X"CB",X"3F",X"28",
		X"13",X"CB",X"59",X"20",X"0C",X"7E",X"FE",X"05",X"30",X"03",X"34",X"18",X"D5",X"36",X"05",X"18",
		X"D1",X"35",X"18",X"CE",X"2A",X"02",X"93",X"CB",X"59",X"20",X"03",X"2B",X"18",X"01",X"23",X"22",
		X"02",X"93",X"3E",X"01",X"32",X"00",X"93",X"18",X"B9",X"36",X"05",X"18",X"B5",X"21",X"E2",X"C0",
		X"11",X"01",X"93",X"06",X"03",X"1A",X"1C",X"CD",X"51",X"01",X"10",X"F9",X"21",X"E2",X"B0",X"3A",
		X"00",X"93",X"06",X"06",X"A7",X"0E",X"04",X"28",X"02",X"0E",X"0C",X"71",X"2D",X"3D",X"10",X"F4",
		X"C9",X"4F",X"E6",X"0F",X"77",X"2D",X"79",X"07",X"07",X"07",X"07",X"E6",X"0F",X"77",X"2D",X"C9",
		X"FD",X"FB",X"F7",X"EF",X"FE",X"3A",X"09",X"04",X"32",X"72",X"85",X"3A",X"FB",X"15",X"32",X"73",
		X"85",X"31",X"80",X"97",X"21",X"00",X"10",X"11",X"00",X"A4",X"01",X"20",X"00",X"ED",X"B0",X"21",
		X"B6",X"01",X"11",X"C0",X"82",X"01",X"40",X"00",X"ED",X"B0",X"21",X"02",X"80",X"7E",X"3D",X"20",
		X"FC",X"77",X"32",X"0A",X"80",X"3A",X"16",X"80",X"CB",X"7F",X"28",X"EE",X"DD",X"21",X"C0",X"82",
		X"06",X"20",X"C5",X"CD",X"AF",X"01",X"C1",X"DD",X"23",X"DD",X"23",X"10",X"F5",X"18",X"DB",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"E9",X"F6",X"01",X"18",X"02",X"8F",X"06",X"8B",X"07",X"27",X"02",
		X"64",X"02",X"CD",X"07",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"A6",X"02",X"1E",X"03",X"21",X"40",X"82",X"11",X"C0",X"87",X"01",X"40",X"00",X"ED",
		X"B0",X"21",X"40",X"83",X"11",X"C0",X"97",X"01",X"40",X"00",X"ED",X"B0",X"21",X"40",X"81",X"11",
		X"C0",X"A7",X"01",X"40",X"00",X"ED",X"B0",X"C9",X"2A",X"0C",X"80",X"7D",X"6C",X"26",X"D0",X"77",
		X"3A",X"0E",X"80",X"32",X"20",X"D0",X"C9",X"3A",X"18",X"80",X"4F",X"3A",X"29",X"80",X"47",X"91",
		X"C8",X"30",X"1B",X"79",X"32",X"29",X"80",X"FE",X"A0",X"C8",X"90",X"27",X"21",X"00",X"A0",X"86",
		X"27",X"77",X"21",X"5D",X"02",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C9",X"27",X"3D",
		X"32",X"22",X"80",X"79",X"32",X"29",X"80",X"3E",X"01",X"32",X"1B",X"80",X"C9",X"30",X"10",X"00",
		X"80",X"FF",X"10",X"10",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"01",X"80",X"1F",X"E6",X"03",X"C6",
		X"25",X"21",X"4F",X"7C",X"06",X"13",X"77",X"2C",X"2C",X"10",X"FB",X"3A",X"01",X"80",X"0F",X"0F",
		X"0F",X"E6",X"07",X"4F",X"21",X"96",X"02",X"D7",X"7E",X"32",X"1C",X"80",X"79",X"21",X"9E",X"02",
		X"D7",X"7E",X"32",X"43",X"80",X"C9",X"07",X"08",X"09",X"0A",X"0B",X"0A",X"09",X"08",X"10",X"11",
		X"12",X"13",X"14",X"13",X"12",X"11",X"3A",X"2A",X"80",X"A7",X"C0",X"CD",X"D4",X"02",X"3A",X"03",
		X"80",X"A7",X"3E",X"40",X"28",X"02",X"3E",X"30",X"2A",X"10",X"80",X"CF",X"29",X"29",X"AF",X"29",
		X"17",X"6C",X"67",X"22",X"0C",X"80",X"3A",X"03",X"80",X"A7",X"3E",X"00",X"28",X"02",X"3E",X"00",
		X"32",X"0E",X"80",X"C9",X"2A",X"10",X"80",X"4C",X"3A",X"14",X"80",X"CF",X"22",X"10",X"80",X"3A",
		X"0F",X"80",X"A7",X"C0",X"7C",X"B9",X"C8",X"FA",X"EC",X"02",X"C6",X"40",X"C6",X"F2",X"6F",X"3A",
		X"03",X"80",X"A7",X"3A",X"13",X"80",X"28",X"02",X"C6",X"FE",X"C6",X"FF",X"67",X"01",X"B8",X"20",
		X"16",X"FE",X"5D",X"22",X"00",X"F0",X"EB",X"E5",X"CD",X"38",X"00",X"3A",X"00",X"F0",X"77",X"3E",
		X"10",X"84",X"67",X"3A",X"01",X"F0",X"77",X"E1",X"EB",X"14",X"24",X"10",X"E5",X"C9",X"21",X"00",
		X"79",X"11",X"00",X"83",X"06",X"40",X"E5",X"CD",X"32",X"03",X"E1",X"2C",X"2C",X"1C",X"1C",X"10",
		X"F5",X"C9",X"7E",X"3D",X"C8",X"E5",X"3C",X"20",X"0C",X"4C",X"24",X"77",X"2C",X"77",X"24",X"77",
		X"2D",X"77",X"3C",X"61",X"77",X"2C",X"4E",X"79",X"12",X"D5",X"24",X"56",X"2D",X"5E",X"EB",X"CD",
		X"B3",X"03",X"FE",X"02",X"38",X"03",X"21",X"00",X"00",X"CD",X"89",X"03",X"E5",X"EB",X"24",X"5E",
		X"2C",X"56",X"EB",X"CD",X"B3",X"03",X"A7",X"28",X"02",X"2E",X"00",X"CD",X"A2",X"03",X"D1",X"E1",
		X"2C",X"72",X"25",X"73",X"2D",X"77",X"25",X"EB",X"E1",X"4C",X"24",X"24",X"24",X"7E",X"12",X"2C",
		X"1C",X"7E",X"12",X"61",X"2D",X"14",X"14",X"1D",X"C9",X"3A",X"03",X"80",X"A7",X"28",X"0F",X"3E",
		X"48",X"CB",X"41",X"20",X"02",X"3E",X"58",X"95",X"6F",X"3E",X"01",X"9C",X"67",X"C9",X"3E",X"08",
		X"D7",X"C9",X"3A",X"03",X"80",X"A7",X"3E",X"EF",X"28",X"07",X"85",X"CB",X"49",X"C0",X"C6",X"10",
		X"C9",X"95",X"C9",X"AF",X"29",X"17",X"29",X"17",X"29",X"17",X"6C",X"67",X"C9",X"0A",X"03",X"21",
		X"D8",X"04",X"CF",X"7E",X"32",X"2B",X"80",X"23",X"7E",X"32",X"2C",X"80",X"ED",X"43",X"85",X"81",
		X"C9",X"3A",X"16",X"80",X"2F",X"07",X"07",X"07",X"E6",X"03",X"21",X"08",X"04",X"D7",X"7E",X"6F",
		X"3A",X"88",X"81",X"85",X"FE",X"80",X"38",X"02",X"D6",X"40",X"32",X"88",X"81",X"18",X"D0",X"21",
		X"88",X"81",X"0A",X"86",X"03",X"FE",X"80",X"38",X"02",X"D6",X"40",X"18",X"C2",X"21",X"00",X"00",
		X"22",X"2B",X"80",X"ED",X"43",X"85",X"81",X"C9",X"02",X"00",X"06",X"10",X"ED",X"43",X"85",X"81",
		X"2A",X"81",X"81",X"3A",X"8B",X"81",X"CD",X"2C",X"04",X"11",X"10",X"00",X"A7",X"ED",X"52",X"19",
		X"38",X"02",X"2E",X"10",X"3A",X"88",X"81",X"85",X"32",X"88",X"81",X"C9",X"C5",X"4F",X"AF",X"06",
		X"10",X"29",X"17",X"38",X"03",X"B9",X"38",X"02",X"91",X"23",X"10",X"F5",X"C1",X"C9",X"0A",X"32",
		X"A0",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A3",X"81",X"03",X"ED",X"43",X"85",
		X"81",X"C9",X"0A",X"32",X"A4",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A2",X"81",
		X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A1",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",
		X"0A",X"32",X"A5",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A6",X"81",X"03",X"ED",
		X"43",X"85",X"81",X"C9",X"0A",X"32",X"A7",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",
		X"B1",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"04",X"0B",X"05",X"0A",X"06",X"09",X"06",X"25",
		X"06",X"5C",X"06",X"29",X"06",X"5E",X"06",X"64",X"06",X"66",X"06",X"72",X"04",X"30",X"04",X"31",
		X"05",X"30",X"06",X"30",X"06",X"3F",X"06",X"48",X"06",X"4B",X"02",X"54",X"03",X"54",X"04",X"54",
		X"02",X"58",X"03",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",
		X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"03",X"01",X"03",X"01",X"03",X"01",X"04",X"01",
		X"04",X"01",X"04",X"01",X"05",X"01",X"05",X"01",X"05",X"01",X"02",X"19",X"02",X"19",X"02",X"19",
		X"04",X"01",X"04",X"01",X"04",X"04",X"04",X"04",X"04",X"05",X"04",X"05",X"05",X"05",X"05",X"05",
		X"06",X"05",X"06",X"05",X"03",X"19",X"03",X"19",X"04",X"19",X"04",X"19",X"05",X"19",X"05",X"19",
		X"03",X"27",X"03",X"27",X"04",X"27",X"04",X"27",X"05",X"27",X"05",X"27",X"03",X"1F",X"03",X"1F",
		X"04",X"1F",X"04",X"1F",X"05",X"1F",X"05",X"1F",X"03",X"13",X"03",X"13",X"04",X"13",X"04",X"13",
		X"05",X"13",X"05",X"13",X"03",X"36",X"03",X"36",X"03",X"37",X"03",X"37",X"04",X"37",X"04",X"37",
		X"03",X"2D",X"03",X"2D",X"04",X"2D",X"04",X"2D",X"05",X"2D",X"05",X"2D",X"04",X"12",X"04",X"12",
		X"04",X"11",X"04",X"11",X"05",X"11",X"05",X"11",X"05",X"17",X"05",X"17",X"06",X"17",X"06",X"17",
		X"02",X"3C",X"03",X"3C",X"03",X"3C",X"04",X"3C",X"04",X"3C",X"05",X"3C",X"05",X"19",X"05",X"19",
		X"06",X"19",X"06",X"19",X"02",X"45",X"03",X"45",X"03",X"45",X"04",X"45",X"04",X"45",X"05",X"45",
		X"05",X"2D",X"05",X"2D",X"06",X"2D",X"06",X"2D",X"04",X"27",X"04",X"27",X"05",X"27",X"05",X"27",
		X"06",X"27",X"06",X"27",X"05",X"0D",X"05",X"0D",X"06",X"0D",X"06",X"0D",X"02",X"6D",X"03",X"6C",
		X"03",X"6C",X"04",X"6C",X"04",X"6C",X"05",X"6C",X"06",X"0D",X"06",X"0D",X"06",X"07",X"06",X"07",
		X"06",X"07",X"06",X"07",X"02",X"4E",X"03",X"4E",X"03",X"4E",X"04",X"4E",X"04",X"4E",X"05",X"4E",
		X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"01",X"54",X"02",X"54",X"06",X"07",X"06",X"07",
		X"06",X"07",X"06",X"07",X"01",X"58",X"02",X"58",X"AF",X"32",X"2D",X"80",X"ED",X"43",X"85",X"81",
		X"C9",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"26",X"7B",X"0A",X"0F",X"0F",X"0F",
		X"5F",X"E6",X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",X"26",X"7D",X"0A",X"77",X"03",X"26",
		X"79",X"CB",X"FD",X"EB",X"60",X"69",X"CF",X"22",X"85",X"81",X"21",X"80",X"93",X"3A",X"42",X"80",
		X"87",X"87",X"87",X"D5",X"EF",X"D1",X"EB",X"72",X"2D",X"73",X"60",X"69",X"01",X"40",X"00",X"ED",
		X"B0",X"3A",X"42",X"80",X"3C",X"FE",X"0C",X"38",X"01",X"AF",X"32",X"42",X"80",X"C9",X"3E",X"31",
		X"32",X"7E",X"7F",X"3C",X"32",X"7C",X"7F",X"AF",X"32",X"2E",X"80",X"ED",X"43",X"85",X"81",X"C9",
		X"3E",X"01",X"32",X"2E",X"80",X"ED",X"43",X"85",X"81",X"C9",X"21",X"1E",X"79",X"36",X"02",X"2C",
		X"36",X"00",X"24",X"36",X"F8",X"24",X"36",X"0E",X"2D",X"36",X"80",X"24",X"36",X"00",X"ED",X"43",
		X"85",X"81",X"AF",X"32",X"2F",X"80",X"21",X"76",X"06",X"11",X"02",X"7F",X"06",X"0F",X"7E",X"12",
		X"1C",X"1C",X"23",X"10",X"F9",X"C9",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"52",
		X"51",X"50",X"4F",X"4A",X"4B",X"ED",X"43",X"85",X"81",X"3E",X"01",X"32",X"2F",X"80",X"C9",X"2A",
		X"85",X"81",X"3A",X"11",X"80",X"BE",X"C0",X"23",X"4D",X"44",X"03",X"7E",X"21",X"A9",X"06",X"D7",
		X"7E",X"21",X"01",X"07",X"CF",X"5E",X"23",X"56",X"EB",X"E9",X"00",X"02",X"03",X"04",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0E",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"06",X"07",X"08",X"09",X"01",
		X"01",X"0A",X"0B",X"0C",X"0D",X"01",X"01",X"0F",X"10",X"11",X"00",X"00",X"12",X"13",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"14",X"15",X"16",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"17",X"31",X"07",X"3F",X"07",X"BD",X"03",X"D1",X"03",X"EF",X"03",X"FD",X"03",X"5D",X"07",X"D8",
		X"05",X"3E",X"04",X"48",X"04",X"8E",X"04",X"52",X"04",X"5C",X"04",X"66",X"04",X"67",X"07",X"E1",
		X"05",X"70",X"04",X"7A",X"04",X"2E",X"06",X"40",X"06",X"4A",X"06",X"85",X"06",X"84",X"04",X"0C",
		X"04",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"ED",X"43",X"85",X"81",X"C9",X"26",
		X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"26",X"7B",X"0A",X"0F",X"0F",X"0F",X"5F",X"E6",
		X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"22",
		X"84",X"03",X"ED",X"43",X"85",X"81",X"C9",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",
		X"26",X"7B",X"0A",X"0F",X"0F",X"0F",X"5F",X"E6",X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",
		X"2D",X"26",X"7E",X"0A",X"77",X"03",X"ED",X"43",X"85",X"81",X"C9",X"F7",X"3A",X"11",X"80",X"FE",
		X"0E",X"C8",X"F7",X"3A",X"11",X"80",X"FE",X"0E",X"C0",X"3A",X"87",X"81",X"3C",X"FE",X"10",X"20",
		X"02",X"3E",X"06",X"32",X"87",X"81",X"4F",X"21",X"BD",X"07",X"D7",X"7E",X"32",X"13",X"80",X"79",
		X"21",X"00",X"10",X"CF",X"5E",X"23",X"56",X"ED",X"53",X"85",X"81",X"18",X"CE",X"24",X"00",X"54",
		X"0E",X"40",X"1A",X"64",X"04",X"2A",X"5C",X"0E",X"04",X"38",X"54",X"1A",X"00",X"3A",X"AD",X"85",
		X"FE",X"00",X"C8",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"0F",X"E6",X"01",X"47",X"21",X"00",X"18",
		X"11",X"00",X"05",X"3A",X"21",X"80",X"A7",X"28",X"01",X"EB",X"4F",X"CD",X"0F",X"08",X"EB",X"3A",
		X"22",X"80",X"A7",X"3E",X"06",X"28",X"07",X"79",X"EE",X"01",X"4F",X"79",X"87",X"81",X"11",X"1F",
		X"08",X"EB",X"D7",X"EB",X"01",X"C0",X"03",X"1A",X"CD",X"28",X"08",X"13",X"10",X"F9",X"C9",X"D5",
		X"C5",X"3A",X"23",X"80",X"A0",X"28",X"02",X"0E",X"02",X"CD",X"FB",X"07",X"C1",X"D1",X"C9",X"01",
		X"1E",X"19",X"02",X"1E",X"19",X"24",X"24",X"24",X"E5",X"F5",X"CD",X"32",X"08",X"F1",X"77",X"E1",
		X"25",X"C9",X"3A",X"03",X"80",X"25",X"A7",X"3E",X"04",X"28",X"03",X"25",X"3E",X"18",X"85",X"E6",
		X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",X"67",X"E6",X"C0",X"B5",X"6F",X"7C",X"E6",X"07",X"81",
		X"67",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"96",
		X"20",X"10",X"C8",X"10",X"AF",X"11",X"3D",X"12",X"CD",X"12",X"A8",X"13",X"73",X"14",X"3F",X"15",
		X"9C",X"16",X"E8",X"16",X"42",X"18",X"24",X"19",X"7A",X"1A",X"29",X"1B",X"77",X"1B",X"F0",X"1C",
		X"0C",X"53",X"00",X"0C",X"FF",X"24",X"0F",X"FF",X"25",X"FF",X"FF",X"28",X"12",X"FF",X"29",X"1F",
		X"FE",X"2A",X"07",X"FE",X"2F",X"1F",X"FE",X"30",X"1F",X"FE",X"2B",X"07",X"FD",X"03",X"EB",X"03",
		X"D7",X"03",X"D6",X"1E",X"04",X"80",X"D6",X"1F",X"06",X"70",X"C3",X"05",X"B7",X"03",X"B6",X"1E",
		X"08",X"80",X"B6",X"26",X"0A",X"70",X"AB",X"1E",X"0C",X"58",X"A9",X"26",X"0E",X"58",X"A1",X"1F",
		X"10",X"40",X"9F",X"26",X"12",X"50",X"9F",X"05",X"9B",X"57",X"9B",X"57",X"93",X"03",X"83",X"03",
		X"7A",X"26",X"14",X"70",X"78",X"1F",X"16",X"70",X"73",X"03",X"69",X"1D",X"18",X"20",X"61",X"2C",
		X"1A",X"5A",X"60",X"25",X"1F",X"5F",X"57",X"5F",X"57",X"5E",X"2C",X"1C",X"5A",X"5B",X"2C",X"1E",
		X"5A",X"5B",X"03",X"53",X"03",X"47",X"03",X"44",X"54",X"00",X"3C",X"1E",X"04",X"60",X"3C",X"26",
		X"06",X"70",X"3B",X"02",X"03",X"27",X"1F",X"08",X"28",X"25",X"26",X"0A",X"38",X"23",X"1F",X"0C",
		X"48",X"23",X"26",X"0E",X"C0",X"21",X"26",X"10",X"58",X"1F",X"1F",X"12",X"68",X"17",X"05",X"17",
		X"1D",X"14",X"D0",X"15",X"2D",X"16",X"68",X"0D",X"FF",X"02",X"01",X"EF",X"05",X"E7",X"2E",X"04",
		X"9C",X"03",X"40",X"00",X"38",X"1C",X"FF",X"18",X"DD",X"26",X"06",X"70",X"DD",X"1E",X"08",X"60",
		X"D3",X"1F",X"0A",X"D0",X"D3",X"26",X"0C",X"C0",X"C9",X"26",X"0E",X"70",X"C9",X"26",X"10",X"60",
		X"C3",X"03",X"BB",X"2E",X"12",X"94",X"03",X"68",X"00",X"20",X"02",X"FF",X"00",X"B3",X"26",X"14",
		X"68",X"B3",X"05",X"A7",X"2E",X"16",X"94",X"03",X"58",X"00",X"C0",X"18",X"FF",X"00",X"A3",X"26",
		X"18",X"70",X"A3",X"1F",X"1A",X"60",X"A3",X"03",X"95",X"26",X"1C",X"68",X"93",X"03",X"83",X"05",
		X"79",X"1F",X"1E",X"D0",X"6F",X"26",X"04",X"70",X"6F",X"1F",X"06",X"60",X"6D",X"1F",X"08",X"70",
		X"6D",X"26",X"0A",X"60",X"67",X"1D",X"0C",X"20",X"67",X"2E",X"0E",X"D8",X"04",X"48",X"1C",X"50",
		X"00",X"20",X"1C",X"FF",X"00",X"5B",X"03",X"4B",X"05",X"47",X"2E",X"10",X"A4",X"04",X"08",X"00",
		X"50",X"08",X"60",X"00",X"C0",X"02",X"44",X"2E",X"12",X"34",X"03",X"78",X"00",X"A8",X"04",X"C0",
		X"06",X"3E",X"1D",X"14",X"70",X"39",X"1F",X"16",X"D0",X"39",X"26",X"18",X"C0",X"33",X"03",X"27",
		X"1E",X"1A",X"90",X"25",X"1F",X"1C",X"80",X"25",X"2E",X"1E",X"60",X"02",X"90",X"04",X"C0",X"08",
		X"23",X"1E",X"04",X"70",X"23",X"05",X"21",X"1F",X"06",X"60",X"1F",X"1E",X"08",X"50",X"1C",X"28",
		X"18",X"1B",X"02",X"01",X"17",X"26",X"0A",X"A0",X"17",X"26",X"0C",X"90",X"15",X"05",X"13",X"1F",
		X"0E",X"B0",X"13",X"1B",X"10",X"A0",X"13",X"1B",X"12",X"90",X"13",X"1F",X"14",X"80",X"0D",X"FF",
		X"22",X"04",X"FF",X"28",X"14",X"EF",X"1F",X"16",X"40",X"E4",X"22",X"02",X"BD",X"26",X"18",X"A0",
		X"BB",X"1F",X"1A",X"A0",X"B8",X"22",X"02",X"A3",X"20",X"1C",X"C0",X"9F",X"1D",X"04",X"E0",X"93",
		X"0F",X"74",X"91",X"26",X"06",X"80",X"8F",X"1E",X"08",X"80",X"8C",X"54",X"00",X"87",X"1E",X"0A",
		X"90",X"87",X"1F",X"0C",X"80",X"83",X"23",X"83",X"57",X"7B",X"03",X"6B",X"1F",X"0E",X"D0",X"6B",
		X"26",X"10",X"A0",X"63",X"05",X"63",X"26",X"12",X"60",X"5B",X"1F",X"14",X"60",X"57",X"36",X"16",
		X"78",X"57",X"03",X"4B",X"57",X"49",X"1F",X"18",X"D0",X"49",X"26",X"1A",X"A0",X"43",X"03",X"36",
		X"1E",X"1C",X"C0",X"36",X"26",X"1E",X"A8",X"36",X"1F",X"04",X"90",X"36",X"1E",X"06",X"78",X"2C",
		X"1F",X"08",X"90",X"2B",X"05",X"1F",X"1F",X"0A",X"80",X"1F",X"26",X"0C",X"60",X"1F",X"1F",X"0E",
		X"40",X"18",X"24",X"03",X"17",X"21",X"10",X"60",X"17",X"1D",X"14",X"20",X"0D",X"FF",X"02",X"01",
		X"F0",X"05",X"ED",X"2E",X"16",X"9C",X"03",X"A0",X"00",X"80",X"10",X"80",X"00",X"E3",X"2E",X"18",
		X"2C",X"02",X"90",X"00",X"80",X"1C",X"DB",X"1E",X"1A",X"60",X"DB",X"1F",X"1C",X"50",X"D1",X"2E",
		X"1E",X"7C",X"03",X"38",X"00",X"80",X"02",X"C0",X"00",X"CB",X"03",X"C5",X"26",X"04",X"B0",X"C5",
		X"1F",X"06",X"A0",X"C5",X"1D",X"08",X"60",X"BD",X"2E",X"0A",X"24",X"03",X"48",X"00",X"28",X"02",
		X"FF",X"00",X"BB",X"05",X"AF",X"1F",X"0C",X"50",X"AD",X"1F",X"0E",X"40",X"AA",X"26",X"10",X"50",
		X"A7",X"26",X"12",X"40",X"A7",X"2E",X"14",X"24",X"04",X"60",X"00",X"D8",X"10",X"28",X"08",X"FF",
		X"02",X"9F",X"03",X"8B",X"05",X"87",X"22",X"01",X"83",X"23",X"73",X"02",X"45",X"73",X"4E",X"2F",
		X"73",X"4C",X"63",X"05",X"5F",X"02",X"45",X"4F",X"05",X"3F",X"22",X"04",X"33",X"23",X"31",X"23",
		X"2B",X"23",X"2B",X"57",X"28",X"03",X"20",X"4D",X"20",X"03",X"10",X"03",X"0D",X"FF",X"24",X"07",
		X"FF",X"2F",X"0F",X"FE",X"30",X"0F",X"FE",X"28",X"1C",X"FD",X"03",X"EF",X"03",X"E3",X"57",X"E3",
		X"05",X"DD",X"1F",X"04",X"A0",X"DD",X"1E",X"06",X"90",X"DB",X"21",X"08",X"70",X"DB",X"1E",X"0C",
		X"A0",X"DB",X"1F",X"0E",X"90",X"D1",X"3D",X"10",X"C0",X"CB",X"03",X"BF",X"3E",X"12",X"A0",X"BB",
		X"03",X"BB",X"3E",X"14",X"60",X"B7",X"3E",X"16",X"A0",X"B3",X"03",X"B3",X"3F",X"18",X"60",X"AF",
		X"3F",X"1A",X"20",X"A7",X"05",X"A5",X"21",X"1C",X"68",X"9B",X"3E",X"04",X"40",X"97",X"3E",X"06",
		X"80",X"95",X"3E",X"08",X"A0",X"93",X"3E",X"0A",X"C0",X"93",X"03",X"7B",X"05",X"7B",X"54",X"00",
		X"71",X"2E",X"0C",X"60",X"0C",X"30",X"00",X"30",X"10",X"30",X"18",X"30",X"08",X"30",X"00",X"30",
		X"10",X"30",X"18",X"30",X"08",X"30",X"00",X"30",X"10",X"30",X"18",X"30",X"08",X"71",X"1D",X"0E",
		X"20",X"70",X"25",X"0F",X"70",X"24",X"0F",X"6B",X"1E",X"10",X"80",X"69",X"26",X"12",X"80",X"67",
		X"1E",X"14",X"80",X"65",X"26",X"16",X"80",X"63",X"03",X"4B",X"05",X"4B",X"1F",X"18",X"C0",X"3F",
		X"03",X"35",X"1F",X"1A",X"80",X"32",X"2E",X"1C",X"D8",X"03",X"C0",X"18",X"18",X"10",X"C0",X"08",
		X"31",X"1D",X"1E",X"40",X"2F",X"05",X"23",X"2E",X"04",X"C0",X"01",X"C0",X"18",X"20",X"2E",X"06",
		X"20",X"01",X"C0",X"08",X"1D",X"2E",X"08",X"C0",X"01",X"C0",X"18",X"17",X"1F",X"0A",X"C0",X"17",
		X"21",X"0C",X"80",X"17",X"1F",X"10",X"40",X"0D",X"FF",X"24",X"07",X"F3",X"26",X"04",X"C0",X"F3",
		X"1E",X"06",X"B0",X"EB",X"2E",X"08",X"3C",X"03",X"C0",X"00",X"C0",X"10",X"C0",X"00",X"DB",X"2E",
		X"0A",X"34",X"02",X"20",X"02",X"FF",X"00",X"D7",X"1F",X"0C",X"C0",X"D5",X"26",X"0E",X"D0",X"D5",
		X"30",X"FF",X"CB",X"2E",X"10",X"1C",X"03",X"98",X"00",X"80",X"02",X"40",X"00",X"BB",X"2E",X"12",
		X"1C",X"01",X"FF",X"00",X"B6",X"1E",X"14",X"C0",X"B6",X"26",X"16",X"D0",X"B4",X"30",X"0F",X"AA",
		X"1F",X"18",X"B0",X"AA",X"1F",X"1A",X"A0",X"9F",X"21",X"1C",X"A0",X"9B",X"03",X"8B",X"1D",X"04",
		X"30",X"83",X"05",X"77",X"2D",X"06",X"C0",X"6F",X"3A",X"10",X"48",X"6B",X"38",X"12",X"60",X"6B",
		X"38",X"14",X"30",X"67",X"38",X"16",X"48",X"5F",X"1F",X"18",X"80",X"5D",X"26",X"1A",X"70",X"56",
		X"2E",X"1C",X"14",X"0B",X"40",X"00",X"38",X"04",X"50",X"06",X"38",X"04",X"3C",X"08",X"30",X"04",
		X"20",X"00",X"20",X"10",X"20",X"00",X"20",X"10",X"20",X"00",X"55",X"26",X"1E",X"70",X"4F",X"26",
		X"04",X"80",X"4F",X"1D",X"06",X"D0",X"48",X"2E",X"08",X"D8",X"03",X"08",X"00",X"58",X"18",X"FF",
		X"00",X"41",X"2E",X"0A",X"48",X"02",X"78",X"00",X"FF",X"08",X"33",X"1F",X"0C",X"70",X"27",X"26",
		X"0E",X"70",X"25",X"26",X"10",X"90",X"23",X"26",X"12",X"B0",X"17",X"21",X"14",X"C0",X"17",X"21",
		X"18",X"A0",X"0D",X"FF",X"22",X"08",X"F1",X"1F",X"04",X"80",X"EF",X"1E",X"06",X"80",X"ED",X"22",
		X"03",X"CA",X"30",X"3F",X"C9",X"2E",X"08",X"70",X"06",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",
		X"1C",X"60",X"00",X"60",X"04",X"C6",X"2E",X"0A",X"58",X"06",X"30",X"04",X"60",X"0C",X"60",X"10",
		X"60",X"14",X"60",X"1C",X"60",X"00",X"C3",X"2E",X"0C",X"40",X"06",X"60",X"04",X"60",X"0C",X"60",
		X"10",X"60",X"14",X"60",X"1C",X"60",X"00",X"C0",X"2E",X"0E",X"40",X"06",X"30",X"00",X"60",X"04",
		X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"BD",X"2E",X"10",X"40",X"06",X"60",X"00",X"60",
		X"04",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"BA",X"2E",X"12",X"58",X"07",X"30",X"1C",
		X"60",X"00",X"60",X"04",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"A7",X"2F",X"07",X"A1",
		X"1E",X"14",X"70",X"9F",X"26",X"16",X"60",X"9E",X"22",X"02",X"9D",X"1F",X"18",X"50",X"9B",X"1E",
		X"1A",X"40",X"83",X"10",X"74",X"81",X"26",X"1C",X"40",X"7B",X"1D",X"1E",X"D8",X"6C",X"23",X"6B",
		X"1E",X"04",X"B0",X"6B",X"1F",X"06",X"80",X"6B",X"1E",X"08",X"50",X"6B",X"1F",X"0A",X"20",X"66",
		X"54",X"00",X"4F",X"22",X"10",X"36",X"1F",X"0C",X"48",X"36",X"1F",X"0E",X"20",X"2B",X"3B",X"10",
		X"C0",X"27",X"3C",X"12",X"A0",X"17",X"11",X"76",X"11",X"1D",X"14",X"20",X"0F",X"23",X"0D",X"F3",
		X"03",X"F3",X"30",X"FF",X"F3",X"57",X"EE",X"2E",X"04",X"14",X"05",X"08",X"00",X"A0",X"08",X"30",
		X"0C",X"FF",X"10",X"FF",X"00",X"EA",X"05",X"E5",X"26",X"06",X"30",X"E5",X"26",X"08",X"C8",X"E2",
		X"1F",X"0A",X"48",X"E2",X"1F",X"0C",X"B0",X"DF",X"26",X"0E",X"60",X"DF",X"26",X"10",X"98",X"CC",
		X"1E",X"12",X"40",X"C8",X"26",X"14",X"60",X"C8",X"26",X"16",X"20",X"C7",X"21",X"18",X"48",X"C3",
		X"1E",X"1C",X"40",X"BB",X"57",X"B3",X"1F",X"1E",X"48",X"A8",X"03",X"A5",X"2E",X"04",X"A0",X"02",
		X"B0",X"02",X"80",X"00",X"A5",X"2E",X"06",X"74",X"04",X"78",X"00",X"50",X"18",X"50",X"08",X"80",
		X"00",X"A5",X"2E",X"08",X"14",X"04",X"78",X"00",X"50",X"08",X"50",X"18",X"80",X"00",X"9B",X"05",
		X"93",X"2E",X"0A",X"7C",X"05",X"A0",X"00",X"F0",X"10",X"30",X"0F",X"30",X"1F",X"80",X"00",X"93",
		X"1F",X"0C",X"50",X"93",X"26",X"0E",X"40",X"93",X"2E",X"10",X"14",X"03",X"AC",X"00",X"FF",X"10",
		X"80",X"00",X"83",X"03",X"7F",X"2E",X"12",X"84",X"07",X"50",X"00",X"C0",X"10",X"50",X"10",X"28",
		X"0B",X"50",X"10",X"70",X"0C",X"60",X"0D",X"77",X"1D",X"14",X"D0",X"73",X"05",X"73",X"26",X"04",
		X"58",X"73",X"1F",X"06",X"48",X"6D",X"2E",X"16",X"14",X"01",X"80",X"00",X"6A",X"2E",X"18",X"14",
		X"01",X"80",X"00",X"67",X"2E",X"1A",X"14",X"01",X"80",X"00",X"64",X"35",X"1C",X"14",X"61",X"35",
		X"1E",X"14",X"47",X"2E",X"08",X"80",X"06",X"08",X"00",X"58",X"08",X"60",X"00",X"60",X"02",X"80",
		X"00",X"60",X"04",X"47",X"2E",X"0A",X"68",X"08",X"08",X"00",X"88",X"08",X"60",X"00",X"60",X"1C",
		X"38",X"00",X"18",X"12",X"A8",X"14",X"80",X"00",X"47",X"2E",X"0C",X"50",X"03",X"08",X"00",X"78",
		X"18",X"80",X"00",X"37",X"1B",X"0E",X"B8",X"37",X"1B",X"10",X"48",X"27",X"2E",X"12",X"50",X"02",
		X"68",X"04",X"E0",X"08",X"24",X"2E",X"14",X"38",X"02",X"98",X"04",X"E0",X"08",X"21",X"2E",X"16",
		X"20",X"02",X"C8",X"04",X"E0",X"08",X"1F",X"2E",X"18",X"90",X"03",X"08",X"1C",X"E0",X"00",X"D0",
		X"08",X"1C",X"2E",X"1A",X"A8",X"03",X"38",X"1C",X"E0",X"00",X"D0",X"08",X"19",X"2E",X"1C",X"C0",
		X"03",X"68",X"1C",X"E0",X"00",X"D0",X"08",X"19",X"1F",X"1E",X"88",X"19",X"1F",X"04",X"68",X"19",
		X"1F",X"06",X"48",X"13",X"1B",X"08",X"88",X"13",X"1B",X"0C",X"48",X"0D",X"FB",X"02",X"1F",X"F5",
		X"1D",X"10",X"A0",X"F3",X"1D",X"12",X"80",X"F1",X"1D",X"14",X"60",X"EF",X"1D",X"16",X"40",X"EB",
		X"05",X"E3",X"02",X"38",X"D5",X"21",X"18",X"50",X"D3",X"05",X"D1",X"57",X"CF",X"03",X"C7",X"03",
		X"C3",X"02",X"6F",X"BF",X"05",X"B3",X"33",X"9F",X"34",X"87",X"18",X"76",X"85",X"4E",X"0F",X"83",
		X"4C",X"73",X"02",X"45",X"63",X"05",X"63",X"57",X"5B",X"02",X"65",X"4B",X"05",X"3F",X"03",X"2F",
		X"03",X"20",X"4D",X"1F",X"03",X"10",X"05",X"0D",X"FF",X"03",X"FF",X"30",X"3F",X"F7",X"05",X"F3",
		X"57",X"EF",X"03",X"E3",X"05",X"DB",X"03",X"CF",X"05",X"C6",X"2E",X"1C",X"D8",X"08",X"60",X"14",
		X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"C6",X"2E",
		X"1E",X"98",X"08",X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"60",
		X"10",X"60",X"00",X"C6",X"2E",X"04",X"58",X"08",X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",X"1C",
		X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",X"1C",X"BE",X"2E",X"06",X"B8",X"08",X"40",X"08",X"60",
		X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"BE",X"2E",X"08",
		X"78",X"08",X"40",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",
		X"60",X"08",X"B8",X"2E",X"0A",X"C8",X"07",X"40",X"1C",X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",
		X"1C",X"60",X"0C",X"60",X"1C",X"B8",X"2E",X"0C",X"98",X"07",X"40",X"00",X"60",X"10",X"60",X"00",
		X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"B8",X"2E",X"0E",X"68",X"07",X"40",X"04",X"60",
		X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"A9",X"1E",X"10",X"B0",X"A9",
		X"1E",X"12",X"90",X"A7",X"1E",X"14",X"A0",X"A5",X"1E",X"16",X"B0",X"A5",X"1E",X"18",X"90",X"9B",
		X"18",X"76",X"91",X"1F",X"1A",X"40",X"8F",X"1F",X"1C",X"40",X"8B",X"18",X"76",X"87",X"1E",X"1E",
		X"50",X"87",X"1E",X"04",X"40",X"7B",X"18",X"76",X"6F",X"1F",X"06",X"C0",X"6F",X"1E",X"08",X"A0",
		X"6F",X"1F",X"0A",X"80",X"64",X"2E",X"0C",X"98",X"10",X"80",X"18",X"80",X"10",X"80",X"09",X"20",
		X"0C",X"40",X"18",X"20",X"1A",X"10",X"18",X"28",X"10",X"10",X"08",X"20",X"06",X"48",X"08",X"18",
		X"0C",X"70",X"18",X"A0",X"13",X"98",X"08",X"80",X"04",X"47",X"1D",X"0E",X"C0",X"47",X"1D",X"10",
		X"A0",X"47",X"1D",X"12",X"80",X"47",X"1D",X"14",X"60",X"43",X"1D",X"16",X"C0",X"43",X"1D",X"18",
		X"A0",X"43",X"1D",X"1A",X"80",X"43",X"1D",X"1C",X"60",X"36",X"1E",X"1E",X"80",X"36",X"26",X"04",
		X"60",X"36",X"1E",X"06",X"40",X"2B",X"1F",X"08",X"50",X"21",X"20",X"0A",X"80",X"1B",X"20",X"0E",
		X"80",X"19",X"1B",X"12",X"D0",X"19",X"1B",X"14",X"20",X"13",X"1B",X"16",X"D0",X"13",X"1B",X"18",
		X"20",X"0D",X"FB",X"11",X"74",X"F3",X"22",X"08",X"E9",X"2D",X"04",X"60",X"E6",X"22",X"08",X"E4",
		X"2E",X"0E",X"9C",X"01",X"80",X"00",X"DC",X"2E",X"10",X"2C",X"02",X"F8",X"00",X"40",X"1C",X"CB",
		X"26",X"12",X"B0",X"CB",X"1F",X"14",X"A0",X"CB",X"2E",X"16",X"2C",X"07",X"70",X"00",X"E8",X"10",
		X"20",X"12",X"B8",X"10",X"B8",X"00",X"20",X"02",X"20",X"00",X"C3",X"23",X"C3",X"35",X"18",X"7C",
		X"BF",X"35",X"1A",X"7C",X"BB",X"35",X"1C",X"7C",X"B7",X"39",X"1E",X"7C",X"AF",X"3B",X"04",X"24",
		X"A7",X"3B",X"06",X"24",X"A3",X"22",X"0C",X"9B",X"03",X"8B",X"05",X"8B",X"1D",X"08",X"70",X"84",
		X"1D",X"0A",X"70",X"84",X"22",X"04",X"77",X"2E",X"0C",X"34",X"09",X"60",X"00",X"A0",X"10",X"28",
		X"0D",X"50",X"10",X"70",X"0C",X"60",X"0D",X"40",X"06",X"30",X"04",X"20",X"08",X"75",X"1F",X"0E",
		X"60",X"73",X"1E",X"10",X"70",X"73",X"23",X"71",X"1F",X"12",X"80",X"6F",X"1E",X"14",X"90",X"6D",
		X"1F",X"16",X"A0",X"6B",X"1E",X"18",X"B0",X"69",X"1F",X"1A",X"C0",X"67",X"1E",X"1C",X"D0",X"67",
		X"57",X"63",X"03",X"63",X"03",X"53",X"22",X"10",X"43",X"03",X"3B",X"05",X"2B",X"2E",X"1E",X"E0",
		X"05",X"08",X"00",X"60",X"18",X"20",X"1C",X"D8",X"18",X"20",X"14",X"27",X"21",X"04",X"68",X"23",
		X"23",X"1E",X"1D",X"08",X"20",X"1D",X"1F",X"0A",X"D0",X"1D",X"1F",X"0C",X"A0",X"1B",X"1D",X"0E",
		X"38",X"18",X"1D",X"10",X"50",X"17",X"1E",X"12",X"D0",X"17",X"1E",X"14",X"A0",X"15",X"1D",X"16",
		X"68",X"13",X"23",X"0D",X"FF",X"30",X"0F",X"FF",X"29",X"0F",X"FF",X"2B",X"03",X"FF",X"2A",X"03",
		X"F3",X"57",X"EE",X"2E",X"04",X"14",X"09",X"08",X"00",X"A0",X"08",X"30",X"0C",X"48",X"10",X"30",
		X"00",X"50",X"10",X"68",X"00",X"30",X"1C",X"20",X"18",X"E5",X"1B",X"06",X"C0",X"E5",X"1F",X"08",
		X"B0",X"E5",X"1F",X"0A",X"48",X"E5",X"1B",X"0C",X"38",X"E3",X"1F",X"0E",X"C0",X"E3",X"1B",X"10",
		X"B0",X"E3",X"1B",X"12",X"48",X"E3",X"1F",X"14",X"38",X"DC",X"2E",X"16",X"7C",X"04",X"08",X"10",
		X"78",X"00",X"50",X"10",X"40",X"00",X"C9",X"35",X"18",X"48",X"C9",X"35",X"1A",X"38",X"C7",X"35",
		X"1C",X"48",X"C7",X"35",X"1E",X"38",X"BD",X"1E",X"04",X"B0",X"BB",X"1E",X"06",X"B0",X"BB",X"1E",
		X"08",X"90",X"B9",X"1E",X"0A",X"90",X"B3",X"2E",X"0C",X"CC",X"01",X"20",X"00",X"A7",X"2E",X"0E",
		X"74",X"04",X"58",X"00",X"A0",X"18",X"A0",X"08",X"20",X"00",X"A3",X"2E",X"10",X"14",X"01",X"20",
		X"00",X"A3",X"57",X"A1",X"2E",X"12",X"14",X"01",X"20",X"00",X"97",X"03",X"93",X"2E",X"14",X"7C",
		X"02",X"98",X"00",X"20",X"02",X"8D",X"1D",X"16",X"E0",X"8D",X"1D",X"18",X"D0",X"8B",X"1D",X"1A",
		X"E0",X"8B",X"1D",X"1C",X"D0",X"87",X"05",X"83",X"03",X"77",X"1E",X"1E",X"60",X"77",X"1F",X"04",
		X"50",X"73",X"05",X"73",X"2E",X"06",X"14",X"04",X"70",X"00",X"E0",X"10",X"A0",X"10",X"20",X"00",
		X"6F",X"1F",X"08",X"60",X"6F",X"1E",X"0A",X"50",X"6B",X"03",X"5B",X"05",X"55",X"1B",X"0C",X"A8",
		X"47",X"2E",X"0E",X"78",X"03",X"08",X"00",X"C8",X"18",X"20",X"00",X"47",X"2E",X"10",X"90",X"03",
		X"08",X"00",X"F8",X"18",X"20",X"00",X"47",X"2E",X"12",X"A8",X"04",X"08",X"00",X"E0",X"18",X"48",
		X"18",X"20",X"00",X"37",X"1F",X"14",X"C0",X"37",X"1F",X"16",X"B0",X"30",X"1B",X"18",X"68",X"2E",
		X"1B",X"1A",X"58",X"2C",X"1B",X"1C",X"48",X"2A",X"1B",X"1E",X"38",X"27",X"36",X"04",X"14",X"23",
		X"36",X"06",X"14",X"1F",X"36",X"08",X"14",X"1B",X"39",X"0A",X"14",X"18",X"2E",X"0C",X"88",X"08",
		X"40",X"00",X"80",X"18",X"80",X"10",X"80",X"08",X"80",X"00",X"80",X"18",X"80",X"10",X"80",X"08",
		X"18",X"2E",X"0E",X"48",X"08",X"40",X"10",X"80",X"08",X"80",X"00",X"80",X"18",X"80",X"10",X"80",
		X"08",X"80",X"00",X"80",X"18",X"17",X"21",X"10",X"70",X"0D",X"F7",X"1B",X"14",X"20",X"F3",X"1B",
		X"16",X"A0",X"F3",X"1B",X"18",X"70",X"ED",X"1F",X"1A",X"A0",X"EB",X"1F",X"1C",X"90",X"E9",X"1F",
		X"1E",X"80",X"E7",X"1F",X"04",X"70",X"E3",X"57",X"DF",X"1B",X"06",X"C0",X"D9",X"1B",X"08",X"C0",
		X"D3",X"03",X"BB",X"05",X"B1",X"21",X"0A",X"B0",X"B1",X"21",X"0E",X"50",X"AB",X"03",X"A1",X"3E",
		X"12",X"90",X"9D",X"3E",X"14",X"70",X"99",X"40",X"16",X"50",X"95",X"3E",X"18",X"30",X"93",X"05",
		X"8D",X"40",X"1A",X"50",X"89",X"3E",X"1C",X"70",X"85",X"3E",X"1E",X"90",X"81",X"3E",X"04",X"B0",
		X"7B",X"03",X"71",X"1F",X"06",X"D0",X"6F",X"26",X"08",X"C0",X"6D",X"1F",X"0A",X"B0",X"6B",X"26",
		X"0C",X"A0",X"69",X"1F",X"0E",X"90",X"63",X"05",X"5F",X"57",X"5B",X"02",X"EC",X"43",X"05",X"40",
		X"1D",X"10",X"30",X"40",X"1D",X"12",X"20",X"3B",X"03",X"36",X"1B",X"14",X"C0",X"25",X"2E",X"16",
		X"E0",X"02",X"C0",X"18",X"C0",X"08",X"25",X"2E",X"18",X"10",X"02",X"C0",X"08",X"C0",X"18",X"23",
		X"2E",X"1A",X"D0",X"02",X"A0",X"18",X"A0",X"08",X"23",X"2E",X"1C",X"20",X"02",X"A0",X"08",X"A0",
		X"18",X"23",X"05",X"1B",X"02",X"E6",X"0E",X"05",X"0D",X"FF",X"02",X"6D",X"F7",X"05",X"F3",X"22",
		X"02",X"E7",X"23",X"E7",X"4E",X"0F",X"E7",X"02",X"F1",X"E3",X"4C",X"DF",X"05",X"DB",X"02",X"34",
		X"D5",X"05",X"CB",X"02",X"49",X"C5",X"05",X"BB",X"02",X"3E",X"BB",X"4D",X"AB",X"05",X"A1",X"33",
		X"8F",X"34",X"7F",X"02",X"46",X"77",X"05",X"73",X"18",X"76",X"67",X"4C",X"67",X"02",X"66",X"65",
		X"05",X"5B",X"02",X"21",X"55",X"05",X"4B",X"03",X"3B",X"05",X"37",X"57",X"33",X"4D",X"33",X"03",
		X"23",X"05",X"1B",X"03",X"1F",X"05",X"0D",X"FF",X"02",X"08",X"F3",X"05",X"EF",X"2E",X"04",X"3C",
		X"05",X"80",X"00",X"80",X"10",X"70",X"00",X"70",X"10",X"70",X"00",X"EE",X"1D",X"06",X"D0",X"EE",
		X"26",X"08",X"80",X"E6",X"2E",X"0A",X"3C",X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"E5",X"1F",
		X"0C",X"80",X"DE",X"2E",X"0E",X"3C",X"03",X"60",X"00",X"60",X"10",X"60",X"00",X"D7",X"1F",X"10",
		X"C0",X"D7",X"2E",X"12",X"26",X"06",X"50",X"02",X"78",X"12",X"18",X"10",X"18",X"00",X"80",X"02",
		X"20",X"00",X"D5",X"1F",X"14",X"D0",X"D2",X"26",X"16",X"50",X"CD",X"2E",X"18",X"1C",X"04",X"40",
		X"00",X"A0",X"10",X"D8",X"00",X"20",X"02",X"C6",X"1F",X"04",X"50",X"C2",X"2E",X"1A",X"1C",X"03",
		X"80",X"00",X"A0",X"00",X"20",X"02",X"BE",X"35",X"1C",X"1C",X"BA",X"3B",X"1E",X"1C",X"B6",X"1F",
		X"06",X"D0",X"B6",X"26",X"08",X"C0",X"B6",X"1D",X"0A",X"50",X"B3",X"03",X"A9",X"1D",X"0C",X"B0",
		X"A3",X"03",X"A0",X"26",X"0E",X"A0",X"A0",X"1F",X"10",X"90",X"93",X"05",X"8B",X"03",X"7B",X"05",
		X"78",X"21",X"12",X"C8",X"76",X"2E",X"16",X"78",X"08",X"50",X"14",X"50",X"04",X"50",X"14",X"50",
		X"04",X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"76",X"2E",X"18",X"18",X"08",X"50",X"0C",
		X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"6B",X"2E",
		X"1A",X"70",X"09",X"40",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",
		X"1C",X"50",X"0C",X"50",X"1C",X"6B",X"2E",X"1C",X"20",X"09",X"40",X"04",X"50",X"14",X"50",X"04",
		X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"61",X"2E",X"1E",X"A4",
		X"07",X"18",X"00",X"10",X"1C",X"60",X"18",X"38",X"14",X"40",X"16",X"60",X"1E",X"20",X"1C",X"5F",
		X"1F",X"04",X"80",X"5B",X"26",X"06",X"60",X"5B",X"1D",X"08",X"20",X"57",X"1F",X"0A",X"40",X"4E",
		X"2E",X"14",X"AC",X"06",X"50",X"00",X"A8",X"10",X"10",X"08",X"E0",X"18",X"A0",X"10",X"C0",X"00",
		X"48",X"2E",X"12",X"D4",X"06",X"08",X"00",X"90",X"18",X"10",X"08",X"A0",X"18",X"E0",X"10",X"C0",
		X"00",X"47",X"2E",X"10",X"44",X"06",X"18",X"00",X"70",X"08",X"70",X"18",X"C0",X"10",X"F0",X"10",
		X"20",X"18",X"3B",X"26",X"16",X"B0",X"37",X"1F",X"18",X"90",X"1F",X"1B",X"1A",X"90",X"1F",X"1B",
		X"1C",X"70",X"1F",X"1B",X"1E",X"50",X"1B",X"1B",X"04",X"70",X"1B",X"35",X"06",X"24",X"1B",X"02",
		X"3F",X"17",X"3B",X"08",X"24",X"15",X"21",X"0A",X"C0",X"13",X"3B",X"0E",X"24",X"0F",X"05",X"0D",
		X"01",X"57",X"FF",X"03",X"F3",X"1D",X"14",X"20",X"EF",X"05",X"E7",X"2E",X"16",X"9C",X"03",X"40",
		X"00",X"38",X"1C",X"40",X"18",X"E5",X"1B",X"18",X"60",X"E1",X"2E",X"1A",X"24",X"03",X"80",X"00",
		X"80",X"10",X"80",X"00",X"DD",X"2E",X"1C",X"9C",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"D7",
		X"1B",X"1E",X"78",X"D7",X"1B",X"04",X"48",X"D7",X"2E",X"06",X"24",X"03",X"80",X"00",X"80",X"10",
		X"80",X"00",X"D3",X"2E",X"08",X"9C",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"D3",X"1B",X"0A",
		X"60",X"CD",X"2E",X"0C",X"24",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"CB",X"26",X"0E",X"C8",
		X"CB",X"26",X"10",X"60",X"C5",X"2E",X"12",X"9C",X"08",X"60",X"00",X"78",X"10",X"20",X"12",X"F8",
		X"10",X"58",X"10",X"50",X"18",X"50",X"08",X"20",X"00",X"C5",X"2E",X"14",X"24",X"08",X"60",X"00",
		X"90",X"10",X"20",X"0C",X"E0",X"10",X"58",X"10",X"50",X"08",X"50",X"18",X"20",X"00",X"C5",X"57",
		X"C3",X"03",X"BB",X"3B",X"16",X"70",X"BB",X"3B",X"18",X"50",X"B7",X"3C",X"1A",X"70",X"B7",X"3B",
		X"1C",X"50",X"B3",X"03",X"A3",X"03",X"95",X"1F",X"1E",X"80",X"93",X"05",X"93",X"1F",X"04",X"70",
		X"91",X"1F",X"06",X"60",X"8F",X"1F",X"08",X"50",X"85",X"03",X"7D",X"26",X"0A",X"E0",X"7D",X"26",
		X"0C",X"88",X"7D",X"26",X"0E",X"50",X"79",X"26",X"10",X"C0",X"79",X"26",X"12",X"6C",X"79",X"26",
		X"14",X"18",X"6F",X"21",X"16",X"80",X"6F",X"3B",X"1A",X"34",X"6B",X"3B",X"1C",X"34",X"6B",X"05",
		X"67",X"1D",X"1E",X"B0",X"65",X"1D",X"04",X"A0",X"63",X"03",X"53",X"05",X"4F",X"26",X"06",X"80",
		X"4C",X"1F",X"08",X"68",X"4B",X"2E",X"0A",X"34",X"02",X"A0",X"04",X"20",X"06",X"44",X"1B",X"0C",
		X"70",X"3E",X"1B",X"0E",X"C0",X"3E",X"1D",X"10",X"70",X"3E",X"1B",X"12",X"18",X"38",X"1B",X"14",
		X"70",X"37",X"2E",X"16",X"A4",X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"37",X"2E",X"04",X"34",
		X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"33",X"02",X"E6",X"23",X"05",X"22",X"2E",X"06",X"48",
		X"02",X"B8",X"04",X"20",X"08",X"22",X"2E",X"08",X"34",X"01",X"20",X"00",X"1B",X"2E",X"0A",X"48",
		X"08",X"30",X"00",X"A0",X"04",X"A0",X"10",X"80",X"0C",X"40",X"10",X"80",X"18",X"A0",X"18",X"20",
		X"00",X"17",X"21",X"18",X"90",X"17",X"21",X"1C",X"70",X"17",X"02",X"7E",X"0F",X"05",X"0F",X"30",
		X"1F",X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"68",
		X"31",X"00",X"A3",X"C3",X"7F",X"00",X"00",X"00",X"87",X"30",X"05",X"24",X"18",X"02",X"00",X"00",
		X"85",X"6F",X"D0",X"24",X"C9",X"00",X"00",X"00",X"77",X"23",X"10",X"FC",X"C9",X"00",X"00",X"00",
		X"3A",X"98",X"A0",X"A7",X"28",X"0B",X"3D",X"28",X"04",X"21",X"90",X"A0",X"C9",X"21",X"8B",X"A0",
		X"C9",X"21",X"86",X"A0",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"3A",X"80",X"A0",X"A7",X"28",X"03",X"F1",X"ED",X"45",
		X"3E",X"01",X"32",X"80",X"A0",X"32",X"22",X"68",X"AF",X"32",X"22",X"68",X"C3",X"9A",X"00",X"3E",
		X"01",X"32",X"22",X"68",X"CD",X"53",X"0A",X"21",X"00",X"A0",X"36",X"00",X"11",X"01",X"A0",X"01",
		X"FF",X"00",X"ED",X"B0",X"AF",X"32",X"22",X"68",X"18",X"FE",X"21",X"81",X"A0",X"36",X"00",X"11",
		X"82",X"A0",X"01",X"0F",X"00",X"ED",X"B0",X"3A",X"94",X"A0",X"A7",X"28",X"0B",X"21",X"00",X"A0",
		X"86",X"77",X"AF",X"32",X"94",X"A0",X"18",X"16",X"3A",X"28",X"80",X"A7",X"28",X"10",X"21",X"01",
		X"A0",X"36",X"00",X"11",X"02",X"A0",X"01",X"26",X"00",X"ED",X"B0",X"C3",X"D2",X"01",X"3A",X"02",
		X"A0",X"A7",X"28",X"0B",X"21",X"95",X"A0",X"36",X"02",X"CD",X"8B",X"02",X"C3",X"D2",X"01",X"3A",
		X"03",X"A0",X"A7",X"28",X"0B",X"21",X"95",X"A0",X"36",X"03",X"CD",X"8B",X"02",X"C3",X"D2",X"01",
		X"3A",X"04",X"A0",X"A7",X"28",X"0B",X"21",X"95",X"A0",X"36",X"04",X"CD",X"8B",X"02",X"C3",X"D2",
		X"01",X"3A",X"0E",X"A0",X"A7",X"28",X"08",X"21",X"95",X"A0",X"36",X"0E",X"CD",X"8B",X"02",X"3A",
		X"0D",X"A0",X"A7",X"28",X"08",X"21",X"95",X"A0",X"36",X"0D",X"CD",X"8B",X"02",X"21",X"95",X"A0",
		X"36",X"05",X"3A",X"05",X"A0",X"A7",X"28",X"09",X"AF",X"32",X"05",X"A0",X"CD",X"14",X"02",X"18",
		X"0A",X"3A",X"19",X"A0",X"A7",X"CA",X"3B",X"01",X"CD",X"48",X"02",X"3A",X"06",X"A0",X"A7",X"28",
		X"0A",X"21",X"95",X"A0",X"36",X"06",X"CD",X"8B",X"02",X"18",X"2E",X"3A",X"07",X"A0",X"A7",X"28",
		X"0A",X"21",X"95",X"A0",X"36",X"07",X"CD",X"8B",X"02",X"18",X"1E",X"3A",X"08",X"A0",X"A7",X"28",
		X"0A",X"21",X"95",X"A0",X"36",X"08",X"CD",X"8B",X"02",X"18",X"0E",X"3A",X"09",X"A0",X"A7",X"28",
		X"08",X"21",X"95",X"A0",X"36",X"09",X"CD",X"8B",X"02",X"21",X"95",X"A0",X"36",X"0A",X"3A",X"0A",
		X"A0",X"A7",X"28",X"09",X"AF",X"32",X"0A",X"A0",X"CD",X"14",X"02",X"18",X"28",X"3A",X"1E",X"A0",
		X"A7",X"28",X"05",X"CD",X"48",X"02",X"18",X"1D",X"21",X"95",X"A0",X"36",X"0B",X"3A",X"0B",X"A0",
		X"A7",X"28",X"09",X"AF",X"32",X"0B",X"A0",X"CD",X"14",X"02",X"18",X"26",X"3A",X"1F",X"A0",X"A7",
		X"28",X"03",X"CD",X"48",X"02",X"21",X"95",X"A0",X"36",X"0C",X"3A",X"0C",X"A0",X"A7",X"28",X"09",
		X"AF",X"32",X"0C",X"A0",X"CD",X"14",X"02",X"18",X"09",X"3A",X"20",X"A0",X"A7",X"28",X"03",X"CD",
		X"48",X"02",X"3A",X"00",X"A0",X"A7",X"28",X"0A",X"21",X"95",X"A0",X"36",X"00",X"CD",X"8B",X"02",
		X"18",X"0E",X"3A",X"01",X"A0",X"A7",X"28",X"08",X"21",X"95",X"A0",X"36",X"01",X"CD",X"8B",X"02",
		X"21",X"81",X"A0",X"11",X"10",X"68",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"91",X"A0",X"32",X"05",
		X"68",X"3A",X"92",X"A0",X"32",X"0A",X"68",X"3A",X"93",X"A0",X"32",X"0F",X"68",X"AF",X"32",X"80",
		X"A0",X"F1",X"ED",X"45",X"21",X"14",X"A0",X"3A",X"95",X"A0",X"D7",X"34",X"21",X"95",X"A0",X"7E",
		X"87",X"86",X"21",X"C0",X"04",X"D7",X"11",X"96",X"A0",X"01",X"03",X"00",X"ED",X"B0",X"21",X"97",
		X"A0",X"46",X"48",X"21",X"54",X"A0",X"3A",X"96",X"A0",X"D7",X"AF",X"DF",X"41",X"21",X"28",X"A0",
		X"3A",X"96",X"A0",X"D7",X"AF",X"DF",X"18",X"12",X"21",X"95",X"A0",X"7E",X"87",X"86",X"21",X"C0",
		X"04",X"D7",X"11",X"96",X"A0",X"01",X"03",X"00",X"ED",X"B0",X"CD",X"07",X"03",X"21",X"97",X"A0",
		X"35",X"28",X"0A",X"21",X"96",X"A0",X"34",X"21",X"98",X"A0",X"34",X"18",X"ED",X"3A",X"99",X"A0",
		X"A7",X"C8",X"AF",X"32",X"99",X"A0",X"21",X"14",X"A0",X"3A",X"95",X"A0",X"D7",X"36",X"00",X"21",
		X"33",X"04",X"3A",X"95",X"A0",X"CF",X"5E",X"23",X"56",X"EB",X"E9",X"21",X"95",X"A0",X"7E",X"87",
		X"86",X"21",X"C0",X"04",X"D7",X"11",X"96",X"A0",X"01",X"03",X"00",X"ED",X"B0",X"21",X"14",X"A0",
		X"3A",X"95",X"A0",X"D7",X"7E",X"A7",X"20",X"19",X"34",X"21",X"97",X"A0",X"46",X"48",X"21",X"54",
		X"A0",X"3A",X"96",X"A0",X"D7",X"AF",X"DF",X"41",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",X"AF",
		X"DF",X"CD",X"07",X"03",X"21",X"97",X"A0",X"35",X"28",X"0A",X"21",X"96",X"A0",X"34",X"21",X"98",
		X"A0",X"34",X"18",X"ED",X"3A",X"99",X"A0",X"A7",X"C8",X"AF",X"32",X"99",X"A0",X"21",X"14",X"A0",
		X"3A",X"95",X"A0",X"D7",X"36",X"00",X"21",X"00",X"A0",X"3A",X"95",X"A0",X"D7",X"3A",X"95",X"A0",
		X"A7",X"28",X"12",X"FE",X"14",X"28",X"0E",X"36",X"00",X"21",X"33",X"04",X"3A",X"95",X"A0",X"CF",
		X"5E",X"23",X"56",X"EB",X"E9",X"35",X"C9",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",X"34",X"3A",
		X"96",X"A0",X"21",X"8A",X"04",X"CF",X"5E",X"23",X"56",X"21",X"54",X"A0",X"3A",X"96",X"A0",X"D7",
		X"7E",X"EB",X"D7",X"22",X"9A",X"A0",X"7E",X"3C",X"C2",X"34",X"03",X"E7",X"36",X"00",X"3E",X"01",
		X"32",X"99",X"A0",X"C9",X"21",X"FC",X"04",X"3A",X"96",X"A0",X"D7",X"7E",X"A7",X"28",X"05",X"11",
		X"82",X"05",X"18",X"03",X"11",X"68",X"05",X"2A",X"9A",X"A0",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"EB",X"CF",X"4E",X"23",X"46",X"EB",X"7E",X"E6",X"0F",X"28",X"07",X"CB",X"38",X"CB",X"19",
		X"3D",X"20",X"F9",X"3A",X"98",X"A0",X"A7",X"28",X"0D",X"3D",X"28",X"05",X"21",X"8C",X"A0",X"18",
		X"08",X"21",X"87",X"A0",X"18",X"03",X"21",X"82",X"A0",X"71",X"7E",X"0F",X"0F",X"0F",X"0F",X"23",
		X"77",X"23",X"70",X"7E",X"0F",X"0F",X"0F",X"0F",X"23",X"77",X"EB",X"E7",X"EB",X"2A",X"9A",X"A0",
		X"7E",X"D6",X"C0",X"28",X"4A",X"3A",X"96",X"A0",X"21",X"32",X"05",X"D7",X"A7",X"28",X"21",X"3D",
		X"28",X"0F",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",X"7E",X"FE",X"06",X"30",X"12",X"2F",X"18",
		X"33",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",X"7E",X"FE",X"08",X"30",X"03",X"87",X"18",X"24",
		X"21",X"4D",X"05",X"3A",X"96",X"A0",X"D7",X"7E",X"A7",X"28",X"17",X"47",X"21",X"28",X"A0",X"3A",
		X"96",X"A0",X"D7",X"7E",X"90",X"38",X"0B",X"D6",X"0A",X"30",X"04",X"ED",X"44",X"18",X"05",X"AF",
		X"18",X"02",X"3E",X"0A",X"12",X"21",X"91",X"A0",X"3A",X"98",X"A0",X"D7",X"EB",X"21",X"17",X"05",
		X"3A",X"96",X"A0",X"D7",X"ED",X"A0",X"21",X"ED",X"04",X"3A",X"95",X"A0",X"D7",X"7E",X"2A",X"9A",
		X"A0",X"23",X"5E",X"16",X"00",X"21",X"00",X"00",X"06",X"08",X"CB",X"3F",X"30",X"01",X"19",X"CB",
		X"23",X"CB",X"12",X"10",X"F5",X"45",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",X"78",X"BE",X"C0",
		X"21",X"54",X"A0",X"3A",X"96",X"A0",X"D7",X"34",X"34",X"21",X"28",X"A0",X"3A",X"96",X"A0",X"D7",
		X"36",X"00",X"C9",X"6F",X"04",X"6F",X"04",X"51",X"04",X"51",X"04",X"6F",X"04",X"51",X"04",X"51",
		X"04",X"60",X"04",X"51",X"04",X"51",X"04",X"67",X"04",X"51",X"04",X"51",X"04",X"52",X"04",X"51",
		X"04",X"C9",X"AF",X"32",X"05",X"A0",X"32",X"19",X"A0",X"AF",X"32",X"09",X"A0",X"32",X"1D",X"A0",
		X"AF",X"32",X"0C",X"A0",X"32",X"20",X"A0",X"AF",X"32",X"0B",X"A0",X"32",X"1F",X"A0",X"C9",X"21",
		X"05",X"A0",X"11",X"06",X"A0",X"01",X"09",X"00",X"36",X"00",X"ED",X"B0",X"21",X"19",X"A0",X"11",
		X"1A",X"A0",X"01",X"09",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"9C",X"05",X"DD",X"05",X"1E",X"06",
		X"65",X"06",X"AC",X"06",X"F5",X"06",X"38",X"07",X"6B",X"07",X"9E",X"07",X"DF",X"07",X"20",X"08",
		X"D9",X"09",X"DB",X"09",X"DD",X"09",X"B3",X"08",X"B9",X"08",X"BF",X"08",X"3D",X"09",X"E1",X"08",
		X"9E",X"09",X"C8",X"08",X"38",X"09",X"3A",X"09",X"47",X"08",X"58",X"08",X"EC",X"09",X"11",X"0A",
		X"00",X"02",X"00",X"02",X"03",X"00",X"05",X"03",X"00",X"08",X"03",X"00",X"0C",X"03",X"00",X"0E",
		X"03",X"00",X"11",X"01",X"01",X"12",X"01",X"01",X"13",X"01",X"02",X"14",X"01",X"02",X"15",X"02",
		X"00",X"17",X"01",X"00",X"18",X"01",X"01",X"19",X"01",X"00",X"1A",X"01",X"00",X"02",X"10",X"0A",
		X"0C",X"10",X"06",X"01",X"05",X"01",X"01",X"06",X"01",X"02",X"04",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"02",X"02",X"05",X"04",X"03",X"07",X"05",X"05",X"05",
		X"05",X"06",X"01",X"01",X"01",X"01",X"05",X"07",X"03",X"03",X"01",X"06",X"01",X"01",X"04",X"01",
		X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"02",X"00",X"00",X"02",X"02",X"00",X"02",X"02",X"02",
		X"00",X"00",X"00",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"04",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"D0",X"5A",X"37",X"60",X"EF",X"65",X"FF",X"6B",
		X"6B",X"72",X"39",X"79",X"6E",X"80",X"11",X"88",X"29",X"90",X"BC",X"98",X"D0",X"A1",X"70",X"AB",
		X"00",X"00",X"11",X"5C",X"8B",X"61",X"58",X"67",X"7D",X"6D",X"00",X"74",X"E6",X"7A",X"35",X"82",
		X"F2",X"89",X"27",X"92",X"D8",X"9A",X"0C",X"A4",X"CE",X"AD",X"00",X"00",X"79",X"01",X"69",X"01",
		X"59",X"01",X"49",X"01",X"39",X"01",X"29",X"01",X"19",X"01",X"09",X"01",X"78",X"01",X"68",X"01",
		X"58",X"01",X"48",X"01",X"38",X"01",X"28",X"01",X"18",X"01",X"08",X"01",X"77",X"01",X"67",X"01",
		X"57",X"01",X"47",X"01",X"37",X"01",X"52",X"01",X"17",X"01",X"07",X"01",X"76",X"01",X"66",X"01",
		X"56",X"01",X"46",X"01",X"36",X"01",X"26",X"01",X"16",X"01",X"06",X"01",X"FF",X"89",X"01",X"79",
		X"01",X"69",X"01",X"59",X"01",X"49",X"01",X"39",X"01",X"29",X"01",X"19",X"01",X"88",X"01",X"78",
		X"01",X"68",X"01",X"58",X"01",X"48",X"01",X"38",X"01",X"28",X"01",X"18",X"01",X"87",X"01",X"77",
		X"01",X"67",X"01",X"57",X"01",X"47",X"01",X"32",X"01",X"27",X"01",X"17",X"01",X"86",X"01",X"76",
		X"01",X"66",X"01",X"56",X"01",X"46",X"01",X"36",X"01",X"26",X"01",X"16",X"01",X"FF",X"56",X"04",
		X"C0",X"01",X"06",X"01",X"56",X"01",X"96",X"01",X"05",X"01",X"96",X"01",X"C0",X"01",X"56",X"01",
		X"76",X"01",X"C0",X"01",X"76",X"01",X"76",X"01",X"C0",X"01",X"26",X"02",X"C0",X"01",X"76",X"01",
		X"56",X"01",X"C0",X"01",X"46",X"01",X"56",X"04",X"C0",X"01",X"06",X"01",X"56",X"01",X"96",X"01",
		X"05",X"01",X"96",X"01",X"C0",X"01",X"56",X"01",X"66",X"01",X"C0",X"01",X"66",X"01",X"66",X"01",
		X"C0",X"01",X"56",X"07",X"FF",X"97",X"04",X"C0",X"01",X"97",X"01",X"97",X"01",X"06",X"01",X"56",
		X"01",X"06",X"01",X"C0",X"01",X"97",X"01",X"A7",X"01",X"C0",X"01",X"A7",X"01",X"A7",X"01",X"C0",
		X"01",X"A7",X"02",X"C0",X"01",X"A7",X"01",X"A7",X"01",X"C0",X"01",X"A7",X"01",X"97",X"04",X"C0",
		X"01",X"97",X"01",X"97",X"01",X"97",X"01",X"97",X"01",X"97",X"01",X"C0",X"01",X"97",X"01",X"A7",
		X"01",X"C0",X"01",X"A7",X"01",X"A7",X"01",X"C0",X"01",X"97",X"07",X"FF",X"59",X"01",X"59",X"01",
		X"59",X"01",X"59",X"01",X"C0",X"02",X"59",X"01",X"59",X"01",X"59",X"01",X"59",X"01",X"C0",X"02",
		X"59",X"01",X"59",X"01",X"59",X"01",X"59",X"01",X"C0",X"02",X"59",X"01",X"59",X"01",X"59",X"01",
		X"59",X"01",X"C0",X"02",X"59",X"01",X"59",X"01",X"59",X"01",X"59",X"01",X"C0",X"02",X"59",X"01",
		X"59",X"01",X"59",X"01",X"59",X"01",X"C0",X"02",X"59",X"01",X"59",X"01",X"59",X"01",X"59",X"01",
		X"C0",X"01",X"59",X"07",X"FF",X"07",X"01",X"07",X"01",X"07",X"02",X"07",X"02",X"07",X"02",X"07",
		X"02",X"07",X"02",X"07",X"02",X"27",X"02",X"47",X"02",X"57",X"02",X"57",X"02",X"57",X"02",X"57",
		X"02",X"57",X"02",X"97",X"02",X"77",X"02",X"57",X"02",X"77",X"02",X"77",X"02",X"77",X"02",X"77",
		X"02",X"77",X"02",X"26",X"02",X"06",X"02",X"A7",X"02",X"97",X"02",X"97",X"02",X"97",X"02",X"97",
		X"02",X"97",X"02",X"A7",X"02",X"06",X"02",X"FF",X"C0",X"02",X"A8",X"02",X"A8",X"02",X"C0",X"04",
		X"A8",X"02",X"A8",X"02",X"C0",X"04",X"98",X"02",X"98",X"02",X"C0",X"04",X"98",X"02",X"98",X"02",
		X"C0",X"04",X"A8",X"02",X"A8",X"02",X"C0",X"04",X"A8",X"02",X"A8",X"02",X"C0",X"04",X"98",X"02",
		X"98",X"02",X"C0",X"04",X"98",X"02",X"98",X"02",X"C0",X"02",X"FF",X"C0",X"02",X"08",X"02",X"08",
		X"02",X"C0",X"04",X"08",X"02",X"08",X"02",X"C0",X"04",X"58",X"02",X"58",X"02",X"C0",X"04",X"58",
		X"02",X"58",X"02",X"C0",X"04",X"08",X"02",X"08",X"02",X"C0",X"04",X"08",X"02",X"08",X"02",X"C0",
		X"04",X"58",X"02",X"58",X"02",X"C0",X"04",X"58",X"02",X"58",X"02",X"C0",X"02",X"FF",X"96",X"04",
		X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",
		X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",
		X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",
		X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"96",X"04",X"FF",X"56",
		X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",
		X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",
		X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",
		X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"56",X"04",X"FF",
		X"58",X"01",X"07",X"01",X"46",X"0D",X"26",X"01",X"16",X"03",X"46",X"01",X"26",X"0C",X"58",X"01",
		X"07",X"01",X"36",X"0D",X"26",X"01",X"36",X"03",X"56",X"01",X"76",X"03",X"56",X"01",X"36",X"03",
		X"26",X"01",X"06",X"03",X"26",X"01",X"FF",X"69",X"01",X"64",X"01",X"79",X"01",X"14",X"01",X"89",
		X"01",X"85",X"01",X"99",X"01",X"35",X"01",X"FF",X"06",X"01",X"16",X"01",X"26",X"01",X"36",X"01",
		X"46",X"01",X"36",X"01",X"26",X"01",X"16",X"01",X"06",X"01",X"B7",X"01",X"A7",X"01",X"97",X"01",
		X"87",X"01",X"77",X"01",X"67",X"01",X"57",X"01",X"47",X"01",X"37",X"01",X"27",X"01",X"17",X"01",
		X"07",X"01",X"B8",X"01",X"A8",X"01",X"98",X"01",X"88",X"01",X"78",X"01",X"68",X"01",X"58",X"01",
		X"48",X"01",X"38",X"01",X"28",X"01",X"18",X"01",X"08",X"01",X"B9",X"01",X"A9",X"01",X"99",X"01",
		X"89",X"01",X"79",X"01",X"69",X"01",X"59",X"01",X"49",X"01",X"39",X"01",X"29",X"01",X"19",X"01",
		X"09",X"01",X"FF",X"04",X"01",X"74",X"01",X"24",X"01",X"94",X"01",X"44",X"01",X"B4",X"01",X"64",
		X"01",X"14",X"01",X"84",X"01",X"34",X"01",X"FF",X"0A",X"01",X"19",X"01",X"0A",X"01",X"19",X"01",
		X"25",X"01",X"34",X"01",X"25",X"01",X"34",X"01",X"43",X"01",X"52",X"01",X"43",X"01",X"52",X"01",
		X"FF",X"09",X"01",X"19",X"01",X"09",X"01",X"29",X"01",X"09",X"01",X"39",X"01",X"09",X"01",X"49",
		X"01",X"09",X"01",X"39",X"01",X"09",X"01",X"29",X"01",X"09",X"01",X"19",X"01",X"09",X"01",X"19",
		X"01",X"09",X"01",X"29",X"01",X"09",X"01",X"39",X"01",X"09",X"01",X"49",X"01",X"09",X"01",X"39",
		X"01",X"09",X"01",X"29",X"01",X"09",X"01",X"19",X"01",X"09",X"01",X"19",X"01",X"09",X"01",X"29",
		X"01",X"09",X"01",X"39",X"01",X"09",X"01",X"49",X"01",X"09",X"01",X"39",X"01",X"09",X"01",X"29",
		X"01",X"09",X"01",X"19",X"01",X"09",X"01",X"FF",X"05",X"01",X"15",X"05",X"FF",X"04",X"01",X"29",
		X"01",X"14",X"01",X"29",X"01",X"04",X"01",X"39",X"01",X"14",X"01",X"39",X"01",X"04",X"01",X"49",
		X"01",X"14",X"01",X"49",X"01",X"04",X"01",X"59",X"01",X"14",X"01",X"59",X"01",X"04",X"01",X"29",
		X"01",X"14",X"01",X"29",X"01",X"04",X"01",X"39",X"01",X"14",X"01",X"39",X"01",X"04",X"01",X"49",
		X"01",X"14",X"01",X"49",X"01",X"04",X"01",X"59",X"01",X"14",X"01",X"59",X"01",X"04",X"01",X"29",
		X"01",X"14",X"01",X"29",X"01",X"04",X"01",X"39",X"01",X"14",X"01",X"39",X"01",X"04",X"01",X"49",
		X"01",X"14",X"01",X"49",X"01",X"04",X"01",X"59",X"01",X"14",X"01",X"59",X"01",X"FF",X"05",X"01",
		X"15",X"01",X"35",X"01",X"65",X"01",X"A5",X"01",X"65",X"01",X"35",X"01",X"25",X"02",X"15",X"02",
		X"05",X"03",X"06",X"03",X"07",X"04",X"08",X"04",X"09",X"08",X"0A",X"08",X"09",X"08",X"0A",X"08",
		X"09",X"08",X"0A",X"08",X"09",X"08",X"0A",X"08",X"09",X"08",X"0A",X"08",X"09",X"08",X"0A",X"08",
		X"09",X"08",X"0A",X"08",X"09",X"08",X"0A",X"08",X"FF",X"05",X"01",X"76",X"01",X"46",X"01",X"06",
		X"01",X"77",X"01",X"06",X"01",X"46",X"01",X"76",X"01",X"05",X"01",X"FF",X"26",X"01",X"56",X"01",
		X"76",X"01",X"96",X"01",X"05",X"01",X"25",X"01",X"26",X"01",X"56",X"01",X"76",X"01",X"96",X"01",
		X"05",X"01",X"25",X"01",X"26",X"01",X"56",X"01",X"76",X"01",X"96",X"01",X"05",X"01",X"25",X"01",
		X"FF",X"06",X"01",X"05",X"01",X"B6",X"01",X"05",X"01",X"45",X"01",X"05",X"01",X"B6",X"01",X"05",
		X"01",X"06",X"01",X"05",X"01",X"A6",X"01",X"05",X"01",X"45",X"01",X"05",X"01",X"A6",X"01",X"05",
		X"01",X"06",X"01",X"05",X"01",X"96",X"01",X"05",X"01",X"45",X"01",X"05",X"01",X"96",X"01",X"05",
		X"01",X"06",X"01",X"05",X"01",X"86",X"01",X"05",X"01",X"45",X"01",X"05",X"01",X"86",X"01",X"05",
		X"01",X"FF",X"E3",X"11",X"71",X"85",X"21",X"00",X"00",X"0E",X"10",X"06",X"00",X"3E",X"01",X"32",
		X"22",X"68",X"78",X"86",X"12",X"23",X"47",X"79",X"BC",X"20",X"F2",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7C",X"82",X"82",X"82",X"FE",X"FE",X"7C",X"00",X"00",X"00",X"FE",X"FE",X"FE",X"80",X"00",X"00",
		X"62",X"F2",X"F2",X"92",X"9E",X"9E",X"8E",X"00",X"6C",X"FE",X"FE",X"92",X"92",X"82",X"44",X"00",
		X"04",X"FE",X"FE",X"FE",X"84",X"44",X"3C",X"00",X"8C",X"9E",X"9E",X"92",X"F2",X"F2",X"F2",X"00",
		X"8C",X"9E",X"9E",X"92",X"F2",X"F2",X"7C",X"00",X"C0",X"F0",X"FE",X"BE",X"8E",X"80",X"C0",X"00",
		X"6C",X"9E",X"9E",X"92",X"F2",X"F2",X"6C",X"00",X"7C",X"9E",X"9E",X"92",X"F2",X"F2",X"62",X"00",
		X"7E",X"FE",X"FE",X"88",X"88",X"88",X"7E",X"00",X"6C",X"92",X"92",X"92",X"FE",X"FE",X"FE",X"00",
		X"82",X"82",X"82",X"82",X"FE",X"FE",X"7C",X"00",X"7C",X"FE",X"FE",X"82",X"82",X"82",X"FE",X"00",
		X"92",X"92",X"92",X"92",X"FE",X"FE",X"FE",X"00",X"90",X"90",X"90",X"90",X"FE",X"FE",X"FE",X"00",
		X"5C",X"DE",X"DE",X"92",X"92",X"82",X"7C",X"00",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"FE",X"00",
		X"00",X"00",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"02",X"02",X"00",
		X"86",X"4E",X"3E",X"18",X"F0",X"F0",X"FE",X"00",X"02",X"02",X"02",X"02",X"FE",X"FE",X"FE",X"00",
		X"7E",X"FE",X"80",X"FE",X"FE",X"80",X"FE",X"00",X"7E",X"FE",X"FE",X"80",X"80",X"80",X"FE",X"00",
		X"7C",X"82",X"82",X"82",X"FE",X"FE",X"7C",X"00",X"70",X"88",X"88",X"88",X"FE",X"FE",X"FE",X"00",
		X"7E",X"8E",X"82",X"82",X"FE",X"FE",X"7C",X"00",X"6E",X"9E",X"9E",X"90",X"F0",X"F0",X"FE",X"00",
		X"4C",X"9E",X"9E",X"92",X"F2",X"F2",X"64",X"00",X"80",X"80",X"FE",X"FE",X"FE",X"80",X"80",X"00",
		X"FC",X"02",X"02",X"02",X"FE",X"FE",X"FC",X"00",X"F0",X"08",X"0C",X"0E",X"FC",X"F8",X"F0",X"00",
		X"FC",X"02",X"FE",X"FE",X"02",X"FE",X"FC",X"00",X"86",X"4E",X"3E",X"38",X"F8",X"E4",X"C2",X"00",
		X"E0",X"10",X"1E",X"1E",X"FE",X"F0",X"E0",X"00",X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"7E",X"D2",X"7E",X"0E",X"06",X"00",
		X"00",X"00",X"00",X"00",X"06",X"07",X"01",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"3C",X"42",X"B9",X"A9",X"BD",X"BD",X"42",X"3C",X"0A",X"44",X"EA",X"F2",X"BE",X"5E",X"0C",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"9A",X"8A",X"80",X"40",X"00",
		X"00",X"60",X"F0",X"FA",X"FA",X"60",X"00",X"00",X"BD",X"BD",X"42",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"A5",X"A5",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"00",X"00",
		X"DB",X"DB",X"DF",X"0E",X"00",X"00",X"7F",X"FF",X"FF",X"00",X"00",X"7F",X"FF",X"FF",X"DB",X"DB",
		X"FF",X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"FF",X"C3",X"C3",X"C3",X"FF",X"7E",X"00",X"00",X"7F",
		X"C3",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"C3",X"00",X"00",X"7E",X"FF",X"C3",X"C3",X"C3",X"C3",
		X"00",X"3E",X"3E",X"2A",X"2A",X"2E",X"00",X"00",X"00",X"3E",X"3E",X"22",X"E2",X"FE",X"00",X"00",
		X"00",X"22",X"22",X"22",X"3E",X"3E",X"00",X"00",X"00",X"FE",X"FE",X"22",X"22",X"3E",X"00",X"00",
		X"00",X"3A",X"3A",X"2A",X"2A",X"3E",X"00",X"00",X"00",X"20",X"A0",X"BE",X"FE",X"20",X"00",X"00",
		X"00",X"27",X"3F",X"25",X"3D",X"3B",X"00",X"00",X"00",X"3E",X"3E",X"20",X"E0",X"FE",X"00",X"00",
		X"00",X"00",X"BE",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"BD",X"01",X"00",X"00",X"00",
		X"00",X"26",X"1E",X"08",X"F8",X"FE",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",
		X"3E",X"3E",X"20",X"3E",X"3E",X"20",X"3E",X"00",X"00",X"3E",X"3E",X"20",X"20",X"3E",X"00",X"00",
		X"00",X"3E",X"3E",X"22",X"22",X"3E",X"00",X"00",X"00",X"3E",X"22",X"22",X"3F",X"3F",X"00",X"00",
		X"00",X"3F",X"23",X"22",X"3E",X"3E",X"00",X"00",X"00",X"00",X"20",X"10",X"3E",X"3E",X"00",X"00",
		X"00",X"2E",X"2E",X"2A",X"3A",X"3A",X"00",X"00",X"00",X"20",X"FE",X"3E",X"20",X"20",X"00",X"00",
		X"00",X"3E",X"02",X"02",X"3E",X"3E",X"00",X"00",X"00",X"38",X"04",X"06",X"3C",X"38",X"00",X"00",
		X"3E",X"02",X"3E",X"3E",X"02",X"3E",X"3E",X"00",X"00",X"26",X"1E",X"08",X"3C",X"32",X"00",X"00",
		X"00",X"3F",X"03",X"02",X"3E",X"3E",X"00",X"00",X"00",X"32",X"3A",X"3E",X"2E",X"26",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"70",X"78",X"7C",X"7E",X"7C",X"78",X"70",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"70",X"78",X"7C",X"7E",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"01",X"07",X"03",X"01",X"00",X"7F",X"7F",X"7F",X"7F",X"78",X"40",X"00",X"00",
		X"00",X"00",X"40",X"78",X"7F",X"7F",X"7F",X"7F",X"7C",X"7E",X"7F",X"7F",X"7F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"60",X"70",X"78",X"70",X"60",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"7F",X"7F",X"7E",X"7C",X"78",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"70",X"78",X"7C",X"7E",X"00",X"00",X"00",X"00",
		X"70",X"3F",X"1F",X"0E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"07",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"FC",X"FF",X"00",X"00",X"00",X"00",X"1F",X"03",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"1F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"01",X"03",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"01",X"03",X"06",X"0C",X"18",X"30",X"60",
		X"38",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"3E",X"3C",
		X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"7F",X"0F",X"01",X"03",X"07",X"0F",X"1F",X"00",X"00",X"00",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"80",X"C0",X"E0",X"F0",
		X"00",X"01",X"03",X"7F",X"3F",X"1F",X"0F",X"07",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"FF",X"FF",X"FF",X"FF",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7E",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",
		X"F0",X"F0",X"F0",X"F0",X"80",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"06",X"78",X"F0",X"F0",
		X"FF",X"3F",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"18",X"3E",X"7F",X"FF",
		X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"F7",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"FF",X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F1",X"F3",X"F7",X"FF",X"FF",X"FF",X"F7",X"F7",X"F6",X"F1",X"F3",X"F7",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"FF",X"FF",X"FF",X"F7",
		X"F0",X"F0",X"F0",X"F7",X"F7",X"F7",X"F7",X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F1",X"F3",X"F7",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F0",
		X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",
		X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"1E",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"0F",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",
		X"F8",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"80",X"C0",X"E0",X"F0",
		X"FF",X"F8",X"C0",X"00",X"80",X"C0",X"E0",X"F0",X"00",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"03",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FC",X"FE",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"03",X"07",X"0F",X"1F",X"BF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"78",X"30",X"01",X"FC",X"FC",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",
		X"FF",X"FF",X"FF",X"7F",X"0F",X"01",X"00",X"01",X"FF",X"FF",X"00",X"00",X"00",X"E0",X"FC",X"FF",
		X"FF",X"FE",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"83",X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"78",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",
		X"C0",X"86",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"7F",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",
		X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"FF",X"FF",X"FF",X"FE",X"F0",X"80",X"00",X"00",
		X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"7F",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"00",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"7F",X"FF",
		X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"3C",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"BC",
		X"FC",X"BC",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",
		X"C3",X"C3",X"C7",X"1F",X"3F",X"3E",X"3C",X"3C",X"03",X"03",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"C3",X"C3",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"3E",X"3F",X"1F",X"07",X"03",X"03",X"03",X"03",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",
		X"7C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FC",X"FE",X"FF",X"FF",X"FE",X"7C",X"38",X"10",
		X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FE",X"3F",X"1F",X"0F",X"07",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"07",X"0F",X"1F",X"3F",X"FE",X"FC",X"F0",X"C0",
		X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"CF",X"C7",X"E1",X"E0",X"E0",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0C",X"0C",X"00",X"81",X"87",X"01",X"07",X"EF",X"E7",X"E1",X"E0",X"0C",X"0C",
		X"8E",X"8C",X"0C",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"EF",X"E0",X"C3",X"C7",
		X"18",X"D8",X"FC",X"3F",X"07",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"07",X"3F",X"FC",X"D8",
		X"FC",X"D8",X"18",X"D8",X"FC",X"3F",X"07",X"00",X"7E",X"38",X"00",X"FF",X"FF",X"00",X"07",X"3F",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"81",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"41",X"41",X"41",X"7F",X"7F",X"3E",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"01",X"00",X"00",
		X"46",X"4F",X"4F",X"49",X"79",X"79",X"71",X"00",X"36",X"7F",X"7F",X"49",X"49",X"41",X"22",X"00",
		X"20",X"7F",X"7F",X"7F",X"21",X"22",X"3C",X"00",X"31",X"79",X"79",X"49",X"4F",X"4F",X"4F",X"00",
		X"31",X"79",X"79",X"49",X"4F",X"4F",X"3E",X"00",X"03",X"0F",X"7F",X"7D",X"71",X"01",X"03",X"00",
		X"36",X"79",X"79",X"49",X"4F",X"4F",X"36",X"00",X"3E",X"79",X"79",X"49",X"4F",X"4F",X"46",X"00",
		X"7E",X"7F",X"7F",X"11",X"11",X"11",X"7E",X"00",X"36",X"49",X"49",X"49",X"7F",X"7F",X"7F",X"00",
		X"41",X"41",X"41",X"41",X"7F",X"7F",X"3E",X"00",X"3E",X"7F",X"7F",X"41",X"41",X"41",X"7F",X"00",
		X"49",X"49",X"49",X"49",X"7F",X"7F",X"7F",X"00",X"09",X"09",X"09",X"09",X"7F",X"7F",X"7F",X"00",
		X"3A",X"7B",X"7B",X"49",X"49",X"41",X"3E",X"00",X"7F",X"08",X"08",X"08",X"7F",X"7F",X"7F",X"00",
		X"00",X"00",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"40",X"40",X"00",
		X"61",X"72",X"7C",X"18",X"0F",X"0F",X"7F",X"00",X"40",X"40",X"40",X"40",X"7F",X"7F",X"7F",X"00",
		X"7E",X"7F",X"01",X"7F",X"7F",X"01",X"7F",X"00",X"7E",X"7F",X"7F",X"01",X"01",X"01",X"7F",X"00",
		X"3E",X"41",X"41",X"41",X"7F",X"7F",X"3E",X"00",X"0E",X"11",X"11",X"11",X"7F",X"7F",X"7F",X"00",
		X"7E",X"71",X"41",X"41",X"7F",X"7F",X"3E",X"00",X"76",X"79",X"79",X"09",X"0F",X"0F",X"7F",X"00",
		X"32",X"79",X"79",X"49",X"4F",X"4F",X"26",X"00",X"01",X"01",X"7F",X"7F",X"7F",X"01",X"01",X"00",
		X"3F",X"40",X"40",X"40",X"7F",X"7F",X"3F",X"00",X"0F",X"10",X"30",X"70",X"3F",X"1F",X"0F",X"00",
		X"3F",X"40",X"7F",X"7F",X"40",X"7F",X"3F",X"00",X"61",X"72",X"7C",X"1C",X"1F",X"27",X"43",X"00",
		X"07",X"08",X"78",X"78",X"7F",X"0F",X"07",X"00",X"43",X"47",X"4F",X"5D",X"79",X"71",X"61",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"7E",X"4B",X"7E",X"70",X"60",X"00",
		X"00",X"00",X"00",X"00",X"60",X"E0",X"80",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"3C",X"42",X"9D",X"95",X"BD",X"BD",X"42",X"3C",X"50",X"22",X"57",X"4F",X"7D",X"7A",X"30",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"59",X"51",X"01",X"02",X"00",
		X"00",X"06",X"0F",X"5F",X"5F",X"06",X"00",X"00",X"BD",X"BD",X"42",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"A5",X"A5",X"03",X"03",X"03",X"03",X"FF",X"FF",X"00",X"00",
		X"DB",X"DB",X"FB",X"70",X"00",X"00",X"FE",X"FF",X"FF",X"00",X"00",X"FE",X"FF",X"FF",X"DB",X"DB",
		X"FF",X"03",X"03",X"FF",X"FF",X"03",X"03",X"FF",X"C3",X"C3",X"C3",X"FF",X"7E",X"00",X"00",X"FE",
		X"C3",X"FF",X"7E",X"00",X"00",X"C3",X"C3",X"C3",X"00",X"00",X"7E",X"FF",X"C3",X"C3",X"C3",X"C3",
		X"00",X"7C",X"7C",X"54",X"54",X"74",X"00",X"00",X"00",X"7C",X"7C",X"44",X"47",X"7F",X"00",X"00",
		X"00",X"44",X"44",X"44",X"7C",X"7C",X"00",X"00",X"00",X"7F",X"7F",X"44",X"44",X"7C",X"00",X"00",
		X"00",X"5C",X"5C",X"54",X"54",X"7C",X"00",X"00",X"00",X"04",X"05",X"7D",X"7F",X"04",X"00",X"00",
		X"00",X"E4",X"FC",X"A4",X"BC",X"DC",X"00",X"00",X"00",X"7C",X"7C",X"04",X"07",X"7F",X"00",X"00",
		X"00",X"00",X"7D",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"BD",X"80",X"00",X"00",X"00",
		X"00",X"64",X"78",X"10",X"1F",X"7F",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"04",X"7C",X"7C",X"04",X"7C",X"00",X"00",X"7C",X"7C",X"04",X"04",X"7C",X"00",X"00",
		X"00",X"7C",X"7C",X"44",X"44",X"7C",X"00",X"00",X"00",X"7C",X"44",X"44",X"FC",X"FC",X"00",X"00",
		X"00",X"FC",X"C4",X"44",X"7C",X"7C",X"00",X"00",X"00",X"00",X"04",X"08",X"7C",X"7C",X"00",X"00",
		X"00",X"74",X"74",X"54",X"5C",X"5C",X"00",X"00",X"00",X"04",X"7F",X"7C",X"04",X"04",X"00",X"00",
		X"00",X"7C",X"40",X"40",X"7C",X"7C",X"00",X"00",X"00",X"1C",X"20",X"60",X"3C",X"1C",X"00",X"00",
		X"7C",X"40",X"7C",X"7C",X"40",X"7C",X"7C",X"00",X"00",X"64",X"78",X"10",X"3C",X"4C",X"00",X"00",
		X"00",X"FC",X"C0",X"40",X"7C",X"7C",X"00",X"00",X"00",X"4C",X"5C",X"7C",X"74",X"64",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"70",X"00",X"00",X"0E",X"1E",X"3E",X"7E",X"3E",X"1E",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"1E",X"3E",X"7E",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"80",X"E0",X"C0",X"80",X"00",X"FE",X"FE",X"FE",X"FE",X"1E",X"02",X"00",X"00",
		X"00",X"00",X"02",X"1E",X"FE",X"FE",X"FE",X"FE",X"3E",X"7E",X"FE",X"FE",X"FE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"06",X"0E",X"1E",X"0E",X"06",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FE",X"7E",X"3E",X"1E",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"0E",X"1E",X"3E",X"7E",X"00",X"00",X"00",X"00",
		X"0E",X"FC",X"F8",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"E0",X"00",X"03",X"03",X"03",X"03",X"03",X"FF",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"3F",X"FF",X"00",X"00",X"00",X"00",X"F8",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"00",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"80",X"C0",X"60",X"30",X"18",X"0C",X"06",
		X"1C",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"7C",X"3C",
		X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FE",X"F0",X"80",X"C0",X"E0",X"F0",X"F8",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"C0",X"80",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"00",X"80",X"C0",X"FE",X"FC",X"F8",X"F0",X"E0",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0F",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"01",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"60",X"1E",X"0F",X"0F",
		X"FF",X"FC",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"18",X"7C",X"FE",X"FF",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CF",X"EF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"FF",X"EF",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"EF",X"EF",X"6F",X"8F",X"CF",X"EF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"FF",X"FF",X"FF",X"EF",
		X"0F",X"0F",X"0F",X"EF",X"EF",X"EF",X"EF",X"EF",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"0F",
		X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",
		X"EF",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"30",X"78",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"F0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"01",X"03",X"07",X"0F",
		X"FF",X"1F",X"03",X"00",X"01",X"03",X"07",X"0F",X"00",X"00",X"C0",X"F8",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"1F",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"3F",X"7F",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"C0",X"E0",X"F0",X"F8",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1E",X"0C",X"80",X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FE",X"F0",X"80",X"00",X"80",X"FF",X"FF",X"00",X"00",X"00",X"07",X"3F",X"FF",
		X"FF",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C1",X"E3",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"C1",X"80",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"3F",X"7F",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"03",X"61",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FE",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",
		X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"FC",X"FF",X"FF",X"FF",X"7F",X"0F",X"01",X"00",X"00",
		X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"7F",X"FF",X"FF",X"FE",X"FC",X"FE",X"FF",
		X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"00",X"FF",X"FF",X"FE",X"FC",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"3C",X"3C",X"3C",X"3D",X"3F",X"3F",X"3F",X"3F",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3D",X"3F",X"3F",X"3F",X"3D",
		X"3F",X"3D",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3D",X"3F",X"3F",X"3F",
		X"C3",X"C3",X"E3",X"F8",X"FC",X"7C",X"3C",X"3C",X"C0",X"C0",X"C3",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"C3",X"C3",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C3",X"C3",X"C3",X"C3",X"C3",
		X"7C",X"FC",X"F8",X"E0",X"C0",X"C0",X"C0",X"C0",X"3C",X"3D",X"3F",X"3F",X"3F",X"3F",X"3F",X"3D",
		X"3E",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"3F",X"7F",X"FF",X"FF",X"7F",X"3E",X"1C",X"08",
		X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"03",X"0F",X"3F",X"7F",X"FC",X"F8",X"F0",X"E0",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"E0",X"F0",X"F8",X"FC",X"7F",X"3F",X"0F",X"03",
		X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F3",X"E3",X"87",X"07",X"07",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"30",X"30",X"00",X"81",X"E1",X"80",X"E0",X"F7",X"E7",X"87",X"07",X"30",X"30",
		X"71",X"31",X"30",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F7",X"07",X"C3",X"E3",
		X"18",X"1B",X"3F",X"FC",X"E0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"E0",X"FC",X"3F",X"1B",
		X"3F",X"1B",X"18",X"1B",X"3F",X"FC",X"E0",X"00",X"7E",X"1C",X"00",X"FF",X"FF",X"00",X"E0",X"FC",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"81",X"E7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"FF",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",
		X"C0",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"1F",X"0F",X"07",X"03",X"03",X"0F",X"0F",
		X"0F",X"07",X"03",X"07",X"06",X"06",X"07",X"07",X"FF",X"FF",X"FF",X"FE",X"FE",X"FB",X"FB",X"FF",
		X"FF",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BB",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EF",X"EF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"9F",X"FF",X"FF",
		X"FF",X"DF",X"DF",X"FF",X"FF",X"FB",X"FB",X"FF",X"3F",X"0F",X"7F",X"FF",X"F0",X"C0",X"80",X"80",
		X"9F",X"BF",X"F0",X"C0",X"80",X"00",X"00",X"00",X"21",X"31",X"69",X"C7",X"1F",X"FF",X"FF",X"DF",
		X"FC",X"7C",X"3E",X"1F",X"07",X"03",X"01",X"00",X"0E",X"0F",X"07",X"03",X"03",X"01",X"01",X"01",
		X"FC",X"76",X"7E",X"3C",X"3E",X"3F",X"1F",X"0F",X"7F",X"9F",X"3F",X"BE",X"1F",X"BF",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FD",X"FD",X"FF",X"FB",X"FB",X"FF",X"FF",X"FF",X"FD",X"BD",X"BF",X"FF",X"F7",X"F7",X"FF",
		X"87",X"CF",X"E7",X"F7",X"FF",X"FF",X"FE",X"FE",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"7C",X"F9",X"FA",X"FA",X"FE",X"7D",X"7E",X"7E",X"3E",X"3E",X"3F",X"1F",X"1F",X"3F",X"7E",X"7C",
		X"F9",X"F3",X"E2",X"F7",X"F6",X"F2",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"9F",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"E3",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"78",X"FF",X"FF",X"3F",X"9F",X"DF",X"CF",X"EF",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F8",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"70",X"F8",X"78",X"78",X"78",X"78",X"7A",X"78",X"78",X"78",X"78",X"70",
		X"78",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"78",X"F0",X"78",X"F0",X"70",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F8",X"F0",X"78",X"F8",X"78",X"F8",X"5A",X"78",X"5A",X"F8",X"78",X"F8",X"78",X"F8",
		X"78",X"F8",X"78",X"F0",X"F8",X"F0",X"F8",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",
		X"F8",X"F8",X"F8",X"F0",X"78",X"F0",X"78",X"F0",X"78",X"F0",X"78",X"F0",X"F8",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"01",X"01",X"09",X"3D",X"3F",X"7F",X"7F",X"1F",X"6F",
		X"FF",X"FF",X"FC",X"F8",X"F8",X"F8",X"F0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"FE",
		X"DF",X"FF",X"7F",X"7F",X"1F",X"07",X"03",X"00",X"00",X"01",X"07",X"07",X"03",X"71",X"7D",X"BD",
		X"FF",X"FF",X"FC",X"F8",X"F8",X"F8",X"F0",X"C0",X"60",X"F0",X"F8",X"FC",X"FC",X"FC",X"F8",X"FE",
		X"FF",X"FF",X"FF",X"FC",X"F9",X"FC",X"D8",X"F7",X"FF",X"FF",X"FF",X"FD",X"78",X"75",X"FB",X"48",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"94",X"D2",X"B9",X"F3",X"E6",X"EC",X"FF",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"78",X"C1",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"6F",X"DF",
		X"F7",X"F7",X"EF",X"FF",X"BF",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"3C",X"E0",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"37",X"EF",
		X"FF",X"7F",X"7F",X"F7",X"EF",X"FE",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C7",X"EF",X"EF",X"FB",X"FB",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"FF",X"FF",X"FF",X"FD",X"F9",X"F9",X"FF",X"DB",X"DF",
		X"FF",X"FF",X"ED",X"DD",X"FD",X"F9",X"F9",X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"EF",X"E7",X"E6",X"E0",X"E0",X"C0",X"C0",X"80",
		X"2F",X"37",X"3F",X"1F",X"1F",X"07",X"01",X"00",X"3F",X"1F",X"3F",X"3F",X"3F",X"0F",X"07",X"03",
		X"00",X"01",X"01",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"0D",X"0B",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"03",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"3F",X"3F",X"E3",X"C0",X"F0",X"F8",X"F8",X"E0",X"C0",X"C0",
		X"04",X"EE",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"18",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"3F",X"1F",X"3F",X"3F",X"3F",X"3F",X"F0",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"C3",X"BD",X"66",X"5E",X"5E",X"66",X"BD",X"C3",X"C0",X"C0",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",
		X"78",X"38",X"3F",X"30",X"30",X"33",X"30",X"30",X"0E",X"06",X"C6",X"06",X"06",X"C6",X"06",X"0E",
		X"00",X"00",X"66",X"66",X"66",X"66",X"66",X"66",X"F0",X"60",X"67",X"67",X"67",X"67",X"60",X"70",
		X"1C",X"18",X"F9",X"F9",X"F9",X"F9",X"18",X"1C",X"07",X"03",X"F3",X"F3",X"F3",X"F3",X"03",X"07",
		X"C3",X"BD",X"46",X"5A",X"46",X"5A",X"9D",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"F8",
		X"00",X"00",X"00",X"CD",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"F0",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FE",X"FE",X"FC",X"F8",X"F8",X"FC",
		X"FF",X"FE",X"F8",X"E0",X"C0",X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FE",X"FE",X"F8",X"C0",X"00",
		X"FE",X"FC",X"E0",X"80",X"00",X"00",X"00",X"00",X"E9",X"EC",X"80",X"05",X"D1",X"89",X"1F",X"7F",
		X"31",X"8B",X"9B",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"13",X"CF",X"87",X"B7",X"1F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"76",X"00",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",X"03",
		X"FF",X"7F",X"0F",X"03",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"03",X"03",
		X"00",X"90",X"08",X"20",X"00",X"C0",X"00",X"00",X"01",X"B4",X"80",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"D0",X"E0",X"F8",X"FA",X"FF",X"FF",X"C0",X"C8",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",
		X"E0",X"B0",X"E0",X"C0",X"D0",X"F8",X"F0",X"C0",X"E0",X"E8",X"F0",X"E0",X"E8",X"F8",X"F0",X"C0",
		X"D0",X"D0",X"E0",X"E0",X"C0",X"E0",X"E8",X"F4",X"FF",X"FE",X"FD",X"F8",X"F8",X"F0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"08",X"A5",X"DF",X"FF",X"CF",X"9C",X"27",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"28",X"DE",X"FF",X"FF",X"65",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"12",X"BA",X"FF",X"FF",X"D5",X"0E",X"05",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"01",X"05",X"0B",X"67",X"FF",X"FF",X"FF",X"C3",X"BD",X"2A",X"02",X"00",X"00",
		X"0F",X"2F",X"5F",X"BF",X"9F",X"FF",X"FF",X"FF",X"0F",X"0F",X"07",X"07",X"1B",X"33",X"23",X"17",
		X"01",X"03",X"07",X"03",X"03",X"01",X"07",X"0B",X"01",X"03",X"07",X"0B",X"0B",X"05",X"05",X"07",
		X"0B",X"07",X"03",X"03",X"01",X"05",X"0F",X"05",X"FF",X"FF",X"BF",X"4F",X"C7",X"37",X"07",X"0B",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"60",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"3C",X"19",X"13",X"07",X"0F",X"FE",X"1F",X"CF",X"E7",X"F7",X"03",X"07",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"18",X"1E",X"1F",X"23",X"73",X"F9",X"E4",X"C2",X"81",X"00",X"00",
		X"00",X"70",X"F8",X"FC",X"FE",X"FF",X"FF",X"DF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"F6",X"76",X"B6",X"D6",X"E6",X"FE",X"FE",X"FE",
		X"06",X"06",X"06",X"06",X"06",X"86",X"C6",X"E6",X"A6",X"46",X"86",X"06",X"06",X"06",X"06",X"06",
		X"F6",X"76",X"B6",X"D6",X"E6",X"F6",X"E6",X"D6",X"E6",X"D6",X"B6",X"66",X"C6",X"86",X"06",X"06",
		X"06",X"06",X"76",X"36",X"D6",X"E6",X"F6",X"F6",X"EC",X"EC",X"88",X"01",X"07",X"07",X"06",X"06",
		X"F8",X"7C",X"8C",X"EC",X"EC",X"EC",X"EC",X"EC",X"EC",X"0C",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"0C",X"EC",X"EC",X"EC",X"EC",X"B7",X"77",X"E1",X"C0",X"80",X"00",X"00",X"00",
		X"06",X"06",X"86",X"C6",X"E6",X"F6",X"E6",X"D6",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"B6",X"76",X"F6",X"E6",X"C6",X"86",X"06",X"06",X"86",X"C6",X"E6",X"F6",X"F6",X"F6",X"E6",X"D6",
		X"2E",X"16",X"06",X"06",X"06",X"06",X"06",X"06",X"E0",X"F0",X"F8",X"FC",X"FE",X"7E",X"BE",X"5E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"FE",X"FF",X"7F",X"3F",X"1F",X"0E",X"04",X"00",
		X"FF",X"7F",X"BF",X"DF",X"EF",X"F7",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6F",X"6F",X"EF",X"EF",X"9F",X"7F",X"FF",X"FF",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",
		X"7F",X"9F",X"EF",X"EF",X"6F",X"6F",X"6F",X"6F",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FF",
		X"1B",X"1A",X"19",X"0F",X"07",X"03",X"01",X"00",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"19",X"1A",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"19",X"1B",
		X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"19",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"19",X"1B",
		X"1A",X"1A",X"1A",X"1A",X"19",X"1B",X"19",X"1A",X"1B",X"1B",X"1B",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"1B",X"1B",X"1B",X"1A",X"19",X"1B",X"19",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1B",
		X"1A",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"81",X"80",X"81",X"83",X"87",X"8F",X"9F",X"BF",
		X"FD",X"FE",X"7F",X"BF",X"9F",X"8F",X"87",X"83",X"81",X"80",X"F8",X"BC",X"5E",X"EF",X"F7",X"FB",
		X"FD",X"FE",X"7F",X"BF",X"9F",X"8F",X"87",X"83",X"FE",X"F0",X"88",X"7C",X"9E",X"6F",X"F7",X"FB",
		X"80",X"80",X"87",X"B8",X"C7",X"3F",X"FF",X"FF",X"87",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"00",X"8F",X"F1",X"FE",X"FF",X"FF",X"3F",X"80",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"BF",X"9F",X"8F",X"87",X"83",X"81",X"80",X"9F",X"BF",X"7F",X"FF",X"FE",X"FD",X"FE",X"FF",
		X"FF",X"80",X"80",X"80",X"81",X"83",X"87",X"8F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",
		X"00",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"82",X"81",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"7F",X"BF",X"DF",X"AF",X"97",X"8B",X"85",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"83",X"83",X"C1",X"C1",X"81",X"85",X"83",
		X"E0",X"F0",X"78",X"B8",X"90",X"80",X"80",X"C0",X"80",X"C0",X"40",X"00",X"00",X"00",X"83",X"C0",
		X"C0",X"C0",X"40",X"80",X"C0",X"C0",X"80",X"80",X"3F",X"3F",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"1C",X"E0",X"00",X"C0",X"80",X"80",X"C0",X"C0",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"03",
		X"C0",X"00",X"E0",X"FC",X"3F",X"C7",X"C0",X"80",X"60",X"20",X"00",X"00",X"E0",X"E0",X"C0",X"80",
		X"B8",X"DC",X"CE",X"C4",X"C0",X"80",X"C0",X"C0",X"8E",X"9E",X"BC",X"78",X"F0",X"E0",X"E0",X"70",
		X"C0",X"00",X"40",X"E0",X"C0",X"80",X"C0",X"C6",X"00",X"80",X"00",X"00",X"80",X"C0",X"00",X"E1",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"BC",X"78",X"00",X"80",X"C0",X"C0",X"80",X"80",
		X"00",X"C0",X"C0",X"81",X"C3",X"C7",X"CF",X"DE",X"00",X"00",X"00",X"01",X"02",X"04",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"30",X"78",X"3C",X"1E",X"0F",X"07",X"03",X"01",X"3F",X"3F",X"1C",X"19",X"02",X"04",X"08",X"10",
		X"0C",X"18",X"31",X"63",X"C7",X"87",X"0F",X"1F",X"CF",X"CF",X"9F",X"3F",X"3C",X"19",X"13",X"06",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C1",X"C3",X"C7",X"0F",X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",
		X"03",X"3C",X"3F",X"1F",X"0F",X"0F",X"77",X"87",X"03",X"00",X"00",X"00",X"80",X"F0",X"FE",X"1F",
		X"38",X"70",X"F0",X"00",X"07",X"3F",X"3F",X"1F",X"1F",X"3F",X"7E",X"79",X"33",X"27",X"0E",X"1C",
		X"7E",X"3F",X"1F",X"0F",X"07",X"07",X"07",X"0F",X"FC",X"00",X"00",X"00",X"00",X"20",X"78",X"7C",
		X"00",X"80",X"00",X"01",X"00",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"20",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"01",X"20",X"01",X"00",X"08",X"00",X"00",X"80",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"F7",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"BE",X"F8",X"D0",X"60",X"C0",X"80",X"80",X"FE",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DB",X"FE",X"1F",X"01",X"00",X"00",X"00",X"00",X"EF",X"BB",X"EF",X"FB",X"1F",X"01",X"00",X"00",
		X"EF",X"FE",X"FF",X"77",X"FD",X"FF",X"1F",X"01",X"EF",X"FE",X"07",X"01",X"00",X"00",X"00",X"00",
		X"EF",X"FE",X"FF",X"B5",X"FF",X"0E",X"03",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E8",X"70",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"FD",X"7F",X"FF",X"DD",X"FF",X"EE",X"BC",X"FC",
		X"E0",X"60",X"C0",X"C0",X"40",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"20",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"01",X"20",X"01",X"00",X"08",X"00",X"00",X"80",X"00",
		X"00",X"80",X"00",X"01",X"00",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"20",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"08",X"00",X"00",X"01",X"20",X"01",X"00",X"08",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"F0",X"B0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"FF",X"DF",X"FE",X"FE",X"FC",X"EC",X"F8",X"F8",
		X"FF",X"FE",X"BC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"FD",X"3F",X"0F",X"03",X"00",X"00",X"00",
		X"FF",X"DF",X"FD",X"F7",X"FF",X"3F",X"0F",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"F8",X"D8",X"F8",X"F8",X"F8",X"F8",X"B8",X"F8",
		X"C0",X"40",X"C0",X"C0",X"80",X"80",X"80",X"80",X"F0",X"D0",X"F0",X"F0",X"E0",X"E0",X"A0",X"E0",
		X"FC",X"BC",X"FC",X"FC",X"F8",X"E8",X"F8",X"F8",X"FF",X"DF",X"FF",X"F7",X"FE",X"FE",X"BE",X"FE",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"EF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"DF",X"FD",X"F7",X"FF",X"FF",X"0F",X"00",
		X"FF",X"EF",X"FB",X"FF",X"00",X"00",X"00",X"00",X"F8",X"18",X"08",X"00",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"F8",X"F0",X"F0",X"F9",X"F1",X"F4",X"F4",X"F0",
		X"F0",X"F4",X"FA",X"FC",X"FE",X"FE",X"FE",X"FE",X"00",X"40",X"44",X"04",X"80",X"C0",X"E0",X"F0",
		X"00",X"10",X"10",X"00",X"00",X"02",X"02",X"00",X"04",X"82",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",
		X"02",X"F9",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"00",X"30",X"00",X"F3",X"FF",X"FF",X"FF",
		X"00",X"00",X"0C",X"60",X"00",X"E0",X"FC",X"FE",X"00",X"00",X"0C",X"00",X"00",X"60",X"00",X"00",
		X"00",X"20",X"20",X"00",X"00",X"04",X"04",X"00",X"C1",X"F7",X"87",X"3F",X"F0",X"C0",X"80",X"80",
		X"67",X"4F",X"30",X"C0",X"80",X"00",X"00",X"00",X"DE",X"CE",X"96",X"39",X"E7",X"1F",X"FF",X"DF",
		X"E3",X"7B",X"39",X"1C",X"06",X"03",X"01",X"00",X"0D",X"0E",X"06",X"03",X"03",X"01",X"01",X"01",
		X"F3",X"79",X"79",X"3B",X"39",X"3E",X"1E",X"0F",X"9F",X"6F",X"C7",X"4E",X"EF",X"47",X"8F",X"8F",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F0",X"FA",X"FA",X"F8",X"FC",X"FC",X"FC",X"FC",
		X"C0",X"E2",X"E2",X"E0",X"E4",X"F4",X"F0",X"F0",X"00",X"02",X"42",X"C0",X"80",X"88",X"C8",X"C0",
		X"87",X"CF",X"E7",X"F6",X"FE",X"F8",X"35",X"F5",X"01",X"07",X"0F",X"0F",X"0E",X"0E",X"0E",X"07",
		X"7B",X"F6",X"E5",X"D5",X"D1",X"52",X"69",X"79",X"31",X"39",X"38",X"18",X"1C",X"3C",X"79",X"73",
		X"E6",X"EC",X"DD",X"C8",X"E9",X"CD",X"C6",X"E0",X"FB",X"FB",X"1F",X"1C",X"8F",X"E7",X"67",X"33",
		X"CF",X"FC",X"3F",X"17",X"81",X"F0",X"1C",X"C7",X"FF",X"CF",X"FB",X"FB",X"FF",X"3F",X"8F",X"C3",
		X"FF",X"FE",X"3E",X"DC",X"DC",X"3C",X"B8",X"B8",X"CF",X"E7",X"E6",X"72",X"3B",X"3B",X"19",X"3D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"7F",X"FF",X"FD",X"FD",X"3B",X"03",X"0E",X"00",X"00",X"0F",X"3F",X"3E",X"7C",X"7E",X"7F",X"7F",
		X"E4",X"EE",X"C4",X"F0",X"F0",X"C0",X"F0",X"00",X"00",X"80",X"C0",X"E0",X"60",X"70",X"F0",X"C0",
		X"FF",X"FF",X"7F",X"7E",X"18",X"03",X"03",X"00",X"00",X"00",X"07",X"07",X"1F",X"7F",X"7F",X"FF",
		X"E4",X"EE",X"C4",X"70",X"F0",X"E0",X"F0",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"C0",
		X"BD",X"BF",X"9F",X"18",X"00",X"00",X"20",X"67",X"FC",X"FC",X"F8",X"30",X"00",X"00",X"B8",X"48",
		X"E7",X"CF",X"8F",X"2F",X"7F",X"FD",X"9F",X"3C",X"B4",X"F2",X"F9",X"F3",X"E7",X"E7",X"E3",X"63",
		X"6F",X"FB",X"FB",X"C8",X"00",X"40",X"60",X"C1",X"FF",X"6F",X"0C",X"40",X"E0",X"4D",X"0C",X"CE",
		X"FF",X"FF",X"FB",X"FB",X"F9",X"FE",X"C7",X"CF",X"EF",X"EF",X"E7",X"E6",X"F0",X"78",X"78",X"B9",
		X"19",X"DD",X"01",X"19",X"FD",X"F2",X"E6",X"FE",X"FC",X"DC",X"8D",X"9D",X"F9",X"F0",X"C3",X"07",
		X"FE",X"FC",X"30",X"00",X"01",X"86",X"CE",X"FC",X"0F",X"5F",X"DE",X"CF",X"EF",X"E7",X"77",X"7B",
		X"7B",X"F9",X"FE",X"E7",X"FC",X"FF",X"73",X"77",X"F7",X"F7",X"73",X"73",X"F8",X"3C",X"FC",X"FC",
		X"B7",X"FD",X"FD",X"64",X"00",X"20",X"30",X"E0",X"FF",X"B7",X"86",X"20",X"70",X"26",X"06",X"E7",
		X"09",X"4E",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"7D",X"FC",X"EE",X"EF",X"6F",X"07",X"DE",
		X"FF",X"7F",X"7F",X"BF",X"FF",X"FF",X"66",X"00",X"FE",X"DE",X"DF",X"8F",X"8F",X"07",X"17",X"1A",
		X"C7",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FC",X"3F",X"F3",X"F7",X"FF",X"FF",X"F7",X"F3",X"F8",
		X"3E",X"FE",X"F7",X"F7",X"B7",X"83",X"EF",X"FF",X"FC",X"7F",X"7F",X"BF",X"FF",X"FF",X"66",X"00",
		X"DB",X"D9",X"C3",X"FE",X"FE",X"BF",X"BF",X"ED",X"78",X"9D",X"F9",X"F1",X"C3",X"E7",X"FE",X"BC",
		X"EC",X"E1",X"FB",X"61",X"00",X"07",X"07",X"FF",X"30",X"00",X"A1",X"39",X"78",X"FC",X"FD",X"FF",
		X"00",X"70",X"FC",X"FC",X"FE",X"FF",X"BF",X"BF",X"DF",X"CF",X"73",X"3B",X"FF",X"B6",X"B0",X"84",
		X"9F",X"1F",X"3F",X"7F",X"FE",X"CC",X"00",X"40",X"AE",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"1F",X"1F",X"06",X"00",X"00",X"01",X"1F",X"3F",X"3F",X"3F",X"0E",X"00",X"03",
		X"01",X"01",X"01",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",X"0F",X"0F",
		X"FF",X"FE",X"F9",X"FB",X"77",X"07",X"1D",X"00",X"38",X"CC",X"E8",X"E8",X"F4",X"F4",X"ED",X"EB",
		X"FF",X"FB",X"FB",X"77",X"07",X"3D",X"30",X"3C",X"83",X"80",X"00",X"20",X"70",X"20",X"80",X"80",
		X"00",X"C8",X"C3",X"FE",X"FE",X"BF",X"BF",X"ED",X"1E",X"7C",X"7E",X"00",X"00",X"00",X"00",X"00",
		X"11",X"33",X"33",X"07",X"07",X"03",X"23",X"37",X"30",X"98",X"EC",X"F6",X"76",X"7A",X"FB",X"F7",
		X"7C",X"CB",X"C3",X"D5",X"CB",X"A5",X"D3",X"7D",X"40",X"7F",X"AD",X"6B",X"E6",X"6F",X"7B",X"72",
		X"68",X"9F",X"A9",X"AF",X"BF",X"D9",X"DF",X"EF",X"0C",X"FB",X"79",X"F3",X"F5",X"73",X"FB",X"F7",
		X"00",X"FF",X"BD",X"9B",X"BD",X"DD",X"B9",X"BB",X"50",X"5F",X"BC",X"BA",X"B5",X"B9",X"D7",X"BF",
		X"14",X"CF",X"DF",X"9F",X"2E",X"9E",X"E7",X"F3",X"04",X"FA",X"CD",X"DD",X"9D",X"3F",X"FD",X"FA",
		X"7C",X"CE",X"85",X"DB",X"C7",X"9B",X"C5",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"02",X"00",
		X"00",X"81",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"F8",
		X"00",X"00",X"00",X"CD",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"F0",X"F9",X"FF",X"FF",X"FF",X"FF",
		X"18",X"10",X"30",X"20",X"60",X"40",X"C0",X"80",X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"0C",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"01",X"01",X"03",X"07",X"07",X"03",
		X"00",X"01",X"07",X"1C",X"30",X"20",X"60",X"C0",X"00",X"00",X"00",X"01",X"01",X"07",X"3C",X"E0",
		X"01",X"03",X"1E",X"70",X"C0",X"00",X"00",X"00",X"E9",X"EC",X"80",X"04",X"D0",X"80",X"00",X"00",
		X"30",X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"77",X"12",X"C0",X"80",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"80",X"40",X"10",X"02",X"40",X"08",X"00",X"00",X"00",X"00",X"80",X"40",X"10",X"44",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"CC",X"80",X"FF",X"FF",X"FF",X"FE",X"CC",X"00",X"00",X"00",
		X"F0",X"B8",X"FC",X"FF",X"CF",X"2F",X"D4",X"EF",X"BC",X"BC",X"B8",X"78",X"D0",X"F0",X"70",X"F0",
		X"B8",X"78",X"FC",X"7C",X"BE",X"FC",X"B8",X"FC",X"B0",X"D8",X"98",X"30",X"D8",X"98",X"50",X"F0",
		X"70",X"F0",X"B0",X"20",X"E0",X"B0",X"D8",X"FC",X"DF",X"EB",X"BF",X"F7",X"E7",X"9C",X"1C",X"B8",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"FF",X"BD",X"D7",X"F9",X"FF",X"FF",X"21",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"1E",X"FF",X"F7",X"BF",X"BB",X"FF",X"F1",X"E0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0E",X"BE",X"E7",X"C9",X"EE",X"FF",X"FF",X"47",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"07",X"1F",X"7E",X"FB",X"FD",X"5E",X"EB",X"FF",X"FF",X"FF",X"03",X"00",X"00",
		X"F9",X"FA",X"F7",X"F3",X"EE",X"5F",X"FD",X"DF",X"19",X"3F",X"1E",X"3C",X"3D",X"3F",X"3F",X"7D",
		X"07",X"06",X"05",X"07",X"0F",X"0E",X"1F",X"1F",X"06",X"07",X"0C",X"0E",X"0F",X"0E",X"07",X"07",
		X"0F",X"0D",X"06",X"05",X"0F",X"0E",X"0F",X"07",X"FF",X"3D",X"C6",X"F3",X"FB",X"FC",X"79",X"1E",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"E0",X"E0",X"40",X"40",X"80",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"C0",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0D",X"1B",X"36",X"6C",X"D8",X"B0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0D",X"1B",X"36",X"6C",X"D8",X"B0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",X"31",X"63",X"C6",X"8C",X"18",X"30",
		X"0C",X"18",X"31",X"63",X"C6",X"8C",X"98",X"70",X"38",X"60",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"38",X"6F",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"00",X"01",X"03",X"06",X"03",X"0C",X"30",X"C0",X"80",X"80",X"80",X"80",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"02",X"01",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"48",X"38",X"08",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"FF",X"00",X"00",X"00",X"FF",
		X"10",X"10",X"08",X"04",X"04",X"02",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"C0",X"A0",X"98",X"84",X"83",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",
		X"8C",X"8A",X"89",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"3F",X"20",X"10",X"08",X"0F",
		X"08",X"08",X"04",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"88",X"88",X"88",X"C8",X"28",X"18",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0C",X"03",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"7F",X"00",X"00",X"00",X"00",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"06",X"40",X"20",X"20",X"1F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"80",X"40",X"40",X"3F",X"88",X"88",X"88",X"88",X"88",X"88",X"68",X"18",
		X"08",X"08",X"08",X"08",X"08",X"06",X"01",X"00",X"00",X"00",X"00",X"E0",X"10",X"10",X"08",X"04",
		X"00",X"00",X"80",X"40",X"30",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"01",X"00",X"00",X"00",X"1F",X"20",X"40",X"80",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"FF",X"11",X"10",X"10",X"10",X"10",X"20",X"40",X"80",
		X"81",X"82",X"84",X"88",X"90",X"A0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"03",X"1C",X"E0",
		X"20",X"20",X"40",X"40",X"40",X"80",X"80",X"80",X"00",X"00",X"01",X"0E",X"70",X"80",X"00",X"00",
		X"07",X"38",X"C0",X"00",X"00",X"01",X"01",X"01",X"E1",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"04",X"08",X"08",X"08",X"10",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"80",X"60",X"18",X"06",
		X"3F",X"00",X"00",X"00",X"3F",X"60",X"18",X"06",X"81",X"60",X"18",X"06",X"01",X"00",X"00",X"E0",
		X"10",X"08",X"08",X"04",X"04",X"82",X"82",X"81",X"11",X"91",X"91",X"51",X"51",X"31",X"20",X"00",
		X"00",X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"C0",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"21",X"26",X"38",X"20",X"01",X"06",X"18",X"60",X"81",X"06",X"18",X"60",
		X"11",X"22",X"22",X"44",X"44",X"88",X"88",X"10",X"10",X"20",X"20",X"40",X"40",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"10",X"10",X"FE",X"01",X"01",X"01",X"FE",X"00",X"00",X"00",
		X"0E",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"A5",X"5A",X"A4",X"59",X"26",X"09",X"16",X"08",
		X"1B",X"24",X"D8",X"21",X"C6",X"19",X"26",X"D8",X"03",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"20",X"C0",X"03",X"1C",X"63",X"8C",X"70",X"00",X"14",X"14",X"28",X"28",X"48",X"51",X"52",X"22",
		X"29",X"51",X"52",X"A5",X"A5",X"4A",X"94",X"94",X"05",X"05",X"02",X"00",X"00",X"00",X"00",X"00",
		X"21",X"52",X"55",X"AA",X"4A",X"15",X"0A",X"05",X"04",X"19",X"66",X"98",X"60",X"80",X"03",X"0C",
		X"C0",X"00",X"01",X"06",X"18",X"E3",X"0C",X"30",X"31",X"C6",X"18",X"E0",X"00",X"03",X"1C",X"E0",
		X"C0",X"00",X"01",X"0E",X"70",X"80",X"00",X"00",X"04",X"08",X"08",X"08",X"10",X"10",X"11",X"21",
		X"24",X"28",X"48",X"50",X"90",X"A0",X"21",X"21",X"21",X"22",X"42",X"44",X"45",X"89",X"8A",X"8A",
		X"42",X"44",X"85",X"8A",X"0A",X"14",X"14",X"28",X"18",X"60",X"87",X"18",X"60",X"80",X"00",X"00",
		X"30",X"C0",X"00",X"00",X"00",X"03",X"1C",X"E0",X"20",X"20",X"40",X"40",X"41",X"81",X"82",X"82",
		X"04",X"04",X"04",X"09",X"09",X"12",X"12",X"24",X"50",X"A1",X"42",X"85",X"0A",X"34",X"48",X"B0",
		X"D0",X"20",X"C1",X"02",X"0C",X"11",X"66",X"88",X"41",X"86",X"09",X"32",X"4C",X"90",X"60",X"83",
		X"30",X"40",X"81",X"06",X"08",X"33",X"CC",X"30",X"24",X"28",X"48",X"50",X"A1",X"A1",X"42",X"44",
		X"24",X"48",X"50",X"90",X"21",X"42",X"45",X"85",X"85",X"8A",X"12",X"14",X"28",X"48",X"51",X"A2",
		X"0A",X"14",X"28",X"50",X"A1",X"A2",X"45",X"8A",X"23",X"C4",X"18",X"20",X"C0",X"00",X"03",X"0C",
		X"00",X"01",X"06",X"18",X"21",X"C6",X"18",X"60",X"11",X"66",X"88",X"30",X"C0",X"00",X"00",X"07",
		X"00",X"00",X"00",X"03",X"0C",X"30",X"C1",X"0E",X"48",X"88",X"90",X"90",X"20",X"20",X"40",X"41",
		X"12",X"24",X"24",X"48",X"48",X"90",X"A0",X"20",X"81",X"82",X"82",X"04",X"09",X"0A",X"12",X"14",
		X"41",X"41",X"82",X"84",X"04",X"09",X"12",X"12",X"63",X"8C",X"30",X"40",X"80",X"00",X"00",X"01",
		X"01",X"01",X"01",X"01",X"06",X"18",X"60",X"80",X"06",X"38",X"C0",X"03",X"1C",X"60",X"80",X"00",
		X"07",X"39",X"C1",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"02",X"02",X"02",X"04",X"04",
		X"0F",X"10",X"10",X"20",X"20",X"40",X"40",X"80",X"08",X"09",X"11",X"12",X"12",X"22",X"24",X"44",
		X"81",X"01",X"02",X"02",X"04",X"05",X"09",X"12",X"28",X"50",X"A0",X"40",X"81",X"02",X"04",X"19",
		X"09",X"32",X"44",X"98",X"20",X"40",X"80",X"01",X"26",X"48",X"90",X"60",X"81",X"02",X"04",X"18",
		X"06",X"08",X"31",X"42",X"8C",X"10",X"60",X"80",X"04",X"09",X"11",X"12",X"24",X"44",X"48",X"90",
		X"81",X"02",X"04",X"09",X"12",X"12",X"24",X"48",X"10",X"21",X"41",X"82",X"84",X"09",X"0A",X"14",
		X"90",X"20",X"41",X"82",X"82",X"05",X"0A",X"14",X"00",X"01",X"02",X"0C",X"10",X"61",X"86",X"08",
		X"43",X"85",X"19",X"21",X"C1",X"01",X"01",X"01",X"30",X"40",X"80",X"00",X"00",X"03",X"0C",X"10",
		X"02",X"04",X"18",X"60",X"83",X"0D",X"31",X"C1",X"F0",X"11",X"22",X"24",X"44",X"48",X"88",X"90",
		X"FF",X"01",X"02",X"04",X"04",X"08",X"11",X"12",X"20",X"20",X"40",X"40",X"81",X"01",X"02",X"04",
		X"22",X"44",X"48",X"88",X"10",X"20",X"20",X"40",X"22",X"44",X"88",X"10",X"20",X"40",X"81",X"02",
		X"02",X"04",X"08",X"10",X"23",X"C5",X"09",X"11",X"04",X"08",X"11",X"62",X"8C",X"10",X"20",X"C0",
		X"61",X"81",X"01",X"01",X"02",X"04",X"18",X"20",X"0F",X"10",X"20",X"40",X"40",X"81",X"01",X"02",
		X"F0",X"11",X"22",X"44",X"88",X"10",X"20",X"20",X"04",X"08",X"11",X"12",X"24",X"48",X"88",X"90",
		X"40",X"81",X"02",X"04",X"08",X"11",X"22",X"44",X"45",X"4A",X"8A",X"14",X"29",X"51",X"A2",X"A5",
		X"14",X"28",X"51",X"A2",X"45",X"4A",X"B4",X"48",X"4A",X"95",X"2A",X"55",X"AA",X"54",X"A9",X"52",
		X"B1",X"46",X"89",X"16",X"28",X"D0",X"23",X"C4",X"28",X"50",X"A0",X"A1",X"42",X"85",X"0A",X"14",
		X"28",X"50",X"A0",X"41",X"82",X"05",X"0A",X"14",X"28",X"50",X"A0",X"41",X"82",X"0D",X"12",X"2C",
		X"20",X"40",X"81",X"02",X"04",X"09",X"12",X"24",X"48",X"90",X"20",X"41",X"82",X"04",X"09",X"12",
		X"FF",X"02",X"04",X"08",X"08",X"11",X"22",X"44",X"0F",X"11",X"21",X"41",X"82",X"04",X"08",X"10",
		X"88",X"10",X"20",X"41",X"82",X"04",X"08",X"11",X"21",X"43",X"85",X"19",X"21",X"41",X"81",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"E1",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"01",X"03",X"07",X"0F",X"FF",X"FE",X"C0",X"E0",X"F0",X"F8",X"04",X"08",X"10",X"20",
		X"00",X"00",X"F0",X"08",X"04",X"02",X"01",X"00",X"70",X"F8",X"FC",X"E6",X"C3",X"81",X"00",X"00",
		X"70",X"F8",X"FC",X"FE",X"FF",X"F9",X"F8",X"F8",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"F9",X"F9",X"79",X"39",X"19",X"01",X"01",X"01",
		X"09",X"09",X"09",X"09",X"09",X"89",X"C9",X"E9",X"69",X"C9",X"89",X"09",X"09",X"09",X"09",X"09",
		X"F9",X"F9",X"79",X"39",X"19",X"09",X"19",X"39",X"19",X"39",X"79",X"E9",X"C9",X"89",X"09",X"09",
		X"09",X"09",X"79",X"F9",X"39",X"19",X"09",X"09",X"1C",X"1C",X"79",X"86",X"08",X"08",X"09",X"09",
		X"F8",X"FC",X"7C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"FC",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"00",X"00",X"00",X"FC",X"1C",X"1C",X"1C",X"1C",X"78",X"F8",X"E6",X"C1",X"80",X"00",X"00",X"00",
		X"09",X"89",X"49",X"29",X"19",X"09",X"19",X"39",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"79",X"F9",X"F9",X"E9",X"C9",X"89",X"09",X"09",X"49",X"29",X"19",X"09",X"09",X"09",X"19",X"39",
		X"31",X"19",X"09",X"09",X"09",X"09",X"09",X"89",X"10",X"08",X"04",X"02",X"01",X"81",X"C1",X"61",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"20",X"01",X"00",X"80",X"40",X"20",X"11",X"0A",X"04",
		X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"9F",X"1F",X"1F",X"7F",X"FF",X"FF",X"FF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"7F",X"1F",X"1F",X"9F",X"9F",X"9F",X"9F",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FF",
		X"27",X"27",X"26",X"10",X"08",X"04",X"02",X"01",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"26",X"24",
		X"27",X"27",X"27",X"27",X"27",X"27",X"26",X"24",X"27",X"27",X"27",X"27",X"27",X"27",X"26",X"24",
		X"27",X"27",X"27",X"27",X"26",X"24",X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"27",X"27",X"26",X"24",X"26",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",X"27",
		X"03",X"04",X"08",X"10",X"20",X"20",X"20",X"26",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"01",X"02",X"04",X"08",X"10",X"20",X"82",X"81",X"82",X"84",X"88",X"90",X"A0",X"C0",
		X"03",X"01",X"80",X"C0",X"A0",X"90",X"88",X"84",X"82",X"81",X"F8",X"FC",X"BE",X"1F",X"0F",X"07",
		X"03",X"01",X"80",X"C0",X"A0",X"90",X"88",X"84",X"01",X"0E",X"78",X"FC",X"FE",X"9F",X"0F",X"07",
		X"80",X"80",X"87",X"BF",X"F8",X"C0",X"00",X"00",X"B8",X"87",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"FF",X"7F",X"0F",X"01",X"00",X"00",X"C0",X"80",X"80",X"80",X"FF",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"A0",X"90",X"88",X"84",X"82",X"81",X"A0",X"C0",X"80",X"00",X"01",X"03",X"01",X"00",
		X"FF",X"80",X"80",X"81",X"82",X"84",X"88",X"90",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"83",X"81",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"01",X"80",X"C0",X"E0",X"B0",X"98",X"8C",X"86",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"02",
		X"C3",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"7F",X"3F",X"3F",X"7F",X"7F",X"67",
		X"E0",X"F1",X"FA",X"7C",X"7A",X"7E",X"7E",X"3C",X"7E",X"3E",X"BC",X"7C",X"39",X"12",X"8F",X"C0",
		X"FD",X"FD",X"FD",X"7D",X"3C",X"3C",X"7C",X"7C",X"FF",X"3F",X"3F",X"31",X"39",X"3D",X"BD",X"FD",
		X"1F",X"FC",X"F2",X"3E",X"7E",X"7C",X"3F",X"38",X"7E",X"3C",X"F0",X"1C",X"03",X"00",X"00",X"03",
		X"3C",X"FF",X"E0",X"FC",X"FF",X"3F",X"37",X"78",X"9E",X"5C",X"3D",X"FF",X"18",X"1E",X"3E",X"7F",
		X"78",X"3C",X"3F",X"3E",X"3C",X"7E",X"3C",X"3C",X"7F",X"7E",X"7C",X"F8",X"F0",X"E0",X"E0",X"F0",
		X"FD",X"7E",X"BE",X"1E",X"3C",X"78",X"34",X"3C",X"FF",X"70",X"FE",X"FE",X"7E",X"3C",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"7C",X"F8",X"FF",X"70",X"3C",X"3E",X"7E",X"7E",
		X"FE",X"3E",X"3D",X"7B",X"3F",X"3F",X"3F",X"3E",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"F0",X"F0",X"60",X"30",X"18",X"0C",X"06",
		X"70",X"F8",X"7C",X"3E",X"1F",X"0F",X"07",X"03",X"80",X"00",X"01",X"03",X"06",X"0C",X"18",X"30",
		X"1C",X"39",X"72",X"E4",X"C8",X"90",X"20",X"40",X"D0",X"E0",X"C0",X"80",X"01",X"03",X"07",X"0E",
		X"C0",X"C0",X"C0",X"C0",X"C1",X"C2",X"C4",X"C8",X"80",X"00",X"00",X"03",X"1C",X"E0",X"00",X"00",
		X"1F",X"03",X"00",X"00",X"80",X"70",X"78",X"F0",X"00",X"FF",X"00",X"00",X"80",X"F0",X"FE",X"FF",
		X"78",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"40",X"80",X"01",X"03",X"07",X"0F",X"1E",X"3C",
		X"01",X"80",X"40",X"20",X"10",X"08",X"10",X"20",X"FC",X"80",X"40",X"20",X"10",X"08",X"04",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"70",X"80",X"F4",X"D7",X"00",X"00",X"81",X"91",X"80",X"07",X"BB",X"BB",
		X"00",X"00",X"0E",X"EE",X"00",X"0E",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"F5",
		X"D7",X"C4",X"F0",X"07",X"03",X"01",X"30",X"00",X"BB",X"BB",X"87",X"78",X"79",X"69",X"F0",X"F0",
		X"FF",X"FE",X"1E",X"F0",X"FE",X"1E",X"F0",X"E0",X"F5",X"FB",X"E0",X"E0",X"C0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"10",X"10",X"77",X"45",X"55",X"00",X"00",X"07",X"77",X"00",X"8F",X"D5",X"DD",
		X"00",X"00",X"0C",X"CC",X"00",X"0C",X"FD",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"EA",
		X"55",X"45",X"77",X"01",X"01",X"00",X"10",X"00",X"DD",X"55",X"8F",X"F0",X"F7",X"87",X"F0",X"70",
		X"FE",X"FD",X"3C",X"F0",X"FC",X"3C",X"F0",X"E0",X"EA",X"E6",X"C0",X"C0",X"C0",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"77",X"00",X"67",X"FA",X"FF",
		X"00",X"00",X"08",X"88",X"00",X"00",X"FB",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"BA",X"E7",X"70",X"77",X"07",X"52",X"30",
		X"F5",X"FB",X"E0",X"E0",X"E8",X"48",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"32",X"00",X"02",X"77",X"76",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E6",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"77",X"34",X"10",X"32",X"21",X"10",X"00",
		X"EA",X"E6",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"12",X"34",X"70",X"83",X"83",
		X"48",X"E0",X"E0",X"E0",X"E0",X"87",X"1E",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C5",X"6B",X"00",X"44",X"62",X"20",X"13",X"10",
		X"5A",X"1E",X"07",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"03",X"44",X"44",X"03",X"07",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"0E",X"0F",X"1E",X"1E",X"1E",X"02",X"80",X"C8",X"00",X"08",X"00",X"80",X"80",X"00",X"20",X"20",
		X"44",X"26",X"33",X"33",X"31",X"10",X"10",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"7F",X"F7",X"73",
		X"C8",X"80",X"22",X"EF",X"EF",X"EF",X"FF",X"EE",X"20",X"20",X"00",X"08",X"08",X"00",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"33",X"FE",X"FD",
		X"00",X"00",X"01",X"01",X"01",X"99",X"D5",X"FB",X"00",X"00",X"08",X"0C",X"0E",X"FF",X"0E",X"0E",
		X"FF",X"7F",X"70",X"70",X"30",X"21",X"10",X"00",X"FD",X"FE",X"D3",X"F0",X"F0",X"F0",X"F0",X"70",
		X"FB",X"F7",X"FD",X"E1",X"E1",X"E1",X"F0",X"F0",X"0E",X"0E",X"FF",X"0E",X"0C",X"08",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"32",X"32",X"00",X"00",X"33",X"CC",X"FF",X"CC",X"88",X"99",
		X"00",X"00",X"CC",X"33",X"DF",X"23",X"11",X"99",X"00",X"00",X"00",X"00",X"88",X"88",X"44",X"44",
		X"32",X"32",X"11",X"11",X"00",X"00",X"00",X"00",X"99",X"88",X"4C",X"BF",X"FC",X"33",X"00",X"00",
		X"99",X"11",X"33",X"FF",X"F3",X"CC",X"00",X"00",X"44",X"44",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"31",X"00",X"00",X"00",X"30",X"C0",X"F4",X"C8",X"91",
		X"00",X"00",X"00",X"C3",X"30",X"D2",X"21",X"98",X"00",X"00",X"00",X"00",X"08",X"80",X"84",X"40",
		X"31",X"31",X"10",X"10",X"00",X"00",X"00",X"00",X"91",X"84",X"C2",X"F0",X"F0",X"30",X"00",X"00",
		X"98",X"10",X"31",X"F0",X"F0",X"C0",X"00",X"00",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"23",X"03",X"00",X"00",X"00",X"00",X"77",X"8F",X"7F",X"9D",
		X"00",X"00",X"00",X"00",X"EE",X"0E",X"CD",X"8A",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"13",X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"08",X"1D",X"0F",X"07",X"00",X"00",X"00",X"00",
		X"EF",X"CF",X"0F",X"0E",X"00",X"00",X"00",X"00",X"0C",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"33",X"00",X"00",X"00",X"00",X"00",X"BF",X"FF",X"B4",
		X"00",X"00",X"00",X"00",X"00",X"6F",X"FF",X"F2",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"B3",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"FE",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"52",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"19",X"3A",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"C3",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",
		X"03",X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"B0",X"00",X"00",X"00",X"00",X"00",X"CC",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"74",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"99",X"77",X"08",X"07",X"00",X"00",X"00",X"00",
		X"88",X"EE",X"10",X"0E",X"00",X"00",X"00",X"00",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"32",X"32",X"00",X"00",X"33",X"FF",X"FF",X"F4",X"88",X"99",
		X"00",X"00",X"CC",X"FF",X"FF",X"F3",X"13",X"99",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",
		X"32",X"31",X"11",X"10",X"00",X"00",X"00",X"00",X"99",X"4C",X"BF",X"FC",X"7B",X"30",X"00",X"00",
		X"99",X"33",X"FD",X"F3",X"FD",X"C0",X"00",X"00",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"30",X"02",X"77",X"10",X"10",X"00",X"77",X"F7",X"F6",X"98",X"FE",X"70",X"F7",
		X"00",X"EE",X"EE",X"6E",X"08",X"4D",X"C3",X"DC",X"00",X"00",X"88",X"88",X"CC",X"08",X"84",X"C8",
		X"10",X"10",X"70",X"03",X"03",X"01",X"00",X"00",X"07",X"F0",X"E1",X"69",X"69",X"78",X"70",X"00",
		X"5C",X"F3",X"62",X"71",X"F9",X"F1",X"E0",X"00",X"FB",X"C4",X"00",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"01",X"00",X"00",X"00",X"77",X"F7",X"F6",X"F6",X"18",X"11",X"00",
		X"00",X"EE",X"EE",X"6E",X"6E",X"08",X"EE",X"FE",X"00",X"00",X"88",X"88",X"00",X"88",X"80",X"EA",
		X"00",X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"F0",X"FF",X"23",X"69",X"69",X"78",X"70",X"00",
		X"FE",X"F8",X"43",X"71",X"F9",X"F1",X"E0",X"00",X"EA",X"C4",X"80",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"77",X"F7",X"F6",X"F6",X"16",X"00",X"33",
		X"00",X"CC",X"89",X"09",X"09",X"3B",X"75",X"FA",X"00",X"00",X"88",X"88",X"00",X"00",X"88",X"80",
		X"00",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"F3",X"00",X"07",X"69",X"69",X"78",X"70",X"00",
		X"FA",X"65",X"43",X"71",X"F9",X"F1",X"E0",X"00",X"80",X"08",X"00",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"77",X"F7",X"F6",X"F6",X"00",X"10",X"F1",
		X"00",X"CC",X"89",X"09",X"09",X"00",X"00",X"C4",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"F1",X"12",X"01",X"69",X"69",X"78",X"70",X"00",
		X"C4",X"C0",X"80",X"71",X"F9",X"F1",X"E0",X"00",X"00",X"00",X"00",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"00",X"00",X"77",X"F7",X"F6",X"F6",X"00",X"44",X"F7",
		X"00",X"EE",X"EE",X"6E",X"6E",X"08",X"88",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"01",X"00",X"00",X"7B",X"37",X"30",X"69",X"69",X"78",X"70",X"00",
		X"88",X"8C",X"06",X"71",X"F9",X"F1",X"E0",X"00",X"00",X"00",X"00",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"00",X"00",X"37",X"00",X"77",X"F7",X"F6",X"F6",X"10",X"10",X"FF",
		X"00",X"EE",X"EE",X"6E",X"6E",X"0B",X"08",X"FF",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"37",X"13",X"01",X"03",X"03",X"01",X"00",X"00",X"11",X"EF",X"E1",X"69",X"69",X"78",X"70",X"00",
		X"88",X"77",X"44",X"71",X"F9",X"F1",X"E0",X"00",X"00",X"00",X"04",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"00",X"10",X"30",X"30",X"01",X"11",X"F6",X"00",X"77",X"F7",X"F6",X"F6",X"18",X"FE",X"F0",
		X"00",X"EE",X"EE",X"6E",X"6E",X"08",X"7F",X"F0",X"00",X"00",X"88",X"88",X"00",X"EE",X"00",X"00",
		X"F3",X"30",X"01",X"03",X"03",X"01",X"00",X"00",X"FE",X"E1",X"67",X"69",X"69",X"78",X"70",X"00",
		X"F7",X"70",X"77",X"71",X"F9",X"F1",X"E0",X"00",X"00",X"00",X"E0",X"CC",X"CC",X"88",X"00",X"00",
		X"00",X"03",X"45",X"66",X"77",X"77",X"77",X"77",X"00",X"0F",X"0F",X"0F",X"07",X"8B",X"CD",X"EE",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"67",X"56",X"34",X"00",X"EF",X"DE",X"BC",X"78",X"F0",X"F0",X"F0",X"00",
		X"88",X"C4",X"E2",X"F1",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"88",X"C4",X"E2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"10",X"00",X"00",X"00",X"00",X"04",X"30",X"32",X"91",X"60",
		X"00",X"00",X"00",X"00",X"00",X"F7",X"23",X"23",X"00",X"00",X"00",X"00",X"EE",X"FF",X"00",X"00",
		X"11",X"01",X"10",X"10",X"00",X"00",X"00",X"00",X"98",X"FE",X"F2",X"F3",X"F1",X"F1",X"70",X"10",
		X"81",X"C1",X"CC",X"88",X"00",X"88",X"88",X"CC",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"70",X"10",X"00",X"00",X"00",X"00",X"24",X"32",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"77",X"C7",X"23",X"23",X"00",X"00",X"00",X"EE",X"CC",X"00",X"00",X"00",
		X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"30",X"FE",X"F3",X"F1",X"F0",X"70",X"70",X"00",
		X"C1",X"E2",X"CC",X"88",X"CC",X"CC",X"E6",X"E6",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"00",X"00",X"00",X"80",X"78",X"77",X"80",
		X"00",X"00",X"00",X"33",X"FF",X"CE",X"23",X"01",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",X"08",
		X"00",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"70",X"98",X"FF",X"F1",X"F0",X"70",X"30",X"00",
		X"C1",X"E2",X"C4",X"88",X"CC",X"E6",X"F3",X"62",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"77",X"00",
		X"00",X"11",X"33",X"77",X"CE",X"CF",X"23",X"01",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"08",
		X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"7F",X"F0",X"70",X"30",X"10",X"00",
		X"E0",X"E2",X"CC",X"CC",X"F7",X"F3",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"11",X"F1",X"E6",X"00",
		X"22",X"33",X"66",X"CC",X"8E",X"47",X"23",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"80",X"FF",X"78",X"70",X"30",X"00",X"00",
		X"E0",X"E2",X"CC",X"FF",X"F3",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"11",X"31",X"E0",X"44",
		X"66",X"66",X"CC",X"CC",X"8E",X"CF",X"23",X"20",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",
		X"00",X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"33",X"54",X"34",X"10",X"00",X"00",
		X"E2",X"E2",X"CC",X"F7",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"CC",X"EE",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"11",X"11",X"33",X"22",X"E0",X"E6",
		X"CC",X"88",X"88",X"08",X"8F",X"CF",X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"34",X"00",X"00",X"00",X"00",X"10",X"60",X"91",X"33",X"34",X"00",X"00",X"00",
		X"E2",X"E2",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"EE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"32",X"75",X"75",X"10",X"03",X"00",X"FF",X"FF",X"F1",X"F0",X"F0",
		X"C0",X"3C",X"03",X"CD",X"CC",X"EE",X"F7",X"F3",X"00",X"80",X"C0",X"68",X"2C",X"24",X"9A",X"9A",
		X"75",X"75",X"32",X"32",X"11",X"00",X"00",X"00",X"F0",X"F0",X"78",X"B4",X"F3",X"FC",X"33",X"00",
		X"F3",X"F1",X"F1",X"F1",X"FD",X"E2",X"CC",X"00",X"9A",X"8A",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"FF",X"66",X"00",X"73",X"00",X"00",X"DD",X"DD",X"33",X"11",X"98",X"7D",
		X"00",X"00",X"00",X"4C",X"6F",X"0F",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"3F",X"E0",X"00",
		X"25",X"30",X"76",X"F7",X"62",X"20",X"10",X"00",X"BD",X"78",X"F1",X"33",X"DD",X"DD",X"30",X"C0",
		X"C0",X"F3",X"0F",X"0F",X"3C",X"C0",X"00",X"00",X"00",X"EE",X"3C",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"33",X"73",X"00",X"11",X"00",X"00",X"DD",X"DD",X"3B",X"00",X"10",X"FD",
		X"00",X"00",X"00",X"4C",X"6E",X"0F",X"10",X"C0",X"00",X"00",X"00",X"00",X"00",X"08",X"E2",X"00",
		X"13",X"21",X"77",X"73",X"21",X"21",X"10",X"00",X"7D",X"F8",X"F0",X"33",X"DD",X"DD",X"38",X"C0",
		X"C0",X"E0",X"0F",X"1E",X"2C",X"C0",X"00",X"00",X"00",X"22",X"6A",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"37",X"BF",X"DF",X"80",X"20",X"3A",
		X"00",X"00",X"08",X"4C",X"6E",X"0F",X"74",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"BA",X"7C",X"70",X"DD",X"BF",X"B7",X"D7",X"70",
		X"C4",X"F7",X"0F",X"1E",X"2C",X"48",X"80",X"00",X"00",X"88",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"76",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"25",X"21",X"01",X"01",X"01",X"01",X"01",
		X"CC",X"C4",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"C0",X"01",
		X"00",X"00",X"46",X"46",X"04",X"08",X"02",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"0F",X"87",X"43",X"21",X"10",X"00",
		X"FF",X"22",X"08",X"00",X"46",X"46",X"04",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"74",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"80",X"03",
		X"00",X"00",X"33",X"33",X"09",X"08",X"03",X"0F",X"00",X"00",X"08",X"08",X"00",X"20",X"08",X"0C",
		X"00",X"44",X"65",X"10",X"00",X"00",X"00",X"00",X"77",X"00",X"0F",X"87",X"43",X"30",X"00",X"00",
		X"FF",X"33",X"08",X"08",X"33",X"33",X"C1",X"22",X"CC",X"88",X"00",X"00",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8B",X"70",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"F7",X"44",
		X"00",X"00",X"BB",X"BB",X"4C",X"7F",X"FC",X"00",X"00",X"00",X"00",X"44",X"EE",X"CC",X"84",X"00",
		X"00",X"77",X"C3",X"30",X"00",X"00",X"00",X"00",X"70",X"FF",X"0F",X"0F",X"C3",X"30",X"00",X"00",
		X"C3",X"FC",X"7F",X"4C",X"BB",X"BB",X"C0",X"30",X"48",X"80",X"CC",X"FF",X"64",X"40",X"80",X"00",
		X"00",X"11",X"33",X"77",X"FF",X"F0",X"F0",X"F0",X"88",X"88",X"88",X"88",X"B8",X"F4",X"71",X"73",
		X"01",X"01",X"01",X"01",X"C1",X"C2",X"F8",X"FC",X"00",X"08",X"8C",X"CE",X"0F",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"0F",X"37",X"13",X"01",X"00",X"73",X"71",X"B4",X"48",X"78",X"78",X"78",X"78",
		X"FC",X"F8",X"E2",X"31",X"F1",X"F1",X"F1",X"F1",X"00",X"00",X"00",X"FF",X"EE",X"CC",X"88",X"00",
		X"00",X"00",X"33",X"22",X"00",X"11",X"32",X"BA",X"00",X"11",X"03",X"00",X"FF",X"F0",X"F2",X"F1",
		X"00",X"08",X"0C",X"07",X"89",X"C4",X"E6",X"F9",X"00",X"00",X"0C",X"84",X"08",X"08",X"0C",X"06",
		X"FA",X"32",X"10",X"11",X"13",X"03",X"00",X"00",X"F1",X"B6",X"96",X"F0",X"F8",X"33",X"10",X"11",
		X"F9",X"F5",X"F1",X"F1",X"E2",X"CC",X"00",X"88",X"26",X"04",X"00",X"00",X"44",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"66",X"44",X"33",X"32",X"32",X"66",X"01",X"03",X"00",X"FF",X"F0",X"F2",X"F1",
		X"00",X"01",X"1E",X"07",X"89",X"C4",X"E6",X"F9",X"00",X"08",X"08",X"00",X"08",X"0A",X"0E",X"04",
		X"32",X"F2",X"D0",X"11",X"00",X"10",X"10",X"00",X"F1",X"B6",X"96",X"F0",X"F8",X"FF",X"80",X"00",
		X"F9",X"F5",X"F1",X"F1",X"E2",X"CC",X"C0",X"66",X"04",X"04",X"04",X"22",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"DD",X"76",X"32",X"44",X"8A",X"03",X"00",X"FF",X"F0",X"F2",X"F1",
		X"00",X"06",X"2C",X"07",X"89",X"C4",X"E6",X"F9",X"00",X"00",X"00",X"00",X"08",X"4A",X"0E",X"04",
		X"32",X"32",X"F6",X"51",X"00",X"00",X"00",X"00",X"F1",X"B6",X"96",X"F0",X"F8",X"77",X"C4",X"40",
		X"F9",X"F5",X"F1",X"F1",X"E2",X"CC",X"77",X"22",X"04",X"06",X"11",X"22",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"99",X"FA",X"72",X"00",X"88",X"07",X"00",X"FF",X"F0",X"F2",X"F1",
		X"00",X"06",X"0C",X"07",X"89",X"C4",X"E6",X"F9",X"00",X"00",X"00",X"06",X"4A",X"0C",X"0C",X"04",
		X"32",X"32",X"32",X"73",X"60",X"00",X"00",X"00",X"F1",X"B6",X"96",X"F0",X"F8",X"33",X"60",X"60",
		X"F9",X"F5",X"F1",X"F1",X"E2",X"EE",X"11",X"00",X"06",X"15",X"11",X"00",X"00",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"32",X"00",X"10",X"43",X"00",X"FF",X"F0",X"F0",X"F0",
		X"00",X"E0",X"3C",X"07",X"89",X"C4",X"E2",X"F1",X"00",X"00",X"80",X"C0",X"48",X"68",X"2C",X"24",
		X"32",X"32",X"10",X"11",X"00",X"00",X"00",X"00",X"F0",X"B4",X"96",X"F0",X"F8",X"33",X"00",X"00",
		X"F1",X"F1",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"24",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"32",X"00",X"10",X"43",X"00",X"FF",X"F0",X"F0",X"F1",
		X"00",X"E0",X"3C",X"07",X"89",X"C4",X"E2",X"F9",X"00",X"00",X"80",X"C0",X"48",X"68",X"2C",X"24",
		X"32",X"32",X"10",X"11",X"00",X"00",X"00",X"00",X"F1",X"B4",X"96",X"F0",X"F8",X"33",X"00",X"00",
		X"F9",X"F1",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"24",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"32",X"00",X"10",X"43",X"00",X"FF",X"F0",X"F1",X"F3",
		X"00",X"E0",X"3C",X"07",X"89",X"C4",X"EA",X"FD",X"00",X"00",X"80",X"C0",X"48",X"68",X"2C",X"24",
		X"32",X"32",X"10",X"11",X"00",X"00",X"00",X"00",X"F3",X"B5",X"96",X"F0",X"F8",X"33",X"00",X"00",
		X"FD",X"F9",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"24",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"32",X"00",X"10",X"43",X"00",X"FF",X"F0",X"F1",X"F3",
		X"00",X"E0",X"3C",X"07",X"89",X"C0",X"E8",X"FD",X"00",X"00",X"80",X"C0",X"48",X"68",X"2C",X"24",
		X"32",X"32",X"10",X"11",X"00",X"00",X"00",X"00",X"F3",X"F1",X"B4",X"F0",X"F8",X"33",X"00",X"00",
		X"FD",X"F9",X"F1",X"F1",X"E2",X"CC",X"00",X"00",X"24",X"04",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"22",X"31",X"30",X"31",X"31",X"31",X"00",X"00",X"00",X"77",X"B8",X"D4",X"62",X"31",
		X"00",X"00",X"00",X"EE",X"C1",X"82",X"14",X"38",X"00",X"00",X"04",X"08",X"00",X"88",X"88",X"88",
		X"31",X"31",X"31",X"30",X"21",X"12",X"00",X"00",X"21",X"52",X"A4",X"48",X"F7",X"F0",X"00",X"00",
		X"B8",X"D4",X"62",X"31",X"FE",X"F0",X"00",X"00",X"88",X"88",X"88",X"00",X"88",X"C4",X"00",X"00",
		X"00",X"00",X"11",X"11",X"11",X"33",X"33",X"33",X"88",X"88",X"BB",X"DC",X"DC",X"2E",X"2E",X"1F",
		X"00",X"00",X"00",X"EE",X"F1",X"E0",X"91",X"67",X"00",X"00",X"00",X"00",X"BB",X"66",X"EE",X"6E",
		X"67",X"77",X"76",X"F1",X"30",X"00",X"00",X"00",X"7E",X"E8",X"80",X"88",X"F7",X"70",X"00",X"00",
		X"8F",X"C7",X"C3",X"73",X"73",X"FD",X"F1",X"10",X"CC",X"CC",X"CC",X"88",X"88",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"67",X"FF",X"11",X"33",X"77",X"DF",X"9F",X"1F",X"1F",X"FF",
		X"08",X"0C",X"4E",X"6B",X"79",X"78",X"78",X"0F",X"00",X"00",X"00",X"00",X"08",X"8C",X"C6",X"0F",
		X"0F",X"37",X"13",X"01",X"00",X"00",X"00",X"00",X"0F",X"EF",X"EF",X"EF",X"6F",X"27",X"03",X"01",
		X"FF",X"8F",X"8F",X"9F",X"BF",X"EE",X"CC",X"88",X"FF",X"6E",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"F7",X"71",X"72",X"62",X"00",X"00",X"77",X"FF",X"8F",X"8F",X"E3",X"71",
		X"11",X"FF",X"EE",X"5D",X"5D",X"B8",X"B8",X"70",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",
		X"31",X"31",X"31",X"10",X"10",X"10",X"00",X"00",X"10",X"31",X"31",X"EB",X"EB",X"F7",X"F7",X"80",
		X"98",X"6E",X"1F",X"1F",X"FF",X"EE",X"00",X"00",X"C4",X"44",X"88",X"FF",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"32",X"EC",X"00",X"11",X"33",X"77",X"FE",X"F8",X"90",X"10",
		X"00",X"00",X"00",X"44",X"88",X"EE",X"9F",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"4C",
		X"62",X"31",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"98",X"D4",X"72",X"30",X"10",X"00",
		X"8F",X"8F",X"9F",X"BF",X"EE",X"CC",X"88",X"00",X"6E",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"EF",X"00",X"11",X"33",X"77",X"DF",X"9F",X"1F",X"1F",
		X"00",X"00",X"00",X"44",X"62",X"71",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"C4",
		X"67",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"9F",X"77",X"11",X"00",X"00",X"00",X"00",
		X"70",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"33",X"67",X"FF",X"11",X"33",X"77",X"DF",X"9F",X"1F",X"1F",X"FF",
		X"08",X"0C",X"4E",X"6B",X"79",X"78",X"78",X"0F",X"00",X"00",X"00",X"00",X"08",X"8C",X"C6",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"67",X"00",X"11",X"33",X"77",X"DF",X"9F",X"1F",X"1F",
		X"00",X"00",X"00",X"44",X"62",X"71",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"C4",
		X"E3",X"31",X"10",X"00",X"00",X"00",X"00",X"00",X"1F",X"9F",X"F7",X"F1",X"72",X"30",X"10",X"00",
		X"70",X"60",X"11",X"77",X"EE",X"CC",X"88",X"00",X"B3",X"44",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"67",X"00",X"00",X"00",X"00",X"11",X"77",X"9F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"EF",X"33",X"11",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"9F",X"DF",X"77",X"33",X"11",X"00",
		X"70",X"70",X"71",X"62",X"44",X"00",X"00",X"00",X"C4",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"37",X"13",X"01",X"00",X"00",X"00",X"00",X"0F",X"EF",X"EF",X"EF",X"6F",X"27",X"03",X"01",
		X"FF",X"8F",X"8F",X"9F",X"BF",X"EE",X"CC",X"88",X"FF",X"6E",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"10",X"FE",X"00",X"22",X"22",X"77",X"F5",X"FA",X"F5",X"F2",
		X"00",X"24",X"24",X"12",X"CD",X"E6",X"FB",X"F5",X"00",X"00",X"00",X"00",X"80",X"68",X"06",X"00",
		X"FE",X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"F2",X"F5",X"7A",X"B4",X"70",X"31",X"31",X"11",
		X"F5",X"FA",X"F5",X"F2",X"E0",X"A8",X"A8",X"88",X"88",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"00",X"00",X"00",X"11",X"33",X"76",X"70",X"70",X"70",X"44",X"EE",X"CC",X"77",X"F8",X"F0",X"F0",
		X"F0",X"02",X"63",X"71",X"8B",X"CD",X"E6",X"F3",X"80",X"C0",X"60",X"38",X"9C",X"D6",X"D0",X"10",
		X"70",X"63",X"73",X"13",X"01",X"00",X"00",X"00",X"F0",X"B4",X"96",X"F0",X"DE",X"7E",X"70",X"00",
		X"F1",X"F1",X"F1",X"E2",X"F1",X"F3",X"E2",X"00",X"10",X"54",X"FE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"76",X"70",X"70",X"70",X"44",X"EE",X"CC",X"77",X"F8",X"F0",X"F0",
		X"F0",X"02",X"63",X"71",X"8B",X"CD",X"E6",X"F3",X"80",X"C0",X"60",X"38",X"9C",X"D6",X"D0",X"10",
		X"70",X"63",X"73",X"13",X"01",X"00",X"00",X"00",X"F0",X"B4",X"96",X"F0",X"DE",X"7E",X"70",X"00",
		X"F1",X"F1",X"F1",X"E2",X"F1",X"F3",X"E2",X"00",X"10",X"54",X"FE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"76",X"70",X"70",X"70",X"44",X"EE",X"CC",X"77",X"F8",X"F0",X"F0",
		X"F0",X"02",X"63",X"71",X"8B",X"CD",X"E6",X"F3",X"80",X"C0",X"60",X"38",X"9C",X"D6",X"D0",X"10",
		X"70",X"63",X"73",X"13",X"01",X"00",X"00",X"00",X"F0",X"B4",X"96",X"F0",X"DE",X"7E",X"70",X"00",
		X"F1",X"F1",X"F1",X"E2",X"F1",X"F3",X"E2",X"00",X"10",X"54",X"FE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"76",X"70",X"70",X"70",X"44",X"EE",X"CC",X"77",X"E8",X"F0",X"B0",
		X"F0",X"02",X"63",X"71",X"8B",X"45",X"E2",X"D1",X"80",X"C0",X"60",X"38",X"9C",X"D6",X"D0",X"10",
		X"70",X"63",X"73",X"13",X"01",X"00",X"00",X"00",X"B0",X"B4",X"86",X"F0",X"DE",X"7E",X"70",X"00",
		X"D1",X"F1",X"71",X"E2",X"F1",X"F3",X"E2",X"00",X"10",X"54",X"FE",X"CC",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"55",X"00",X"00",X"00",X"00",X"0F",X"7F",X"0F",X"55",
		X"00",X"00",X"00",X"00",X"0F",X"9F",X"0F",X"55",X"00",X"00",X"00",X"00",X"0F",X"EF",X"0F",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"00",X"00",X"00",X"00",X"0F",X"7F",X"0F",X"55",X"00",X"00",X"00",X"00",X"0F",X"9F",X"0F",X"55",
		X"00",X"00",X"00",X"00",X"0F",X"EF",X"0F",X"55",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"AA",X"F0",X"F7",X"F0",X"00",X"00",X"00",X"00",
		X"AA",X"F0",X"F9",X"F0",X"00",X"00",X"00",X"00",X"AA",X"F0",X"FE",X"F0",X"00",X"00",X"00",X"00",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",
		X"AA",X"F0",X"F7",X"F0",X"00",X"00",X"00",X"00",X"AA",X"F0",X"F9",X"F0",X"00",X"00",X"00",X"00",
		X"AA",X"F0",X"FE",X"F0",X"00",X"00",X"00",X"00",X"AA",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",
		X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"FF",X"FB",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"FF",
		X"11",X"00",X"00",X"30",X"F0",X"F0",X"F0",X"F0",X"FF",X"FE",X"F7",X"F1",X"F3",X"F3",X"F7",X"F7",
		X"F7",X"FE",X"FC",X"F9",X"F2",X"F0",X"F4",X"F4",X"F0",X"F3",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"80",X"E0",X"F0",X"E1",X"C3",X"87",X"8F",X"EF",
		X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"F0",X"FC",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F7",X"F3",X"F9",X"F4",X"F0",X"F2",X"F2",
		X"0F",X"8F",X"9E",X"FC",X"CC",X"CC",X"EE",X"EE",X"48",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"01",X"F7",X"F7",X"F3",X"F3",X"33",X"17",X"1F",X"0F",
		X"F4",X"F4",X"F0",X"F2",X"F9",X"FC",X"FE",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F3",X"F0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"7F",X"1F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"FF",X"FF",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"FC",X"F0",X"F2",X"F2",X"F0",X"F4",X"F9",X"F3",X"F7",X"FE",
		X"EE",X"EE",X"CC",X"CC",X"FC",X"FE",X"F7",X"FF",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C8",
		X"FF",X"FF",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"FD",X"F7",X"F7",X"F3",X"91",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8F",X"F8",X"F8",X"F8",X"F8",X"FA",X"FA",X"FA",X"0F",X"F0",X"F7",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"E0",X"E0",X"E0",X"E0",X"E4",X"E4",X"E4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FA",X"FA",X"F8",X"F8",X"F8",X"F8",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"DE",X"BC",X"78",X"EF",X"DE",X"BC",X"78",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"E4",X"E4",X"E4",X"E0",X"E0",X"E0",X"E0",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"88",X"C4",X"E2",X"F1",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"88",X"C4",X"E2",X"F1",
		X"00",X"00",X"13",X"54",X"36",X"00",X"72",X"72",X"00",X"00",X"F1",X"F0",X"FC",X"CC",X"DD",X"DD",
		X"00",X"00",X"F1",X"F0",X"B0",X"0F",X"F8",X"FC",X"00",X"00",X"84",X"82",X"C4",X"08",X"04",X"CC",
		X"72",X"72",X"30",X"54",X"52",X"21",X"00",X"00",X"DD",X"DD",X"FC",X"FC",X"F0",X"E1",X"00",X"00",
		X"FC",X"F8",X"F0",X"F4",X"F0",X"E1",X"00",X"00",X"CC",X"04",X"88",X"82",X"C4",X"C4",X"00",X"00",
		X"00",X"00",X"12",X"54",X"36",X"00",X"72",X"72",X"00",X"00",X"F2",X"F0",X"FC",X"CC",X"DD",X"DD",
		X"00",X"00",X"F2",X"F0",X"70",X"0F",X"F8",X"FC",X"00",X"00",X"84",X"82",X"44",X"08",X"04",X"CC",
		X"72",X"72",X"30",X"54",X"52",X"30",X"00",X"00",X"DD",X"DD",X"FC",X"FC",X"F0",X"D2",X"00",X"00",
		X"FC",X"F8",X"F0",X"F8",X"F0",X"D2",X"00",X"00",X"CC",X"04",X"88",X"8A",X"C4",X"C4",X"00",X"00",
		X"00",X"00",X"12",X"54",X"26",X"00",X"72",X"72",X"00",X"00",X"F4",X"F0",X"EC",X"CC",X"DD",X"DD",
		X"00",X"00",X"F4",X"F0",X"E0",X"0F",X"F8",X"FC",X"00",X"00",X"84",X"82",X"C4",X"08",X"04",X"CC",
		X"72",X"72",X"30",X"55",X"52",X"30",X"00",X"00",X"DD",X"DD",X"FC",X"FD",X"F0",X"B4",X"00",X"00",
		X"FC",X"F8",X"F0",X"F1",X"F0",X"B4",X"00",X"00",X"CC",X"04",X"88",X"82",X"C4",X"C4",X"00",X"00",
		X"00",X"00",X"12",X"54",X"36",X"00",X"72",X"72",X"00",X"00",X"F8",X"F0",X"DC",X"CC",X"DD",X"DD",
		X"00",X"00",X"F8",X"F0",X"D0",X"0F",X"F8",X"FC",X"00",X"00",X"8C",X"82",X"C4",X"08",X"04",X"CC",
		X"72",X"72",X"30",X"54",X"52",X"30",X"00",X"00",X"DD",X"DD",X"FC",X"FE",X"F0",X"78",X"00",X"00",
		X"FC",X"F8",X"F0",X"F2",X"F0",X"78",X"00",X"00",X"CC",X"04",X"88",X"82",X"C4",X"4C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"C9",X"00",X"00",X"00",X"00",X"FF",X"01",X"FF",X"3C",
		X"33",X"77",X"FF",X"00",X"FF",X"0F",X"FF",X"F0",X"EE",X"0E",X"F0",X"00",X"EE",X"0C",X"DF",X"D1",
		X"C8",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"0F",X"4F",X"5E",X"01",X"00",X"00",X"00",
		X"F0",X"0F",X"0F",X"F0",X"F8",X"7C",X"37",X"03",X"D0",X"1E",X"0C",X"E0",X"00",X"0F",X"EE",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"87",X"F0",X"F0",X"F0",X"F0",X"E1",X"87",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"C3",X"2D",X"1E",X"0F",X"0F",X"F1",X"F7",X"3F",X"97",X"4B",X"2D",X"96",X"4A",
		X"47",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"8F",X"47",X"23",X"11",X"00",
		X"0F",X"0F",X"0E",X"1C",X"28",X"43",X"87",X"0F",X"1C",X"28",X"C1",X"07",X"0F",X"0F",X"0F",X"0F",
		X"6F",X"BF",X"DF",X"FF",X"EE",X"5C",X"30",X"F0",X"DF",X"EF",X"9B",X"71",X"F0",X"F0",X"F0",X"F0",
		X"D2",X"E9",X"FC",X"FE",X"FF",X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"D2",X"E9",X"FC",X"FE",
		X"F0",X"F8",X"7C",X"3E",X"1F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"7C",X"3E",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"D1",X"A3",X"93",X"DF",X"B7",X"A3",X"77",X"FF",X"BF",X"DF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"1E",X"2C",X"49",X"1C",X"28",X"49",X"43",X"83",X"07",X"0F",X"0F",
		X"43",X"2D",X"96",X"4B",X"2D",X"1E",X"0F",X"0F",X"BF",X"7E",X"3E",X"B4",X"78",X"78",X"F0",X"F0",
		X"47",X"23",X"11",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"8F",X"47",X"23",X"11",X"00",
		X"0F",X"1E",X"1E",X"3C",X"3C",X"78",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"E0",X"80",X"00",X"00",X"30",X"37",X"E0",X"80",X"10",X"31",X"50",X"A1",X"43",X"87",
		X"66",X"77",X"FE",X"FC",X"FE",X"F7",X"7B",X"3D",X"70",X"F0",X"F0",X"E0",X"E2",X"F7",X"FF",X"CC",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"F7",X"F3",X"F1",X"CB",X"ED",X"FE",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"1E",X"2C",X"58",X"A0",X"C8",X"C8",X"08",X"00",X"C8",X"90",X"10",X"30",X"30",X"70",X"70",X"F0",
		X"0E",X"0C",X"08",X"00",X"00",X"00",X"01",X"9A",X"11",X"00",X"01",X"12",X"24",X"58",X"A1",X"43",
		X"F1",X"F8",X"F0",X"FC",X"F6",X"7B",X"3D",X"1E",X"80",X"C8",X"C0",X"E0",X"E0",X"F0",X"F8",X"B8",
		X"EC",X"FF",X"FF",X"FF",X"F7",X"F1",X"F0",X"F0",X"87",X"CB",X"ED",X"FE",X"FE",X"FF",X"F7",X"F1",
		X"3C",X"68",X"D0",X"B0",X"74",X"FE",X"DF",X"8F",X"70",X"ED",X"C7",X"C1",X"C1",X"E0",X"E8",X"7E",
		X"81",X"E8",X"F8",X"7C",X"7C",X"3E",X"7F",X"EE",X"1E",X"34",X"F6",X"E2",X"D0",X"B0",X"61",X"C3",
		X"E0",X"F0",X"70",X"FC",X"F6",X"7B",X"3D",X"1E",X"00",X"80",X"E0",X"F2",X"F1",X"F0",X"F8",X"FA",
		X"FE",X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"F0",X"87",X"CB",X"ED",X"FE",X"EE",X"FE",X"FF",X"FF",
		X"2C",X"58",X"A1",X"42",X"84",X"08",X"00",X"88",X"95",X"08",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"10",X"10",X"30",X"30",X"70",X"70",X"E2",X"F0",X"F0",X"F1",X"F1",X"D0",X"A1",X"43",X"87",
		X"F7",X"FF",X"F7",X"FB",X"FD",X"F6",X"7B",X"3D",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"F7",X"FA",
		X"F1",X"C8",X"CC",X"88",X"88",X"00",X"00",X"11",X"CB",X"ED",X"76",X"33",X"11",X"10",X"74",X"FE",
		X"1E",X"2C",X"58",X"B0",X"70",X"F8",X"E0",X"80",X"FC",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"03",X"03",X"07",X"04",X"04",X"07",X"00",X"09",X"08",X"0C",X"0F",X"25",X"25",X"0F",
		X"00",X"0C",X"0F",X"0F",X"09",X"00",X"09",X"0B",X"00",X"00",X"00",X"08",X"0C",X"0C",X"4A",X"4A",
		X"07",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"09",X"09",X"0B",X"0F",X"C2",X"0F",X"01",X"00",
		X"0E",X"4A",X"0E",X"03",X"01",X"07",X"08",X"00",X"0E",X"06",X"0C",X"0C",X"0C",X"08",X"00",X"00",
		X"C0",X"86",X"07",X"07",X"02",X"00",X"86",X"00",X"00",X"10",X"01",X"33",X"53",X"CB",X"8E",X"CE",
		X"02",X"03",X"07",X"06",X"8A",X"11",X"33",X"11",X"10",X"02",X"06",X"04",X"04",X"00",X"16",X"16",
		X"00",X"0F",X"0F",X"11",X"01",X"03",X"07",X"06",X"00",X"11",X"19",X"33",X"00",X"0E",X"00",X"00",
		X"02",X"06",X"21",X"BA",X"11",X"08",X"08",X"80",X"00",X"00",X"00",X"8C",X"04",X"0E",X"07",X"02",
		X"00",X"12",X"12",X"70",X"70",X"E1",X"F0",X"34",X"16",X"F0",X"F0",X"E1",X"F0",X"78",X"F0",X"F0",
		X"A4",X"C3",X"F0",X"78",X"F0",X"F0",X"B4",X"96",X"00",X"00",X"C0",X"86",X"E0",X"F0",X"F0",X"C3",
		X"3C",X"F0",X"F0",X"34",X"16",X"10",X"01",X"00",X"F0",X"96",X"F0",X"F0",X"F0",X"E1",X"F0",X"70",
		X"F0",X"F0",X"E1",X"F0",X"78",X"F0",X"E1",X"C2",X"F0",X"F0",X"E0",X"E0",X"C2",X"A4",X"80",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"32",X"00",X"00",X"73",X"FC",X"FF",X"FF",X"FB",X"F7",
		X"00",X"00",X"CC",X"FF",X"FF",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"88",X"80",X"80",X"CC",X"CC",
		X"33",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F3",X"F7",X"77",X"00",X"00",
		X"FB",X"F3",X"FF",X"FF",X"FC",X"C8",X"00",X"00",X"C8",X"C8",X"CC",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"50",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"61",X"10",X"01",X"01",
		X"1E",X"87",X"8C",X"9D",X"1E",X"D2",X"0E",X"6E",X"18",X"1E",X"72",X"F9",X"FC",X"A1",X"C3",X"8F",
		X"00",X"00",X"00",X"00",X"10",X"10",X"21",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"60",
		X"00",X"00",X"00",X"00",X"00",X"10",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"25",X"0F",X"08",X"33",X"3B",X"0B",X"DE",X"5E",X"D2",X"87",X"89",X"DD",X"11",X"C1",X"83",X"1A",
		X"80",X"80",X"08",X"0C",X"88",X"00",X"78",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"E1",X"10",X"61",X"10",X"30",X"01",X"10",
		X"C4",X"1D",X"84",X"6E",X"C2",X"1F",X"1B",X"A5",X"FC",X"BC",X"8F",X"61",X"61",X"C9",X"C9",X"8F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"40",X"80",X"00",X"00",X"00",X"00",X"00",
		X"2D",X"68",X"C0",X"80",X"00",X"00",X"00",X"00",X"0F",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"1E",X"34",X"76",X"0D",X"B7",X"E6",X"B3",X"0E",X"3C",X"E6",X"F7",X"6E",X"C0",X"60",X"07",
		X"08",X"E0",X"00",X"00",X"0C",X"84",X"C0",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"87",X"82",X"82",X"00",X"00",X"00",X"00",X"00",X"69",X"3C",X"10",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"00",X"00",X"30",X"10",X"00",X"00",X"80",X"C0",X"E0",X"70",X"30",X"96",X"D2",
		X"40",X"60",X"60",X"30",X"B4",X"F0",X"87",X"0F",X"10",X"10",X"10",X"30",X"B0",X"3C",X"3C",X"1E",
		X"00",X"00",X"00",X"00",X"70",X"30",X"01",X"00",X"70",X"70",X"25",X"25",X"2D",X"E1",X"C3",X"0F",
		X"0D",X"08",X"28",X"18",X"18",X"0F",X"3C",X"F0",X"4B",X"69",X"3C",X"3C",X"87",X"E0",X"68",X"0E",
		X"20",X"20",X"20",X"68",X"68",X"69",X"4B",X"C3",X"00",X"10",X"30",X"60",X"61",X"E1",X"69",X"0F",
		X"00",X"00",X"00",X"10",X"30",X"F0",X"C0",X"80",X"00",X"60",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"86",X"0C",X"0F",X"C3",X"70",X"34",X"03",X"03",X"01",X"01",X"21",X"C3",X"92",X"92",X"0B",X"01",
		X"81",X"F0",X"87",X"0E",X"86",X"3C",X"0E",X"E1",X"80",X"00",X"00",X"00",X"E0",X"80",X"00",X"08",
		X"00",X"30",X"40",X"00",X"01",X"30",X"60",X"00",X"61",X"E1",X"07",X"3C",X"F0",X"E1",X"30",X"61",
		X"18",X"09",X"0D",X"85",X"87",X"A5",X"4B",X"0F",X"78",X"F0",X"C3",X"0F",X"2D",X"78",X"78",X"69",
		X"00",X"10",X"00",X"10",X"30",X"70",X"C0",X"00",X"D0",X"30",X"70",X"C0",X"90",X"10",X"30",X"00",
		X"84",X"0C",X"4A",X"E0",X"C3",X"00",X"00",X"00",X"69",X"4B",X"43",X"0F",X"96",X"90",X"10",X"00",
		X"E1",X"3C",X"0F",X"0F",X"0F",X"87",X"01",X"01",X"01",X"03",X"A4",X"68",X"C2",X"E1",X"69",X"1E",
		X"F0",X"78",X"07",X"34",X"61",X"2D",X"3C",X"78",X"E0",X"08",X"08",X"80",X"C0",X"00",X"00",X"80",
		X"03",X"12",X"42",X"4A",X"C2",X"80",X"80",X"80",X"0F",X"3C",X"B0",X"90",X"00",X"00",X"00",X"00",
		X"18",X"08",X"80",X"80",X"C0",X"40",X"20",X"00",X"C0",X"60",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"03",X"34",X"F0",X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"12",X"34",X"34",X"F0",X"F0",X"F0",X"F0",
		X"C3",X"D2",X"96",X"78",X"F0",X"F0",X"F0",X"3C",X"C3",X"87",X"78",X"F0",X"F0",X"F0",X"E1",X"C3",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"78",X"96",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"F0",X"F0",X"C3",X"C3",X"E1",X"F0",X"78",X"D2",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"E1",
		X"80",X"E0",X"E0",X"E0",X"E0",X"78",X"78",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F0",X"78",X"3C",X"34",X"34",X"30",X"30",
		X"3C",X"78",X"78",X"F0",X"F0",X"E1",X"E1",X"F0",X"C3",X"F0",X"F0",X"F0",X"F0",X"78",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"3C",X"12",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"78",X"F0",X"78",X"87",X"C3",X"F0",X"F0",X"F0",X"E1",X"F0",X"F0",X"F0",X"F0",X"E1",X"D2",X"F0",
		X"E0",X"F0",X"E1",X"C2",X"86",X"86",X"84",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"C3",X"86",X"00",X"00",X"00",X"00",X"F0",X"78",X"08",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"44",X"22",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"22",X"AA",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"8C",X"DF",X"FF",X"EE",X"77",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",
		X"33",X"01",X"10",X"30",X"00",X"00",X"00",X"00",X"DD",X"77",X"7F",X"B7",X"55",X"88",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"00",X"CC",X"88",X"88",X"44",X"88",X"CC",X"66",X"11",
		X"00",X"00",X"00",X"02",X"23",X"11",X"08",X"88",X"04",X"00",X"00",X"10",X"02",X"30",X"09",X"12",
		X"00",X"00",X"09",X"81",X"00",X"02",X"01",X"08",X"00",X"00",X"08",X"00",X"00",X"08",X"00",X"66",
		X"88",X"30",X"00",X"10",X"00",X"02",X"00",X"00",X"20",X"03",X"83",X"82",X"00",X"00",X"00",X"02",
		X"0F",X"0F",X"38",X"02",X"00",X"10",X"00",X"00",X"04",X"00",X"00",X"02",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"33",X"76",X"0C",X"00",X"CC",X"00",X"00",X"00",X"E8",X"80",X"00",X"44",X"00",
		X"33",X"44",X"08",X"00",X"00",X"00",X"00",X"00",X"F1",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"F0",X"80",X"C4",X"37",X"31",X"10",X"00",X"00",X"C4",X"00",X"00",X"88",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"44",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"33",X"76",X"0C",X"00",X"CC",X"00",X"00",X"00",X"E8",X"80",X"00",X"44",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F1",X"12",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"F0",X"80",X"C4",X"37",X"31",X"10",X"00",X"00",X"C4",X"00",X"00",X"88",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"08",X"09",X"00",X"00",
		X"08",X"00",X"00",X"04",X"00",X"00",X"80",X"00",X"11",X"00",X"00",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"04",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"42",X"60",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F8",X"FF",X"1F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FF",X"3F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"FF",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"7F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"C0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"70",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",X"F0",X"B0",X"D0",X"F0",
		X"FF",X"FF",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F8",X"FF",X"FF",X"3F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F8",X"FF",X"FF",X"7F",X"1F",X"3D",X"35",X"F0",X"D0",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",X"0F",X"0F",X"0F",X"0F",X"3F",X"FF",X"FF",X"F8",
		X"70",X"70",X"73",X"F0",X"F0",X"F0",X"F0",X"F0",X"3F",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"3F",X"FF",X"FF",X"FE",X"F0",X"F0",X"3F",X"7F",X"FF",X"FF",X"FC",X"F0",X"F0",X"F0",
		X"35",X"35",X"9A",X"CD",X"E2",X"F0",X"F0",X"F0",X"7F",X"7F",X"7F",X"7F",X"7E",X"F8",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F7",X"F0",X"F0",X"F0",X"F0",X"F1",X"E7",X"FF",X"4F",
		X"F0",X"F0",X"F1",X"D5",X"DD",X"BB",X"FC",X"F8",X"F1",X"D5",X"BA",X"FC",X"E9",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"27",X"00",X"00",X"01",X"03",X"07",X"0F",X"0F",X"0F",
		X"80",X"48",X"48",X"3C",X"2C",X"1E",X"1E",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"80",
		X"5B",X"2D",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"4F",X"A7",X"79",X"5A",X"6D",X"ED",
		X"0F",X"0F",X"1E",X"2D",X"4B",X"96",X"E1",X"69",X"80",X"C0",X"48",X"68",X"A4",X"3E",X"7E",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"10",X"01",X"03",X"07",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"A7",X"5B",X"2D",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"FF",X"B7",X"5A",X"2D",
		X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"C3",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"96",X"F0",X"F0",X"F0",X"F0",X"F0",X"5A",X"96",X"2D",X"4B",X"F1",X"F0",X"F0",X"E0",
		X"1F",X"3F",X"7E",X"ED",X"CB",X"87",X"0F",X"0F",X"CB",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"BF",X"E7",X"A3",X"F1",X"68",X"3C",X"38",X"32",
		X"0F",X"C3",X"6D",X"FE",X"BF",X"E3",X"60",X"F0",X"0F",X"0F",X"0F",X"0F",X"86",X"EA",X"F7",X"F0",
		X"0E",X"0C",X"08",X"00",X"10",X"30",X"61",X"D2",X"10",X"30",X"61",X"D2",X"F0",X"F0",X"F0",X"F0",
		X"E1",X"F0",X"F0",X"F1",X"E2",X"F3",X"B3",X"DD",X"D1",X"F6",X"BA",X"FC",X"FC",X"70",X"70",X"F0",
		X"F0",X"F1",X"F1",X"E3",X"E0",X"F1",X"F0",X"F0",X"FF",X"FF",X"FF",X"0F",X"7B",X"34",X"8B",X"CC",
		X"FF",X"7E",X"DE",X"FC",X"7C",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F1",X"F1",X"F1",X"F3",X"F3",X"F3",X"FF",X"FF",X"EF",X"CF",X"CF",X"CF",X"8F",X"8F",
		X"EE",X"FF",X"FF",X"0F",X"FF",X"D3",X"1F",X"07",X"B8",X"30",X"30",X"38",X"FC",X"FC",X"FC",X"FE",
		X"F0",X"B0",X"F0",X"E0",X"D0",X"F0",X"F0",X"F0",X"78",X"F0",X"F0",X"F0",X"F0",X"B0",X"F0",X"B0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FE",X"FE",X"7E",X"7F",X"7F",X"3F",X"3F",X"3F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"B0",X"E0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",
		X"F7",X"F7",X"E7",X"EF",X"CF",X"CF",X"8F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F3",X"E3",X"E3",X"F4",X"F4",X"F0",X"80",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"7C",X"7E",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",
		X"7E",X"3E",X"3E",X"3F",X"F1",X"F1",X"F1",X"11",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"D2",X"F0",X"78",X"F0",X"F4",X"FE",X"DF",X"87",X"F0",X"ED",X"C7",X"C1",X"C1",X"E0",X"E8",X"7E",
		X"FE",X"08",X"08",X"0C",X"0C",X"0E",X"0E",X"87",X"0F",X"0F",X"87",X"87",X"87",X"00",X"00",X"00",
		X"0F",X"69",X"FC",X"77",X"3F",X"0F",X"0F",X"0F",X"1E",X"0F",X"87",X"E1",X"F8",X"78",X"78",X"78",
		X"0E",X"0D",X"0B",X"07",X"3C",X"70",X"31",X"31",X"F0",X"78",X"F0",X"F3",X"CC",X"8B",X"16",X"35",
		X"0F",X"0F",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"F7",X"11",X"11",X"33",X"33",X"77",X"77",X"EE",
		X"F0",X"C8",X"CC",X"88",X"88",X"00",X"00",X"11",X"B4",X"F0",X"61",X"30",X"10",X"10",X"74",X"EE",
		X"F1",X"F1",X"F0",X"FC",X"33",X"1D",X"86",X"CA",X"FF",X"FF",X"FF",X"FF",X"F3",X"F0",X"F8",X"F8",
		X"77",X"FF",X"EE",X"88",X"10",X"01",X"01",X"01",X"FF",X"99",X"11",X"10",X"C3",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"3C",X"F0",X"78",X"79",X"7F",X"78",X"78",X"78",X"F0",X"F1",X"F7",X"FF",X"9E",
		X"31",X"31",X"70",X"74",X"FF",X"FF",X"FF",X"FF",X"35",X"16",X"8B",X"CC",X"F3",X"F0",X"D8",X"00",
		X"EE",X"FF",X"FE",X"F4",X"F2",X"79",X"F0",X"D2",X"70",X"F0",X"F0",X"E0",X"E2",X"F7",X"FF",X"F7",
		X"F7",X"7E",X"7E",X"FC",X"FC",X"F8",X"F8",X"1E",X"F0",X"F0",X"F0",X"87",X"87",X"87",X"0F",X"0F",
		X"CA",X"86",X"1D",X"33",X"FC",X"F0",X"A1",X"01",X"F8",X"F8",X"F0",X"D2",X"0E",X"0D",X"0B",X"07",
		X"01",X"01",X"01",X"10",X"08",X"0E",X"0F",X"87",X"0F",X"0F",X"0F",X"C3",X"10",X"11",X"19",X"1F",
		X"F0",X"F0",X"F0",X"1F",X"1F",X"1F",X"0F",X"0F",X"1E",X"87",X"87",X"C3",X"CB",X"E9",X"ED",X"CF",
		X"81",X"E8",X"F8",X"7C",X"7C",X"3E",X"7F",X"F6",X"1E",X"34",X"F6",X"F2",X"F0",X"E1",X"F0",X"B4",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"80",X"80",X"C4",X"E6",X"F3",X"73",X"73",X"71",
		X"00",X"00",X"00",X"00",X"0F",X"8F",X"CF",X"EF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"71",X"31",X"30",X"30",X"30",X"10",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"F7",X"0F",X"8F",X"CF",X"EF",X"DF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",
		X"10",X"10",X"10",X"10",X"3C",X"2C",X"2C",X"68",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"1E",
		X"68",X"48",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C8",X"48",X"EC",X"E4",X"70",X"F0",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"F3",X"F3",X"F3",X"F1",X"F1",X"71",X"70",X"70",X"DF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",
		X"B0",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E1",X"80",X"C0",X"C0",X"E0",X"60",X"B0",X"F0",X"F0",
		X"70",X"30",X"31",X"20",X"30",X"31",X"31",X"90",X"CC",X"8B",X"34",X"7B",X"F0",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",X"FF",X"3C",X"BC",X"FC",X"B8",X"98",X"89",X"01",X"01",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"20",X"71",X"70",X"B0",
		X"33",X"0C",X"C2",X"ED",X"F0",X"FF",X"FF",X"FF",X"01",X"02",X"02",X"02",X"C0",X"C8",X"C8",X"80",
		X"00",X"10",X"10",X"30",X"20",X"70",X"70",X"B0",X"90",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"78",
		X"F0",X"F0",X"F0",X"F0",X"B4",X"68",X"C0",X"80",X"B4",X"68",X"C0",X"80",X"00",X"01",X"03",X"07",
		X"B0",X"F8",X"12",X"07",X"0F",X"0F",X"0F",X"0F",X"FF",X"67",X"A3",X"F1",X"78",X"3C",X"0F",X"0F",
		X"C4",X"67",X"E5",X"F2",X"53",X"73",X"E1",X"A1",X"0F",X"0F",X"0F",X"0F",X"87",X"CB",X"ED",X"AD",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"3D",X"0F",X"0F",X"1E",X"3D",X"7B",X"E7",X"CF",X"8F",
		X"E8",X"7E",X"CF",X"9E",X"2D",X"C3",X"D2",X"69",X"00",X"80",X"E0",X"3C",X"4B",X"87",X"0F",X"0F",
		X"00",X"00",X"00",X"80",X"68",X"1E",X"0F",X"0F",X"80",X"80",X"80",X"80",X"80",X"80",X"68",X"1E",
		X"3D",X"D2",X"FC",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"4F",X"A7",X"5B",X"2D",X"1E",X"0F",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"88",X"08",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"3C",X"4B",X"96",X"2D",X"C3",X"87",X"87",X"C3",
		X"7B",X"B7",X"5B",X"3D",X"2D",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"4F",X"A7",X"4B",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C3",X"C3",X"E1",X"E1",X"E1",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"00",X"2C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",X"00",X"0E",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"78",X"E0",X"D0",X"E0",X"80",X"F0",X"F0",X"B0",X"D0",X"E0",X"80",X"00",X"00",
		X"E2",X"70",X"E0",X"80",X"00",X"00",X"00",X"00",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"70",X"F6",X"FE",X"FE",X"FE",X"FE",X"01",X"0E",X"00",X"00",X"3B",X"95",X"CA",X"CA",
		X"1E",X"00",X"00",X"33",X"FF",X"FF",X"EF",X"FF",X"F0",X"F0",X"47",X"EF",X"FF",X"FF",X"EF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"C3",
		X"00",X"00",X"00",X"00",X"10",X"F0",X"87",X"0F",X"80",X"80",X"80",X"00",X"F0",X"00",X"00",X"00",
		X"E1",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"F6",X"70",X"00",X"80",X"CA",X"CA",X"95",X"3B",X"74",X"F0",X"10",X"00",
		X"FF",X"EF",X"FF",X"FF",X"F3",X"F0",X"F0",X"10",X"FF",X"EF",X"FF",X"FF",X"FF",X"F7",X"F0",X"F0",
		X"E0",X"F0",X"D0",X"E0",X"78",X"F0",X"F0",X"F0",X"00",X"80",X"E0",X"F0",X"B0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"80",X"E0",X"70",X"71",X"E0",X"10",X"00",X"00",X"00",X"00",X"80",X"E8",X"7E",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"CF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"F3",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F7",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"F0",X"00",X"80",X"80",X"80",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"A3",X"03",X"47",X"07",X"8F",
		X"00",X"88",X"4C",X"2E",X"1F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"88",X"4C",X"0C",
		X"00",X"10",X"11",X"21",X"30",X"61",X"63",X"D3",X"8F",X"0F",X"87",X"4B",X"2D",X"96",X"4B",X"2C",
		X"0F",X"0F",X"0E",X"0C",X"0D",X"19",X"31",X"70",X"09",X"03",X"07",X"0F",X"0F",X"0F",X"8F",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"97",X"D7",X"FF",X"CE",X"4C",X"EC",X"F3",X"8C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",
		X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"F3",X"F1",X"70",X"30",X"10",X"00",X"00",
		X"F7",X"F3",X"79",X"B4",X"F0",X"F0",X"F0",X"F0",X"88",X"CC",X"EE",X"FF",X"F7",X"F3",X"79",X"B4",
		X"00",X"00",X"00",X"00",X"88",X"D9",X"B7",X"E7",X"00",X"00",X"23",X"77",X"BF",X"6F",X"CF",X"F8",
		X"0F",X"0F",X"8F",X"CF",X"E7",X"C0",X"81",X"03",X"0F",X"0E",X"0C",X"09",X"03",X"07",X"0F",X"0F",
		X"00",X"00",X"4C",X"2E",X"1F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"88",X"4C",X"2E",
		X"25",X"96",X"4B",X"2D",X"9E",X"FC",X"E0",X"80",X"0F",X"0F",X"87",X"5B",X"6C",X"80",X"00",X"00",
		X"0F",X"0F",X"2E",X"88",X"00",X"00",X"00",X"00",X"2E",X"88",X"00",X"80",X"80",X"80",X"80",X"80",
		X"00",X"01",X"00",X"00",X"00",X"30",X"30",X"77",X"07",X"F0",X"77",X"77",X"77",X"08",X"80",X"FF",
		X"08",X"E0",X"00",X"00",X"00",X"08",X"08",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"77",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"70",X"F0",X"77",X"67",X"47",X"07",X"F0",
		X"FF",X"F8",X"88",X"00",X"00",X"00",X"08",X"E0",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"33",X"33",X"00",X"77",X"77",X"47",X"F7",X"00",X"07",X"88",X"00",X"FF",
		X"00",X"88",X"E0",X"00",X"00",X"08",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"77",X"37",X"30",X"30",X"00",X"00",X"01",X"00",X"FF",X"F8",X"E7",X"47",X"70",X"40",X"F0",X"70",
		X"11",X"7F",X"88",X"00",X"00",X"80",X"E0",X"00",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"77",X"00",X"00",X"70",X"30",X"38",X"00",X"80",X"F8",
		X"00",X"00",X"00",X"00",X"06",X"88",X"88",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"77",X"04",X"20",X"21",X"00",X"00",X"00",X"00",X"C8",X"40",X"40",X"F0",X"40",X"70",X"00",X"00",
		X"F7",X"F0",X"80",X"E0",X"80",X"00",X"00",X"00",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"66",X"00",X"00",X"00",X"77",X"47",X"4F",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"04",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"76",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"47",X"C7",X"47",X"77",X"00",X"00",X"00",
		X"F1",X"F8",X"88",X"88",X"00",X"00",X"00",X"00",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"23",X"00",X"77",X"00",X"00",X"77",X"30",X"00",X"C7",X"47",X"CF",
		X"00",X"00",X"00",X"00",X"00",X"E8",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"77",X"04",X"30",X"21",X"00",X"00",X"00",X"00",X"FF",X"70",X"F0",X"C7",X"47",X"77",X"00",X"00",
		X"77",X"F8",X"88",X"E8",X"88",X"00",X"00",X"00",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"03",X"03",X"00",X"74",X"00",X"00",X"B0",X"00",X"77",X"0F",X"00",X"F7",
		X"00",X"00",X"60",X"00",X"00",X"08",X"08",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"8A",
		X"77",X"34",X"33",X"33",X"00",X"00",X"01",X"00",X"FF",X"F0",X"F8",X"67",X"47",X"00",X"C7",X"66",
		X"FF",X"F8",X"88",X"00",X"00",X"00",X"E8",X"00",X"8A",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"11",X"30",X"10",X"00",X"00",X"02",X"F8",X"C3",X"C5",X"D0",X"E3",
		X"00",X"00",X"04",X"F3",X"E4",X"3C",X"5A",X"2D",X"00",X"00",X"00",X"00",X"08",X"00",X"84",X"80",
		X"32",X"30",X"11",X"01",X"00",X"00",X"00",X"00",X"D3",X"E0",X"F0",X"FC",X"B0",X"31",X"00",X"00",
		X"57",X"1C",X"1E",X"E1",X"D1",X"C4",X"00",X"00",X"0C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"11",X"30",X"10",X"00",X"00",X"02",X"F8",X"C3",X"85",X"D0",X"E3",
		X"00",X"00",X"04",X"F3",X"E0",X"3C",X"5A",X"2D",X"00",X"00",X"00",X"00",X"08",X"00",X"84",X"80",
		X"32",X"30",X"11",X"01",X"00",X"00",X"00",X"00",X"D3",X"E0",X"F0",X"F8",X"B0",X"31",X"00",X"00",
		X"46",X"1C",X"1E",X"E1",X"D1",X"C4",X"00",X"00",X"0C",X"4C",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"70",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"71",
		X"00",X"00",X"10",X"30",X"F0",X"70",X"34",X"18",X"00",X"00",X"C0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"12",X"10",X"00",X"00",X"00",X"00",X"00",
		X"88",X"C4",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"66",X"E6",X"F1",
		X"00",X"10",X"70",X"F0",X"30",X"16",X"06",X"08",X"70",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"96",X"16",X"30",X"00",X"00",X"00",X"00",
		X"88",X"E6",X"E6",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"00",X"44",X"EE",X"E6",X"F1",
		X"30",X"70",X"F0",X"30",X"12",X"07",X"06",X"08",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"60",X"40",
		X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"96",X"1E",X"34",X"30",X"00",X"00",X"00",
		X"88",X"E6",X"F7",X"E2",X"C0",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"70",X"00",X"00",X"00",X"10",X"30",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"31",X"30",X"30",X"00",X"10",X"00",X"CC",X"CC",X"EE",X"E6",X"F1",
		X"70",X"F0",X"10",X"03",X"03",X"07",X"06",X"08",X"F0",X"F0",X"F0",X"F0",X"78",X"38",X"30",X"20",
		X"30",X"30",X"21",X"01",X"00",X"00",X"00",X"00",X"E1",X"96",X"1E",X"3C",X"3C",X"70",X"00",X"00",
		X"88",X"E6",X"F7",X"F3",X"F3",X"E0",X"00",X"00",X"20",X"00",X"88",X"88",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"00",X"00",X"30",X"70",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"30",X"F0",X"F0",
		X"00",X"10",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"80",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"71",X"70",X"70",X"30",X"00",X"88",X"CC",X"CC",X"EE",X"E6",X"F1",
		X"F0",X"10",X"01",X"03",X"03",X"07",X"06",X"08",X"F0",X"F0",X"F0",X"78",X"3C",X"18",X"10",X"10",
		X"70",X"70",X"61",X"03",X"01",X"00",X"00",X"00",X"E1",X"96",X"1E",X"3C",X"3C",X"78",X"70",X"00",
		X"88",X"E6",X"F7",X"F3",X"F3",X"F1",X"E0",X"00",X"10",X"10",X"88",X"CC",X"88",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"FA",X"B6",X"FF",X"F2",
		X"00",X"00",X"00",X"CC",X"E6",X"F7",X"FF",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"00",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"FF",X"FF",X"66",X"22",X"00",X"00",X"00",
		X"E6",X"FF",X"CC",X"45",X"4C",X"00",X"00",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"FE",X"B6",X"F2",X"F7",
		X"00",X"00",X"00",X"CC",X"E6",X"F7",X"F7",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FB",X"FF",X"EE",X"33",X"00",X"00",X"00",
		X"F7",X"CC",X"CC",X"77",X"CC",X"00",X"00",X"00",X"88",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"FA",X"B7",X"FE",X"F2",
		X"00",X"00",X"00",X"CC",X"E6",X"FF",X"F7",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"FF",X"FF",X"66",X"22",X"00",X"00",X"00",
		X"E6",X"FF",X"CC",X"45",X"4C",X"00",X"00",X"00",X"88",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"33",X"FE",X"B6",X"F2",X"FA",
		X"00",X"00",X"00",X"CC",X"F7",X"F7",X"F7",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"FB",X"FF",X"66",X"33",X"00",X"00",X"00",
		X"EE",X"CC",X"CC",X"67",X"CC",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"30",X"10",X"10",X"10",X"07",X"39",X"00",X"00",X"80",X"F0",X"A7",X"D7",X"C7",X"C7",
		X"03",X"37",X"4F",X"87",X"E1",X"AD",X"5E",X"3E",X"0E",X"EE",X"00",X"2E",X"2E",X"CC",X"E3",X"A1",
		X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A7",X"D3",X"70",X"54",X"00",X"00",X"00",X"00",
		X"3E",X"9E",X"F6",X"E1",X"98",X"44",X"33",X"00",X"B1",X"B3",X"80",X"C0",X"E2",X"40",X"EC",X"00",
		X"10",X"00",X"00",X"40",X"21",X"01",X"00",X"01",X"00",X"80",X"C0",X"05",X"3B",X"05",X"0A",X"01",
		X"00",X"31",X"34",X"3C",X"9E",X"4F",X"27",X"03",X"00",X"88",X"C4",X"88",X"00",X"00",X"78",X"48",
		X"00",X"03",X"D1",X"32",X"74",X"33",X"00",X"00",X"0A",X"00",X"00",X"01",X"80",X"8C",X"80",X"80",
		X"0A",X"04",X"0B",X"05",X"38",X"74",X"32",X"11",X"C4",X"C4",X"00",X"00",X"80",X"C8",X"A0",X"88",
		X"00",X"01",X"12",X"35",X"71",X"35",X"7B",X"7B",X"03",X"3C",X"F3",X"FF",X"DF",X"0F",X"88",X"8B",
		X"0C",X"C2",X"EF",X"FE",X"33",X"1D",X"AC",X"F8",X"00",X"00",X"0C",X"C2",X"CA",X"CA",X"CA",X"ED",
		X"7B",X"7B",X"7B",X"24",X"35",X"12",X"12",X"01",X"F9",X"BC",X"AD",X"DC",X"FF",X"FE",X"E1",X"0E",
		X"FD",X"4E",X"1D",X"F5",X"FF",X"F3",X"78",X"07",X"ED",X"ED",X"ED",X"CA",X"0C",X"84",X"0C",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"11",X"44",X"21",X"51",X"32",
		X"00",X"00",X"00",X"00",X"04",X"98",X"80",X"01",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"B3",X"4F",X"23",X"88",X"00",X"00",X"00",X"00",
		X"84",X"82",X"00",X"44",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"00",X"00",X"01",X"01",X"10",X"1E",
		X"3D",X"7B",X"EE",X"88",X"88",X"88",X"88",X"CD",X"FF",X"11",X"00",X"44",X"E8",X"00",X"00",X"80",
		X"00",X"00",X"00",X"08",X"08",X"09",X"8B",X"FE",X"00",X"00",X"04",X"04",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"11",X"00",X"00",X"20",X"08",X"4C",X"88",X"88",X"CB",X"ED",X"22",X"22",X"33",X"B3",X"5D",
		X"0C",X"08",X"00",X"00",X"00",X"00",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"11",X"00",X"00",X"00",X"01",X"01",X"00",
		X"98",X"99",X"88",X"CC",X"62",X"7B",X"33",X"11",X"00",X"00",X"20",X"24",X"16",X"00",X"CC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"01",X"02",X"06",X"0C",X"08",X"00",X"00",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"64",X"00",X"00",X"00",X"99",X"FF",X"44",X"11",X"33",X"33",X"77",X"EF",X"ED",X"8B",
		X"88",X"CA",X"CB",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"4A",X"04",X"04",X"06",X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"4C",X"8D",X"1A",
		X"00",X"04",X"27",X"47",X"07",X"0F",X"0F",X"0F",X"00",X"00",X"05",X"1A",X"25",X"1A",X"78",X"F7",
		X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"34",X"78",X"4B",X"0F",X"0F",X"0F",X"1F",X"1B",
		X"1F",X"0F",X"87",X"0F",X"0F",X"0F",X"0F",X"0F",X"88",X"07",X"0F",X"0F",X"6E",X"EE",X"0F",X"0F",
		X"00",X"00",X"04",X"4A",X"A5",X"5A",X"E1",X"F8",X"00",X"00",X"00",X"08",X"85",X"5A",X"A5",X"5A",
		X"00",X"01",X"06",X"0C",X"8C",X"08",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"76",X"3B",X"00",X"0F",X"0F",X"2F",X"6F",X"E1",X"F0",X"F8",X"30",X"1C",X"0E",X"0F",X"0F",
		X"84",X"4A",X"A5",X"D2",X"A5",X"96",X"A5",X"1E",X"00",X"06",X"44",X"08",X"00",X"08",X"00",X"00",
		X"00",X"00",X"23",X"26",X"09",X"00",X"00",X"00",X"1D",X"1B",X"1F",X"1B",X"07",X"0B",X"07",X"0B",
		X"0B",X"84",X"C3",X"F8",X"FC",X"7F",X"3F",X"1F",X"0D",X"12",X"2D",X"E1",X"C3",X"8F",X"8F",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"01",X"13",X"03",X"02",X"04",X"08",
		X"0F",X"0F",X"07",X"8A",X"00",X"00",X"00",X"00",X"78",X"0F",X"0D",X"0A",X"05",X"00",X"00",X"00",
		X"2F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4B",X"69",X"3C",X"78",X"7C",X"6F",X"CF",
		X"0F",X"2F",X"2F",X"0F",X"0F",X"0E",X"0C",X"0E",X"00",X"4E",X"44",X"08",X"00",X"00",X"00",X"00",
		X"87",X"0B",X"05",X"0A",X"05",X"02",X"22",X"01",X"0F",X"0F",X"0F",X"0A",X"00",X"00",X"00",X"00",
		X"26",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"04",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"8C",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"01",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"40",X"40",X"01",X"92",X"92",X"12",
		X"09",X"12",X"21",X"4B",X"87",X"3F",X"7F",X"7D",X"C3",X"0F",X"0F",X"7F",X"FF",X"DF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"20",X"00",X"08",X"C3",X"00",X"00",X"00",X"00",X"00",X"40",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3C",X"0F",X"0F",X"EF",X"FF",X"BF",X"FF",X"FF",X"09",X"84",X"48",X"2D",X"1E",X"CF",X"EF",X"EB",
		X"40",X"40",X"20",X"20",X"08",X"94",X"94",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"92",X"92",X"01",X"40",X"40",X"20",X"20",
		X"7D",X"7F",X"3F",X"87",X"4B",X"21",X"12",X"09",X"FF",X"FF",X"DF",X"FF",X"7F",X"0F",X"0F",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"3C",X"01",X"00",X"40",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"BF",X"FF",X"EF",X"0F",X"0F",X"3C",X"EB",X"EF",X"CF",X"1E",X"2D",X"48",X"84",X"09",
		X"84",X"94",X"94",X"08",X"20",X"20",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"08",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"30",X"40",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"88",
		X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"88",X"88",X"80",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"08",X"0C",X"0E",X"F0",X"0F",
		X"03",X"03",X"03",X"03",X"30",X"0F",X"80",X"0F",X"0E",X"0F",X"0F",X"0F",X"F0",X"0F",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"E0",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"0F",X"00",X"00",X"00",X"01",X"00",X"00",X"FF",X"0F",X"00",X"00",X"08",X"04",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"08",
		X"0F",X"0F",X"0F",X"0F",X"07",X"34",X"43",X"0C",X"00",X"0C",X"0E",X"0F",X"78",X"87",X"0C",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"48",X"87",X"0C",X"33",X"FF",X"00",X"00",X"00",X"00",X"08",X"22",X"33",X"CC",
		X"00",X"00",X"00",X"00",X"77",X"77",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"3C",X"C3",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"B7",X"3F",X"6F",X"06",X"00",X"00",X"00",X"00",X"FF",X"CF",X"0C",X"00",X"00",X"05",X"04",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"01",X"01",X"00",X"00",
		X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"1E",X"61",X"00",X"00",X"08",X"0F",X"3C",X"E1",X"86",X"19",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"83",X"0C",X"2A",X"77",X"EF",X"00",X"00",X"00",X"00",X"77",X"CC",X"8C",X"08",
		X"11",X"66",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3C",X"43",X"0E",X"08",X"00",
		X"06",X"19",X"B3",X"FF",X"07",X"02",X"00",X"00",X"77",X"FF",X"CF",X"0C",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8E",X"08",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"07",X"01",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"1E",X"2D",X"4A",X"84",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"84",X"08",X"33",X"77",X"EF",X"11",X"33",X"33",X"66",X"CC",X"8C",X"08",X"00",
		X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1E",X"10",
		X"1E",X"25",X"02",X"04",X"61",X"C3",X"84",X"08",X"19",X"13",X"37",X"6F",X"CE",X"8C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CE",X"8C",X"08",X"00",X"00",X"05",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"80",X"40",X"20",X"10",X"01",
		X"00",X"00",X"00",X"00",X"0F",X"50",X"1E",X"A1",X"00",X"00",X"00",X"20",X"48",X"80",X"08",X"CC",
		X"FF",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"11",X"10",X"20",X"40",X"80",X"00",X"00",
		X"C1",X"F5",X"FE",X"55",X"FF",X"00",X"00",X"00",X"CC",X"CC",X"88",X"80",X"C8",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"40",X"40",X"4B",X"50",X"4B",X"49",X"00",X"00",X"00",X"00",X"08",X"00",X"08",X"CC",
		X"FE",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"FB",X"FB",X"51",X"FB",X"40",X"40",X"00",X"F0",X"CC",X"88",X"00",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"17",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"EE",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"33",X"22",X"22",X"33",X"33",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"23",X"23",X"23",X"03",X"01",X"01",X"01",
		X"43",X"43",X"43",X"00",X"08",X"00",X"80",X"04",X"00",X"08",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"52",X"70",X"70",X"30",X"70",X"70",X"00",X"00",X"5A",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"5A",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"70",X"31",X"70",X"40",X"52",X"00",X"00",X"00",X"F0",X"F8",X"FF",X"00",X"5A",X"00",X"00",X"00",
		X"F3",X"E6",X"FF",X"10",X"5A",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"25",X"34",X"70",X"30",X"70",X"70",X"00",X"00",X"A5",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"A5",X"E1",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"E0",
		X"70",X"31",X"70",X"04",X"25",X"00",X"00",X"00",X"F0",X"F8",X"FF",X"00",X"A5",X"00",X"00",X"00",
		X"F3",X"E6",X"FF",X"01",X"A5",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"03",X"03",X"03",X"03",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",
		X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",
		X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"4B",X"00",X"00",X"FF",X"FF",X"48",X"48",X"48",X"48",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"03",X"03",X"03",X"30",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",
		X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",
		X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",
		X"4B",X"4B",X"4B",X"F0",X"00",X"00",X"FF",X"FF",X"48",X"48",X"48",X"C0",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"27",X"12",
		X"00",X"00",X"00",X"00",X"00",X"40",X"E4",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"72",X"20",X"00",X"00",X"00",X"00",X"00",
		X"84",X"4E",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"35",
		X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"12",X"01",X"00",X"00",X"00",X"00",X"00",
		X"CA",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"75",X"23",
		X"00",X"00",X"00",X"00",X"00",X"04",X"4A",X"8C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"13",X"25",X"02",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"EA",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"36",
		X"00",X"00",X"00",X"00",X"00",X"08",X"8C",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"36",X"13",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C6",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"57",X"73",X"EF",
		X"00",X"00",X"00",X"00",X"44",X"EE",X"FB",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"9B",X"55",X"33",X"00",X"00",X"00",X"00",
		X"F7",X"DF",X"C8",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"93",X"33",
		X"00",X"00",X"00",X"00",X"00",X"A8",X"C4",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"23",X"15",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"C9",X"88",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"04",X"00",X"33",
		X"00",X"00",X"00",X"00",X"10",X"08",X"88",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"27",X"11",X"10",X"08",X"00",X"00",X"00",X"00",
		X"44",X"88",X"20",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"04",X"00",X"00",X"00",X"08",X"22",X"45",X"31",
		X"00",X"00",X"00",X"00",X"00",X"04",X"64",X"88",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"11",X"04",X"64",X"00",X"00",X"00",X"00",X"00",
		X"AE",X"80",X"88",X"10",X"00",X"00",X"00",X"20",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"44",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"30",X"C3",X"96",X"F0",X"F0",
		X"00",X"00",X"00",X"C0",X"C3",X"F0",X"78",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"96",X"E1",X"F0",X"30",X"00",X"00",X"00",
		X"F0",X"E1",X"F0",X"F0",X"0C",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F4",X"72",X"30",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"F0",X"E1",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"F4",X"72",X"30",X"00",X"00",X"00",X"00",
		X"78",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"21",X"30",X"00",X"00",X"30",X"D2",X"5A",X"A5",X"5A",X"B4",
		X"00",X"00",X"C0",X"B4",X"A5",X"5A",X"A5",X"D2",X"00",X"00",X"00",X"00",X"80",X"80",X"48",X"C0",
		X"30",X"21",X"10",X"10",X"00",X"00",X"00",X"00",X"B4",X"5A",X"AD",X"5E",X"D2",X"30",X"00",X"00",
		X"D2",X"A5",X"5A",X"A5",X"B4",X"C0",X"00",X"00",X"C0",X"48",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"30",X"40",X"40",X"00",X"00",X"00",X"45",X"00",X"11",X"00",X"01",X"00",X"01",X"00",X"04",
		X"00",X"88",X"00",X"08",X"00",X"08",X"00",X"02",X"00",X"C0",X"20",X"20",X"00",X"00",X"00",X"2A",
		X"45",X"00",X"00",X"00",X"40",X"40",X"30",X"00",X"04",X"00",X"01",X"00",X"01",X"00",X"11",X"00",
		X"02",X"00",X"08",X"00",X"08",X"00",X"88",X"00",X"2A",X"00",X"00",X"00",X"20",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"AE",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"A4",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AE",X"4E",X"AE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A4",X"4A",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"44",X"26",X"44",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"40",X"24",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"11",X"00",X"02",X"00",X"00",X"00",X"08",X"44",X"00",X"02",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"08",X"40",X"00",X"20",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"02",X"00",X"11",X"00",X"00",
		X"08",X"00",X"11",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"01",X"00",X"00",X"20",
		X"00",X"00",X"04",X"00",X"00",X"10",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"52",X"25",
		X"00",X"00",X"00",X"00",X"00",X"48",X"A4",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"52",X"21",X"00",X"00",X"00",X"00",X"00",
		X"4A",X"A4",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"12",X"25",
		X"00",X"00",X"00",X"00",X"00",X"08",X"84",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"12",X"01",X"00",X"00",X"00",X"00",X"00",
		X"4A",X"84",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"70",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"06",X"04",X"04",X"07",X"03",X"00",X"00",X"06",X"0F",X"09",X"09",X"0B",X"02",X"00",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",
		X"00",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"0F",
		X"00",X"00",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"88",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"01",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"88",X"00",X"00",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"2E",X"2E",X"2E",X"2E",X"2E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"34",X"34",X"34",X"34",X"34",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",
		X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"34",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"34",X"34",X"34",X"34",X"34",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"88",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"88",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"88",X"88",X"CC",X"CC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"03",X"03",X"03",X"03",X"03",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"88",X"00",X"00",
		X"FF",X"FF",X"EE",X"88",X"00",X"00",X"00",X"00",X"CC",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",
		X"EE",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"01",
		X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"03",X"03",
		X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"05",X"03",X"07",
		X"00",X"00",X"00",X"00",X"02",X"04",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"02",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"09",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"05",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"04",X"0B",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"05",X"03",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"01",X"01",X"00",X"00",X"00",X"00",
		X"08",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0B",X"07",
		X"00",X"00",X"00",X"08",X"08",X"04",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"02",X"02",X"00",X"00",X"00",X"00",
		X"0B",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0F",X"03",
		X"00",X"00",X"00",X"04",X"08",X"08",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"02",X"04",X"00",X"00",X"00",X"00",
		X"0E",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"07",X"03",
		X"00",X"00",X"00",X"00",X"04",X"08",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"F0",X"F0",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",
		X"90",X"E3",X"F1",X"F3",X"F7",X"F7",X"F0",X"F2",X"3F",X"8F",X"8F",X"EE",X"FF",X"FF",X"F4",X"F4",
		X"0E",X"0F",X"8F",X"31",X"9F",X"EF",X"F1",X"F0",X"00",X"08",X"0C",X"0C",X"0E",X"4E",X"AC",X"EE",
		X"F2",X"F3",X"F0",X"F7",X"F3",X"F1",X"70",X"F0",X"F4",X"F4",X"F0",X"F8",X"F8",X"F8",X"70",X"F0",
		X"F0",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"FC",X"F0",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"71",X"70",X"71",X"71",X"70",X"70",X"70",X"F7",X"7F",X"FF",X"F8",X"FF",X"F7",X"F2",X"F2",
		X"FE",X"7F",X"FF",X"F3",X"FF",X"FF",X"C3",X"01",X"F0",X"78",X"F8",X"FC",X"CC",X"0C",X"08",X"0C",
		X"70",X"71",X"40",X"01",X"F1",X"E0",X"E0",X"E0",X"C2",X"0A",X"00",X"70",X"F0",X"F0",X"F0",X"F0",
		X"01",X"03",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"0C",X"78",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"70",X"C0",X"00",X"00",X"00",X"00",X"00",X"C3",X"07",X"07",X"00",X"07",X"09",X"01",X"70",
		X"F8",X"FC",X"7C",X"36",X"1E",X"0E",X"7C",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"80",X"F0",X"F5",X"F0",X"F0",X"E0",X"90",X"00",X"B0",
		X"FE",X"FC",X"E0",X"A0",X"20",X"40",X"00",X"00",X"E0",X"A0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"01",X"07",X"01",X"01",
		X"08",X"08",X"08",X"08",X"0C",X"0C",X"08",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"08",X"00",X"00",X"00",X"10",X"30",X"70",X"00",X"10",X"30",X"70",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"50",X"01",X"13",X"33",X"77",X"F7",X"F7",X"F7",X"F7",
		X"FC",X"FE",X"FE",X"EE",X"FE",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F3",X"71",X"B7",X"D3",X"C1",X"E1",X"B0",X"10",
		X"FF",X"FF",X"EF",X"DE",X"BE",X"6E",X"1E",X"94",X"F0",X"70",X"F0",X"B0",X"70",X"D0",X"90",X"20",
		X"00",X"01",X"01",X"03",X"03",X"13",X"33",X"73",X"07",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"DF",X"EF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"F0",X"78",X"08",X"CE",X"EA",X"FA",
		X"93",X"E1",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"3F",X"81",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"6D",X"01",X"81",X"E1",X"F0",X"F0",X"BA",X"6A",X"DE",X"B8",X"08",X"00",X"80",X"F0",
		X"E0",X"C1",X"83",X"13",X"37",X"77",X"F0",X"F0",X"37",X"7F",X"FF",X"FF",X"FF",X"FC",X"F1",X"F3",
		X"CF",X"CF",X"EF",X"FF",X"FF",X"F6",X"FA",X"FC",X"40",X"1C",X"58",X"0C",X"9E",X"C0",X"CF",X"CF",
		X"F0",X"F0",X"B0",X"10",X"40",X"10",X"90",X"00",X"F3",X"F1",X"F0",X"F0",X"F0",X"70",X"10",X"00",
		X"FC",X"F8",X"F0",X"F1",X"E1",X"C1",X"80",X"00",X"EF",X"CF",X"80",X"0E",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"40",X"20",X"20",X"10",X"50",X"33",X"30",X"F0",X"F0",X"F1",
		X"F0",X"F0",X"F0",X"FC",X"D2",X"C1",X"C0",X"88",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"38",
		X"00",X"90",X"30",X"30",X"B0",X"70",X"70",X"F0",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"88",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",X"10",X"30",X"30",X"70",X"50",
		X"F0",X"F0",X"F0",X"F0",X"F1",X"F0",X"F2",X"F0",X"70",X"F0",X"F3",X"FC",X"F3",X"F0",X"F0",X"F1",
		X"00",X"C0",X"8C",X"D3",X"EC",X"E2",X"E1",X"F8",X"00",X"00",X"00",X"00",X"08",X"40",X"04",X"48",
		X"F0",X"F0",X"F0",X"B0",X"F0",X"F0",X"F0",X"B0",X"F1",X"F4",X"F3",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F8",X"F2",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",X"48",X"98",X"80",X"C0",X"D0",X"E0",X"E0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",X"81",
		X"00",X"00",X"10",X"10",X"30",X"31",X"72",X"79",X"F0",X"F0",X"F0",X"D0",X"F0",X"F8",X"F4",X"D0",
		X"F0",X"F0",X"F0",X"F0",X"10",X"F0",X"F0",X"F0",X"87",X"82",X"90",X"10",X"30",X"30",X"70",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F8",X"F0",X"F0",X"D0",X"F0",X"F0",X"F0",X"00",
		X"F0",X"F0",X"F0",X"B0",X"F0",X"F0",X"F1",X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F4",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F9",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"FC",
		X"F0",X"F0",X"F0",X"B0",X"F0",X"F0",X"F0",X"00",X"F6",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"10",X"F0",X"F0",X"F0",X"F0",X"80",X"F0",X"F0",X"F0",
		X"00",X"00",X"10",X"30",X"70",X"70",X"30",X"70",X"00",X"10",X"B0",X"F0",X"F0",X"F0",X"F7",X"F0",
		X"10",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"D0",X"D0",X"D0",X"F0",X"F0",X"F0",X"F4",
		X"F1",X"F0",X"30",X"80",X"C0",X"F0",X"80",X"F0",X"F2",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",
		X"F4",X"F0",X"F0",X"F0",X"C0",X"80",X"C0",X"C0",X"FC",X"A0",X"00",X"00",X"30",X"70",X"F0",X"F0",
		X"F0",X"B0",X"A0",X"A0",X"E0",X"F0",X"F3",X"F3",X"00",X"E0",X"E0",X"C0",X"C0",X"8F",X"8E",X"1C",
		X"00",X"30",X"30",X"70",X"70",X"FF",X"F1",X"E1",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"8C",X"1C",
		X"F0",X"50",X"00",X"00",X"C0",X"E0",X"F0",X"F0",X"0F",X"80",X"C2",X"E0",X"30",X"10",X"30",X"10",
		X"8F",X"00",X"14",X"70",X"E0",X"F0",X"F0",X"F0",X"00",X"68",X"E0",X"E0",X"30",X"F0",X"10",X"F0",
		X"F0",X"80",X"F0",X"F0",X"F0",X"F1",X"F3",X"F2",X"F0",X"F0",X"F0",X"F0",X"F7",X"FF",X"F4",X"F8",
		X"C0",X"C0",X"80",X"80",X"8E",X"CF",X"E3",X"F1",X"F0",X"F0",X"70",X"30",X"00",X"08",X"2C",X"FC",
		X"73",X"01",X"10",X"30",X"10",X"00",X"00",X"00",X"F5",X"F8",X"F7",X"F0",X"D0",X"90",X"10",X"00",
		X"FB",X"F1",X"FE",X"F0",X"F0",X"F0",X"F0",X"F0",X"FC",X"F8",X"F0",X"F0",X"D0",X"D0",X"D0",X"F0",
		X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"50",X"F0",X"10",X"30",X"10",X"30",X"F0",X"F0",X"F4",X"F1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"10",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"E0",X"A0",X"A0",X"B0",X"F0",X"F1",X"F0",X"F0",X"F0",X"70",X"70",X"30",X"30",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"00",X"E0",X"C0",X"80",X"C0",X"C0",X"80",X"00",X"00",
		X"F0",X"F0",X"F0",X"10",X"F3",X"F0",X"F2",X"F2",X"00",X"70",X"30",X"10",X"06",X"80",X"88",X"80",
		X"00",X"F0",X"F1",X"F9",X"FF",X"7B",X"33",X"13",X"00",X"F0",X"F8",X"FC",X"D0",X"F8",X"FC",X"FF",
		X"F2",X"F2",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"88",X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",
		X"03",X"00",X"09",X"08",X"00",X"00",X"00",X"00",X"DC",X"78",X"38",X"10",X"08",X"08",X"00",X"00",
		X"00",X"F0",X"F0",X"F0",X"B0",X"F3",X"F1",X"F1",X"00",X"F0",X"F0",X"F0",X"F0",X"FE",X"FE",X"FF",
		X"10",X"F0",X"F1",X"F9",X"F9",X"FF",X"F1",X"F1",X"F0",X"F0",X"F8",X"8C",X"FC",X"F0",X"FC",X"FC",
		X"B1",X"F1",X"F3",X"F0",X"B0",X"70",X"30",X"10",X"F0",X"F0",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F1",X"F0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"FC",X"F8",X"F0",X"F0",X"F8",X"F8",X"F0",X"F0",
		X"F0",X"70",X"F0",X"30",X"30",X"90",X"10",X"C1",X"E0",X"F0",X"F0",X"F0",X"F0",X"F6",X"F3",X"FC",
		X"00",X"02",X"07",X"0F",X"0F",X"8C",X"8A",X"87",X"00",X"00",X"08",X"0C",X"0C",X"00",X"00",X"00",
		X"41",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"F0",X"73",X"76",X"30",X"B0",X"50",X"10",X"00",
		X"87",X"CA",X"C8",X"D8",X"C0",X"E0",X"E0",X"F0",X"30",X"70",X"F0",X"F0",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"F0",X"70",X"30",X"70",X"70",X"71",X"F3",X"F3",
		X"F0",X"F2",X"F7",X"FF",X"FF",X"F8",X"FC",X"F8",X"F0",X"E0",X"E8",X"CC",X"DC",X"80",X"80",X"40",
		X"C0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"F3",X"F1",X"F0",X"F0",X"30",X"30",X"30",X"70",
		X"F8",X"E0",X"E0",X"C8",X"D0",X"80",X"80",X"40",X"60",X"00",X"00",X"80",X"08",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"00",X"10",X"30",X"70",X"F0",X"F3",X"F3",X"F0",
		X"40",X"00",X"E1",X"F9",X"F9",X"FE",X"F4",X"F4",X"00",X"90",X"58",X"0C",X"8C",X"C0",X"F0",X"F0",
		X"70",X"B0",X"30",X"10",X"A0",X"80",X"10",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"70",
		X"F4",X"F4",X"FE",X"F8",X"F0",X"F0",X"E0",X"C0",X"F0",X"F0",X"E0",X"C0",X"88",X"18",X"30",X"70",
		X"70",X"90",X"30",X"60",X"D0",X"31",X"23",X"90",X"F0",X"F0",X"70",X"D0",X"B0",X"7E",X"FE",X"F0",
		X"F0",X"F0",X"F1",X"F9",X"F9",X"FF",X"FF",X"F0",X"70",X"70",X"78",X"7C",X"7C",X"FC",X"F8",X"F8",
		X"C0",X"60",X"30",X"70",X"F0",X"F0",X"F0",X"F0",X"FE",X"70",X"B0",X"D0",X"E0",X"F0",X"F0",X"F0",
		X"F7",X"F8",X"FB",X"F8",X"E0",X"40",X"80",X"00",X"E8",X"C8",X"8C",X"00",X"08",X"08",X"00",X"00",
		X"00",X"80",X"80",X"C0",X"C0",X"E1",X"E2",X"F0",X"D0",X"B0",X"60",X"D0",X"30",X"7E",X"70",X"30",
		X"80",X"C0",X"E1",X"E9",X"F9",X"FF",X"F8",X"F0",X"F0",X"F0",X"F8",X"7C",X"7C",X"B0",X"DC",X"FC",
		X"F0",X"F0",X"F1",X"F0",X"00",X"F0",X"F0",X"F0",X"30",X"B0",X"98",X"D0",X"50",X"E0",X"E0",X"F0",
		X"F0",X"F8",X"F8",X"F8",X"E0",X"C0",X"80",X"00",X"EC",X"CC",X"80",X"00",X"08",X"08",X"00",X"00",
		X"F0",X"F7",X"F3",X"F1",X"E0",X"C0",X"80",X"00",X"E0",X"CF",X"8F",X"0F",X"0F",X"07",X"03",X"01",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"0E",X"06",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"17",X"21",X"10",X"70",X"00",X"00",X"40",X"23",X"10",X"78",X"F6",X"F1",
		X"10",X"80",X"1F",X"7F",X"FF",X"F0",X"FF",X"FF",X"10",X"70",X"F0",X"FE",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"F6",X"F0",X"F0",X"F0",X"C0",X"E0",X"F0",X"F0",
		X"F7",X"F3",X"FF",X"CF",X"08",X"00",X"00",X"00",X"F8",X"F8",X"B8",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F7",X"F0",X"F0",X"F0",X"F0",X"F1",X"F7",X"F1",X"F0",X"FF",X"F1",
		X"F0",X"F6",X"FF",X"FF",X"F8",X"F3",X"FF",X"FF",X"70",X"70",X"7C",X"F0",X"F0",X"E0",X"E0",X"E0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"20",X"10",X"F4",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",
		X"F3",X"F3",X"FF",X"F6",X"F0",X"F0",X"E0",X"F0",X"E8",X"E8",X"E8",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"FF",X"F0",X"F0",X"F0",X"E3",X"C7",X"87",X"00",X"E8",X"F7",
		X"00",X"0F",X"0F",X"0C",X"00",X"06",X"0F",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"70",X"10",X"20",X"10",X"00",X"00",X"00",X"00",X"F0",X"F6",X"70",X"10",X"40",X"00",X"00",X"00",
		X"F3",X"F3",X"F7",X"F6",X"70",X"90",X"80",X"10",X"E8",X"F8",X"F0",X"F0",X"F0",X"F0",X"70",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"60",X"33",X"17",X"0F",X"00",X"00",X"0F",
		X"F0",X"EE",X"FC",X"F8",X"F2",X"77",X"3F",X"1F",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E8",
		X"00",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"07",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"01",X"03",X"07",X"E2",X"F0",X"F0",X"F0",X"F0",X"E8",X"60",X"20",X"00",X"F0",X"70",X"70",X"70",
		X"F0",X"F0",X"F0",X"00",X"F0",X"F1",X"F0",X"F0",X"F0",X"E3",X"F7",X"5F",X"FE",X"B0",X"F1",X"77",
		X"04",X"0C",X"88",X"C0",X"E6",X"FF",X"FF",X"FD",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"E8",
		X"FF",X"E0",X"E0",X"D0",X"C0",X"90",X"90",X"20",X"78",X"F7",X"70",X"B0",X"D0",X"60",X"B0",X"D0",
		X"F1",X"F3",X"F6",X"F0",X"F0",X"E0",X"C0",X"80",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"30",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"07",X"07",X"0F",X"0E",X"0C",X"01",X"03",
		X"08",X"08",X"00",X"00",X"06",X"0F",X"0F",X"0D",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"01",X"87",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"0E",X"00",X"00",X"02",X"00",X"80",X"C0",X"E0",
		X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"20",X"00",X"31",X"B1",X"11",X"00",X"71",X"B7",X"7E",X"FE",X"FC",X"FD",X"F1",X"F1",
		X"C0",X"E0",X"F0",X"F8",X"FF",X"FF",X"FD",X"F9",X"10",X"00",X"00",X"80",X"C0",X"E8",X"F8",X"F8",
		X"00",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"76",X"39",X"12",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"F3",X"F0",X"F0",X"70",X"20",X"40",X"10",X"F0",X"F0",X"D0",X"80",X"40",X"90",X"30",X"00",
		X"F0",X"F0",X"70",X"31",X"12",X"30",X"71",X"F1",X"F1",X"F3",X"FF",X"F3",X"F0",X"F0",X"F0",X"F0",
		X"0C",X"8F",X"8F",X"CF",X"E3",X"F1",X"F0",X"F0",X"00",X"08",X"0C",X"0E",X"0E",X"0E",X"8F",X"CF",
		X"D1",X"61",X"B0",X"D0",X"60",X"00",X"10",X"70",X"F0",X"F0",X"70",X"A0",X"93",X"70",X"F0",X"F0",
		X"F0",X"F0",X"D0",X"70",X"FC",X"F1",X"F0",X"F0",X"DF",X"7E",X"F4",X"74",X"78",X"70",X"70",X"70",
		X"10",X"01",X"02",X"04",X"00",X"01",X"43",X"00",X"FC",X"03",X"0C",X"0C",X"00",X"FE",X"77",X"0B",
		X"E0",X"00",X"0C",X"0B",X"09",X"8F",X"FC",X"8E",X"00",X"00",X"00",X"00",X"0C",X"0C",X"C0",X"60",
		X"00",X"30",X"30",X"00",X"00",X"00",X"10",X"00",X"07",X"81",X"00",X"00",X"1C",X"3C",X"F0",X"00",
		X"8E",X"00",X"0F",X"0F",X"0C",X"00",X"E0",X"00",X"60",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"03",X"03",X"04",X"00",X"73",X"02",X"0C",X"BB",X"0C",X"7C",X"78",X"7F",X"FF",X"03",
		X"00",X"60",X"0C",X"0A",X"09",X"8F",X"FE",X"8E",X"00",X"00",X"00",X"00",X"08",X"0E",X"C0",X"60",
		X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"0B",X"01",X"10",X"38",X"0C",X"BC",X"08",X"00",
		X"EE",X"81",X"0F",X"0E",X"0C",X"60",X"00",X"00",X"60",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"11",X"30",X"70",X"00",X"07",X"0A",X"0E",X"76",X"F2",X"F7",X"FF",X"0F",
		X"00",X"08",X"0C",X"8A",X"E9",X"EF",X"F8",X"88",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"60",
		X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"37",X"B2",X"B8",X"02",X"36",X"06",X"02",X"00",
		X"08",X"00",X"6F",X"0E",X"0C",X"08",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"10",X"01",X"01",X"01",X"01",X"31",X"B3",X"73",X"F3",
		X"08",X"08",X"08",X"08",X"08",X"08",X"FC",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",
		X"00",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"03",X"B2",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"01",X"70",X"00",X"00",X"01",X"03",X"77",X"FF",X"3F",X"B3",X"33",
		X"0E",X"0F",X"0F",X"8F",X"EF",X"0F",X"7F",X"0F",X"00",X"00",X"00",X"08",X"08",X"00",X"C0",X"60",
		X"00",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"0F",X"37",X"33",X"01",X"00",X"00",
		X"80",X"8D",X"EF",X"0F",X"0F",X"0F",X"0F",X"06",X"60",X"00",X"00",X"08",X"08",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"31",X"37",X"70",X"00",X"70",X"F0",X"73",X"77",X"0F",X"FF",X"F7",X"07",
		X"03",X"ED",X"8B",X"0B",X"0D",X"8F",X"FF",X"8F",X"00",X"08",X"0C",X"0C",X"0E",X"0C",X"CC",X"6C",
		X"00",X"03",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"0F",X"0F",X"17",X"33",X"F0",X"30",X"10",
		X"80",X"8C",X"0F",X"0D",X"0B",X"EB",X"01",X"01",X"60",X"04",X"0E",X"0E",X"0C",X"0C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"13",X"07",X"10",X"30",X"00",X"00",X"33",X"0F",X"3F",X"FF",X"A0",X"93",
		X"03",X"0C",X"C3",X"03",X"58",X"C8",X"A3",X"DF",X"00",X"08",X"04",X"02",X"81",X"82",X"4C",X"4E",
		X"10",X"10",X"03",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FF",X"7F",X"73",X"00",X"00",X"00",
		X"B0",X"E0",X"E8",X"F8",X"E3",X"03",X"00",X"00",X"C2",X"84",X"02",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"10",X"00",X"10",X"30",X"07",X"07",X"37",X"07",X"34",X"F3",X"AF",X"9F",
		X"0F",X"0F",X"CF",X"0F",X"13",X"CD",X"AE",X"DE",X"00",X"08",X"0C",X"0E",X"8F",X"8F",X"4F",X"4F",
		X"10",X"10",X"00",X"00",X"03",X"01",X"00",X"00",X"EF",X"FF",X"F7",X"73",X"70",X"00",X"00",X"00",
		X"BE",X"EE",X"ED",X"FC",X"E0",X"00",X"00",X"00",X"CF",X"8F",X"0F",X"80",X"0C",X"08",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"04",X"01",X"00",X"03",X"0F",X"00",X"00",X"03",X"03",
		X"08",X"08",X"0C",X"0F",X"07",X"03",X"CD",X"CC",X"00",X"00",X"0C",X"0C",X"08",X"08",X"0C",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"01",X"00",X"08",X"00",X"0D",X"0C",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"07",X"03",X"0F",X"00",X"00",X"13",X"03",
		X"00",X"01",X"0F",X"0F",X"77",X"F3",X"FD",X"EC",X"00",X"08",X"08",X"00",X"08",X"0B",X"0F",X"0E",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"0C",X"00",X"00",X"01",X"00",X"02",X"00",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"06",X"07",X"0F",X"00",X"10",X"13",X"03",
		X"02",X"07",X"1E",X"3F",X"F7",X"F3",X"FD",X"FC",X"00",X"00",X"C0",X"C0",X"CA",X"8F",X"0E",X"0C",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"02",X"00",
		X"6C",X"0C",X"00",X"00",X"01",X"02",X"00",X"00",X"0C",X"0E",X"0E",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"0F",X"1F",X"30",X"10",X"13",X"03",
		X"06",X"1E",X"7C",X"FF",X"F7",X"F3",X"FD",X"FC",X"70",X"F0",X"F0",X"E6",X"EE",X"CC",X"CC",X"8C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"01",X"00",
		X"7C",X"1C",X"00",X"00",X"01",X"01",X"00",X"00",X"8E",X"0E",X"0A",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"08",X"00",X"10",X"70",X"F0",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"01",
		X"00",X"0E",X"0F",X"0F",X"07",X"03",X"01",X"08",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"70",X"F0",X"F0",X"E0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"17",X"3F",X"30",X"10",X"11",X"03",
		X"30",X"7E",X"FF",X"FF",X"F7",X"F3",X"F9",X"FC",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"EE",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"18",X"00",X"00",X"01",X"00",X"00",X"00",X"CE",X"8C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"80",X"01",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"03",X"07",X"07",
		X"00",X"0E",X"0F",X"0F",X"07",X"0F",X"0F",X"0E",X"00",X"00",X"08",X"0C",X"0C",X"0E",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"0C",X"00",X"01",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"0F",X"0F",X"07",X"03",X"09",X"0C",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"01",X"03",X"07",X"00",X"00",X"00",
		X"07",X"03",X"09",X"0C",X"0E",X"00",X"10",X"70",X"0C",X"0C",X"0C",X"1C",X"34",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"07",X"07",X"0B",X"0B",X"0D",X"0D",X"3E",
		X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0E",X"89",X"00",X"00",X"00",X"0C",X"0C",X"08",X"04",X"0C",
		X"03",X"32",X"70",X"F1",X"F0",X"F0",X"F0",X"F0",X"F8",X"F1",X"F7",X"FF",X"E7",X"E0",X"C0",X"80",
		X"87",X"83",X"03",X"09",X"09",X"0C",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"10",X"72",X"36",X"3E",X"1E",X"1E",X"00",
		X"78",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"EF",
		X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"00",X"00",
		X"70",X"17",X"07",X"07",X"06",X"04",X"00",X"00",X"E0",X"CC",X"48",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"E0",X"E0",X"C1",X"80",X"82",X"03",X"80",X"00",X"00",X"07",X"0F",X"07",X"01",X"08",
		X"00",X"00",X"0D",X"0B",X"0B",X"07",X"07",X"0F",X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",X"0C",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"0E",X"0C",X"0C",X"09",X"09",X"03",X"00",X"00",
		X"07",X"09",X"0E",X"0F",X"0E",X"00",X"00",X"00",X"0E",X"0E",X"06",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"02",X"00",X"00",X"06",X"0E",
		X"00",X"08",X"0C",X"0E",X"07",X"01",X"06",X"07",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"0B",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"06",X"02",X"00",X"00",X"10",
		X"07",X"07",X"07",X"06",X"04",X"30",X"70",X"F0",X"0C",X"08",X"30",X"70",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"13",X"00",X"00",X"00",X"02",X"16",X"3E",X"FE",X"FE",
		X"00",X"18",X"3C",X"FE",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"E0",X"C8",X"8C",X"8F",
		X"71",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FE",X"F6",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"FF",X"EF",X"CE",X"C8",X"80",X"00",X"00",X"00",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"30",X"70",X"72",X"36",X"3E",X"1E",X"1E",X"00",
		X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"60",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C1",X"83",X"C0",X"C0",X"80",X"02",X"06",X"0E",X"0E",X"0E",
		X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"06",X"00",X"00",X"02",X"00",X"00",X"00",
		X"0F",X"0F",X"0E",X"08",X"04",X"00",X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"20",X"20",X"20",X"F6",X"2E",
		X"00",X"00",X"00",X"40",X"58",X"4E",X"FF",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"8E",
		X"03",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"FE",X"2E",X"B6",X"32",X"00",X"00",X"00",
		X"5F",X"FF",X"7F",X"FF",X"CE",X"0C",X"08",X"00",X"8F",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"60",X"20",X"20",X"70",
		X"00",X"00",X"00",X"C0",X"70",X"40",X"40",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"10",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"A0",X"20",X"20",X"F8",X"34",X"02",X"00",X"00",
		X"50",X"77",X"77",X"F7",X"C6",X"04",X"00",X"00",X"80",X"8C",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"10",X"01",X"01",X"01",X"20",X"20",X"33",X"E7",X"27",
		X"08",X"0E",X"0E",X"4F",X"53",X"CD",X"7E",X"5E",X"00",X"00",X"00",X"00",X"08",X"0E",X"8E",X"8F",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"27",X"E7",X"33",X"B0",X"30",X"00",X"00",X"00",
		X"5E",X"7E",X"FC",X"F0",X"C0",X"06",X"06",X"00",X"87",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"1A",X"05",X"0A",X"05",X"3A",X"E5",X"2A",X"25",X"AA",
		X"05",X"0A",X"05",X"CA",X"75",X"4A",X"45",X"5A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"8A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"75",X"2A",X"25",X"FA",X"35",X"0A",X"05",X"0A",
		X"F5",X"7A",X"75",X"FA",X"C5",X"0A",X"05",X"0A",X"85",X"8A",X"05",X"0A",X"05",X"0A",X"05",X"0A",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"07",X"03",X"05",X"0B",X"08",X"00",X"00",X"00",
		X"0F",X"0E",X"0F",X"0F",X"07",X"03",X"01",X"00",X"08",X"0C",X"06",X"0B",X"0D",X"0F",X"0F",X"0F",
		X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"00",X"00",
		X"00",X"00",X"00",X"01",X"07",X"06",X"00",X"00",X"0F",X"0B",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"07",X"03",X"05",X"0B",X"08",X"00",X"00",X"01",
		X"0F",X"0E",X"0F",X"0F",X"07",X"03",X"01",X"08",X"08",X"0C",X"06",X"0B",X"0D",X"0F",X"0F",X"0F",
		X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"08",X"04",X"00",X"00",
		X"08",X"00",X"00",X"01",X"07",X"06",X"00",X"00",X"0F",X"0B",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"07",X"03",X"05",X"0B",X"08",X"00",X"01",X"03",
		X"0F",X"0E",X"0F",X"0F",X"07",X"03",X"09",X"0C",X"08",X"0C",X"06",X"0B",X"0D",X"0F",X"0F",X"0F",
		X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"08",X"04",X"00",X"00",
		X"0C",X"08",X"00",X"01",X"07",X"06",X"00",X"00",X"0F",X"0B",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"07",X"03",X"05",X"0B",X"08",X"01",X"03",X"07",
		X"0F",X"0E",X"0F",X"0F",X"07",X"0B",X"0D",X"0E",X"08",X"0C",X"06",X"0B",X"0D",X"0F",X"0F",X"0F",
		X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"08",X"04",X"00",X"00",
		X"0E",X"0C",X"08",X"01",X"07",X"06",X"00",X"00",X"0F",X"0B",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"7F",X"FA",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0A",
		X"30",X"70",X"F0",X"70",X"1F",X"1F",X"0F",X"0A",X"E0",X"E0",X"F0",X"E0",X"EF",X"CF",X"FF",X"7A",
		X"F5",X"7A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"85",X"EA",X"15",X"0A",X"05",X"0A",
		X"05",X"0A",X"05",X"0A",X"E5",X"FA",X"75",X"3A",X"75",X"7A",X"45",X"2A",X"25",X"BA",X"C5",X"EA",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"1A",X"00",X"00",X"00",X"30",X"CF",X"FF",X"FF",X"FA",
		X"00",X"10",X"30",X"F0",X"7F",X"BF",X"DF",X"FA",X"00",X"80",X"C0",X"80",X"0C",X"0E",X"0F",X"0A",
		X"15",X"1A",X"15",X"3A",X"75",X"3A",X"05",X"0A",X"F5",X"FA",X"F5",X"FA",X"F5",X"8A",X"05",X"0A",
		X"F5",X"FA",X"E5",X"EA",X"F5",X"7A",X"35",X"1A",X"C5",X"CA",X"05",X"0A",X"05",X"8A",X"85",X"8A",
		X"05",X"0A",X"05",X"0A",X"45",X"0A",X"05",X"1A",X"05",X"0A",X"45",X"0A",X"05",X"DA",X"75",X"7A",
		X"05",X"0A",X"65",X"0A",X"C5",X"2A",X"B5",X"FA",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"2A",
		X"05",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"F5",X"F0",X"67",X"30",X"00",X"40",X"00",X"00",
		X"F5",X"70",X"29",X"A0",X"00",X"C0",X"00",X"00",X"05",X"00",X"4E",X"00",X"80",X"00",X"00",X"00",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"15",X"0A",X"05",X"0A",X"05",X"1A",X"45",X"AA",X"25",X"0A",
		X"05",X"0A",X"05",X"0A",X"05",X"0A",X"25",X"8A",X"05",X"0A",X"25",X"0A",X"05",X"0A",X"05",X"0A",
		X"05",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"A5",X"A0",X"89",X"00",X"00",X"00",X"00",X"00",
		X"05",X"80",X"0E",X"40",X"00",X"20",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"10",
		X"00",X"00",X"0F",X"07",X"03",X"01",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"30",X"10",X"10",X"08",X"0C",X"00",X"00",X"00",X"E0",
		X"80",X"81",X"13",X"77",X"7F",X"7F",X"7F",X"2F",X"0F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"8F",X"8F",X"93",X"30",X"00",X"08",X"0E",X"4F",X"4F",X"8F",X"8F",X"07",X"01",
		X"00",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",
		X"0F",X"EF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"00",X"38",X"1C",X"CE",X"CF",X"CF",X"CF",X"6F",
		X"CF",X"87",X"07",X"03",X"03",X"03",X"41",X"01",X"0C",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"7F",X"7F",X"7F",X"3F",X"17",X"83",X"01",X"00",X"FF",X"FF",X"FF",X"BF",X"9F",X"FF",X"3F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"0F",X"FF",X"EF",X"CF",X"CF",X"8E",X"0C",X"18",X"30",
		X"01",X"21",X"33",X"03",X"03",X"01",X"00",X"80",X"0F",X"0F",X"CF",X"0F",X"0C",X"0C",X"0C",X"04",
		X"00",X"A0",X"40",X"40",X"60",X"20",X"20",X"00",X"10",X"00",X"08",X"0C",X"08",X"08",X"00",X"00",
		X"C0",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"07",X"03",X"C1",X"60",X"20",X"10",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"87",X"D3",X"A1",X"40",
		X"0F",X"4F",X"6F",X"4F",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",X"AF",X"5F",X"AF",X"5F",X"0F",X"0F",
		X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"87",X"7F",X"8F",X"0F",X"0F",X"7F",X"FF",X"0F",X"0F",
		X"0F",X"0F",X"AF",X"5F",X"AF",X"5F",X"2F",X"0F",X"0F",X"0F",X"0F",X"4F",X"AF",X"5F",X"AF",X"5F",
		X"0F",X"1F",X"6F",X"CF",X"CF",X"0F",X"8F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"8F",X"4F",X"FF",X"0F",X"0F",X"2F",X"6F",X"2F",X"1F",X"0F",X"CF",X"2F",X"1F",X"0F",X"0F",
		X"AF",X"5F",X"AF",X"5F",X"2F",X"1F",X"2F",X"1F",X"0F",X"6F",X"CF",X"0F",X"8F",X"0F",X"8F",X"0F",
		X"00",X"10",X"20",X"70",X"80",X"00",X"00",X"00",X"20",X"40",X"20",X"40",X"A0",X"50",X"A0",X"50",
		X"C7",X"77",X"37",X"07",X"07",X"07",X"87",X"40",X"3F",X"EF",X"DF",X"1F",X"2F",X"4F",X"4F",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"30",X"30",X"20",X"40",X"80",
		X"A0",X"50",X"A0",X"90",X"00",X"00",X"00",X"00",X"80",X"50",X"A0",X"50",X"80",X"00",X"00",X"00",
		X"2F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"2F",X"2F",X"0F",X"0F",X"1F",X"2F",X"0F",X"0F",X"6F",X"CF",X"0F",X"8F",X"0F",X"0F",X"0F",
		X"00",X"40",X"A0",X"50",X"A0",X"40",X"20",X"10",X"00",X"00",X"00",X"50",X"80",X"00",X"00",X"00",
		X"A7",X"33",X"81",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"8F",X"4F",X"47",X"23",X"01",X"00",
		X"00",X"00",X"02",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"0E",X"07",X"0F",X"0F",X"02",X"02",
		X"00",X"00",X"0E",X"07",X"0F",X"0F",X"07",X"03",X"00",X"00",X"0C",X"46",X"0A",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"02",X"02",X"0C",X"0F",X"07",X"0E",X"00",X"00",
		X"03",X"07",X"00",X"0B",X"07",X"0E",X"00",X"00",X"00",X"0C",X"04",X"0E",X"02",X"08",X"00",X"80",
		X"00",X"00",X"03",X"02",X"01",X"03",X"00",X"00",X"00",X"00",X"0D",X"0E",X"0F",X"0F",X"02",X"02",
		X"00",X"00",X"0D",X"0E",X"0F",X"0F",X"07",X"03",X"00",X"40",X"8C",X"0E",X"0A",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"03",X"00",X"01",X"00",X"00",X"02",X"02",X"0C",X"0F",X"0E",X"0D",X"00",X"00",
		X"03",X"07",X"00",X"07",X"0E",X"0D",X"00",X"00",X"00",X"0C",X"04",X"06",X"0A",X"08",X"00",X"00",
		X"00",X"00",X"03",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"0B",X"0D",X"0F",X"0F",X"42",X"02",
		X"00",X"00",X"0B",X"0D",X"0F",X"0F",X"07",X"03",X"00",X"00",X"0C",X"0E",X"0A",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"02",X"01",X"11",X"00",X"00",X"02",X"02",X"0C",X"0E",X"0D",X"8B",X"00",X"00",
		X"03",X"07",X"00",X"0E",X"0D",X"0B",X"00",X"00",X"00",X"0C",X"04",X"1E",X"0A",X"08",X"00",X"00",
		X"00",X"00",X"03",X"03",X"01",X"03",X"00",X"00",X"00",X"00",X"07",X"0B",X"0F",X"0F",X"02",X"02",
		X"00",X"00",X"07",X"0B",X"0F",X"0F",X"07",X"03",X"00",X"00",X"04",X"0E",X"0A",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"03",X"41",X"01",X"00",X"00",X"02",X"12",X"0C",X"0D",X"0B",X"07",X"00",X"00",
		X"03",X"07",X"00",X"0D",X"0B",X"07",X"00",X"00",X"00",X"0C",X"04",X"0E",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"01",X"04",X"0F",X"00",X"0E",
		X"00",X"03",X"04",X"0F",X"00",X"0F",X"00",X"01",X"00",X"0E",X"00",X"0E",X"00",X"0C",X"02",X"02",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"04",X"04",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"08",X"04",X"03",X"00",X"02",X"02",X"00",X"00",X"0E",X"00",X"0E",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FE",X"FB",X"FD",X"FE",X"FF",X"FF",X"0E",X"08",X"0C",X"06",X"0B",X"0D",X"06",X"0B",
		X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F9",X"F4",X"F2",X"F0",X"F1",X"FB",X"FF",X"FF",X"02",X"01",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"08",X"0C",X"0E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FE",X"0E",X"0C",X"0D",X"08",X"00",X"04",X"02",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FB",X"FD",X"F6",X"FB",X"FD",X"FE",X"FF",X"FF",X"84",X"09",X"0D",X"07",X"0B",X"0F",X"07",X"0F",
		X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FE",X"F8",X"F0",X"F0",X"F3",X"F6",X"0E",X"08",X"01",X"03",X"06",X"0C",X"08",X"00",
		X"F7",X"F0",X"71",X"F3",X"F9",X"F4",X"F2",X"F1",X"0F",X"0F",X"0F",X"0F",X"0D",X"09",X"01",X"00",
		X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"FF",X"00",X"08",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"70",X"F1",X"F3",X"F6",X"74",X"FC",X"F8",X"F0",X"0C",X"09",X"01",X"03",X"03",X"07",X"07",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",
		X"70",X"F0",X"F8",X"F8",X"F4",X"F2",X"F1",X"F0",X"8F",X"07",X"07",X"03",X"03",X"01",X"01",X"0C",
		X"F7",X"F3",X"F0",X"F0",X"F8",X"FE",X"FF",X"FF",X"00",X"00",X"08",X"04",X"03",X"01",X"08",X"0E",
		X"F1",X"F3",X"F7",X"FF",X"FF",X"F7",X"F3",X"F7",X"08",X"01",X"0B",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F1",X"0E",X"0C",X"08",X"0D",X"0F",X"0E",X"0C",X"08",
		X"77",X"F1",X"F8",X"F8",X"F4",X"F2",X"F1",X"F0",X"8F",X"0F",X"07",X"01",X"00",X"00",X"00",X"0C",
		X"73",X"F9",X"F8",X"FC",X"7C",X"FE",X"7E",X"FF",X"00",X"00",X"08",X"04",X"03",X"03",X"81",X"00",
		X"71",X"F3",X"F7",X"FF",X"7F",X"FF",X"FF",X"7F",X"0E",X"0F",X"0F",X"0F",X"0F",X"8F",X"8F",X"8F",
		X"7F",X"7E",X"7E",X"7C",X"FC",X"F8",X"F9",X"F3",X"80",X"80",X"82",X"83",X"86",X"0C",X"88",X"00",
		X"70",X"F0",X"F0",X"F0",X"F8",X"F4",X"F2",X"F1",X"87",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F1",X"F3",X"F3",X"F7",X"F7",X"FF",X"FF",X"FE",X"00",X"08",X"0C",X"0E",X"0F",X"0E",X"08",X"00",
		X"F0",X"F1",X"F3",X"F6",X"FC",X"F8",X"F1",X"F7",X"08",X"0C",X"00",X"00",X"01",X"07",X"0F",X"0F",
		X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0D",X"0D",X"0F",
		X"00",X"08",X"0D",X"0F",X"0F",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"08",X"0C",X"0C",X"8A",X"CA",
		X"05",X"04",X"03",X"33",X"13",X"00",X"00",X"10",X"0F",X"0F",X"0F",X"8F",X"C3",X"EF",X"F7",X"F0",
		X"3F",X"2B",X"3F",X"3F",X"3F",X"7F",X"F8",X"F0",X"6E",X"BE",X"7C",X"FC",X"F4",X"F0",X"F0",X"F0",
		X"00",X"06",X"07",X"07",X"03",X"01",X"07",X"01",X"00",X"00",X"01",X"0C",X"0A",X"03",X"07",X"03",
		X"00",X"02",X"07",X"0F",X"07",X"0E",X"0C",X"0E",X"00",X"02",X"06",X"04",X"0C",X"08",X"0E",X"0E",
		X"03",X"07",X"83",X"C0",X"E1",X"F3",X"F7",X"F0",X"0F",X"0E",X"0E",X"0C",X"0F",X"8E",X"F0",X"20",
		X"0F",X"0F",X"0D",X"04",X"0E",X"0C",X"FC",X"70",X"08",X"08",X"08",X"04",X"0C",X"0E",X"04",X"C0",
		X"00",X"03",X"13",X"07",X"07",X"0F",X"0F",X"07",X"F7",X"EF",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"7E",X"7F",X"3F",X"3F",X"3F",X"2F",X"3F",X"7F",X"F0",X"F0",X"FC",X"FE",X"7E",X"BF",X"6F",X"CF",
		X"0F",X"0F",X"0F",X"07",X"07",X"01",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"7F",X"7F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"8F",X"0F",X"0E",X"0E",X"0E",X"0E",X"08",X"00",
		X"F0",X"F0",X"E0",X"C0",X"81",X"01",X"03",X"03",X"F0",X"C0",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"08",X"08",X"08",X"0C",X"0C",
		X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"31",
		X"00",X"00",X"00",X"00",X"00",X"00",X"82",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"13",X"11",X"00",X"00",X"03",X"01",X"01",X"81",
		X"FF",X"DF",X"A7",X"E6",X"7E",X"7F",X"7F",X"79",X"09",X"CF",X"E9",X"F6",X"F3",X"FF",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"0F",X"CC",X"FC",X"FF",X"F3",X"FB",X"0F",X"0F",X"07",X"02",X"BE",X"EB",X"3F",X"CF",
		X"08",X"08",X"08",X"6C",X"F0",X"70",X"8E",X"0C",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"10",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"F3",X"F7",X"F1",X"73",X"71",X"E1",X"C1",X"01",
		X"FB",X"FE",X"7F",X"39",X"1F",X"1E",X"0E",X"0F",X"F3",X"F5",X"F7",X"FF",X"FF",X"A7",X"B3",X"D7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"FF",X"E4",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"FF",X"EF",X"E9",X"CF",X"8C",X"89",X"0C",X"CF",X"0F",X"09",X"00",X"09",X"0F",X"0D",X"0F",
		X"08",X"0C",X"00",X"08",X"0C",X"0C",X"0C",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0A",X"02",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"01",X"00",X"00",X"03",X"01",X"00",X"00",X"08",X"0C",X"0E",X"07",X"03",X"0F",X"0F",
		X"04",X"06",X"06",X"03",X"0F",X"0F",X"0F",X"0F",X"01",X"01",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"01",X"01",X"01",X"07",X"03",X"01",X"01",X"0F",X"7F",X"7F",X"7F",X"1F",X"1F",X"0F",X"0F",
		X"0F",X"CF",X"FF",X"9F",X"5F",X"FF",X"FF",X"7F",X"0F",X"0F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"02",X"02",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"01",X"03",X"0E",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"01",X"03",X"0F",X"0E",X"0E",X"00",X"06",X"0C",X"08",X"08",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"BF",X"FF",X"EF",X"FF",X"FF",X"0F",X"1F",X"3F",X"CF",X"7F",X"CF",X"CF",X"8F",
		X"1F",X"EF",X"EF",X"CF",X"0F",X"0F",X"0F",X"0F",X"08",X"00",X"00",X"08",X"0E",X"08",X"08",X"08",
		X"01",X"03",X"35",X"11",X"01",X"03",X"06",X"00",X"0F",X"0F",X"EF",X"FF",X"7F",X"FF",X"BF",X"1F",
		X"7F",X"7F",X"FF",X"FF",X"9F",X"8F",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"7F",X"7F",
		X"00",X"01",X"00",X"01",X"03",X"07",X"0C",X"00",X"3F",X"33",X"07",X"0C",X"09",X"01",X"03",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"1F",X"0F",X"09",X"01",X"00",
		X"FF",X"FF",X"FF",X"EF",X"EF",X"6F",X"6F",X"4F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"08",X"08",X"08",X"0C",X"00",X"00",X"08",
		X"CF",X"CF",X"CF",X"0F",X"0E",X"08",X"08",X"08",X"0F",X"0F",X"0F",X"09",X"00",X"00",X"00",X"00",
		X"09",X"08",X"08",X"08",X"0C",X"04",X"02",X"00",X"0C",X"06",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"37",X"7F",X"FF",X"7F",X"1F",
		X"0F",X"0F",X"0F",X"FF",X"5F",X"FF",X"5F",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"3F",X"FF",X"EF",X"FF",X"FF",X"FF",X"7F",X"FF",X"BF",X"6F",X"CF",X"CF",X"8F",X"8F",
		X"88",X"8E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"07",X"0F",X"0F",X"0F",X"07",X"F7",X"F3",X"13",
		X"FF",X"7F",X"3F",X"3F",X"7F",X"EF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"6F",X"63",X"60",X"40",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"AF",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"0E",X"0F",X"0F",X"0E",X"0E",X"0E",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"7F",X"7F",X"2E",X"00",X"00",X"00",X"00",X"8F",X"8F",X"08",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"82",X"0A",X"2F",X"1F",X"0F",
		X"00",X"00",X"00",X"04",X"03",X"5B",X"1E",X"AF",X"00",X"00",X"00",X"28",X"00",X"80",X"00",X"C0",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"1F",X"27",X"05",X"89",X"00",X"00",
		X"4F",X"EF",X"13",X"0F",X"0F",X"0D",X"08",X"00",X"CC",X"CC",X"08",X"80",X"08",X"2C",X"06",X"01",
		X"00",X"00",X"00",X"02",X"01",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"0D",X"06",
		X"00",X"00",X"48",X"01",X"40",X"56",X"47",X"48",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"C0",
		X"12",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"70",X"03",X"00",X"02",X"08",X"00",X"00",X"00",
		X"F5",X"63",X"48",X"42",X"40",X"03",X"40",X"00",X"D4",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"F0",X"00",X"03",X"00",
		X"00",X"01",X"02",X"24",X"C8",X"2C",X"0F",X"02",X"00",X"0F",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"84",X"F3",X"80",X"00",X"00",X"00",X"00",X"04",X"10",X"E8",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"20",X"20",X"30",X"73",X"F0",
		X"00",X"01",X"82",X"84",X"88",X"8C",X"CF",X"E2",X"00",X"0F",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"10",X"30",X"70",X"60",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"30",X"10",X"10",X"30",X"50",
		X"F2",X"F0",X"F4",X"83",X"00",X"00",X"80",X"40",X"00",X"84",X"C0",X"C8",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"70",X"00",X"00",X"10",X"00",X"00",X"00",X"F0",X"F0",X"00",X"70",X"C0",X"80",
		X"00",X"00",X"F0",X"F0",X"00",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"20",
		X"10",X"00",X"00",X"70",X"70",X"00",X"00",X"00",X"80",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"70",X"70",X"00",X"00",X"10",X"00",X"00",X"00",X"F0",X"F0",X"00",X"70",X"C0",X"80",
		X"00",X"00",X"F0",X"F0",X"00",X"90",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"10",X"00",X"00",X"70",X"70",X"00",X"00",X"00",X"80",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F1",X"F1",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"80",X"80",X"00",X"80",X"00",X"80",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"00",X"00",X"30",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F4",X"F0",
		X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"90",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"30",X"30",X"30",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C4",X"C0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"F0",X"F0",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
