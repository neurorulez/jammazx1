-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "FFFFFFFFFFF0FFF01000FD40FFFFFFFF0000017F000000003C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF00000000005F7FFFFFFF003FFFFFFFFFFF7CFFFF";
    attribute INIT_03 of inst : label is "57FFBFFFFFFDFFFFF500FFFF4000FD000000E000000F00002FFF00BFC6832558";
    attribute INIT_04 of inst : label is "283F83FF0002340000001FF0000000000FFF42FF0000001F00000000FFFDFFFF";
    attribute INIT_05 of inst : label is "FBFF003C000F17D0000000000082003400000000003CFF1F0D020BF0C0FF703F";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "FFFFFFFF4400980050002000000000240000000A0F0003402F5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "3FA00000FFFFFFFF0000FC3D00000000000F000F01F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "800300000E00C00303703FC30000000C1C003E00C0003FC0000AC00000000000";
    attribute INIT_0D of inst : label is "BAFF00FCFDFFFFFF0000401F0FC000B0001E0780000004030000000000D40008";
    attribute INIT_0E of inst : label is "000001D0A000000050023C00FFFF02FF00003540000000000200000000F003C0";
    attribute INIT_0F of inst : label is "0F8FFFE000C00407E3F2C0030003000FD7F0FFF000000000C000FC00FF80F800";
    attribute INIT_10 of inst : label is "0000000001010000020200000000000000000000F01F007FFFECFF0003FF3FFF";
    attribute INIT_11 of inst : label is "0000000000000360000000000000028000000000000001010000020200000000";
    attribute INIT_12 of inst : label is "0360000000000000028000000000000000000000000000000000000000000110";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000110000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "67899006CF532418C003275801D82498071029C001500A240000000000000000";
    attribute INIT_16 of inst : label is "00006789241800000000CF53082000000550CFA3000000001BE4CA0300000000";
    attribute INIT_17 of inst : label is "3D4C90600F50000005F00000CFA3082000000550CA03000000001BE490060000";
    attribute INIT_18 of inst : label is "4C00600000CF00245300180000330009D4C00600000C0002F530418000030000";
    attribute INIT_19 of inst : label is "2C2038E603049EB40204298C33D40906C00000000CF5024130008000033D0090";
    attribute INIT_1A of inst : label is "000001FF0FFF0FFF00000000F5500000FFFF00000AFF0000000A00000033A498";
    attribute INIT_1B of inst : label is "02400240D4000F0F00170F0F0000FF40FFF0FFF000000000057E000000000000";
    attribute INIT_1C of inst : label is "02400240D4000F0F00170F0F0000F0F000000000BFFE382C024002401414A41A";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "3D01800A2BDF0A00FFFEFDE04540BC003D010142500F0A00FFFEFDE04540BC00";
    attribute INIT_21 of inst : label is "000142FA7FDF0A00FFFEFDE04540BC003D0102AA7FDF0A00FFFEFDE04540BC00";
    attribute INIT_22 of inst : label is "F07F0142500F282AFFF6FC554540A000200182FA7FDF0000FFFEFDE04540BC00";
    attribute INIT_23 of inst : label is "3DF5800A2BDF0A28FFFEFDE04540BC003DF50142500F0A28FFFEFDE04540BC00";
    attribute INIT_24 of inst : label is "007542FA7FDF0A28FFFEFDE04540BC003DF502AA7FDF0A28FFFEFDE04540BC00";
    attribute INIT_25 of inst : label is "FF7F0142500F2AAAFFF6FC554540A000200582FA7FDF0028FFFEFDE04540BC00";
    attribute INIT_26 of inst : label is "3D01800A2BDF0A00FFFEFD784540BC003D010142502F0A00FFFEFD784540BC00";
    attribute INIT_27 of inst : label is "000142FA7FDF0A00FFFEFD784540BC003D0102AA7FDF0A00FFFEFD784540BC00";
    attribute INIT_28 of inst : label is "200182FA7FDF0000FFFEFD784540BC00200182FA7FDF0000FFFEFD784540BC00";
    attribute INIT_29 of inst : label is "3D0102AA7FDF0A00FFFEFD784540BC00000142FA7FDF0A00FFFEFD784540BC00";
    attribute INIT_2A of inst : label is "3D010142502F0A00FFFEFD784540BC003D01800A2BDF0A00FFFEFD784540BC00";
    attribute INIT_2B of inst : label is "F07F0142500F282AFFF6FC7D4540A000F07F0142500F282AFFF6FC7D4540A000";
    attribute INIT_2C of inst : label is "082000000000000A0855BD2A3C00AF60820800000000000A0855BD2A3C0CAF60";
    attribute INIT_2D of inst : label is "820800000000000A0855BD2A3C00AF60208200000000000A086ABD3F3C0CAF60";
    attribute INIT_2E of inst : label is "208200000000000A0855BD2A3C00AF60082000000000000A087FBD153C0CAF60";
    attribute INIT_2F of inst : label is "082000000080000A0855BD2A3C00AF60820800000080000A0855BD2A3C0CAF60";
    attribute INIT_30 of inst : label is "820800000080000A0855BD2A3C00AF60208200000080000A0855BD2A3C0CAF60";
    attribute INIT_31 of inst : label is "208200000080000A0855BD2A3C00AF60082000000080000A0855BD2A3C0CAF60";
    attribute INIT_32 of inst : label is "0000010000000000400080104000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "00BA02DA00130080FE0072E0D4480000012300A900040000B040D34000000000";
    attribute INIT_34 of inst : label is "000033330000000000003335000000001FBFE7C81BE70028FEF48BDDFC102000";
    attribute INIT_35 of inst : label is "0000333300000000000033170000000000003333000000000000351700000000";
    attribute INIT_36 of inst : label is "0000033300000000000030C00000000000003333000000000000330C00000000";
    attribute INIT_37 of inst : label is "0028006800000000290021000000000000680048000000002800290000000000";
    attribute INIT_38 of inst : label is "5002400240404D41155350504D44464E18BF01C8D04364EC400637400D2C437C";
    attribute INIT_39 of inst : label is "5F595A4A5D4B5F4B0A1F0E5F4B343972949591D545454554C5C4C58410515045";
    attribute INIT_3A of inst : label is "D5430141E11B4151E81141547401151000961300545400CC44ED444F41150145";
    attribute INIT_3B of inst : label is "15410740F1104954F1104D5454143F014445E1074350114951115039011414F4";
    attribute INIT_3C of inst : label is "ADD96DF8B0A6A022F8F5F0B4C2F6F3F004AA0400025E020E009B00000E5B0E1A";
    attribute INIT_3D of inst : label is "0F0F0F0F343F3C2F0B020A042FDB0FFAAF0F2FCBFDAFBF2FFAF2FAFD2FFACBFA";
    attribute INIT_3E of inst : label is "00F54140007D5414007D541400571501007E5414009010050094150104E04445";
    attribute INIT_3F of inst : label is "007D5414005715010057150100DD414000D7150100C5414000C54140007F5414";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "FFFCFFFFFFFCFFF00000FC001FFFFFFF0000000F0000000005540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF00000000000501FFFFFFAAFFFFFFFFFFFC00FFFD";
    attribute INIT_03 of inst : label is "01FFFFFFFFFEFFFF5000FFD50000F00000004000003F00023FFF0BFF1AA4C943";
    attribute INIT_04 of inst : label is "BC3F50FF00030000000005D0000000003FFF0FFF000000010000000BFFFEFFFF";
    attribute INIT_05 of inst : label is "FFFF80B0000F0003000000000BFF00100000000002F4D42D3C2F0FD002FF30FF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "FFFFFFFF01006400C0007800002400370010003B00000B001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "FFFC0000FCFFFFFF0000100000030000000F000F2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "C00300003F000001003B1FF3C00200050F003D00C000DF40000F400000000000";
    attribute INIT_0D of inst : label is "FFFF00FCD07FFFFF000000003D0003F00C07007000000000000000008003000C";
    attribute INIT_0E of inst : label is "00000000F8000000003F3C007FFF2FFF00000000000000000300000000F003C0";
    attribute INIT_0F of inst : label is "8FCF5FFCCCFB00C3F1CBC0010003000701F8FFF000000000E000F0003FE0FF00";
    attribute INIT_10 of inst : label is "0000020200000000000000000101000002020000F807E03FFFFFFF8000FF07FF";
    attribute INIT_11 of inst : label is "0000000000000000000000000000011000000360000000000000000000000101";
    attribute INIT_12 of inst : label is "0000000000000000011000000000000003600000000000000280000000000000";
    attribute INIT_13 of inst : label is "00000000000036000000000000000D8000000000000000000000028000000000";
    attribute INIT_14 of inst : label is "00000036000000000000000D000080000000000300006000000000000000D800";
    attribute INIT_15 of inst : label is "0550CFA31BE4CA031AA4C1030620376400842DD810C03B78000000D800000000";
    attribute INIT_16 of inst : label is "00000550CA03000000001BE49006000000006789241800000000CF5308200000";
    attribute INIT_17 of inst : label is "6F90280C03C00A0003C000A06789900600000000CF53241800000000CFA30820";
    attribute INIT_18 of inst : label is "90000C00001B00CAE400030000060032F90080C00001000CBE40A03000000003";
    attribute INIT_19 of inst : label is "00826D68104136D9001011B406F932800000C00001BE0CA040003000006F0328";
    attribute INIT_1A of inst : label is "000000000FFF0FFF02AFFFFFFFE80AAFFFFFAAA0FFFF0000AAFF000006203764";
    attribute INIT_1B of inst : label is "02400240C000E0000003000B00000000FFF0FFF0FA80FFFF2BFFFA80FFEA0000";
    attribute INIT_1C of inst : label is "02400240C000E0000003000B000000000000000003C00FF00240024094168412";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "5E8280BF0FFA0B03FE1778000000FDE0DE82400B02FA0B03FE1778000000FDE0";
    attribute INIT_21 of inst : label is "5002EFFF0FFA0303FE1778000000FDE08002EFFF0FFA0B03FE1778000000FDE0";
    attribute INIT_22 of inst : label is "DE87400B02FA2CFFFFAD780000007FEA8002EFFF0FFA0003FE1778000000FDE0";
    attribute INIT_23 of inst : label is "5E8280BF0FFA0BB7FE1778000000FDE0DE82400B02FA0BB7FE1778000000FDE0";
    attribute INIT_24 of inst : label is "5002EFFF0FFA03B7FE1778000000FDE08002EFFF0FFA0BB7FE1778000000FDE0";
    attribute INIT_25 of inst : label is "DE87400B02FA2FFFFFAD780000007FEA8002EFFF0FFA0037FE1778000000FDE0";
    attribute INIT_26 of inst : label is "5E8280BF0FFA0B03FEB7797C0000FDE0DE82400B02FA0B03FEB7797C0000FDE0";
    attribute INIT_27 of inst : label is "5002EFFF0FFA0303FEB7797C0000FDE08002EFFF0FFA0B03FEB7797C0000FDE0";
    attribute INIT_28 of inst : label is "8002EFFF0FFA0003FEB7797C0000FDE08002EFFF0FFA0003FEB7797C0000FDE0";
    attribute INIT_29 of inst : label is "8002EFFF0FFA0B03FEB7797C0000FDE05002EFFF0FFA0303FEB7797C0000FDE0";
    attribute INIT_2A of inst : label is "DE82400B02FA0B03FEB7797C0000FDE05E8280BF0FFA0B03FEB7797C0000FDE0";
    attribute INIT_2B of inst : label is "DE87400B02FA2CFFFFAD787C00007FEADE87400B02FA2CFFFFAD787C00007FEA";
    attribute INIT_2C of inst : label is "82080000000200003F3F3D15BC0017AA20820000000200003F3F3D15BC0017AA";
    attribute INIT_2D of inst : label is "20820000000200003F3F3D15BC0017AA08200000000200003F153D00BC0017AA";
    attribute INIT_2E of inst : label is "08200000000200003F3F3D15BC0017AA82080000000200003F2A3D15BC001780";
    attribute INIT_2F of inst : label is "8208000002C200003F3F3D15BC0017AA2082000002C200003F3F3D15BC0017AA";
    attribute INIT_30 of inst : label is "2082000002C200003F3F3D15BC0017AA0820000002C200003F3F3D15BC0017AA";
    attribute INIT_31 of inst : label is "0820000002C200003F3F3D15BC0017AA8208000002C200003F3F3D15BC0017AA";
    attribute INIT_32 of inst : label is "0000000400000000840000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "06E508BD00001000CDF08FA0000000040199008E000000080C409C8000000000";
    attribute INIT_34 of inst : label is "373715150000000037351515000000003F68BDDF044108758FA7DFF04100F9A0";
    attribute INIT_35 of inst : label is "3737151500000000373515150000000037371515000000001735151500000000";
    attribute INIT_36 of inst : label is "037301510000000070E05150000000003737151500000000370E151500000000";
    attribute INIT_37 of inst : label is "0048000800000000280025000000000000280058000000002100200000000000";
    attribute INIT_38 of inst : label is "A0228282A29A0881A6A2A0A28A838B0AA5A287ACA03287AC05276441A8A22248";
    attribute INIT_39 of inst : label is "A5A4AF8DACAD870727A78DAD8D9034B3787AD29ADACA7A683A329898E0A2A09A";
    attribute INIT_3A of inst : label is "42838280E22B22A8C0202AA830080A20020A2882202A200E82C28227C680A808";
    attribute INIT_3B of inst : label is "8A800380F2082CA8F22824A828023E02822AF20323A0002EA022203C082820B8";
    attribute INIT_3C of inst : label is "0A12C2820A080ACA222A8E0A1A2A8888080A0800A0A8A2A200A00020A2A8AAAA";
    attribute INIT_3D of inst : label is "0808020207082302000C000F081032800272C830210208C88084202342803020";
    attribute INIT_3E of inst : label is "80D88228283EA802283EA80202832A80283CA802084220880042288282CA882A";
    attribute INIT_3F of inst : label is "283EA80202C32A8002C32A8080E8822802832A8080F8822880F88228283DA802";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "FFFEFE001F4FFFFF0000000000000000FFFFFE8000003FF13C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF7FFCFFFF00000000";
    attribute INIT_03 of inst : label is "57FFFFFE00020000F50000BFBFFF02FF007FFFFFFFFFFFFFD000FFFFC6832558";
    attribute INIT_04 of inst : label is "C03F03FFFEFF00BFFFFFE00FFC50FFFF0FFF02FFFFFFFFE0FF40FFFF00020000";
    attribute INIT_05 of inst : label is "000003C0F1F4E8007FE0FC3CD082FE00001F0FFFFFC000E04002C00000FF803F";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "FFFFFFFFC400FE00D400F8000024002F004C002F0C5400002F5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "3FA01FFFFFFFFFFF0000FC3D07FF0FFF0FF000F001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "7FFCFFFFF1FF3FFCFC80C0000FF1FFF0E3F0C1C037F0C03CFCF534BC3FFFFC3F";
    attribute INIT_0D of inst : label is "BAFFF0FCFDFFFFFF0000401FF03FFF4FFFE1F87FFFFFFBFCFFF3FFFF0F007FE0";
    attribute INIT_0E of inst : label is "FFFFFE2F5FFFFFFFA542C3FFFFFF02FF3F40356847933FF74203C0C7E0F003C0";
    attribute INIT_0F of inst : label is "0000001F073C0BC0E000C3FCFFC0FC00280000000000005C3FF303FF007F07FA";
    attribute INIT_10 of inst : label is "0000000051050000A20A00000000000000000000F0000000FFECFF00FC00C000";
    attribute INIT_11 of inst : label is "0000000000003FFC0000000001502FF807F40AA0000051050000A20A00000000";
    attribute INIT_12 of inst : label is "3FFC0000000000002FF80000000001500AA00000000007F40000000000001FFC";
    attribute INIT_13 of inst : label is "000000007F40AA00000000001FD02A8000000000000000001FFC000000000000";
    attribute INIT_14 of inst : label is "007F00AA40000000001F002AD00080000007000AF400A00000010002FD00A800";
    attribute INIT_15 of inst : label is "078003000F5003400F50034033D83FFE1758BFF84DD72FFC01FD02A800000000";
    attribute INIT_16 of inst : label is "000007800340000000000F500280000000000FA00000000001400B0000000000";
    attribute INIT_17 of inst : label is "3D400D000F50034005F001C00FA00280000000000B0000000000014003000000";
    attribute INIT_18 of inst : label is "40000000000F00035000400000030000D400D00000000000F500340000000000";
    attribute INIT_19 of inst : label is "2C68BFFE0B87BFFE0664AFAE03D400D00000000000F5003400000000003D000D";
    attribute INIT_1A of inst : label is "00003FFFFFFFFFFFFFFFFFFF0AAF02AF000002A8F500000000A500003233BFFE";
    attribute INIT_1B of inst : label is "00000000D400FFFF0017FFFF0000FFFCFFFFFFFFFFFFFFFFFA81FA80FFA00000";
    attribute INIT_1C of inst : label is "00000000D400FFFF0017FFFF0000FFFFBFFE382CBFFE382C000000001FF4A28A";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "00007FF55400340000000000000000000000FEBDAFD034000000000000000000";
    attribute INIT_21 of inst : label is "BF80BD050000340000000000000000008000FD55000034000000000000000000";
    attribute INIT_22 of inst : label is "0000FEBDAFD0D00000AB0000000000005FF07D0500001F000000000000000000";
    attribute INIT_23 of inst : label is "00F57FF554003428000000000000000000F5FEBDAFD034280000000000000000";
    attribute INIT_24 of inst : label is "BFF5BD0500003428000000000000000080F5FD55000034280000000000000000";
    attribute INIT_25 of inst : label is "0F54FEBDAFD0D28000AB0000000000005FF57D0500001F280000000000000000";
    attribute INIT_26 of inst : label is "00007FF55400340000000038009600000000FEBDAFD034000000003800960000";
    attribute INIT_27 of inst : label is "BF80BD050000340000000038003400008000FD55000034000000003800960000";
    attribute INIT_28 of inst : label is "5FF07D0500001F0000000038009600005FF07D0500001F000000003800340000";
    attribute INIT_29 of inst : label is "8000FD55000034000000003800340000BF80BD05000034000000003800960000";
    attribute INIT_2A of inst : label is "0000FEBDAFD03400000000380034000000007FF5540034000000003800340000";
    attribute INIT_2B of inst : label is "0000FEBDAFD0D00000AB0028003400000000FEBDAFD0D00000AB002800960000";
    attribute INIT_2C of inst : label is "0820000000000000543FA83F000000008208000000000000543FA83F003F0000";
    attribute INIT_2D of inst : label is "8208000000000000543FA83F000000002082000000000000543FA83F003F0000";
    attribute INIT_2E of inst : label is "2082000000000000543FA83F000000000820000000000000543FA83F003F0000";
    attribute INIT_2F of inst : label is "082003C000D00000543FA83F00000000820803C000D00000543FA83F003F0000";
    attribute INIT_30 of inst : label is "820803C000D00000543FA83F00000000208203C000D00000543FA83F003F0000";
    attribute INIT_31 of inst : label is "208203C000D00000543FA83F00000000082003C000D00000543FA83F003F0000";
    attribute INIT_32 of inst : label is "0020010400000000420084104000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "00000027000400800420780000080100010A005B00C00000C840F70810000000";
    attribute INIT_34 of inst : label is "0000333300000000000033350000000005020832060000000180C40102042020";
    attribute INIT_35 of inst : label is "0000333300000000000033170000000000003333000000000000351700000000";
    attribute INIT_36 of inst : label is "0000033300000000000030C00000000000003333000000000000330C00000000";
    attribute INIT_37 of inst : label is "002B006F00000000E900F10000000000006B004F00000000E800F90000000000";
    attribute INIT_38 of inst : label is "0083008FAE9CAC020D0300030D0C018CDCFA01BEDBCF39C7323B3280BD3F0FAF";
    attribute INIT_39 of inst : label is "0808080808A828A8880280029863682C2B202CA000300003A0AAA2AB0F0C0F00";
    attribute INIT_3A of inst : label is "00032800C0030000E800000238008002028802220080008C02E80A0BE4808080";
    attribute INIT_3B of inst : label is "00082300E0020800E00200000000BE000000E0030B00200808800038800002B0";
    attribute INIT_3C of inst : label is "02820A222A0B0A0B028A022A8B0B2B0BFB75FBFFAFA7ADA5FF65FFEFA5A5A5A7";
    attribute INIT_3D of inst : label is "820000080022080002000000008208200008008288002200200800880820A200";
    attribute INIT_3E of inst : label is "00C40002003D0080003D008000430028003E008000000A200002022B08E00002";
    attribute INIT_3F of inst : label is "003D0080004300280043002800D400020043002800D4000200D40002003C0080";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "FFFFFFE000017FFF00000000E0000000FFFFFFF00000074005540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF00D4FFFF00000000";
    attribute INIT_03 of inst : label is "01FFFFFF002F00005000E3D5FFFF0FFF003D43FFFFFFFFFFC000F4551AA4C943";
    attribute INIT_04 of inst : label is "403FA0FFFFFF20FFFFFFFA2FD000FFFC3FFF0FFFFFFFFFFEF400FFFF002F0000";
    attribute INIT_05 of inst : label is "00000040FCF0FFF000F0FF04CBFFFD00000101FFF5002BD0002FC00002FFC0FF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "FFFFFFFF4900FD00C400FE000024007F003200FF03C008001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "FFFC0017FCFFFFFF0000100000FC0FFF0FF008F02ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "3FFCFFFFC0DFFFFEFFC0E000C5421FF2F0F0C2C0304020B0FC70B0FF3FFF7CFF";
    attribute INIT_0D of inst : label is "FFFF40FCD07FFFFF00000000C2FFFC0FF3F8FF8FFFFFFFFFFFCBFFFF80033FF0";
    attribute INIT_0E of inst : label is "FFFFFFFF07FFFFFFC03FC3FD7FFF2FFF0100AFF001CF9FF30303C003F0F0C3C0";
    attribute INIT_0F of inst : label is "80000003C3040F30F000C3FCFFF0FF80F4000000000000011FF10FF7C01F00FF";
    attribute INIT_10 of inst : label is "0000A20A000000000000000051050000A20A0000F800E000FFFFFF80FF00F800";
    attribute INIT_11 of inst : label is "0AA00000000007F40000000000001FFC00003FFC000000000000000000005105";
    attribute INIT_12 of inst : label is "07F40AA0000000001FFC0000000000003FFC0000000000002FF8000000000150";
    attribute INIT_13 of inst : label is "000000030000FFC0000000000000FFF0000000000000000001502FF800000000";
    attribute INIT_14 of inst : label is "000003FF0000C000000000FF0000F0000000003F0000FC000000000F0000FF00";
    attribute INIT_15 of inst : label is "00000FA001400B0001400B0006A07FFD0CA4BFFE32C4FFFE00000FFF00000000";
    attribute INIT_16 of inst : label is "000000000B0000000000014003000000000007800340000000000F5002800000";
    attribute INIT_17 of inst : label is "05002C0003C00B0003C000E007800300000000000F500340000000000FA00280";
    attribute INIT_18 of inst : label is "000000000001000B40000000000000025000C000000000001400B00000000000";
    attribute INIT_19 of inst : label is "0CE27FFD30657FFD001057FD005002C000000000001400B0000000000005002C";
    attribute INIT_1A of inst : label is "000005FFFFFFFFFFFFFF00000017F5500000555F0000AAFF5500000006A47F7D";
    attribute INIT_1B of inst : label is "00000000C000E0000003000B0000FF50FFFFFFFFFFFF0000D400057E00158000";
    attribute INIT_1C of inst : label is "00000000C000E0000003000B0000000003C00FF003C00FF00000000097D68FF2";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "A0207F400000000001E00000000008002020BFF4BD00000001E0000000000800";
    attribute INIT_21 of inst : label is "AFFC10000000A80001E00000000008007FE810000000000001E0000000000800";
    attribute INIT_22 of inst : label is "2020BFF4BD000002005F0000000000007FFC100000001FC001E0000000000800";
    attribute INIT_23 of inst : label is "A0787F40000000B401E00000000008002078BFF4BD0000B401E0000000000800";
    attribute INIT_24 of inst : label is "AFFC10000000A8B401E00000000008007FF81000000000B401E0000000000800";
    attribute INIT_25 of inst : label is "2170BFF4BD000B42005F0000000000007FFC100000001FF401E0000000000800";
    attribute INIT_26 of inst : label is "A0207F400000000001E0017C014108002020BFF4BD00000001E0017C01410800";
    attribute INIT_27 of inst : label is "AFFC10000000A80001E0017C005008007FE810000000000001E0017C01410800";
    attribute INIT_28 of inst : label is "7FFC100000001FC001E0017C014108007FFC100000001FC001E0017C00500800";
    attribute INIT_29 of inst : label is "7FE810000000000001E0017C00500800AFFC10000000A80001E0017C01410800";
    attribute INIT_2A of inst : label is "2020BFF4BD00000001E0017C00500800A0207F400000000001E0017C00500800";
    attribute INIT_2B of inst : label is "2020BFF4BD000002005F007C005000002020BFF4BD000002005F007C01410000";
    attribute INIT_2C of inst : label is "D75D00000000000040FF00150000E82A75D700000000000040FF0015000CE82A";
    attribute INIT_2D of inst : label is "75D700000000000040FF00150000E82A5D7500000000000040FF0015000CE82A";
    attribute INIT_2E of inst : label is "5D7500000000000040FF00150000E82AD75D00000000000040FF0015000CE82A";
    attribute INIT_2F of inst : label is "D75D0AF002C0000040FF00150000E82A75D70AF002C0000040FF0015000CE82A";
    attribute INIT_30 of inst : label is "75D70AF002C0000040FF00150000E82A5D750AF002C0000040FF0015000CE82A";
    attribute INIT_31 of inst : label is "5D750AF002C0000040FF00150000E82AD75D0AF002C0000040FF0015000CE82A";
    attribute INIT_32 of inst : label is "0004002400000000840006000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "8029084702001200FA08740004004004084F001F00000008BF80D18000000400";
    attribute INIT_34 of inst : label is "373715150000000037351515000000004819C02000002880920C310000000400";
    attribute INIT_35 of inst : label is "3737151500000000373515150000000037371515000000001735151500000000";
    attribute INIT_36 of inst : label is "037301510000000070E05150000000003737151500000000370E151500000000";
    attribute INIT_37 of inst : label is "004F000100000000F800450000000000002F005100000000F100400000000000";
    attribute INIT_38 of inst : label is "A0E0B0AC5C005187E4A0A1A0818888004C059D4C1480AE047F4EC1D7130060D3";
    attribute INIT_39 of inst : label is "AAAFAFBBA3558154EAEDAEA9003B72AD5F0A1ECA5A3A4A2BDA8F9ACB6FAEAF8A";
    attribute INIT_3A of inst : label is "14170140D4470110E945001471510004519601055005464C14E54103B0155545";
    attribute INIT_3B of inst : label is "11104745E0500101E0400D1154403D144001C457030144401010457111114474";
    attribute INIT_3C of inst : label is "01218100000700C3C005380433C60233F7EBF7FF0E5A0E0EFFDEFFCF0F5E0F1E";
    attribute INIT_3D of inst : label is "90535C507A40434C5058505A433060000CE08320030C00830038C003800020C0";
    attribute INIT_3E of inst : label is "55F94000557C1400557C140055970100557E1400509502015594000150E04401";
    attribute INIT_3F of inst : label is "557C1400555701005557010055C540005557010055E9400055E94000557F1400";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
