-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "000F000FF000F000000000000000000000030003C000C00000FA02FF00000000";
    attribute INIT_01 of inst : label is "000F000FF000F000000000000000000000030003C000C000EBC0FFE000000000";
    attribute INIT_02 of inst : label is "C003C003C003C00300000000D0030003C003D557C007C000D000000000070000";
    attribute INIT_03 of inst : label is "C000C00000030003C3C3C3C3000303C3C000C3C003C30003C3C0C000FAAFF55F";
    attribute INIT_04 of inst : label is "01800000FFF4782FFFFF5FF51FFFF82DFFFFF82FFFFFF82F03F0004000000000";
    attribute INIT_05 of inst : label is "2FFFAAA0000003C00BE0AAAAFFF80AAAFFFFF82FFFFFF82F1FFFFFFD00000000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0018180000F400E009D818C907C002C009000009014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC6832558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "000015552FFFAAA0FFF80AAAFFF47FFF00000000201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "60C0FFFC05432DE1C00052CF0001FE01000000000000000000000000FFFFFFFF";
    attribute INIT_0E of inst : label is "037D07F8707DB4BE0FFCFAB41D3C0A0BF8B800002F813A0000003F800000BC00";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000FFFF0000FFFFFFFF000FFFFFF000FFFF0000FFFF0000000FFFFFF000FFFF";
    attribute INIT_11 of inst : label is "0000FFFF0000FFFFFFFF000FFFFFF000FFFF0000FFFF0000000FFFFFF000FFFF";
    attribute INIT_12 of inst : label is "3E00000057D0FF000054003E003C0000FF00E0000000FD00000001F50BFF002F";
    attribute INIT_13 of inst : label is "F000C0000000FC000000003F000F00003FFC0BE000000FF40000000000000000";
    attribute INIT_14 of inst : label is "0000000000000400000000080020002008000000000066000000001800030000";
    attribute INIT_15 of inst : label is "E0000000D400FE00005F02FF002F0003FC0000000000FF0000000000000700FA";
    attribute INIT_16 of inst : label is "FFC0FE00800000000000000003FF00BFFFC0E8000000D000007400410FFF00BF";
    attribute INIT_17 of inst : label is "FFE0BE00C000FFFC00000FFF03FF002F810055500000CC00000000CC010A1555";
    attribute INIT_18 of inst : label is "002F0003000700FA002000200054003EFF00E0000000FD00000001F50BFF002F";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000010A1555002F00000FFF00BF";
    attribute INIT_1A of inst : label is "005F02FF0000000000000008000000180000003F000000000054003E000001F5";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000CC14000FFF00740041";
    attribute INIT_1C of inst : label is "00003FC000000400000066000000FC0000000FF457D0FF000000FD0000000000";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000000CC000000FD000000D000D400FE00";
    attribute INIT_1E of inst : label is "FC0000000000000008000000F000C0003FFC0BE03E000000FF00E00000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000081005550FF000280FFF0FA00E0000000";
    attribute INIT_20 of inst : label is "0FF501FF000002FFD7FCFFD00000FFE000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0FFF03F4003F02BFFFF0C7C0FF00FAA03FF507FF00002FFFD7FFFFF40000FFFE";
    attribute INIT_22 of inst : label is "0000FFF51FFF00000000F5FFFFF400000FFF03FC001F7800A8003D7FFFFC0000";
    attribute INIT_23 of inst : label is "07FF00000000FF57FFF400000000D5FF000A1FFF00FF0000BFFF5C3CFFF0002C";
    attribute INIT_24 of inst : label is "0FFF3FEA07FF000AFFFCEAFFFFF4A8001FF503FF003F2FFFD7FCFFD0C000FAA8";
    attribute INIT_25 of inst : label is "0000000000000008001000000000A880003F03F02FFF0000FFC0C3FCFFFF0000";
    attribute INIT_26 of inst : label is "0000000000000000FF00FF00000000000003000000020000F000400020000000";
    attribute INIT_27 of inst : label is "00000000000000000B0004000000000000000000000000000F000F0000000000";
    attribute INIT_28 of inst : label is "01010000000000D7D01000000000F5C0000000D40A0000800000351E00181201";
    attribute INIT_29 of inst : label is "005F024605002580FD40E46000140096005E024611001580AD40E46000110095";
    attribute INIT_2A of inst : label is "002F1A4100000294FE00D069000005A00078003D030026000B40DF0040300026";
    attribute INIT_2B of inst : label is "000258D4020B20044000350409060600007E003C00601580AF40CF0002400095";
    attribute INIT_2C of inst : label is "000F000D00FD0FFFFC009C001FC0FFFC02F900000000001FBE0000000000D000";
    attribute INIT_2D of inst : label is "0007000000002FBFFFE02EEC7474F0F0000F000D3FF40FFFFC009C0007FFFFFC";
    attribute INIT_2E of inst : label is "07FA0141003F3F0002A87FA0EFD400007DFF00010003002FFFD07F7CEFD04028";
    attribute INIT_2F of inst : label is "0002FFFF01F40000BF8053BB3FD00F00FFE0BF55000B00000BFF57DEFFD00000";
    attribute INIT_30 of inst : label is "005B0000000008DF940000000000DC805800500C0900118060340304B0800C06";
    attribute INIT_31 of inst : label is "008701B7001E01C9F480F790ED0060D03C030003000501C9F00F7000540060D0";
    attribute INIT_32 of inst : label is "0780241F240FC000C280BAA8FFC00000000E3000000000C3B6FF7F40FF544000";
    attribute INIT_33 of inst : label is "ADEB27FF030000280C30FF00FF543CF05FE000BD3000000000FC57EA17E00028";
    attribute INIT_34 of inst : label is "000F0B4D07952E25C000C7805B4042E020ED617F10000D0238B4FF00FFFC8A00";
    attribute INIT_35 of inst : label is "000D0000000000021C0000000000A000200C5400424801808040002A0C16002B";
    attribute INIT_36 of inst : label is "00000002001F00140000A000FD00050000000002001F00140000A000FD000500";
    attribute INIT_37 of inst : label is "00000000000000000203000000000000000000000000A0000203000000000028";
    attribute INIT_38 of inst : label is "0000000000000800000000000000000800000000000000F00203000000003C00";
    attribute INIT_39 of inst : label is "CC93CCCF33333274C3C00F1DC3E0F5F000000000000000004000000080000000";
    attribute INIT_3A of inst : label is "3C301F4300010F83A004E0C0D3F2FFFC3FF800070000FC010003C0000000F4CF";
    attribute INIT_3B of inst : label is "07FE0E03BFFF38000000F838FCDF0000D0000000C0003C000FC0000000003F00";
    attribute INIT_3C of inst : label is "C3C3F0FFFC00BCBCC30F03FF0F000FA02F3F3F3C0C0F000BC0700FFC0000FABC";
    attribute INIT_3D of inst : label is "003EE00F1FD0000003C000FC00070F0708023C33EE0C0000263F330F0000003F";
    attribute INIT_3E of inst : label is "0000000000000000000B000F003F000000030000E000FD03F000F800FC00C540";
    attribute INIT_3F of inst : label is "FE0303C303C30000D078C00FC02D0000F5F400F300000AF83C023C3D3C300800";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "000F000FF000F000000000000000000000030003C000C000001F03F500000000";
    attribute INIT_01 of inst : label is "FFFF000FFFFFF000FFFC00003FFF0000FFFF0003FFFFC000FD00D7F0FFFF0000";
    attribute INIT_02 of inst : label is "4001C0034001C003000000000003E003EAABC003C000C00B0000E0000000000B";
    attribute INIT_03 of inst : label is "4000C00000010003C3C3C3C3FFFFFFC3FFFFC3FFC3C3FFC3C3C3C3FFFFFFF00F";
    attribute INIT_04 of inst : label is "0040000000002FFF00000BE00000FFF8F41FFFFFF41FFFFF004000C000000000";
    attribute INIT_05 of inst : label is "F41F7FFE00000000FFFF5FF5F41FBFFDFFFFFFFFFFFFFFFF0000FFF8FFFF0000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0001018000402AFE10412BFA00402FEA100000900000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C943";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "00000000FFFF7FFEFFFFBFFD00002FFF00000000155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "537B588400013EB20000000100001FFE000000000000000000000000FFFFFFFF";
    attribute INIT_0E of inst : label is "0F00C30F3C00C0C382A048700C0F3F3FFCDFA000FD7F017F0000074040005000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "00000000000000000000000F0000F000000F0000F0000000000F000FF000F000";
    attribute INIT_11 of inst : label is "FFFC00003FFF0000FFFC000F3FFFF000FFFF0000FFFF0000FFFF000FFFFFF000";
    attribute INIT_12 of inst : label is "FC00800000001E00000002F8000F000FFFC0FC0000000000000000000FFF02FF";
    attribute INIT_13 of inst : label is "F800C0000000F4000000001F002F00031FFC2FFC000001D00000000000000000";
    attribute INIT_14 of inst : label is "00000000000040000000000000200020880000000000AD000000000104810004";
    attribute INIT_15 of inst : label is "F000C0000000FF00000003FF003F000FFF00E00000007C00000000000001001F";
    attribute INIT_16 of inst : label is "FF00FFC0400000000002000000FF03CFFF40FF00000040000000000907FF03FF";
    attribute INIT_17 of inst : label is "F0F8FF8040005FD0000B01FD0FFF00FF164068800000440000000044065008A5";
    attribute INIT_18 of inst : label is "003F000F0001001F00200020000002F8FFC0FC0000000000000000000FFF02FF";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000065008A502FF000007FF03FF";
    attribute INIT_1A of inst : label is "000003FF0000000000000000000000010000001F00000000000002F800000000";
    attribute INIT_1B of inst : label is "00000000000000000000000000000000000000000000004400003F1700000009";
    attribute INIT_1C of inst : label is "00001F00000040000000AD000000F400000001D000001E000000000000000000";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000000440000005000000040000000FF00";
    attribute INIT_1E of inst : label is "FF00E0000000000088000000F800C0001FFC2FFCFC008000FFC0FC0000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000016406880FD00BFC0FFD0FFC0F000C000";
    attribute INIT_20 of inst : label is "03FA001700000FFFEBF0F5000000FFFC00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "07FF00F800070FFFFFD0CB40FC00FFFC0FFA017F00003FFFEBFCFF500000FFFF";
    attribute INIT_22 of inst : label is "FFEA3FF0017F0000BFAFF0FDFF40000003FF00FE00001FA0FFFFBC3F55500000";
    attribute INIT_23 of inst : label is "005F000000003FABFD4000000000EAFDABFF03FF00170000FFFFAFFCFF4002FF";
    attribute INIT_24 of inst : label is "2FD51FFF001502FFD5FEFFFD5500FFE00FF0007F00073FFFC3F4F500F000FFFF";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000FF0FFF3D57000BFFF0FFFEFFFFFE00";
    attribute INIT_26 of inst : label is "0000000000000000FF001400010028000003000300000002F000F0000000E000";
    attribute INIT_27 of inst : label is "00000000000000000F0000000100000000000000000000000F00010001000200";
    attribute INIT_28 of inst : label is "00000000000002A9000000000000DAA0105C00541400001017B0150080000000";
    attribute INIT_29 of inst : label is "003D0C00000003A0DF00400C000002B0003D0C00000003A0DF00400C000002B0";
    attribute INIT_2A of inst : label is "003C0400000006BECF0000040000AFA4001F009601A00380FD00E580029000B0";
    attribute INIT_2B of inst : label is "00DC0054240618243700952024038389002F00C1000D0380FE00D0C01C0000B0";
    attribute INIT_2C of inst : label is "000B00BF00F4053FF8007F8007C0FF14005000000000000D140000000000C000";
    attribute INIT_2D of inst : label is "0000000000001F7F1F7CFCFC0000EBC0000B0ABF0540053FF8007FA80054FF14";
    attribute INIT_2E of inst : label is "0FFF002A00071E80FF540D9CFD000000001F00000001BEBFFFE00EECFD00C2FC";
    attribute INIT_2F of inst : label is "02BF02F800000000FFDE0AF43D003E000FFF7D0000070000FF800BBBF5000000";
    attribute INIT_30 of inst : label is "000000000000060E000000000000C240238C0054900000380300151AD0103004";
    attribute INIT_31 of inst : label is "0B13002B00000079F138BA0000008B4007AB003D000000EAFAB4DF000000EAC0";
    attribute INIT_32 of inst : label is "02FD1801400578006B40FA8FF800A0000A57069000000079E3D0AFFC0540E028";
    attribute INIT_33 of inst : label is "00F21815A400023AAED0AFFC05400C30017F09000680BE00FFD03FFF0000003F";
    attribute INIT_34 of inst : label is "00AF0CF700F011EFE8007CC03C00AD10CCFA18010000078387C05FA85F80350F";
    attribute INIT_35 of inst : label is "000000000000000000000000000040008500A90309242040000B0000000010B0";
    attribute INIT_36 of inst : label is "0000002C0001000000000E00500000000000002C0001000000000E0050000000";
    attribute INIT_37 of inst : label is "000000000000000003D00000000000000000000000007C0003D0000000000054";
    attribute INIT_38 of inst : label is "000000000002040000000000A0000004000000000000000003D0000000000000";
    attribute INIT_39 of inst : label is "CCCFCC631B1A33330F2EC3C0F0F0C3D002000203000000000200000100000000";
    attribute INIT_3A of inst : label is "3EF3000300003DF044C032C0011D7FFC07FF00000000FF000000C0000000034F";
    attribute INIT_3B of inst : label is "005F3FE0FD1F1F80E000FCFEFCCF0000000000000000FC000100000000003FC0";
    attribute INIT_3C of inst : label is "C3C3F0143C00F2FFC30F03140F0003FE3F3F0C3C0C0F0B2F08300FD4C2A0FFF0";
    attribute INIT_3D of inst : label is "000FFEBD0000000001F0003F00000F803C331C35017A0000383F0501AA00003F";
    attribute INIT_3E of inst : label is "0000000000000000000F003F003F00020003000070000003F000FC000000C000";
    attribute INIT_3F of inst : label is "4F0303C30F432803C01CC00FFAF4AFE0C0F20FFF0000FFFC3C0B3C343E3E3C00";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "000F000FF000F00000030003C000C000000000000000000000E002FF00000000";
    attribute INIT_01 of inst : label is "000F000FF000F00000030003C000C000000000000000000082C0FFE000000000";
    attribute INIT_02 of inst : label is "C003C003FFFFEAAB00000000FC00A000C003D557003F000AFC00A000003F000A";
    attribute INIT_03 of inst : label is "C000C00000030003000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "01800000000000000000000000000000000000000000000003F0004000000000";
    attribute INIT_05 of inst : label is "00000000000003C0000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0018180000F400E009D818C907C002C009000009014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC0032558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "0000155500000000000000000000000000000000201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "C000C000F000F000FC00FC00FF00FF00FFC0FFC0FFF0FFF0FFFCFFFCFFFFFFFF";
    attribute INIT_0D of inst : label is "0000FFFC00000001000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "037D07F8707DB4BE0FFCFAB4003C000B000000000000000000003F800000BC00";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0003FFFFC000FFFFFFFF000FFFFFF000FFFF0003FFFFC000000FFFFFF000FFFF";
    attribute INIT_11 of inst : label is "0003FFFFC000FFFFFFFF000FFFFFF000FFFF0003FFFFC000000FFFFFF000FFFF";
    attribute INIT_12 of inst : label is "FC00C000000048000003003D003F000380000000680000000024000A00400002";
    attribute INIT_13 of inst : label is "F000C0006900FC00007D003F000F0000CFBCF6C00000F3D000000005F7FF00AA";
    attribute INIT_14 of inst : label is "000000000000240000000018003000303FC0E0000A40002C000000002FE0002F";
    attribute INIT_15 of inst : label is "00000000D400FE00005F02FF0000000080000000D00020000003000000000020";
    attribute INIT_16 of inst : label is "FFC0FE005000FC000000001F03FF00BFFFC0E800F400FFC0000002FF0FFF00BF";
    attribute INIT_17 of inst : label is "FFE0BE001F80FFFC00000FFF03FF002FFFC0AA800000CC00000000CC0FFF0AAA";
    attribute INIT_18 of inst : label is "0010000C00000020003000300003003D80000000680000000024000A00400002";
    attribute INIT_19 of inst : label is "00000000000000000000000000000000000000000FFF0AAA03FF00020FFF00BF";
    attribute INIT_1A of inst : label is "005F02FF000300000000001800000000007D003F000000050003003D0024000A";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000CC15002FFF000002FF";
    attribute INIT_1C of inst : label is "F4000800000024000A40002C6900FC000000F3D0000048006800000000000000";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000000CC000000FD00F400FFC0D400FE00";
    attribute INIT_1E of inst : label is "80000000000000003FC0E000F000C000CFBCF6C0FC00C0008000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFC0AA80FF00BFC0FFF0FA0000000000";
    attribute INIT_20 of inst : label is "0FC001FA000002FF00FCEBD00000FFE000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0FF703F0003F02BFF7F003C0FF00FAA03FC007FA00002FFF00FFEBF40000FFFE";
    attribute INIT_22 of inst : label is "0000FF401FEA00000000407FEAF400000FFF03C0001F7800A800101FFABC0000";
    attribute INIT_23 of inst : label is "07AB00000000FF57EAF400000000D5FF000A1FFC00FF0000BFFF000CAFF0002C";
    attribute INIT_24 of inst : label is "0FD53F0007FF000AD5FC003FFFF4A8001FD003FA003F2FFF41FCEBD0C000FAA8";
    attribute INIT_25 of inst : label is "00000000000056AB000000000000ABAA003F03C02FFF0000FFC000FCFFFF0000";
    attribute INIT_26 of inst : label is "000F001F0001000FFF00FFD0FFFF43D0008F0057003D01F3FC80F540DF00F3D0";
    attribute INIT_27 of inst : label is "000F001F00011E8FFF00FFD0FFFF43D0000F000300012A00FF00FF00FFFFF400";
    attribute INIT_28 of inst : label is "01010000000000D7D0100000000075C001025FD40A4C06821242356430181009";
    attribute INIT_29 of inst : label is "005F0247050025807D40F46000140096005E0247110015802D40F46000110095";
    attribute INIT_2A of inst : label is "002F1A4100000294BE00D069000005A00078003F030026000B40FF0040300026";
    attribute INIT_2B of inst : label is "280258D4020B20004000350009060600007E003F00601580AF40FF0002400095";
    attribute INIT_2C of inst : label is "0000000200300000000020000300000000A40000000000006800000000000000";
    attribute INIT_2D of inst : label is "00000000000000000010011010100C08000000020B4000000000200000780000";
    attribute INIT_2E of inst : label is "000400000007002F00000000802800000000000000000090002D0000822C0000";
    attribute INIT_2F of inst : label is "0000000000000000000000440B6C00D0001E00000000000000000000A92D0000";
    attribute INIT_30 of inst : label is "00000000000000000000000000000000000050000000018000000004B0000000";
    attribute INIT_31 of inst : label is "0000000000100000000000000100000000000000000000000000800000000000";
    attribute INIT_32 of inst : label is "00000000000D000000000000000000000000000000000000002B0040E0800000";
    attribute INIT_33 of inst : label is "000000000000000000000000E08000005E00000000000000002C000014100000";
    attribute INIT_34 of inst : label is "00000002000000000000000000000000000000000000000000000000D0000000";
    attribute INIT_35 of inst : label is "0013000000000009F100690000005800200C00DC40080100800037280802C000";
    attribute INIT_36 of inst : label is "00FF1FFD00E20028FFC05FFD22C00A0003FF2FFD00E20028FFF05FFE22C00A00";
    attribute INIT_37 of inst : label is "0FFF3015000003CAFDFC500000008F000FFF0615000000FAFDFC500000008F00";
    attribute INIT_38 of inst : label is "03FF2FFF00FF02A8FFF0FFFEFFC00AA00FFF24150000280AFDFC5000000080A8";
    attribute INIT_39 of inst : label is "00000000000000000000000000000000584018DC9530200E040ADCA0020600D0";
    attribute INIT_3A of inst : label is "0000000000000003000400000000FFFC00000000000000000000000000000000";
    attribute INIT_3B of inst : label is "00000000000000000000000000000000D000000000003C000FC0000000003F00";
    attribute INIT_3C of inst : label is "C3C3F0FFFC00BCBCC30F03FF0F000FA0003F003C000F000BC0700FFC0000FABC";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000008023C33EE0C00002600330000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "000F000FF000F00000030003C000C0000000000000000000001F03D000000000";
    attribute INIT_01 of inst : label is "000F000FF000F00000030003C000C0000000000000000000FD0041F000000000";
    attribute INIT_02 of inst : label is "4001C0034001FFFF000000005000FC00EAABC0030005003F5000FC000005003F";
    attribute INIT_03 of inst : label is "4000C00000010003000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "004000000000000000000000000000000000000000000000004000C000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0001018000402AFE10412BFA00402FEA100000900000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C003";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "C000C000F000F000FC00FC00FF00FF00FFC0FFC0FFF0FFF0FFFCFFFCFFFFFFFF";
    attribute INIT_0D of inst : label is "0000000400000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0F00C30F3C00C0C382A04870000F003F00000000000000000000074000005000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "00030003C000C0000003000FC000F000000F0003F000C000000F000FF000F000";
    attribute INIT_11 of inst : label is "00030003C000C0000003000FC000F000000F0003F000C000000F000FF000F000";
    attribute INIT_12 of inst : label is "3FC03C00000014000000000300FF000F080020000000D6000000025701080000";
    attribute INIT_13 of inst : label is "F800C0000000F4000000021F002F0003E7F4DB700000064000000000007FBFFF";
    attribute INIT_14 of inst : label is "080000000000400000000001003000300500DA0000000010000000001F50001F";
    attribute INIT_15 of inst : label is "000000000000FF00000003FF0000000020000000000080000000000000000002";
    attribute INIT_16 of inst : label is "FF00FFC00000FC000000000700FF03FFFF40FF000000D0000000005207FF03FF";
    attribute INIT_17 of inst : label is "FFF8FF800000BFD0000001FD0FFF00FFFFC0FFC00000CC00000000CC0FFF0FFF";
    attribute INIT_18 of inst : label is "0000FFF0000000020030003000000003080020000000D6000000025701080000";
    attribute INIT_19 of inst : label is "00000000000000000000000000000000000000000FFF0FFF0FFD00BF07FF03FF";
    attribute INIT_1A of inst : label is "000003FF0000000000000001000000000000021F000000000000000300000257";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000CC00003FFF00000052";
    attribute INIT_1C of inst : label is "0000200000004000000000100000F40000000640000014000000D60000000000";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000000CC00000050000000D0000000FF00";
    attribute INIT_1E of inst : label is "20000000080000000500DA00F800C000E7F4DB703FC03C000800200000000000";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFC0FFC02D00FFC0FFD0FFC000000000";
    attribute INIT_20 of inst : label is "03C0001700000FF500F0F5000000D7FC00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "07F000F800070FFF43D08B40FC00FFFC0FC0017F00003FF500FCFF500000D7FF";
    attribute INIT_22 of inst : label is "FFEA3F00017F0000BFAF003DFF40000003F500E000001FA07FFF200F55500000";
    attribute INIT_23 of inst : label is "005F000000003C00FD4000000000003DABFF03FC00170000541F002CFF4002FF";
    attribute INIT_24 of inst : label is "2F001FEA001502FF003EEAFD5500FFE00FC0007F00073FFF00F4F500F000FFFF";
    attribute INIT_25 of inst : label is "000000000000001500000000000055EA00D00FE03D57000B41F082FEFFFFFE00";
    attribute INIT_26 of inst : label is "00A30003000017AFFF28FD007C01EF4001CF000B0007007FFCD0F8007400FF40";
    attribute INIT_27 of inst : label is "00A300030000007BFF28FD007C01EF40000300030000017BFF00FD007C01FE00";
    attribute INIT_28 of inst : label is "00000000000002AB000000000000FAA00ADD845C14301831177015018C01E004";
    attribute INIT_29 of inst : label is "003F0C00000003A0FF00400C000002B0003F0C00000003A0FF00400C000002B0";
    attribute INIT_2A of inst : label is "003F0400000006BEFF0000040000AFA4001F009701A003807D00F580029000B0";
    attribute INIT_2B of inst : label is "00DC0054240618243740952024438389002F00C1000D0380BE00D0C01C0000B0";
    attribute INIT_2C of inst : label is "0000000C0010000000000C000100000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000030300000103400000024000000000000060000000000";
    attribute INIT_2E of inst : label is "000000000000003C00A0022052D0000000000000000001400010011056D00003";
    attribute INIT_2F of inst : label is "00000000000000000000008B04F401C00000000000002AA0005400444AD00000";
    attribute INIT_30 of inst : label is "00000000000000010000000000000000200000000000003800020000D0020000";
    attribute INIT_31 of inst : label is "0000002000000000000042000000000000000030000000000000030000000000";
    attribute INIT_32 of inst : label is "00000000000500000000000004000000000000000000000000D0A00000000000";
    attribute INIT_33 of inst : label is "00000000000000000000A000000000000100000000008000001034000000000B";
    attribute INIT_34 of inst : label is "000000C00000000000000C000000000000000000000000000000000050400000";
    attribute INIT_35 of inst : label is "000100000000003ED80000000000AF0085DCA95700240800370B150003803000";
    attribute INIT_36 of inst : label is "08FF0001004000BFFFC8D0000040FF8001FF0401005000BFFFD0D0040140FF80";
    attribute INIT_37 of inst : label is "0DFFC00000000BFFFC1000000000FFE009FF6900000003FFFC1000000000FFA0";
    attribute INIT_38 of inst : label is "01FF042F005101FFFFD0FE045140FFD00BFF680000001FFFFC1000000000FFF0";
    attribute INIT_39 of inst : label is "00000000000000000000000000000000000C005400C006030C50542030600841";
    attribute INIT_3A of inst : label is "00000000000000000000000000007FFC00000000000000000000000000000000";
    attribute INIT_3B of inst : label is "00000000000000000000000000000000000000000000FC000100000000003FC0";
    attribute INIT_3C of inst : label is "C3C3F0143C00F2FFC30F03140F0003FE003F003C000F002F08300FD4C2A0FFF0";
    attribute INIT_3D of inst : label is "000000000000000000000000000000003C331C35017A000038000500AA000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
