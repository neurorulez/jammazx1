library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity travusa_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of travusa_cpu is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"F3",X"31",X"00",X"E8",X"ED",X"56",X"3A",X"04",X"D0",X"A7",X"F2",X"D0",X"05",X"DD",
		X"21",X"75",X"07",X"CD",X"94",X"06",X"A7",X"C2",X"3C",X"00",X"C3",X"9B",X"56",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"80",X"56",X"F3",X"76",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F3",X"76",X"72",X"00",X"81",X"00",X"95",X"00",X"A5",X"00",
		X"B3",X"00",X"4B",X"06",X"BA",X"BB",X"00",X"B6",X"B7",X"B8",X"B9",X"00",X"10",X"B6",X"10",X"BC",
		X"01",X"4B",X"06",X"BA",X"BB",X"00",X"B6",X"B7",X"B8",X"B9",X"00",X"10",X"B6",X"B7",X"B8",X"B9",
		X"00",X"06",X"BA",X"BB",X"01",X"4B",X"04",X"BA",X"BB",X"00",X"B7",X"BD",X"BE",X"BF",X"00",X"C0",
		X"C0",X"C1",X"10",X"BF",X"01",X"4B",X"B6",X"10",X"BC",X"00",X"B6",X"B7",X"B8",X"B9",X"00",X"06",
		X"BA",X"BB",X"01",X"5B",X"C0",X"C0",X"C1",X"10",X"BF",X"00",X"10",X"B7",X"BD",X"BE",X"BF",X"00",
		X"04",X"BA",X"BB",X"01",X"01",X"02",X"03",X"05",X"06",X"07",X"09",X"0A",X"0C",X"0E",X"0F",X"10",
		X"E0",X"00",X"0C",X"01",X"22",X"01",X"39",X"01",X"4F",X"01",X"6A",X"01",X"7D",X"01",X"96",X"01",
		X"40",X"01",X"C1",X"A1",X"C1",X"A1",X"E1",X"A1",X"C1",X"A1",X"C1",X"14",X"05",X"E1",X"A1",X"C1",
		X"A1",X"C1",X"C1",X"A1",X"C1",X"15",X"0E",X"1D",X"06",X"A1",X"C1",X"A1",X"C1",X"14",X"0E",X"1D",
		X"0B",X"A1",X"C1",X"A1",X"C1",X"15",X"0E",X"1C",X"10",X"A1",X"C1",X"00",X"40",X"1D",X"4D",X"86",
		X"41",X"1E",X"C1",X"A1",X"C1",X"49",X"22",X"49",X"23",X"A1",X"49",X"25",X"C1",X"A1",X"4D",X"28",
		X"A1",X"00",X"44",X"2A",X"A1",X"C1",X"81",X"81",X"C1",X"15",X"05",X"48",X"30",X"A1",X"48",X"90",
		X"41",X"32",X"4D",X"33",X"A1",X"4E",X"35",X"C1",X"00",X"40",X"37",X"C1",X"4A",X"39",X"81",X"48",
		X"3B",X"A1",X"C1",X"A1",X"49",X"3F",X"4D",X"94",X"41",X"40",X"52",X"9A",X"41",X"0E",X"00",X"40",
		X"41",X"49",X"42",X"81",X"C1",X"A1",X"48",X"8B",X"41",X"46",X"C1",X"41",X"8E",X"49",X"91",X"44",
		X"C8",X"4A",X"95",X"44",X"49",X"52",X"90",X"41",X"4A",X"00",X"44",X"4B",X"A1",X"52",X"4D",X"81",
		X"49",X"4F",X"49",X"50",X"A1",X"4D",X"52",X"A1",X"52",X"9B",X"44",X"54",X"00",X"40",X"55",X"49",
		X"56",X"81",X"C1",X"81",X"81",X"49",X"5B",X"49",X"92",X"41",X"0E",X"4D",X"96",X"41",X"8E",X"1C",
		X"0B",X"41",X"5C",X"52",X"5D",X"00",X"40",X"5E",X"49",X"5F",X"49",X"60",X"81",X"81",X"49",X"63",
		X"4D",X"06",X"41",X"64",X"4E",X"65",X"52",X"EC",X"00",X"35",X"03",X"44",X"4D",X"43",X"03",X"44",
		X"4D",X"48",X"03",X"44",X"C3",X"4B",X"03",X"34",X"C3",X"E1",X"01",X"A8",X"80",X"16",X"02",X"48",
		X"80",X"3B",X"02",X"88",X"80",X"67",X"02",X"78",X"80",X"9D",X"02",X"8B",X"80",X"E8",X"02",X"7B",
		X"80",X"54",X"03",X"44",X"CD",X"61",X"03",X"44",X"CD",X"69",X"03",X"44",X"CD",X"77",X"03",X"44",
		X"CD",X"81",X"A9",X"66",X"AE",X"82",X"AF",X"A8",X"08",X"29",X"B2",X"81",X"B1",X"29",X"B6",X"81",
		X"B5",X"29",X"B6",X"81",X"B9",X"29",X"B6",X"81",X"BC",X"23",X"B6",X"82",X"C4",X"C3",X"24",X"B6",
		X"81",X"BF",X"23",X"A6",X"82",X"C6",X"C5",X"24",X"A6",X"81",X"C2",X"23",X"B6",X"82",X"C8",X"C7",
		X"24",X"B6",X"19",X"81",X"BF",X"00",X"90",X"B0",X"AF",X"AB",X"AA",X"B4",X"B3",X"B2",X"B2",X"B8",
		X"B7",X"B6",X"B6",X"BB",X"BA",X"B6",X"B6",X"8E",X"BE",X"BD",X"B6",X"B6",X"B4",X"C1",X"C0",X"B6",
		X"B8",X"CA",X"C9",X"A6",X"BB",X"CB",X"19",X"82",X"C0",X"B6",X"00",X"66",X"D1",X"81",X"A8",X"08",
		X"27",X"B2",X"81",X"B1",X"27",X"B6",X"81",X"B5",X"27",X"B6",X"81",X"B9",X"27",X"B6",X"84",X"BC",
		X"B6",X"C4",X"C3",X"24",X"B6",X"84",X"BF",X"A6",X"C6",X"C5",X"24",X"A6",X"84",X"C2",X"B6",X"C8",
		X"C7",X"24",X"B6",X"19",X"81",X"BF",X"00",X"62",X"D5",X"63",X"CF",X"62",X"D3",X"83",X"D6",X"B4",
		X"B3",X"24",X"B6",X"83",X"D7",X"B8",X"B7",X"24",X"B6",X"83",X"D8",X"BB",X"BA",X"24",X"B6",X"83",
		X"D9",X"BE",X"BD",X"24",X"B6",X"84",X"D6",X"B4",X"C1",X"C0",X"23",X"B6",X"84",X"D7",X"B8",X"CA",
		X"C9",X"23",X"A6",X"83",X"D8",X"BB",X"CB",X"19",X"81",X"C0",X"23",X"B6",X"00",X"66",X"D1",X"81",
		X"A8",X"08",X"63",X"DD",X"64",X"DD",X"9F",X"EC",X"EE",X"ED",X"B6",X"EE",X"ED",X"B6",X"E6",X"EC",
		X"F0",X"EF",X"B6",X"F0",X"EF",X"B6",X"E7",X"EC",X"F2",X"F1",X"B6",X"F2",X"F1",X"B6",X"E8",X"EC",
		X"C3",X"B6",X"B6",X"C4",X"C3",X"B6",X"92",X"E9",X"EC",X"C5",X"F7",X"F7",X"F3",X"C5",X"F7",X"EA",
		X"EC",X"F4",X"F6",X"F6",X"F5",X"F4",X"F6",X"EB",X"EC",X"26",X"F6",X"82",X"F8",X"EC",X"26",X"F6",
		X"82",X"F9",X"EC",X"27",X"FA",X"81",X"EC",X"00",X"62",X"D5",X"63",X"CF",X"62",X"D3",X"84",X"D6",
		X"B4",X"DE",X"DB",X"63",X"DD",X"87",X"D7",X"B8",X"DF",X"B6",X"EE",X"ED",X"B6",X"87",X"D8",X"BB",
		X"E0",X"E2",X"F0",X"EF",X"B6",X"87",X"D9",X"BE",X"E1",X"E3",X"F2",X"F1",X"B6",X"87",X"D6",X"B4",
		X"E1",X"E4",X"B6",X"B6",X"C4",X"87",X"D7",X"B8",X"E1",X"E5",X"F7",X"F7",X"F3",X"83",X"D8",X"BB",
		X"E1",X"23",X"F6",X"84",X"F5",X"D9",X"BE",X"E1",X"24",X"F6",X"83",X"D6",X"B4",X"E1",X"24",X"F6",
		X"63",X"FD",X"24",X"FA",X"00",X"88",X"5A",X"5E",X"63",X"64",X"66",X"6C",X"70",X"74",X"44",X"7C",
		X"44",X"81",X"00",X"47",X"85",X"49",X"8D",X"00",X"50",X"A0",X"00",X"46",X"D8",X"08",X"42",X"DF",
		X"08",X"42",X"E2",X"00",X"44",X"F0",X"14",X"84",X"66",X"6C",X"70",X"74",X"44",X"7C",X"44",X"81",
		X"00",X"44",X"F4",X"14",X"43",X"89",X"49",X"8D",X"00",X"44",X"F0",X"14",X"84",X"66",X"6C",X"70",
		X"74",X"44",X"7C",X"1C",X"44",X"F8",X"00",X"44",X"F4",X"14",X"43",X"89",X"45",X"8D",X"1C",X"44",
		X"FC",X"00",X"8C",X"03",X"FA",X"03",X"5D",X"04",X"C2",X"04",X"38",X"05",X"84",X"18",X"00",X"18",
		X"18",X"00",X"69",X"6A",X"00",X"6B",X"6C",X"6D",X"6E",X"00",X"6F",X"70",X"71",X"72",X"00",X"F1",
		X"6F",X"70",X"F1",X"73",X"F1",X"72",X"00",X"6B",X"6C",X"F1",X"74",X"F1",X"6E",X"F1",X"00",X"75",
		X"76",X"00",X"77",X"78",X"00",X"79",X"7A",X"7B",X"7C",X"00",X"7D",X"7E",X"7F",X"80",X"00",X"81",
		X"82",X"83",X"84",X"00",X"18",X"85",X"00",X"86",X"87",X"88",X"00",X"89",X"8A",X"8B",X"8C",X"00",
		X"8D",X"8E",X"00",X"8F",X"90",X"91",X"00",X"F1",X"8D",X"F1",X"92",X"93",X"00",X"94",X"95",X"96",
		X"00",X"97",X"98",X"99",X"9A",X"00",X"F1",X"97",X"F1",X"9B",X"9C",X"9D",X"00",X"9E",X"9F",X"A0",
		X"A1",X"00",X"A2",X"A3",X"A4",X"A5",X"00",X"18",X"7C",X"00",X"85",X"01",X"00",X"02",X"03",X"04",
		X"00",X"02",X"05",X"01",X"01",X"00",X"06",X"02",X"02",X"02",X"00",X"07",X"08",X"5A",X"5A",X"00",
		X"09",X"0A",X"0B",X"0C",X"00",X"02",X"0D",X"0E",X"00",X"0F",X"10",X"11",X"12",X"00",X"02",X"13",
		X"14",X"00",X"15",X"16",X"00",X"17",X"14",X"00",X"19",X"01",X"00",X"19",X"02",X"1A",X"00",X"1B",
		X"02",X"1C",X"00",X"15",X"F1",X"06",X"01",X"01",X"F1",X"00",X"17",X"06",X"02",X"02",X"00",X"02",
		X"5A",X"5A",X"5A",X"00",X"15",X"01",X"00",X"17",X"02",X"16",X"00",X"06",X"02",X"14",X"00",X"01",
		X"08",X"00",X"02",X"0A",X"16",X"00",X"1B",X"15",X"14",X"00",X"15",X"17",X"00",X"85",X"2F",X"3A",
		X"3A",X"00",X"31",X"5A",X"5A",X"00",X"09",X"2F",X"00",X"3A",X"31",X"00",X"2A",X"55",X"00",X"2A",
		X"04",X"00",X"09",X"38",X"38",X"00",X"2F",X"3A",X"3A",X"00",X"31",X"5A",X"5A",X"00",X"38",X"38",
		X"00",X"3A",X"3A",X"38",X"38",X"00",X"39",X"39",X"3A",X"3A",X"00",X"5A",X"5A",X"F4",X"66",X"F4",
		X"5A",X"00",X"2A",X"F4",X"E9",X"67",X"F4",X"00",X"2F",X"F4",X"6D",X"6E",X"F4",X"00",X"31",X"F4",
		X"71",X"72",X"7A",X"F4",X"00",X"2A",X"F4",X"7B",X"7C",X"7F",X"F4",X"00",X"2F",X"38",X"38",X"00",
		X"31",X"3A",X"3A",X"00",X"09",X"2F",X"5A",X"00",X"3A",X"31",X"00",X"5A",X"55",X"00",X"2F",X"00",
		X"31",X"00",X"85",X"1D",X"1E",X"03",X"04",X"00",X"01",X"1F",X"20",X"21",X"22",X"23",X"00",X"02",
		X"24",X"25",X"26",X"27",X"28",X"00",X"29",X"00",X"1E",X"2A",X"00",X"29",X"2B",X"2C",X"00",X"2E",
		X"2D",X"2D",X"00",X"01",X"2F",X"5A",X"00",X"02",X"31",X"00",X"2F",X"32",X"1E",X"03",X"00",X"31",
		X"29",X"5A",X"33",X"00",X"34",X"1E",X"1E",X"2A",X"35",X"00",X"36",X"36",X"36",X"00",X"2C",X"2C",
		X"37",X"00",X"2D",X"2D",X"38",X"38",X"38",X"00",X"2F",X"07",X"3A",X"3A",X"3A",X"00",X"31",X"5A",
		X"5A",X"5A",X"33",X"00",X"02",X"2A",X"35",X"00",X"01",X"3B",X"38",X"38",X"00",X"02",X"3C",X"3D",
		X"3E",X"3F",X"40",X"41",X"00",X"42",X"43",X"44",X"45",X"46",X"30",X"F1",X"41",X"F1",X"00",X"1D",
		X"03",X"04",X"00",X"5A",X"33",X"00",X"2A",X"00",X"86",X"3A",X"3A",X"3A",X"00",X"47",X"5A",X"5A",
		X"00",X"48",X"49",X"00",X"4A",X"F1",X"4B",X"F1",X"4C",X"00",X"4D",X"47",X"4E",X"4F",X"F2",X"4F",
		X"F2",X"00",X"50",X"4B",X"4F",X"47",X"5A",X"00",X"51",X"4B",X"4A",X"33",X"00",X"52",X"4B",X"4D",
		X"00",X"3A",X"39",X"4E",X"4F",X"4F",X"49",X"53",X"00",X"07",X"38",X"38",X"38",X"5A",X"33",X"00",
		X"4B",X"4A",X"3A",X"3A",X"00",X"4B",X"4D",X"39",X"51",X"4B",X"4C",X"00",X"F2",X"4F",X"F2",X"56",
		X"4F",X"47",X"5A",X"33",X"00",X"47",X"5C",X"5C",X"57",X"4B",X"4C",X"54",X"00",X"38",X"38",X"38",
		X"5A",X"5A",X"33",X"00",X"4A",X"3A",X"3A",X"00",X"4D",X"58",X"5A",X"00",X"59",X"5D",X"00",X"F2",
		X"4F",X"F2",X"5D",X"00",X"4E",X"4F",X"49",X"00",X"47",X"5E",X"5F",X"60",X"61",X"62",X"63",X"00",
		X"A7",X"64",X"65",X"66",X"67",X"68",X"00",X"4A",X"5D",X"00",X"4D",X"5D",X"00",X"C0",X"CC",X"A0",
		X"D8",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AF",X"32",X"00",X"90",X"32",X"00",X"A0",X"FD",X"21",X"EC",X"05",X"3E",X"01",X"57",X"06",X"08",
		X"21",X"00",X"E0",X"7A",X"77",X"5E",X"BB",X"28",X"03",X"C3",X"76",X"07",X"2C",X"20",X"F4",X"24",
		X"10",X"F1",X"7A",X"07",X"30",X"E7",X"3E",X"55",X"4F",X"06",X"08",X"21",X"00",X"E0",X"77",X"EE",
		X"FF",X"2C",X"20",X"FA",X"24",X"10",X"F7",X"FD",X"21",X"19",X"06",X"79",X"06",X"08",X"21",X"00",
		X"E0",X"57",X"5E",X"BB",X"28",X"03",X"C3",X"76",X"07",X"EE",X"FF",X"2C",X"20",X"F3",X"24",X"10",
		X"F0",X"79",X"EE",X"FF",X"FE",X"55",X"20",X"D0",X"31",X"00",X"E8",X"3E",X"01",X"57",X"06",X"10",
		X"21",X"00",X"80",X"7A",X"77",X"CD",X"D5",X"07",X"2C",X"20",X"F8",X"24",X"10",X"F5",X"7A",X"07",
		X"30",X"EB",X"3E",X"55",X"4F",X"06",X"10",X"21",X"00",X"80",X"77",X"EE",X"FF",X"2C",X"20",X"FA",
		X"24",X"10",X"F7",X"79",X"06",X"10",X"21",X"00",X"80",X"57",X"CD",X"D5",X"07",X"EE",X"FF",X"2C",
		X"20",X"F7",X"24",X"10",X"F4",X"79",X"EE",X"FF",X"FE",X"55",X"20",X"D8",X"CD",X"29",X"08",X"21",
		X"9E",X"0D",X"CD",X"24",X"07",X"DD",X"21",X"75",X"07",X"CD",X"94",X"06",X"CD",X"17",X"08",X"3E",
		X"FF",X"32",X"FF",X"E0",X"FB",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"3E",X"03",X"32",X"01",
		X"E7",X"C3",X"3E",X"08",X"DD",X"E5",X"DD",X"21",X"75",X"07",X"11",X"00",X"00",X"AF",X"32",X"00",
		X"E7",X"32",X"EF",X"E7",X"CD",X"BB",X"06",X"D1",X"CD",X"BB",X"06",X"D1",X"CD",X"BB",X"06",X"D1",
		X"CD",X"BB",X"06",X"D1",X"3A",X"EF",X"E7",X"DD",X"E1",X"DD",X"E9",X"21",X"00",X"00",X"06",X"20",
		X"1A",X"85",X"30",X"01",X"24",X"6F",X"1C",X"20",X"F7",X"14",X"10",X"F4",X"C1",X"D5",X"C5",X"C3",
		X"D2",X"06",X"E5",X"3A",X"00",X"E7",X"21",X"40",X"47",X"87",X"85",X"6F",X"5E",X"23",X"56",X"E1",
		X"7A",X"BC",X"20",X"09",X"7B",X"BD",X"20",X"05",X"21",X"BC",X"0D",X"18",X"0A",X"3A",X"EF",X"E7",
		X"3C",X"32",X"EF",X"E7",X"21",X"CB",X"0D",X"11",X"82",X"E0",X"01",X"20",X"00",X"ED",X"B0",X"3A",
		X"00",X"E7",X"87",X"87",X"4F",X"3E",X"36",X"91",X"6F",X"26",X"82",X"22",X"80",X"E0",X"FD",X"21",
		X"8C",X"E0",X"3A",X"00",X"E7",X"C6",X"30",X"32",X"85",X"E0",X"21",X"00",X"E7",X"34",X"21",X"80",
		X"E0",X"C3",X"28",X"07",X"DD",X"21",X"75",X"07",X"5E",X"23",X"56",X"23",X"EB",X"01",X"80",X"00",
		X"1A",X"13",X"FE",X"01",X"EB",X"28",X"F1",X"EB",X"38",X"21",X"77",X"09",X"18",X"F2",X"DD",X"21",
		X"75",X"07",X"06",X"02",X"4F",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",
		X"02",X"C6",X"07",X"77",X"11",X"80",X"00",X"19",X"79",X"10",X"EE",X"DD",X"E9",X"F5",X"0F",X"0F",
		X"0F",X"0F",X"CD",X"66",X"07",X"F1",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",
		X"FD",X"77",X"00",X"FD",X"23",X"C9",X"08",X"D9",X"DD",X"21",X"7F",X"07",X"C3",X"2D",X"08",X"21",
		X"A9",X"0D",X"DD",X"21",X"89",X"07",X"C3",X"28",X"07",X"D9",X"7C",X"D9",X"21",X"BA",X"87",X"DD",
		X"21",X"96",X"07",X"C3",X"42",X"07",X"D9",X"7D",X"D9",X"DD",X"21",X"A0",X"07",X"C3",X"42",X"07",
		X"19",X"D9",X"7A",X"D9",X"DD",X"21",X"AB",X"07",X"C3",X"42",X"07",X"19",X"D9",X"7B",X"D9",X"DD",
		X"21",X"B6",X"07",X"C3",X"42",X"07",X"3A",X"00",X"D0",X"CB",X"4F",X"CA",X"75",X"06",X"CB",X"47",
		X"20",X"F4",X"01",X"00",X"20",X"10",X"FE",X"0D",X"20",X"FB",X"3A",X"00",X"D0",X"CB",X"47",X"28",
		X"F4",X"08",X"D9",X"FD",X"E9",X"5E",X"BB",X"C8",X"08",X"D9",X"0E",X"01",X"CD",X"F0",X"07",X"FD",
		X"21",X"E6",X"07",X"C3",X"7F",X"07",X"D9",X"08",X"0E",X"00",X"CD",X"F0",X"07",X"D9",X"08",X"C9",
		X"21",X"20",X"80",X"11",X"00",X"E3",X"CD",X"12",X"08",X"06",X"20",X"7E",X"12",X"36",X"00",X"23",
		X"13",X"10",X"F8",X"CD",X"12",X"08",X"D5",X"11",X"60",X"00",X"19",X"D1",X"7C",X"FE",X"90",X"38",
		X"E5",X"C9",X"0C",X"0D",X"C0",X"EB",X"C9",X"DD",X"21",X"75",X"07",X"21",X"00",X"E0",X"06",X"07",
		X"36",X"00",X"2C",X"20",X"FB",X"24",X"10",X"F8",X"C9",X"DD",X"21",X"75",X"07",X"21",X"00",X"80",
		X"06",X"10",X"7D",X"E6",X"01",X"77",X"2C",X"20",X"F9",X"24",X"10",X"F6",X"DD",X"E9",X"CD",X"29",
		X"08",X"21",X"59",X"10",X"CD",X"24",X"07",X"3A",X"01",X"E7",X"06",X"05",X"CD",X"42",X"0C",X"3A",
		X"00",X"D0",X"CB",X"47",X"20",X"14",X"3A",X"01",X"E7",X"07",X"4F",X"06",X"00",X"DD",X"21",X"DA",
		X"0D",X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"DD",X"21",X"02",X"E7",X"CD",X"17",
		X"0C",X"47",X"E6",X"55",X"FE",X"55",X"28",X"09",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"13",X"18",
		X"CE",X"DD",X"36",X"00",X"55",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"01",X"CD",X"A3",X"08",
		X"18",X"BD",X"DD",X"36",X"00",X"AA",X"DD",X"36",X"01",X"03",X"DD",X"36",X"02",X"FF",X"CD",X"A3",
		X"08",X"18",X"AC",X"DD",X"56",X"00",X"1E",X"02",X"CD",X"02",X"0C",X"28",X"0E",X"CD",X"BF",X"08",
		X"DD",X"56",X"00",X"1E",X"01",X"CD",X"02",X"0C",X"20",X"F3",X"C9",X"CD",X"BF",X"08",X"C9",X"3A",
		X"01",X"E7",X"DD",X"BE",X"01",X"C8",X"06",X"01",X"CD",X"42",X"0C",X"DD",X"86",X"02",X"32",X"01",
		X"E7",X"06",X"05",X"CD",X"42",X"0C",X"C9",X"CD",X"29",X"08",X"21",X"EC",X"0D",X"CD",X"24",X"07",
		X"3A",X"03",X"D0",X"21",X"B2",X"85",X"CD",X"05",X"09",X"3A",X"04",X"D0",X"21",X"AE",X"85",X"CD",
		X"05",X"09",X"21",X"42",X"09",X"CD",X"12",X"09",X"CD",X"BD",X"09",X"3A",X"00",X"D0",X"CB",X"4F",
		X"20",X"DE",X"C3",X"3E",X"08",X"06",X"08",X"0E",X"30",X"0F",X"38",X"01",X"0C",X"71",X"24",X"10",
		X"F6",X"C9",X"7E",X"3C",X"C8",X"3D",X"11",X"03",X"D0",X"FE",X"10",X"38",X"03",X"11",X"04",X"D0",
		X"E6",X"07",X"47",X"1A",X"28",X"03",X"1F",X"10",X"FD",X"2F",X"23",X"A6",X"87",X"23",X"8E",X"5F",
		X"23",X"3E",X"00",X"8E",X"23",X"E5",X"67",X"6B",X"5E",X"23",X"56",X"EB",X"CD",X"24",X"07",X"E1",
		X"18",X"D0",X"00",X"03",X"57",X"09",X"02",X"01",X"77",X"09",X"03",X"01",X"87",X"09",X"11",X"01",
		X"97",X"09",X"13",X"01",X"AF",X"09",X"FF",X"5F",X"09",X"65",X"09",X"6B",X"09",X"71",X"09",X"26",
		X"8A",X"4C",X"4F",X"57",X"00",X"26",X"8A",X"4D",X"45",X"44",X"00",X"26",X"8A",X"48",X"49",X"20",
		X"00",X"26",X"8A",X"4D",X"41",X"58",X"00",X"7B",X"09",X"81",X"09",X"1E",X"8A",X"4C",X"4F",X"57",
		X"00",X"1E",X"8A",X"48",X"49",X"20",X"00",X"8B",X"09",X"91",X"09",X"1A",X"8A",X"4E",X"4F",X"20",
		X"00",X"1A",X"8A",X"59",X"45",X"53",X"00",X"9B",X"09",X"A5",X"09",X"0A",X"89",X"54",X"41",X"42",
		X"4C",X"45",X"20",X"20",X"00",X"0A",X"89",X"55",X"50",X"52",X"49",X"47",X"48",X"54",X"00",X"B3",
		X"09",X"B8",X"09",X"16",X"8A",X"5E",X"5F",X"00",X"16",X"8A",X"5B",X"5C",X"00",X"CD",X"52",X"0A",
		X"3A",X"04",X"D0",X"CB",X"57",X"CA",X"F6",X"09",X"CD",X"3F",X"0A",X"CD",X"34",X"0A",X"FE",X"08",
		X"30",X"12",X"FE",X"06",X"30",X"18",X"C6",X"31",X"32",X"82",X"E0",X"D6",X"31",X"28",X"46",X"21",
		X"87",X"E0",X"18",X"3F",X"E6",X"07",X"FE",X"07",X"28",X"44",X"FE",X"05",X"38",X"2D",X"06",X"0D",
		X"21",X"12",X"89",X"C3",X"49",X"0A",X"CD",X"34",X"0A",X"E6",X"03",X"FE",X"03",X"28",X"2C",X"CD",
		X"D6",X"09",X"21",X"7E",X"0A",X"CD",X"24",X"07",X"CD",X"34",X"0A",X"1F",X"1F",X"E6",X"03",X"FE",
		X"02",X"DE",X"FF",X"CD",X"52",X"0A",X"21",X"80",X"E0",X"36",X"0E",X"C6",X"32",X"32",X"89",X"E0",
		X"21",X"8E",X"E0",X"36",X"53",X"21",X"80",X"E0",X"C3",X"24",X"07",X"CD",X"3F",X"0A",X"21",X"6E",
		X"0A",X"C3",X"24",X"07",X"3A",X"03",X"D0",X"1F",X"1F",X"1F",X"1F",X"2F",X"E6",X"0F",X"C9",X"21",
		X"92",X"87",X"36",X"00",X"21",X"0E",X"82",X"06",X"1B",X"11",X"80",X"00",X"36",X"00",X"19",X"10",
		X"FB",X"C9",X"21",X"5E",X"0A",X"11",X"80",X"E0",X"01",X"10",X"00",X"ED",X"B0",X"C9",X"12",X"89",
		X"31",X"43",X"4F",X"49",X"4E",X"20",X"20",X"31",X"50",X"4C",X"41",X"59",X"20",X"00",X"12",X"89",
		X"20",X"46",X"52",X"45",X"45",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"92",X"87",
		X"41",X"01",X"0E",X"82",X"43",X"4F",X"49",X"4E",X"20",X"4D",X"4F",X"44",X"45",X"20",X"20",X"42",
		X"00",X"AF",X"32",X"0F",X"E7",X"67",X"6F",X"22",X"0D",X"E7",X"CD",X"29",X"08",X"21",X"7E",X"0E",
		X"CD",X"24",X"07",X"3A",X"00",X"D0",X"21",X"B2",X"85",X"CD",X"05",X"09",X"3A",X"01",X"D0",X"21",
		X"AE",X"85",X"CD",X"05",X"09",X"3A",X"02",X"D0",X"21",X"AA",X"85",X"CD",X"05",X"09",X"CD",X"E9",
		X"0A",X"3A",X"0D",X"E7",X"21",X"26",X"86",X"CD",X"3E",X"07",X"3A",X"0E",X"E7",X"CD",X"3E",X"07",
		X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"CC",X"3A",X"01",X"D0",X"CB",X"4F",X"20",X"C5",X"CD",X"29",
		X"08",X"3E",X"01",X"CD",X"58",X"0C",X"C3",X"3E",X"08",X"21",X"0F",X"E7",X"3A",X"22",X"E0",X"E6",
		X"C0",X"BE",X"C8",X"32",X"0F",X"E7",X"3A",X"0E",X"E7",X"C6",X"01",X"27",X"32",X"0E",X"E7",X"D0",
		X"3A",X"0D",X"E7",X"C6",X"01",X"27",X"32",X"0D",X"E7",X"C9",X"2A",X"AD",X"0E",X"22",X"06",X"E7",
		X"21",X"C2",X"0E",X"FD",X"21",X"AF",X"0E",X"CD",X"1D",X"0B",X"C3",X"3E",X"08",X"FD",X"22",X"0B",
		X"E7",X"E5",X"CD",X"29",X"08",X"E1",X"CD",X"24",X"07",X"DD",X"21",X"08",X"E7",X"3E",X"01",X"32",
		X"05",X"E7",X"06",X"05",X"CD",X"49",X"0C",X"3E",X"01",X"0E",X"40",X"CD",X"5A",X"0C",X"CD",X"CF",
		X"0B",X"CD",X"D2",X"0B",X"3E",X"FF",X"32",X"11",X"E7",X"3A",X"00",X"D0",X"CB",X"4F",X"28",X"4A",
		X"CD",X"2C",X"0C",X"E6",X"AA",X"FE",X"2A",X"28",X"13",X"CD",X"17",X"0C",X"47",X"E6",X"55",X"FE",
		X"55",X"28",X"11",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"1D",X"18",X"DD",X"CD",X"CF",X"0B",X"CD",
		X"D2",X"0B",X"18",X"D5",X"DD",X"36",X"00",X"55",X"3A",X"06",X"E7",X"DD",X"77",X"01",X"DD",X"36",
		X"02",X"01",X"CD",X"AC",X"0B",X"18",X"C2",X"DD",X"36",X"00",X"AA",X"3A",X"07",X"E7",X"DD",X"77",
		X"01",X"DD",X"36",X"02",X"FF",X"CD",X"AC",X"0B",X"18",X"AF",X"CD",X"CF",X"0B",X"3E",X"01",X"0E",
		X"20",X"CD",X"5A",X"0C",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"9E",X"C9",X"CD",X"CF",X"0B",X"DD",
		X"56",X"00",X"1E",X"02",X"CD",X"02",X"0C",X"28",X"0F",X"CD",X"EA",X"0B",X"DD",X"56",X"00",X"1E",
		X"01",X"CD",X"02",X"0C",X"20",X"F3",X"18",X"03",X"CD",X"EA",X"0B",X"CD",X"D2",X"0B",X"C9",X"AF",
		X"18",X"0F",X"3A",X"05",X"E7",X"4F",X"06",X"00",X"FD",X"2A",X"0B",X"E7",X"FD",X"09",X"FD",X"7E",
		X"00",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"C9",X"3A",X"05",X"E7",X"DD",X"BE",X"01",
		X"C8",X"06",X"01",X"CD",X"49",X"0C",X"DD",X"86",X"02",X"32",X"05",X"E7",X"06",X"05",X"CD",X"49",
		X"0C",X"C9",X"0E",X"00",X"06",X"0C",X"CD",X"1C",X"0C",X"A2",X"C8",X"10",X"F9",X"0D",X"20",X"F4",
		X"1D",X"20",X"EF",X"3E",X"FF",X"A2",X"C9",X"CD",X"1C",X"0C",X"18",X"1F",X"21",X"10",X"E7",X"3A",
		X"01",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",X"FF",X"C9",X"21",X"11",X"E7",X"3A",
		X"00",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",X"FF",X"F5",X"AF",X"3D",X"20",X"FD",
		X"F1",X"C9",X"4F",X"D6",X"03",X"07",X"3C",X"18",X"01",X"4F",X"87",X"2F",X"D6",X"C8",X"6F",X"26",
		X"82",X"70",X"C6",X"80",X"6F",X"70",X"79",X"C9",X"0E",X"00",X"06",X"00",X"10",X"FE",X"0D",X"20",
		X"F9",X"3D",X"20",X"F4",X"C9",X"C5",X"0E",X"00",X"06",X"00",X"10",X"FE",X"F5",X"3A",X"00",X"D0",
		X"CB",X"4F",X"28",X"09",X"F1",X"0D",X"20",X"F0",X"3D",X"20",X"EB",X"C1",X"C9",X"F1",X"C1",X"06",
		X"01",X"C9",X"CD",X"29",X"08",X"11",X"C0",X"E1",X"21",X"39",X"10",X"01",X"10",X"00",X"ED",X"B0",
		X"11",X"60",X"E1",X"21",X"49",X"10",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"00",X"D0",X"CB",X"4F",
		X"20",X"F9",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"7F",X"01",X"ED",X"B0",X"C3",
		X"3E",X"08",X"AF",X"32",X"11",X"E7",X"18",X"15",X"3A",X"00",X"D0",X"CB",X"4F",X"CA",X"3E",X"08",
		X"CD",X"2C",X"0C",X"E6",X"AA",X"FE",X"2A",X"20",X"EF",X"3A",X"12",X"E7",X"3C",X"32",X"12",X"E7",
		X"FE",X"05",X"30",X"DE",X"21",X"B8",X"0C",X"E5",X"3D",X"28",X"26",X"3D",X"28",X"4B",X"3D",X"28",
		X"56",X"3D",X"28",X"57",X"CD",X"29",X"08",X"21",X"AE",X"81",X"06",X"1A",X"3E",X"41",X"CD",X"F8",
		X"0C",X"21",X"9E",X"81",X"06",X"0A",X"3E",X"30",X"11",X"80",X"00",X"77",X"3C",X"19",X"10",X"FB",
		X"C9",X"21",X"00",X"80",X"E5",X"7C",X"E6",X"0E",X"4F",X"7D",X"E6",X"30",X"B1",X"CB",X"3F",X"6F",
		X"26",X"00",X"11",X"4D",X"0D",X"19",X"7E",X"E1",X"4F",X"87",X"3E",X"1C",X"CE",X"00",X"77",X"23",
		X"79",X"E6",X"0F",X"77",X"CD",X"3F",X"0D",X"18",X"DB",X"0E",X"00",X"21",X"00",X"80",X"36",X"1C",
		X"23",X"71",X"CD",X"3F",X"0D",X"18",X"F7",X"0E",X"01",X"18",X"F0",X"0E",X"0A",X"18",X"EC",X"23",
		X"CB",X"75",X"C8",X"11",X"40",X"00",X"19",X"7C",X"FE",X"90",X"D8",X"E1",X"C9",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"88",X"00",X"01",X"09",X"0A",X"0B",X"81",X"89",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0E",X"A2",X"21",
		X"00",X"80",X"3E",X"03",X"A9",X"4F",X"FE",X"A3",X"20",X"01",X"AF",X"77",X"23",X"36",X"01",X"23",
		X"CB",X"75",X"3E",X"02",X"28",X"EE",X"11",X"40",X"00",X"19",X"7C",X"FE",X"90",X"38",X"E3",X"21",
		X"1E",X"88",X"36",X"A4",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"C3",X"3E",X"08",X"3A",X"82",
		X"52",X"41",X"4D",X"20",X"20",X"20",X"4F",X"4B",X"00",X"3A",X"82",X"52",X"41",X"4D",X"20",X"20",
		X"20",X"4E",X"47",X"20",X"20",X"3A",X"20",X"20",X"20",X"20",X"3A",X"00",X"52",X"4F",X"4D",X"20",
		X"20",X"20",X"4F",X"4B",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"52",X"4F",X"4D",X"20",X"20",
		X"20",X"4E",X"47",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D7",X"08",X"91",X"0A",X"0A",X"0B",X"82",X"0C",X"B2",X"0C",X"6D",X"0D",X"36",X"82",X"44",X"49",
		X"50",X"20",X"53",X"57",X"20",X"31",X"20",X"32",X"20",X"33",X"20",X"34",X"20",X"35",X"20",X"36",
		X"20",X"37",X"20",X"38",X"01",X"32",X"83",X"44",X"53",X"57",X"31",X"01",X"2E",X"83",X"44",X"53",
		X"57",X"32",X"01",X"2A",X"81",X"46",X"55",X"45",X"4C",X"20",X"43",X"4F",X"4E",X"53",X"55",X"4D",
		X"50",X"54",X"49",X"4F",X"4E",X"20",X"41",X"54",X"20",X"43",X"4F",X"4C",X"4C",X"49",X"53",X"49",
		X"4F",X"4E",X"01",X"22",X"81",X"46",X"55",X"45",X"4C",X"20",X"43",X"4F",X"4E",X"53",X"55",X"4D",
		X"50",X"54",X"49",X"4F",X"4E",X"20",X"49",X"4E",X"20",X"52",X"55",X"4E",X"4E",X"49",X"4E",X"47",
		X"01",X"1A",X"81",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"49",X"54",X"59",X"01",X"16",X"81",
		X"53",X"50",X"45",X"45",X"44",X"01",X"12",X"82",X"43",X"4F",X"49",X"4E",X"20",X"4D",X"4F",X"44",
		X"45",X"01",X"0A",X"82",X"42",X"4F",X"44",X"59",X"20",X"54",X"59",X"50",X"45",X"00",X"B6",X"85",
		X"31",X"20",X"32",X"20",X"33",X"20",X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"20",X"38",X"01",
		X"B2",X"82",X"4B",X"45",X"59",X"30",X"01",X"AE",X"82",X"4B",X"45",X"59",X"31",X"01",X"AA",X"82",
		X"4B",X"45",X"59",X"32",X"01",X"A6",X"82",X"54",X"49",X"4D",X"4E",X"47",X"00",X"12",X"01",X"00",
		X"01",X"16",X"17",X"19",X"15",X"13",X"14",X"1F",X"1C",X"1B",X"1D",X"1E",X"1A",X"18",X"20",X"21",
		X"12",X"11",X"3C",X"83",X"53",X"20",X"4F",X"20",X"55",X"20",X"4E",X"20",X"44",X"20",X"53",X"01",
		X"34",X"82",X"30",X"31",X"20",X"48",X"4F",X"52",X"4E",X"20",X"53",X"4F",X"55",X"4E",X"44",X"20",
		X"01",X"32",X"82",X"30",X"32",X"20",X"42",X"52",X"41",X"4B",X"45",X"20",X"53",X"4F",X"55",X"4E",
		X"44",X"01",X"30",X"82",X"30",X"33",X"20",X"53",X"50",X"49",X"4E",X"4E",X"49",X"4E",X"47",X"20",
		X"53",X"4F",X"55",X"4E",X"44",X"01",X"2E",X"82",X"30",X"34",X"20",X"50",X"41",X"53",X"53",X"49",
		X"4E",X"47",X"20",X"53",X"4F",X"55",X"4E",X"44",X"20",X"31",X"01",X"2C",X"82",X"30",X"35",X"20",
		X"43",X"4F",X"55",X"4E",X"54",X"44",X"4F",X"57",X"4E",X"20",X"53",X"4F",X"55",X"4E",X"44",X"01",
		X"2A",X"82",X"30",X"36",X"20",X"41",X"44",X"44",X"2E",X"20",X"46",X"55",X"45",X"4C",X"20",X"53",
		X"4F",X"55",X"4E",X"44",X"01",X"28",X"82",X"30",X"37",X"20",X"4A",X"55",X"4D",X"50",X"49",X"4E",
		X"47",X"20",X"53",X"4F",X"55",X"4E",X"44",X"01",X"26",X"82",X"30",X"38",X"20",X"43",X"4F",X"4C",
		X"4C",X"49",X"53",X"49",X"4F",X"4E",X"20",X"53",X"4F",X"55",X"4E",X"44",X"01",X"24",X"82",X"30",
		X"39",X"20",X"4F",X"50",X"45",X"4E",X"49",X"4E",X"47",X"20",X"4D",X"55",X"53",X"49",X"43",X"01",
		X"22",X"82",X"31",X"30",X"20",X"45",X"4E",X"44",X"49",X"4E",X"47",X"20",X"4D",X"55",X"53",X"49",
		X"43",X"01",X"20",X"82",X"31",X"31",X"20",X"41",X"52",X"52",X"49",X"56",X"41",X"4C",X"20",X"4D",
		X"55",X"53",X"49",X"43",X"01",X"1E",X"82",X"31",X"32",X"20",X"46",X"49",X"4E",X"41",X"4C",X"20",
		X"47",X"4F",X"41",X"4C",X"20",X"4D",X"55",X"53",X"49",X"43",X"01",X"1C",X"82",X"31",X"33",X"20",
		X"43",X"48",X"45",X"43",X"4B",X"50",X"4F",X"49",X"4E",X"54",X"20",X"4D",X"55",X"53",X"49",X"43",
		X"01",X"1A",X"82",X"31",X"34",X"20",X"42",X"47",X"4D",X"20",X"31",X"20",X"20",X"20",X"53",X"54",
		X"52",X"45",X"45",X"54",X"01",X"18",X"82",X"31",X"35",X"20",X"42",X"47",X"4D",X"20",X"32",X"20",
		X"20",X"20",X"52",X"4F",X"55",X"47",X"48",X"20",X"57",X"41",X"59",X"01",X"16",X"82",X"31",X"36",
		X"20",X"42",X"47",X"4D",X"20",X"33",X"20",X"20",X"20",X"48",X"49",X"47",X"48",X"57",X"41",X"59",
		X"01",X"14",X"82",X"31",X"37",X"20",X"57",X"41",X"52",X"4E",X"49",X"4E",X"47",X"20",X"53",X"4F",
		X"55",X"4E",X"44",X"01",X"12",X"82",X"31",X"38",X"20",X"50",X"41",X"53",X"53",X"49",X"4E",X"47",
		X"20",X"53",X"4F",X"55",X"4E",X"44",X"20",X"32",X"00",X"A8",X"C1",X"7C",X"60",X"A8",X"81",X"7C",
		X"98",X"90",X"41",X"7C",X"60",X"90",X"01",X"7C",X"98",X"68",X"C1",X"7C",X"60",X"68",X"81",X"7C",
		X"98",X"50",X"41",X"7C",X"60",X"50",X"01",X"7C",X"98",X"34",X"82",X"30",X"31",X"20",X"20",X"44",
		X"49",X"50",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"01",X"30",X"82",X"30",X"32",X"20",X"20",
		X"49",X"3D",X"4F",X"20",X"50",X"4F",X"41",X"54",X"01",X"2C",X"82",X"30",X"33",X"20",X"20",X"53",
		X"4F",X"55",X"4E",X"44",X"53",X"01",X"28",X"82",X"30",X"34",X"20",X"20",X"43",X"48",X"41",X"52",
		X"41",X"43",X"54",X"45",X"52",X"01",X"24",X"82",X"30",X"35",X"20",X"20",X"43",X"4F",X"4C",X"4F",
		X"52",X"01",X"20",X"82",X"30",X"36",X"20",X"20",X"43",X"52",X"4F",X"53",X"53",X"20",X"48",X"41",
		X"54",X"43",X"48",X"20",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"A2",X"8C",X"A3",X"8C",X"96",X"00",X"02",X"A2",X"8C",X"96",X"C1",X"0C",X"00",X"8C",X"96",
		X"01",X"CC",X"00",X"C2",X"2F",X"01",X"8C",X"00",X"42",X"0C",X"C2",X"2F",X"00",X"0E",X"A5",X"8E",
		X"A5",X"0E",X"92",X"8E",X"92",X"00",X"0E",X"A5",X"0E",X"92",X"00",X"02",X"0D",X"82",X"2F",X"00",
		X"02",X"0D",X"42",X"2F",X"00",X"02",X"0D",X"C2",X"21",X"00",X"22",X"24",X"42",X"28",X"9B",X"2A",
		X"00",X"22",X"25",X"52",X"29",X"B2",X"28",X"00",X"0A",X"2A",X"92",X"2A",X"A2",X"25",X"00",X"32",
		X"2A",X"AC",X"2B",X"27",X"26",X"66",X"26",X"00",X"22",X"26",X"5C",X"2B",X"C7",X"27",X"00",X"0C",
		X"2B",X"A2",X"29",X"06",X"27",X"00",X"32",X"25",X"52",X"29",X"C2",X"22",X"00",X"22",X"15",X"99",
		X"10",X"00",X"0A",X"2A",X"82",X"26",X"C2",X"24",X"00",X"32",X"15",X"62",X"11",X"C2",X"16",X"00",
		X"52",X"28",X"92",X"25",X"00",X"52",X"12",X"A2",X"0F",X"00",X"22",X"13",X"52",X"17",X"C2",X"13",
		X"00",X"02",X"11",X"32",X"17",X"99",X"10",X"00",X"08",X"10",X"C7",X"10",X"00",X"06",X"10",X"00",
		X"32",X"15",X"C2",X"0D",X"00",X"02",X"12",X"72",X"11",X"A2",X"0D",X"00",X"08",X"10",X"92",X"16",
		X"C2",X"12",X"00",X"12",X"24",X"42",X"28",X"9B",X"2A",X"00",X"42",X"12",X"82",X"16",X"00",X"42",
		X"27",X"92",X"2A",X"00",X"32",X"25",X"52",X"29",X"C2",X"22",X"00",X"0A",X"2A",X"82",X"28",X"C2",
		X"24",X"00",X"82",X"2F",X"00",X"02",X"06",X"82",X"2A",X"00",X"12",X"07",X"00",X"12",X"14",X"00",
		X"22",X"12",X"A2",X"16",X"A2",X"21",X"00",X"52",X"26",X"92",X"29",X"00",X"12",X"25",X"B2",X"26",
		X"C2",X"16",X"00",X"02",X"24",X"62",X"10",X"92",X"14",X"00",X"02",X"08",X"82",X"2A",X"00",X"02",
		X"08",X"00",X"8E",X"A5",X"00",X"42",X"2F",X"00",X"8E",X"92",X"00",X"45",X"21",X"B5",X"22",X"24",
		X"15",X"B5",X"14",X"00",X"15",X"21",X"A5",X"22",X"35",X"14",X"C5",X"16",X"00",X"34",X"22",X"B4",
		X"21",X"24",X"15",X"B4",X"16",X"00",X"04",X"23",X"B4",X"21",X"44",X"16",X"84",X"15",X"00",X"15",
		X"21",X"65",X"24",X"C5",X"23",X"25",X"16",X"75",X"15",X"C5",X"15",X"00",X"15",X"21",X"74",X"22",
		X"B5",X"21",X"04",X"16",X"65",X"15",X"B5",X"16",X"00",X"04",X"23",X"54",X"23",X"B4",X"22",X"24",
		X"15",X"74",X"16",X"C4",X"17",X"00",X"44",X"21",X"84",X"20",X"C4",X"20",X"04",X"16",X"44",X"13",
		X"84",X"15",X"00",X"05",X"21",X"45",X"22",X"85",X"20",X"C5",X"23",X"05",X"16",X"45",X"17",X"85",
		X"16",X"C5",X"16",X"00",X"05",X"22",X"45",X"21",X"85",X"24",X"C5",X"23",X"05",X"14",X"45",X"13",
		X"85",X"14",X"C5",X"14",X"00",X"04",X"23",X"44",X"24",X"84",X"23",X"C4",X"23",X"04",X"14",X"44",
		X"15",X"84",X"13",X"C4",X"15",X"00",X"04",X"20",X"44",X"23",X"84",X"20",X"C4",X"21",X"04",X"17",
		X"44",X"17",X"84",X"13",X"C4",X"15",X"00",X"15",X"21",X"75",X"22",X"15",X"17",X"55",X"16",X"B5",
		X"14",X"00",X"14",X"21",X"65",X"22",X"C4",X"21",X"45",X"16",X"A4",X"16",X"00",X"24",X"21",X"84",
		X"23",X"64",X"16",X"00",X"24",X"21",X"24",X"16",X"00",X"25",X"21",X"95",X"21",X"25",X"15",X"85",
		X"15",X"C5",X"16",X"00",X"05",X"21",X"64",X"22",X"B5",X"21",X"04",X"17",X"45",X"14",X"A5",X"16",
		X"00",X"24",X"22",X"84",X"24",X"C4",X"21",X"14",X"14",X"B4",X"15",X"00",X"44",X"24",X"A4",X"21",
		X"04",X"16",X"54",X"12",X"A4",X"14",X"00",X"03",X"27",X"43",X"28",X"73",X"24",X"C3",X"25",X"00",
		X"03",X"25",X"43",X"26",X"93",X"24",X"B3",X"28",X"00",X"75",X"24",X"34",X"17",X"00",X"24",X"23",
		X"A4",X"24",X"05",X"16",X"85",X"17",X"00",X"F4",X"20",X"F5",X"AF",X"30",X"4A",X"00",X"90",X"78",
		X"FE",X"A8",X"1A",X"FE",X"AB",X"1A",X"A0",X"00",X"A0",X"00",X"FC",X"90",X"79",X"10",X"5A",X"78",
		X"90",X"00",X"FF",X"F0",X"00",X"20",X"20",X"1F",X"1D",X"1C",X"18",X"14",X"10",X"0C",X"08",X"04",
		X"02",X"00",X"F5",X"AF",X"F1",X"09",X"67",X"65",X"5F",X"5C",X"58",X"58",X"58",X"00",X"F6",X"78",
		X"F7",X"AF",X"09",X"4A",X"00",X"E4",X"09",X"07",X"05",X"02",X"03",X"4B",X"79",X"07",X"4A",X"00",
		X"E3",X"09",X"0C",X"0A",X"C3",X"4B",X"08",X"06",X"03",X"83",X"00",X"05",X"4A",X"00",X"E3",X"09",
		X"0C",X"0A",X"C2",X"4B",X"08",X"0B",X"86",X"00",X"03",X"4A",X"78",X"E3",X"10",X"0E",X"0A",X"C2",
		X"4B",X"08",X"0B",X"88",X"00",X"83",X"79",X"E3",X"11",X"0F",X"0B",X"98",X"00",X"82",X"78",X"8E",
		X"00",X"FC",X"82",X"78",X"FC",X"88",X"00",X"E3",X"29",X"08",X"75",X"8B",X"00",X"E3",X"29",X"08",
		X"0B",X"87",X"00",X"82",X"78",X"84",X"00",X"81",X"2A",X"89",X"00",X"FC",X"82",X"78",X"FC",X"99",
		X"00",X"C5",X"4F",X"09",X"07",X"23",X"7A",X"7A",X"89",X"00",X"E3",X"26",X"24",X"22",X"84",X"7B",
		X"89",X"00",X"E2",X"27",X"25",X"85",X"7B",X"89",X"00",X"E1",X"28",X"FC",X"86",X"7A",X"FC",X"02",
		X"4B",X"78",X"8E",X"00",X"FC",X"82",X"78",X"4E",X"5B",X"00",X"90",X"79",X"10",X"5A",X"78",X"10",
		X"5A",X"00",X"F5",X"57",X"F6",X"78",X"F7",X"AF",X"FE",X"A8",X"1A",X"FE",X"E2",X"17",X"FC",X"90",
		X"7A",X"60",X"5B",X"00",X"FE",X"DA",X"13",X"F5",X"57",X"F6",X"78",X"F2",X"09",X"79",X"7C",X"80",
		X"84",X"86",X"88",X"88",X"00",X"F7",X"AF",X"F3",X"09",X"B2",X"B6",X"BA",X"BD",X"BE",X"BE",X"BE",
		X"00",X"FE",X"A8",X"1A",X"FE",X"E2",X"17",X"08",X"6D",X"78",X"E2",X"01",X"04",X"86",X"00",X"88",
		X"7B",X"C1",X"6F",X"A0",X"01",X"2F",X"EF",X"C2",X"6D",X"07",X"09",X"84",X"00",X"8B",X"7B",X"E5",
		X"22",X"0E",X"10",X"78",X"78",X"40",X"5B",X"00",X"88",X"79",X"E3",X"11",X"0F",X"0B",X"85",X"00",
		X"08",X"5A",X"78",X"E2",X"10",X"0E",X"C6",X"5B",X"0A",X"08",X"06",X"03",X"00",X"00",X"0A",X"5A",
		X"00",X"E4",X"09",X"07",X"05",X"02",X"02",X"5B",X"79",X"F5",X"57",X"F6",X"88",X"F7",X"BF",X"FE",
		X"A8",X"1A",X"FE",X"E2",X"17",X"FE",X"C6",X"1A",X"A0",X"00",X"A0",X"00",X"10",X"5B",X"79",X"FF",
		X"F5",X"BF",X"F7",X"BF",X"F1",X"00",X"57",X"57",X"5A",X"5F",X"00",X"F2",X"00",X"88",X"88",X"85",
		X"80",X"00",X"FE",X"A8",X"1A",X"40",X"4F",X"00",X"E4",X"7A",X"7A",X"2B",X"2C",X"FE",X"C6",X"14",
		X"01",X"4F",X"2D",X"FC",X"FE",X"C6",X"14",X"01",X"4F",X"2E",X"8C",X"00",X"03",X"5D",X"00",X"01",
		X"5F",X"2E",X"8C",X"00",X"03",X"5D",X"00",X"01",X"5F",X"2D",X"8C",X"00",X"E4",X"7A",X"7A",X"2B",
		X"2C",X"12",X"4F",X"00",X"84",X"78",X"84",X"00",X"82",X"78",X"FC",X"86",X"00",X"84",X"78",X"84",
		X"00",X"82",X"78",X"FE",X"68",X"14",X"82",X"00",X"84",X"78",X"84",X"00",X"82",X"78",X"03",X"4D",
		X"00",X"FF",X"F5",X"BF",X"FE",X"A8",X"1A",X"FE",X"AB",X"1A",X"FE",X"AB",X"1A",X"FE",X"68",X"14",
		X"FA",X"00",X"F5",X"BF",X"F1",X"0C",X"BD",X"BB",X"B7",X"B4",X"00",X"FE",X"A8",X"1A",X"FE",X"AB",
		X"1A",X"40",X"6B",X"00",X"82",X"78",X"84",X"00",X"84",X"78",X"86",X"00",X"FC",X"82",X"78",X"84",
		X"00",X"84",X"78",X"B4",X"00",X"E2",X"16",X"06",X"8B",X"00",X"E4",X"03",X"06",X"13",X"15",X"C1",
		X"7A",X"05",X"0B",X"7B",X"79",X"C5",X"7A",X"18",X"05",X"12",X"14",X"04",X"FA",X"00",X"F1",X"00",
		X"B1",X"AD",X"A8",X"A3",X"A2",X"9F",X"9C",X"99",X"97",X"94",X"92",X"91",X"90",X"8F",X"8F",X"8F",
		X"00",X"FE",X"A8",X"1A",X"FE",X"AB",X"1A",X"48",X"7B",X"00",X"E5",X"16",X"06",X"13",X"1D",X"1F",
		X"83",X"79",X"85",X"00",X"E4",X"16",X"06",X"13",X"15",X"C4",X"7A",X"05",X"1A",X"1C",X"1E",X"83",
		X"78",X"83",X"7B",X"C3",X"7B",X"0B",X"13",X"15",X"C4",X"7A",X"05",X"12",X"14",X"04",X"86",X"00",
		X"01",X"7B",X"00",X"E2",X"0B",X"08",X"C4",X"7A",X"0A",X"12",X"14",X"04",X"89",X"00",X"01",X"7B",
		X"08",X"C3",X"7A",X"0A",X"0C",X"09",X"89",X"00",X"C3",X"7C",X"30",X"7A",X"7A",X"C2",X"7A",X"07",
		X"09",X"86",X"00",X"C8",X"7C",X"25",X"21",X"1A",X"1C",X"1E",X"2F",X"26",X"00",X"85",X"7B",X"E5",
		X"25",X"21",X"12",X"14",X"04",X"86",X"00",X"F5",X"8F",X"FE",X"A8",X"1A",X"FE",X"AB",X"1A",X"FE",
		X"26",X"13",X"90",X"00",X"10",X"5C",X"7A",X"A0",X"00",X"FA",X"00",X"F0",X"0D",X"02",X"05",X"07",
		X"00",X"F5",X"8F",X"FE",X"DC",X"15",X"FE",X"A8",X"1A",X"FE",X"F1",X"14",X"FA",X"00",X"F0",X"00",
		X"0A",X"0E",X"11",X"17",X"1A",X"1E",X"22",X"25",X"29",X"2C",X"2D",X"2F",X"30",X"30",X"30",X"30",
		X"00",X"F5",X"8F",X"FE",X"DC",X"15",X"FE",X"A8",X"1A",X"FE",X"37",X"15",X"F9",X"00",X"20",X"4C",
		X"00",X"90",X"7A",X"A0",X"7B",X"10",X"4A",X"78",X"FF",X"F4",X"30",X"F5",X"8F",X"FE",X"DE",X"15",
		X"FE",X"A8",X"1A",X"FE",X"26",X"13",X"FE",X"A2",X"15",X"F0",X"00",X"30",X"30",X"30",X"30",X"2F",
		X"2D",X"2B",X"29",X"27",X"25",X"23",X"21",X"1F",X"00",X"F5",X"8F",X"F1",X"0B",X"90",X"92",X"00",
		X"FF",X"FA",X"00",X"F9",X"00",X"FE",X"F9",X"15",X"F0",X"0D",X"70",X"73",X"75",X"00",X"F1",X"0D",
		X"95",X"98",X"9B",X"00",X"F2",X"0D",X"1D",X"1B",X"18",X"00",X"F3",X"0D",X"6D",X"6A",X"67",X"00",
		X"FE",X"50",X"16",X"FA",X"00",X"FE",X"F9",X"15",X"F0",X"0D",X"1D",X"1B",X"18",X"00",X"F1",X"0D",
		X"6D",X"6A",X"67",X"00",X"F2",X"0D",X"70",X"73",X"75",X"00",X"F3",X"0D",X"95",X"98",X"9B",X"00",
		X"20",X"4C",X"00",X"8E",X"7A",X"C2",X"4A",X"50",X"55",X"8B",X"00",X"E5",X"60",X"59",X"58",X"5F",
		X"54",X"87",X"00",X"E5",X"60",X"59",X"58",X"62",X"61",X"84",X"7B",X"84",X"78",X"E5",X"59",X"6A",
		X"68",X"67",X"65",X"87",X"7B",X"03",X"4B",X"79",X"E4",X"6E",X"6D",X"6B",X"69",X"97",X"00",X"C2",
		X"7B",X"06",X"13",X"8D",X"00",X"C1",X"3B",X"EE",X"C1",X"7B",X"6F",X"8A",X"00",X"C1",X"4B",X"6F",
		X"C1",X"0B",X"EE",X"0B",X"4B",X"00",X"E4",X"6F",X"71",X"13",X"06",X"86",X"00",X"82",X"78",X"84",
		X"00",X"E2",X"72",X"16",X"88",X"00",X"02",X"5B",X"78",X"8D",X"00",X"01",X"7B",X"25",X"8D",X"00",
		X"E1",X"57",X"C1",X"7F",X"3F",X"C1",X"7D",X"14",X"0D",X"7B",X"00",X"C1",X"6B",X"25",X"C2",X"6D",
		X"21",X"12",X"20",X"5B",X"00",X"88",X"79",X"C2",X"4B",X"5B",X"5C",X"86",X"00",X"09",X"7A",X"78",
		X"C5",X"5A",X"1E",X"1C",X"1A",X"21",X"25",X"82",X"7B",X"8C",X"00",X"E4",X"04",X"14",X"12",X"21",
		X"8F",X"00",X"E1",X"04",X"10",X"5C",X"7A",X"20",X"0C",X"00",X"FA",X"00",X"F9",X"00",X"F4",X"90",
		X"F0",X"00",X"78",X"7A",X"7D",X"7F",X"82",X"85",X"87",X"8A",X"8C",X"8E",X"8F",X"00",X"F5",X"AF",
		X"F1",X"00",X"9F",X"A2",X"A6",X"AD",X"AD",X"AD",X"AE",X"00",X"F6",X"08",X"F2",X"00",X"14",X"12",
		X"10",X"0E",X"0C",X"0B",X"0A",X"00",X"F7",X"57",X"F3",X"00",X"64",X"61",X"5F",X"5C",X"5A",X"58",
		X"00",X"FE",X"59",X"17",X"FA",X"00",X"F4",X"08",X"F0",X"00",X"14",X"12",X"10",X"0E",X"0C",X"0B",
		X"0A",X"00",X"F5",X"57",X"F1",X"00",X"64",X"61",X"5F",X"5C",X"5A",X"58",X"00",X"F6",X"90",X"F2",
		X"00",X"78",X"7A",X"7D",X"7F",X"82",X"85",X"87",X"8A",X"8C",X"8E",X"8F",X"00",X"F7",X"AF",X"F3",
		X"00",X"9F",X"A2",X"A6",X"AD",X"AD",X"AD",X"AE",X"00",X"06",X"7F",X"7B",X"81",X"30",X"89",X"7A",
		X"E8",X"7B",X"25",X"21",X"1A",X"1C",X"1E",X"2F",X"26",X"88",X"00",X"01",X"4A",X"56",X"C2",X"7F",
		X"78",X"04",X"33",X"6F",X"00",X"84",X"78",X"84",X"00",X"82",X"78",X"C2",X"7D",X"16",X"72",X"04",
		X"7F",X"00",X"84",X"78",X"84",X"00",X"82",X"78",X"E2",X"71",X"6F",X"40",X"7D",X"7B",X"E4",X"25",
		X"21",X"1A",X"1C",X"8A",X"78",X"E4",X"21",X"12",X"14",X"04",X"9C",X"00",X"C2",X"6D",X"14",X"04",
		X"8E",X"00",X"E5",X"25",X"21",X"12",X"14",X"04",X"8B",X"00",X"83",X"7B",X"E5",X"25",X"21",X"12",
		X"14",X"04",X"88",X"00",X"86",X"7B",X"E5",X"25",X"21",X"1A",X"1C",X"1E",X"85",X"78",X"10",X"5A",
		X"7B",X"81",X"25",X"8F",X"7B",X"E3",X"14",X"12",X"22",X"8D",X"7B",X"02",X"5C",X"7A",X"C2",X"5A",
		X"5D",X"56",X"02",X"6F",X"78",X"E2",X"2F",X"26",X"88",X"00",X"86",X"7B",X"81",X"30",X"89",X"7A",
		X"90",X"7B",X"A0",X"00",X"A0",X"00",X"10",X"4F",X"7A",X"A0",X"7B",X"FF",X"F9",X"08",X"10",X"5F",
		X"7B",X"F4",X"90",X"F5",X"AF",X"F6",X"08",X"F7",X"57",X"FE",X"11",X"18",X"F9",X"00",X"F4",X"90",
		X"F5",X"AF",X"F6",X"08",X"F7",X"57",X"FE",X"11",X"18",X"F4",X"08",X"F5",X"57",X"F6",X"90",X"F7",
		X"AF",X"10",X"5F",X"7A",X"FC",X"FE",X"AB",X"1A",X"FE",X"E2",X"17",X"30",X"5F",X"7B",X"90",X"7A",
		X"FE",X"E2",X"17",X"FB",X"08",X"FE",X"2A",X"18",X"F9",X"08",X"F6",X"08",X"F7",X"27",X"FE",X"C7",
		X"18",X"10",X"4D",X"00",X"90",X"78",X"40",X"4F",X"00",X"8E",X"7A",X"C2",X"5F",X"36",X"3B",X"FE",
		X"96",X"18",X"FA",X"00",X"FE",X"C7",X"18",X"F5",X"AF",X"4F",X"5F",X"7B",X"C1",X"5D",X"46",X"8E",
		X"00",X"C1",X"5D",X"46",X"C1",X"5F",X"47",X"FE",X"E4",X"18",X"41",X"4F",X"00",X"90",X"7A",X"90",
		X"7B",X"F9",X"08",X"10",X"5F",X"7B",X"F4",X"60",X"F5",X"AF",X"7F",X"5F",X"7B",X"B1",X"7B",X"90",
		X"7A",X"FC",X"FE",X"AB",X"1A",X"FE",X"E2",X"17",X"FA",X"00",X"FE",X"87",X"18",X"FB",X"08",X"FE",
		X"84",X"18",X"F9",X"08",X"10",X"5F",X"7B",X"FE",X"C7",X"18",X"4F",X"5D",X"00",X"E1",X"46",X"8E",
		X"00",X"E1",X"46",X"C1",X"5F",X"47",X"FE",X"E4",X"18",X"01",X"5F",X"46",X"0E",X"5D",X"7B",X"01",
		X"5F",X"46",X"01",X"5D",X"47",X"8D",X"7B",X"E3",X"43",X"44",X"45",X"8B",X"7B",X"E3",X"40",X"41",
		X"42",X"82",X"00",X"87",X"7B",X"C2",X"5F",X"76",X"35",X"C3",X"5D",X"37",X"38",X"39",X"84",X"00",
		X"87",X"78",X"E2",X"32",X"34",X"97",X"00",X"F4",X"60",X"F0",X"06",X"5F",X"5D",X"5A",X"56",X"52",
		X"4D",X"46",X"3E",X"36",X"2E",X"00",X"F5",X"AF",X"F1",X"08",X"AE",X"AC",X"AA",X"A7",X"A3",X"9E",
		X"9A",X"93",X"00",X"FF",X"8D",X"7B",X"C1",X"5D",X"46",X"C2",X"5F",X"47",X"45",X"8C",X"7B",X"C1",
		X"5D",X"46",X"C3",X"5F",X"47",X"45",X"00",X"8B",X"7B",X"C1",X"5D",X"46",X"C4",X"5F",X"47",X"45",
		X"00",X"00",X"8A",X"7B",X"E3",X"43",X"44",X"45",X"83",X"00",X"88",X"7B",X"E3",X"40",X"41",X"42",
		X"85",X"00",X"86",X"7A",X"E3",X"37",X"38",X"39",X"86",X"00",X"FC",X"E1",X"52",X"8E",X"00",X"E2",
		X"52",X"77",X"8E",X"00",X"E1",X"53",X"9A",X"00",X"E1",X"49",X"86",X"00",X"82",X"78",X"84",X"00",
		X"E4",X"4E",X"4C",X"4B",X"4A",X"86",X"00",X"FC",X"82",X"78",X"84",X"00",X"C2",X"4F",X"4F",X"4D",
		X"87",X"00",X"FF",X"FA",X"00",X"F0",X"00",X"08",X"08",X"08",X"08",X"09",X"0B",X"0D",X"10",X"14",
		X"19",X"1D",X"24",X"2A",X"2D",X"2D",X"2B",X"00",X"F1",X"00",X"27",X"27",X"27",X"28",X"2A",X"2D",
		X"31",X"36",X"3B",X"41",X"4C",X"A8",X"A4",X"A0",X"9B",X"94",X"00",X"F2",X"00",X"60",X"60",X"60",
		X"60",X"60",X"60",X"5F",X"5D",X"5A",X"56",X"52",X"00",X"F3",X"00",X"AF",X"AF",X"AF",X"AF",X"AF",
		X"AF",X"AF",X"AF",X"AE",X"AD",X"AB",X"00",X"FE",X"D6",X"19",X"FB",X"08",X"FE",X"91",X"19",X"F9",
		X"08",X"10",X"4D",X"00",X"F0",X"00",X"60",X"60",X"60",X"60",X"60",X"60",X"5F",X"5D",X"5A",X"56",
		X"52",X"24",X"2A",X"2D",X"2D",X"2B",X"00",X"F1",X"00",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",
		X"AF",X"AE",X"AD",X"AB",X"A8",X"A4",X"A0",X"9B",X"94",X"00",X"F2",X"00",X"08",X"08",X"08",X"08",
		X"09",X"0B",X"0D",X"10",X"14",X"19",X"1D",X"00",X"F3",X"00",X"27",X"27",X"27",X"28",X"2A",X"2D",
		X"31",X"36",X"3B",X"41",X"4C",X"00",X"03",X"4D",X"78",X"E2",X"32",X"34",X"8B",X"00",X"83",X"7B",
		X"C2",X"4F",X"76",X"35",X"C3",X"4D",X"37",X"38",X"39",X"88",X"00",X"87",X"7B",X"E3",X"40",X"41",
		X"42",X"86",X"00",X"89",X"7B",X"E3",X"43",X"44",X"45",X"84",X"00",X"8A",X"7B",X"C1",X"4F",X"46",
		X"C2",X"4D",X"47",X"3C",X"82",X"00",X"FD",X"81",X"3C",X"03",X"4F",X"7A",X"E3",X"37",X"38",X"39",
		X"85",X"00",X"E1",X"46",X"C2",X"4D",X"3D",X"3E",X"FD",X"E2",X"3E",X"3D",X"05",X"4F",X"7B",X"E3",
		X"40",X"41",X"42",X"88",X"00",X"87",X"7B",X"E3",X"43",X"44",X"45",X"86",X"00",X"88",X"7B",X"C1",
		X"4D",X"46",X"C2",X"4F",X"47",X"45",X"85",X"00",X"89",X"7B",X"C1",X"4D",X"46",X"C1",X"4F",X"3A",
		X"85",X"00",X"88",X"7B",X"FC",X"E3",X"40",X"41",X"42",X"85",X"00",X"86",X"7A",X"E3",X"37",X"38",
		X"39",X"06",X"4F",X"00",X"E1",X"52",X"8E",X"00",X"E2",X"52",X"77",X"8E",X"00",X"E1",X"53",X"9A",
		X"00",X"E1",X"49",X"86",X"00",X"82",X"78",X"84",X"00",X"E4",X"4E",X"4C",X"4B",X"4A",X"86",X"00",
		X"FC",X"82",X"78",X"84",X"00",X"FC",X"E2",X"4F",X"4D",X"87",X"00",X"01",X"5F",X"46",X"8E",X"00",
		X"01",X"5F",X"46",X"01",X"5D",X"47",X"8D",X"7B",X"E3",X"43",X"44",X"45",X"8B",X"7B",X"E3",X"40",
		X"41",X"42",X"82",X"00",X"87",X"7B",X"C2",X"5F",X"76",X"35",X"C3",X"5D",X"37",X"38",X"39",X"84",
		X"00",X"87",X"78",X"E2",X"32",X"34",X"97",X"00",X"10",X"4B",X"79",X"A0",X"00",X"A0",X"00",X"82",
		X"78",X"84",X"00",X"84",X"78",X"84",X"00",X"82",X"78",X"FC",X"82",X"78",X"84",X"00",X"84",X"78",
		X"84",X"00",X"82",X"78",X"FC",X"FF",X"A0",X"7B",X"10",X"5F",X"7A",X"A0",X"00",X"FF",X"F9",X"F7",
		X"FE",X"D5",X"1A",X"FB",X"F7",X"F0",X"0E",X"09",X"09",X"00",X"09",X"4D",X"00",X"E1",X"AD",X"C3",
		X"7F",X"B5",X"AA",X"A9",X"C3",X"4B",X"B3",X"B0",X"B0",X"FE",X"6A",X"1B",X"C2",X"7B",X"00",X"2A",
		X"89",X"00",X"C5",X"7D",X"AC",X"AB",X"AA",X"A9",X"78",X"C2",X"7B",X"08",X"29",X"87",X"00",X"FE",
		X"33",X"1B",X"FA",X"00",X"F0",X"0E",X"08",X"08",X"00",X"0D",X"4D",X"00",X"E3",X"B4",X"78",X"78",
		X"89",X"00",X"E1",X"AD",X"C3",X"7F",X"B5",X"AA",X"A9",X"C3",X"4D",X"B3",X"AC",X"7B",X"FE",X"6A",
		X"1B",X"E3",X"29",X"08",X"75",X"88",X"00",X"C5",X"7D",X"AC",X"AB",X"AA",X"A9",X"78",X"01",X"4B",
		X"0B",X"88",X"00",X"C4",X"7D",X"AC",X"AF",X"AE",X"AD",X"83",X"00",X"87",X"7B",X"E4",X"AC",X"AF",
		X"AE",X"AD",X"85",X"00",X"85",X"7B",X"E4",X"AC",X"AF",X"AE",X"AD",X"87",X"00",X"83",X"7B",X"E4",
		X"AC",X"AF",X"AE",X"AD",X"89",X"00",X"E1",X"7B",X"E4",X"AC",X"AF",X"AE",X"AD",X"8B",X"00",X"E3",
		X"AF",X"AE",X"AD",X"8D",X"00",X"E1",X"AD",X"7F",X"4D",X"00",X"F0",X"00",X"37",X"33",X"2F",X"2B",
		X"27",X"23",X"1F",X"1B",X"17",X"13",X"0F",X"0D",X"0B",X"09",X"00",X"F1",X"00",X"8D",X"89",X"85",
		X"81",X"7D",X"79",X"75",X"71",X"6D",X"69",X"65",X"61",X"5E",X"5B",X"59",X"58",X"00",X"07",X"4D",
		X"00",X"E4",X"AD",X"AE",X"AF",X"AC",X"85",X"7B",X"85",X"00",X"E4",X"AD",X"AE",X"AF",X"AC",X"87",
		X"7B",X"83",X"00",X"E4",X"AD",X"AE",X"AF",X"AC",X"89",X"7B",X"E5",X"00",X"AD",X"AE",X"AF",X"AC",
		X"89",X"7B",X"02",X"4F",X"78",X"C3",X"4D",X"AE",X"AF",X"AC",X"8B",X"7B",X"02",X"5F",X"78",X"01",
		X"4D",X"AC",X"07",X"4F",X"00",X"C3",X"4B",X"29",X"08",X"75",X"8B",X"00",X"E3",X"29",X"08",X"0B",
		X"8D",X"00",X"81",X"2A",X"99",X"00",X"FF",X"FA",X"00",X"FE",X"C7",X"1C",X"C7",X"4F",X"9C",X"9F",
		X"97",X"80",X"E9",X"A1",X"A1",X"09",X"0F",X"BC",X"C7",X"4F",X"9D",X"96",X"C6",X"D0",X"A8",X"A0",
		X"00",X"09",X"0F",X"BC",X"C1",X"4F",X"9E",X"86",X"00",X"09",X"0F",X"BC",X"FE",X"1B",X"1C",X"FE",
		X"1B",X"1C",X"FE",X"1B",X"1C",X"FE",X"1B",X"1C",X"82",X"00",X"C5",X"7F",X"F5",X"F1",X"EE",X"EB",
		X"A1",X"09",X"0F",X"BC",X"C2",X"7F",X"FB",X"F8",X"FE",X"45",X"1D",X"87",X"00",X"09",X"0F",X"BC",
		X"87",X"00",X"89",X"BC",X"FF",X"FA",X"00",X"F0",X"00",X"58",X"58",X"58",X"58",X"58",X"58",X"57",
		X"55",X"53",X"51",X"4D",X"4A",X"47",X"44",X"40",X"3D",X"00",X"F1",X"00",X"A7",X"A7",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A6",X"A4",X"A2",X"A1",X"9E",X"9B",X"98",X"95",X"92",X"00",X"6D",X"4F",X"7B",
		X"E3",X"FE",X"99",X"9B",X"09",X"4F",X"7B",X"E7",X"F2",X"F6",X"F9",X"FC",X"FF",X"9A",X"F8",X"07",
		X"4F",X"7B",X"E8",X"EC",X"EF",X"F3",X"F7",X"FA",X"FD",X"98",X"F5",X"81",X"00",X"EC",X"D1",X"D2",
		X"D3",X"D2",X"D3",X"D2",X"EA",X"ED",X"F0",X"F4",X"F8",X"FB",X"84",X"00",X"86",X"A1",X"E4",X"EB",
		X"EE",X"F1",X"F5",X"5E",X"7F",X"00",X"A5",X"00",X"E3",X"F5",X"98",X"FD",X"8B",X"00",X"E3",X"9E",
		X"F8",X"9A",X"C2",X"0F",X"F3",X"F5",X"07",X"7F",X"00",X"E4",X"A8",X"D0",X"C6",X"96",X"C5",X"0F",
		X"F3",X"F5",X"F6",X"F7",X"F4",X"07",X"5F",X"A1",X"C6",X"0F",X"F2",X"F3",X"F5",X"F6",X"F7",X"F4",
		X"03",X"5F",X"7B",X"E7",X"D1",X"D2",X"D3",X"D2",X"D3",X"D2",X"D3",X"C3",X"0F",X"F1",X"F7",X"F4",
		X"16",X"4F",X"7B",X"F4",X"30",X"F5",X"7F",X"04",X"4E",X"7B",X"C5",X"0E",X"E8",X"E2",X"DC",X"D6",
		X"BF",X"87",X"BC",X"05",X"4E",X"7B",X"C4",X"0E",X"E3",X"DD",X"D7",X"C4",X"87",X"BC",X"04",X"4E",
		X"7B",X"C5",X"0E",X"E9",X"E4",X"DE",X"D8",X"C8",X"87",X"BC",X"04",X"4E",X"7B",X"C5",X"0E",X"EA",
		X"E5",X"DF",X"D9",X"D0",X"87",X"BC",X"03",X"4E",X"7B",X"81",X"8C",X"C4",X"0E",X"D2",X"E6",X"E0",
		X"DA",X"88",X"BC",X"FF",X"C5",X"4F",X"9C",X"9F",X"97",X"80",X"E9",X"8B",X"A1",X"E6",X"9D",X"96",
		X"C6",X"D0",X"A8",X"A0",X"8A",X"00",X"E1",X"9E",X"FF",X"C4",X"7F",X"F5",X"F1",X"EE",X"EB",X"8A",
		X"A1",X"FF",X"C4",X"0F",X"FA",X"FD",X"FE",X"FF",X"C4",X"1E",X"D2",X"E6",X"E0",X"DA",X"86",X"BC",
		X"FF",X"FA",X"00",X"FE",X"C3",X"1C",X"FE",X"04",X"1D",X"51",X"7F",X"00",X"40",X"7F",X"00",X"FE",
		X"19",X"1D",X"E2",X"FB",X"F8",X"FE",X"22",X"1D",X"01",X"7F",X"FA",X"C3",X"0E",X"F8",X"FB",X"FC",
		X"FE",X"92",X"1D",X"E3",X"F6",X"F7",X"F9",X"03",X"4E",X"7B",X"C5",X"1E",X"E9",X"E4",X"DE",X"D8",
		X"C8",X"85",X"BC",X"07",X"4E",X"7B",X"C4",X"1E",X"EA",X"DD",X"D7",X"C4",X"85",X"BC",X"06",X"4E",
		X"7B",X"C5",X"1E",X"E8",X"E2",X"DC",X"D6",X"BF",X"85",X"BC",X"06",X"4E",X"7B",X"C5",X"1E",X"E7",
		X"E1",X"DB",X"D5",X"BE",X"85",X"BC",X"06",X"4E",X"7B",X"C5",X"1E",X"E9",X"E4",X"DE",X"D8",X"C8",
		X"85",X"BC",X"02",X"4E",X"7B",X"C5",X"1E",X"EA",X"E5",X"DF",X"D9",X"D0",X"05",X"0E",X"BC",X"FF",
		X"FA",X"00",X"FE",X"C3",X"1C",X"FE",X"04",X"1D",X"2F",X"4F",X"00",X"81",X"E3",X"8F",X"00",X"81",
		X"E5",X"8F",X"00",X"81",X"E7",X"8F",X"00",X"81",X"CF",X"8F",X"00",X"E2",X"C7",X"E3",X"8E",X"00",
		X"E2",X"C8",X"E5",X"8E",X"00",X"E2",X"C9",X"CA",X"FE",X"19",X"1D",X"C2",X"4F",X"DF",X"CB",X"FE",
		X"22",X"1D",X"C2",X"4F",X"E1",X"CC",X"C2",X"0E",X"FB",X"FC",X"FE",X"92",X"1D",X"C2",X"4F",X"D6",
		X"CD",X"01",X"0E",X"F9",X"FE",X"57",X"1D",X"FA",X"00",X"6D",X"4F",X"7B",X"E3",X"D6",X"D9",X"DA",
		X"89",X"7B",X"85",X"D6",X"E2",X"DB",X"DC",X"87",X"7B",X"87",X"D6",X"E2",X"DD",X"DE",X"E5",X"D1",
		X"D2",X"D3",X"D2",X"D4",X"89",X"D6",X"E2",X"DF",X"E0",X"84",X"A1",X"E1",X"D5",X"89",X"D6",X"E2",
		X"E1",X"E2",X"84",X"00",X"E1",X"D7",X"8A",X"D6",X"E1",X"E4",X"84",X"00",X"E1",X"D8",X"8A",X"D6",
		X"E1",X"E6",X"84",X"00",X"E1",X"D8",X"8A",X"D6",X"E1",X"E8",X"84",X"00",X"E1",X"D8",X"8A",X"D6",
		X"E1",X"E1",X"FE",X"54",X"1E",X"FE",X"54",X"1E",X"FE",X"5A",X"1E",X"84",X"00",X"FC",X"E1",X"D7",
		X"8B",X"D6",X"84",X"A1",X"E1",X"D5",X"88",X"D6",X"83",X"7B",X"E5",X"D1",X"D2",X"D3",X"D2",X"D4",
		X"85",X"D6",X"96",X"7B",X"84",X"00",X"E1",X"D8",X"8B",X"D6",X"84",X"00",X"E1",X"D8",X"8B",X"D6",
		X"FF",X"F4",X"30",X"F5",X"7F",X"50",X"07",X"BC",X"10",X"4F",X"A1",X"60",X"4F",X"00",X"40",X"0F",
		X"00",X"10",X"5F",X"A1",X"70",X"07",X"BC",X"F0",X"04",X"08",X"0C",X"00",X"F0",X"0B",X"10",X"14",
		X"08",X"00",X"F1",X"02",X"B0",X"AC",X"AC",X"B0",X"00",X"F1",X"0B",X"A8",X"A4",X"B0",X"00",X"FE",
		X"92",X"1E",X"60",X"07",X"BC",X"60",X"07",X"BC",X"F0",X"01",X"08",X"0C",X"00",X"F0",X"0A",X"10",
		X"14",X"08",X"00",X"F1",X"03",X"A8",X"A4",X"B0",X"00",X"F1",X"0A",X"B8",X"B4",X"00",X"FE",X"8F",
		X"1E",X"F0",X"03",X"10",X"14",X"14",X"10",X"00",X"F0",X"0B",X"08",X"0C",X"0C",X"08",X"00",X"F1",
		X"02",X"B0",X"AC",X"AC",X"B0",X"00",X"F1",X"0B",X"B8",X"B4",X"B4",X"B8",X"00",X"FE",X"8F",X"1E",
		X"F0",X"00",X"18",X"1C",X"1C",X"18",X"00",X"F0",X"0B",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"04",
		X"B8",X"B4",X"B4",X"B8",X"B0",X"AC",X"AC",X"B0",X"00",X"FE",X"8F",X"1E",X"F0",X"01",X"08",X"0C",
		X"00",X"F0",X"06",X"20",X"24",X"18",X"00",X"F0",X"0C",X"18",X"1C",X"10",X"00",X"F1",X"02",X"B8",
		X"B4",X"00",X"F1",X"07",X"B0",X"AC",X"B8",X"00",X"F1",X"0C",X"B0",X"AC",X"B8",X"00",X"FE",X"8F",
		X"1E",X"F0",X"01",X"08",X"0C",X"00",X"F0",X"07",X"10",X"14",X"14",X"10",X"08",X"0C",X"00",X"F1",
		X"00",X"B8",X"B4",X"B4",X"B8",X"BF",X"BF",X"B0",X"AC",X"B8",X"BF",X"BF",X"B8",X"B4",X"00",X"FE",
		X"8F",X"1E",X"F0",X"00",X"18",X"1C",X"1C",X"18",X"01",X"18",X"1C",X"1C",X"18",X"01",X"01",X"10",
		X"14",X"14",X"10",X"00",X"F1",X"02",X"B0",X"AC",X"AC",X"B0",X"BF",X"B8",X"B4",X"B4",X"B8",X"BF",
		X"BF",X"BC",X"BC",X"00",X"FE",X"8F",X"1E",X"F0",X"08",X"0C",X"0C",X"08",X"01",X"04",X"04",X"01",
		X"01",X"04",X"04",X"00",X"F1",X"00",X"B8",X"B4",X"B4",X"B8",X"A0",X"9C",X"9C",X"A0",X"B0",X"AC",
		X"AC",X"B0",X"00",X"FE",X"8F",X"1E",X"F0",X"00",X"08",X"0C",X"01",X"01",X"10",X"14",X"08",X"01",
		X"01",X"04",X"01",X"01",X"18",X"1C",X"10",X"00",X"F1",X"00",X"B8",X"B4",X"BF",X"BF",X"BF",X"BC",
		X"BF",X"BF",X"B8",X"B4",X"BF",X"BF",X"B8",X"B4",X"00",X"FE",X"8F",X"1E",X"F0",X"00",X"10",X"14",
		X"08",X"01",X"08",X"0C",X"01",X"01",X"20",X"24",X"18",X"01",X"18",X"1C",X"10",X"00",X"F1",X"00",
		X"A8",X"A4",X"B0",X"BF",X"A0",X"9C",X"A8",X"BF",X"A8",X"A4",X"B0",X"BF",X"A8",X"A4",X"B0",X"00",
		X"FE",X"8F",X"1E",X"F0",X"00",X"18",X"1C",X"1C",X"18",X"20",X"24",X"24",X"20",X"18",X"1C",X"1C",
		X"18",X"18",X"1C",X"1C",X"18",X"00",X"F1",X"00",X"A8",X"A4",X"A4",X"A8",X"B0",X"AC",X"AC",X"B0",
		X"A0",X"9C",X"9C",X"A0",X"B0",X"AC",X"AC",X"B0",X"00",X"F0",X"01",X"04",X"04",X"01",X"18",X"1C",
		X"1C",X"18",X"01",X"04",X"04",X"01",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"01",X"BC",X"BC",X"BF",
		X"BF",X"BC",X"BC",X"BF",X"A0",X"9C",X"9C",X"A0",X"B0",X"AC",X"AC",X"B0",X"00",X"FE",X"8F",X"1E",
		X"F0",X"01",X"08",X"0C",X"00",X"F0",X"07",X"10",X"14",X"08",X"00",X"F1",X"02",X"BC",X"BF",X"BF",
		X"B8",X"BC",X"00",X"F1",X"0B",X"A8",X"A4",X"B0",X"00",X"FE",X"8F",X"1E",X"F0",X"01",X"08",X"0C",
		X"0C",X"08",X"01",X"10",X"14",X"08",X"01",X"01",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"04",X"B8",
		X"B4",X"00",X"F1",X"0A",X"B8",X"B4",X"B4",X"B8",X"00",X"FE",X"8F",X"1E",X"F0",X"02",X"08",X"0C",
		X"0C",X"08",X"01",X"01",X"18",X"1C",X"1C",X"18",X"00",X"F1",X"06",X"B8",X"B4",X"B4",X"B8",X"00",
		X"FE",X"8F",X"1E",X"F0",X"02",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"02",X"B8",X"B4",X"B4",X"B8",
		X"00",X"F1",X"0A",X"B8",X"B4",X"B4",X"B8",X"00",X"FE",X"8F",X"1E",X"F0",X"02",X"08",X"0C",X"00",
		X"F0",X"09",X"08",X"0C",X"00",X"F1",X"02",X"B0",X"AC",X"B8",X"00",X"F1",X"08",X"B0",X"AC",X"B8",
		X"BF",X"B8",X"B4",X"00",X"FE",X"8F",X"1E",X"F0",X"00",X"08",X"0C",X"00",X"F0",X"06",X"10",X"14",
		X"14",X"10",X"01",X"08",X"0C",X"00",X"F1",X"01",X"BC",X"BC",X"BF",X"A8",X"A4",X"B0",X"BF",X"BF",
		X"BF",X"B8",X"B4",X"00",X"FE",X"8F",X"1E",X"F0",X"02",X"10",X"14",X"14",X"10",X"01",X"01",X"20",
		X"24",X"24",X"20",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"01",X"A8",X"A4",X"A4",X"A8",X"00",X"F1",
		X"0B",X"B0",X"AC",X"AC",X"B0",X"00",X"FE",X"8F",X"1E",X"F0",X"04",X"20",X"24",X"24",X"20",X"01",
		X"01",X"08",X"0C",X"0C",X"08",X"00",X"F1",X"00",X"B8",X"B4",X"B4",X"B8",X"BF",X"98",X"94",X"94",
		X"98",X"BF",X"A8",X"A4",X"A4",X"A8",X"00",X"FE",X"8F",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"21",X"00",X"E3",X"3E",X"1D",X"32",X"0C",X"E0",X"DD",X"7E",X"00",X"E6",X"7F",X"D6",X"02",
		X"FA",X"17",X"21",X"21",X"26",X"21",X"EF",X"11",X"10",X"00",X"DD",X"19",X"21",X"0C",X"E0",X"35",
		X"20",X"E7",X"CD",X"0B",X"2B",X"C9",X"18",X"25",X"37",X"25",X"97",X"25",X"F1",X"25",X"00",X"00",
		X"00",X"00",X"27",X"26",X"3B",X"26",X"F7",X"24",X"0D",X"25",X"00",X"00",X"00",X"00",X"4A",X"26",
		X"63",X"26",X"94",X"26",X"C0",X"26",X"14",X"27",X"66",X"27",X"8E",X"27",X"A1",X"27",X"F7",X"24",
		X"33",X"28",X"24",X"29",X"24",X"29",X"06",X"29",X"6C",X"2A",X"20",X"2F",X"09",X"30",X"46",X"30",
		X"84",X"30",X"70",X"31",X"00",X"00",X"44",X"32",X"BD",X"32",X"CE",X"32",X"76",X"33",X"D4",X"33",
		X"0D",X"34",X"0D",X"35",X"CD",X"15",X"22",X"CD",X"BF",X"21",X"18",X"1E",X"F5",X"CD",X"15",X"22",
		X"CD",X"BF",X"21",X"18",X"07",X"F5",X"CD",X"EE",X"21",X"CD",X"B0",X"21",X"F1",X"A7",X"28",X"0A",
		X"11",X"64",X"00",X"1F",X"38",X"03",X"11",X"9C",X"FF",X"19",X"DD",X"5E",X"04",X"DD",X"56",X"05",
		X"19",X"7C",X"FE",X"0C",X"38",X"03",X"FE",X"F5",X"D8",X"DD",X"75",X"04",X"DD",X"74",X"05",X"C9",
		X"3A",X"04",X"E7",X"47",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"29",X"29",X"7C",X"18",X"0A",X"3A",
		X"04",X"E7",X"47",X"2A",X"08",X"E3",X"29",X"29",X"7C",X"C6",X"28",X"10",X"02",X"D6",X"08",X"6F",
		X"26",X"00",X"29",X"29",X"EB",X"DD",X"7E",X"05",X"87",X"87",X"38",X"0C",X"C6",X"38",X"CD",X"98",
		X"22",X"EB",X"21",X"00",X"00",X"ED",X"52",X"C9",X"2F",X"C6",X"35",X"C3",X"98",X"22",X"F5",X"DD",
		X"6E",X"04",X"DD",X"66",X"05",X"29",X"29",X"DD",X"56",X"09",X"14",X"DD",X"5E",X"08",X"CB",X"3A",
		X"CB",X"1B",X"CB",X"3A",X"CB",X"1B",X"D5",X"7C",X"87",X"18",X"27",X"11",X"55",X"01",X"29",X"29",
		X"6C",X"9F",X"67",X"18",X"2C",X"F5",X"2A",X"04",X"E3",X"29",X"ED",X"5B",X"08",X"E3",X"7A",X"FE",
		X"02",X"38",X"07",X"20",X"E6",X"7B",X"FE",X"AA",X"30",X"E1",X"CB",X"3A",X"CB",X"1B",X"D5",X"7C",
		X"29",X"84",X"CB",X"7C",X"28",X"5D",X"2F",X"CD",X"98",X"22",X"11",X"00",X"00",X"EB",X"ED",X"52",
		X"D1",X"F1",X"A7",X"28",X"07",X"ED",X"52",X"1F",X"30",X"02",X"19",X"19",X"DD",X"5E",X"02",X"DD",
		X"56",X"03",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"DD",
		X"7E",X"05",X"A7",X"FA",X"67",X"22",X"2F",X"3C",X"28",X"0D",X"87",X"87",X"FE",X"E0",X"30",X"03",
		X"87",X"C6",X"20",X"EB",X"CD",X"98",X"22",X"DD",X"7E",X"00",X"FE",X"17",X"30",X"03",X"22",X"86",
		X"E2",X"DD",X"5E",X"0A",X"DD",X"56",X"0B",X"19",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"D0",X"DD",
		X"34",X"0C",X"C9",X"CD",X"98",X"22",X"18",X"A8",X"4F",X"06",X"00",X"C5",X"60",X"68",X"CB",X"3B",
		X"30",X"01",X"09",X"28",X"06",X"CB",X"21",X"CB",X"10",X"18",X"F3",X"C1",X"6C",X"60",X"CB",X"3A",
		X"30",X"01",X"09",X"C8",X"CB",X"21",X"CB",X"10",X"18",X"F4",X"3A",X"04",X"D0",X"E6",X"40",X"C8",
		X"DD",X"7E",X"07",X"A7",X"C0",X"3A",X"0D",X"E3",X"FE",X"0F",X"D0",X"87",X"5F",X"16",X"00",X"21",
		X"6B",X"23",X"19",X"06",X"00",X"FD",X"21",X"90",X"46",X"FD",X"09",X"3A",X"D8",X"E2",X"A7",X"28",
		X"0B",X"3D",X"28",X"0D",X"3A",X"D9",X"E2",X"FE",X"10",X"D0",X"18",X"05",X"CD",X"51",X"23",X"38",
		X"07",X"23",X"3E",X"24",X"CD",X"53",X"23",X"D0",X"F5",X"79",X"FE",X"2C",X"28",X"3E",X"FE",X"40",
		X"28",X"3A",X"F1",X"87",X"FD",X"BE",X"01",X"3E",X"10",X"30",X"03",X"04",X"3E",X"18",X"32",X"0D",
		X"E3",X"3E",X"01",X"32",X"0F",X"E3",X"3E",X"04",X"32",X"00",X"E3",X"AF",X"32",X"D8",X"E2",X"3E",
		X"1F",X"CD",X"B6",X"5E",X"3E",X"17",X"CD",X"B6",X"5E",X"3A",X"0C",X"E3",X"D6",X"02",X"30",X"01",
		X"AF",X"21",X"25",X"E7",X"BE",X"30",X"01",X"7E",X"23",X"77",X"37",X"C9",X"21",X"00",X"E3",X"3E",
		X"0B",X"BE",X"28",X"06",X"77",X"3E",X"17",X"CD",X"B6",X"5E",X"F1",X"3E",X"04",X"32",X"0F",X"E3",
		X"C9",X"3E",X"30",X"DD",X"96",X"06",X"FD",X"86",X"02",X"FD",X"BE",X"03",X"D0",X"3A",X"03",X"E3",
		X"86",X"DD",X"96",X"03",X"FD",X"86",X"00",X"FD",X"BE",X"01",X"C9",X"FA",X"02",X"FC",X"00",X"00",
		X"00",X"04",X"00",X"06",X"FE",X"FE",X"FE",X"FF",X"FF",X"00",X"00",X"01",X"01",X"02",X"02",X"FE",
		X"FE",X"FF",X"FF",X"00",X"00",X"01",X"01",X"02",X"02",X"19",X"EB",X"DD",X"7E",X"06",X"C6",X"18",
		X"6F",X"CB",X"3F",X"CB",X"3F",X"85",X"2F",X"CD",X"98",X"22",X"EB",X"DD",X"6E",X"05",X"DD",X"66",
		X"06",X"C9",X"DD",X"CB",X"0E",X"7E",X"28",X"07",X"EB",X"21",X"FF",X"FF",X"A7",X"ED",X"52",X"DD",
		X"5E",X"02",X"DD",X"56",X"03",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"DD",X"7E",X"06",X"11",
		X"00",X"00",X"D6",X"30",X"F8",X"1C",X"D6",X"20",X"D8",X"1C",X"D6",X"18",X"D8",X"CB",X"3F",X"CB",
		X"3F",X"C6",X"03",X"5F",X"C9",X"CD",X"9D",X"24",X"DD",X"7E",X"03",X"FD",X"BE",X"01",X"38",X"2E",
		X"47",X"FD",X"7E",X"03",X"B8",X"38",X"58",X"FD",X"96",X"02",X"FE",X"04",X"18",X"31",X"CD",X"A7",
		X"24",X"DD",X"7E",X"03",X"C6",X"0E",X"4F",X"D6",X"1C",X"30",X"01",X"AF",X"47",X"FD",X"7E",X"01",
		X"FD",X"96",X"00",X"FE",X"24",X"38",X"2B",X"FD",X"7E",X"01",X"B9",X"38",X"07",X"78",X"FD",X"BE",
		X"00",X"3E",X"00",X"C9",X"FD",X"7E",X"03",X"B9",X"38",X"25",X"FD",X"96",X"02",X"FE",X"24",X"38",
		X"1E",X"FD",X"7E",X"02",X"B8",X"3F",X"D0",X"FD",X"86",X"01",X"1F",X"DD",X"BE",X"03",X"9F",X"3C",
		X"37",X"C9",X"FD",X"7E",X"03",X"B9",X"38",X"07",X"78",X"FD",X"BE",X"02",X"3E",X"00",X"C9",X"3E",
		X"01",X"C9",X"DD",X"21",X"00",X"E3",X"3A",X"04",X"E7",X"1F",X"38",X"0E",X"CD",X"9D",X"24",X"FD",
		X"7E",X"01",X"FD",X"86",X"00",X"1F",X"DD",X"77",X"03",X"C9",X"CD",X"D0",X"2E",X"82",X"18",X"F5",
		X"3A",X"04",X"E7",X"1F",X"38",X"23",X"CD",X"9D",X"24",X"CD",X"71",X"24",X"D0",X"FD",X"23",X"FD",
		X"23",X"FD",X"7E",X"01",X"FD",X"96",X"00",X"FE",X"4A",X"D8",X"DE",X"2A",X"4F",X"ED",X"5F",X"87",
		X"B9",X"3F",X"D8",X"FD",X"86",X"00",X"C6",X"15",X"C9",X"CD",X"D0",X"2E",X"5F",X"7A",X"93",X"D8",
		X"FE",X"88",X"30",X"D2",X"57",X"ED",X"5F",X"87",X"BA",X"3F",X"D8",X"83",X"C9",X"DD",X"7E",X"0C",
		X"1F",X"DD",X"7E",X"0B",X"1F",X"18",X"14",X"E5",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"29",X"DD",
		X"7E",X"0C",X"1F",X"DD",X"7E",X"0B",X"1F",X"84",X"C6",X"28",X"E1",X"E6",X"FC",X"4F",X"06",X"00",
		X"FD",X"21",X"00",X"E5",X"FD",X"09",X"C9",X"EB",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"19",X"DD",
		X"75",X"0A",X"DD",X"74",X"0B",X"30",X"03",X"DD",X"34",X"0C",X"CB",X"12",X"30",X"03",X"DD",X"35",
		X"0C",X"6C",X"DD",X"66",X"0C",X"ED",X"5B",X"0B",X"E3",X"A7",X"ED",X"52",X"11",X"30",X"00",X"19",
		X"DD",X"74",X"07",X"DD",X"75",X"06",X"C9",X"2A",X"08",X"E3",X"11",X"F6",X"FF",X"19",X"30",X"03",
		X"22",X"08",X"E3",X"DD",X"7E",X"00",X"FE",X"0A",X"28",X"49",X"C3",X"66",X"26",X"DD",X"35",X"0F",
		X"28",X"3A",X"CD",X"B6",X"27",X"AF",X"18",X"3E",X"3A",X"1E",X"E7",X"A7",X"28",X"3B",X"3E",X"01",
		X"CD",X"B9",X"27",X"2A",X"08",X"E3",X"25",X"20",X"2A",X"7D",X"FE",X"A0",X"38",X"25",X"DD",X"34",
		X"00",X"AF",X"32",X"1A",X"E2",X"18",X"1C",X"2A",X"D8",X"E2",X"7D",X"A7",X"28",X"12",X"25",X"20",
		X"02",X"2E",X"00",X"22",X"D8",X"E2",X"3D",X"28",X"C9",X"AF",X"18",X"0A",X"DD",X"36",X"00",X"03",
		X"CD",X"B6",X"27",X"3A",X"1F",X"E0",X"CD",X"7C",X"21",X"3A",X"D8",X"E2",X"0E",X"02",X"A7",X"20",
		X"1D",X"CD",X"1D",X"28",X"3A",X"04",X"E7",X"1F",X"38",X"14",X"2A",X"08",X"E3",X"29",X"7C",X"FE",
		X"05",X"38",X"0B",X"06",X"0A",X"FE",X"07",X"30",X"02",X"06",X"05",X"78",X"81",X"4F",X"DD",X"71",
		X"0D",X"3A",X"04",X"D0",X"CB",X"77",X"CA",X"C0",X"40",X"CD",X"D5",X"23",X"D2",X"C0",X"40",X"87",
		X"87",X"87",X"C6",X"10",X"C3",X"0E",X"23",X"DD",X"7E",X"00",X"FE",X"04",X"28",X"07",X"DD",X"35",
		X"0F",X"C0",X"C3",X"86",X"57",X"2A",X"86",X"E2",X"11",X"F0",X"FF",X"19",X"38",X"03",X"21",X"00",
		X"00",X"22",X"86",X"E2",X"ED",X"5B",X"0A",X"E3",X"19",X"30",X"03",X"DD",X"34",X"0C",X"22",X"0A",
		X"E3",X"DD",X"35",X"0F",X"C0",X"DD",X"7E",X"0D",X"3C",X"47",X"E6",X"07",X"20",X"0B",X"78",X"D6",
		X"08",X"47",X"2A",X"86",X"E2",X"7C",X"B5",X"28",X"0F",X"DD",X"70",X"0D",X"2A",X"86",X"E2",X"3E",
		X"09",X"94",X"DD",X"77",X"0F",X"C3",X"C0",X"40",X"DD",X"36",X"0F",X"20",X"DD",X"36",X"00",X"84",
		X"C9",X"2A",X"08",X"E3",X"11",X"E8",X"FF",X"19",X"38",X"03",X"21",X"00",X"00",X"22",X"08",X"E3",
		X"DD",X"35",X"0F",X"20",X"12",X"DD",X"36",X"0F",X"50",X"DD",X"36",X"00",X"08",X"3E",X"0F",X"CD",
		X"B6",X"5E",X"3E",X"1F",X"CD",X"B6",X"5E",X"AF",X"2A",X"04",X"E3",X"CD",X"15",X"22",X"CD",X"1D",
		X"28",X"DD",X"71",X"0D",X"C3",X"C0",X"40",X"21",X"00",X"00",X"22",X"86",X"E2",X"DD",X"36",X"0D",
		X"26",X"CD",X"C0",X"40",X"DD",X"35",X"0F",X"C0",X"C3",X"86",X"57",X"CD",X"C0",X"40",X"DD",X"35",
		X"0F",X"C0",X"DD",X"35",X"00",X"DD",X"36",X"0F",X"50",X"C9",X"3E",X"01",X"CD",X"B9",X"27",X"2A",
		X"08",X"E3",X"7C",X"FE",X"01",X"38",X"0F",X"20",X"05",X"7D",X"FE",X"D0",X"38",X"08",X"DD",X"34",
		X"00",X"18",X"03",X"CD",X"B6",X"27",X"3A",X"1F",X"E0",X"CD",X"7C",X"21",X"CD",X"1D",X"28",X"79",
		X"C6",X"20",X"DD",X"77",X"0D",X"3A",X"04",X"D0",X"E6",X"40",X"CA",X"C0",X"40",X"3A",X"03",X"E3",
		X"D6",X"06",X"FE",X"B5",X"DA",X"C0",X"40",X"3E",X"2B",X"DD",X"CB",X"03",X"7E",X"28",X"02",X"3E",
		X"2F",X"C3",X"DC",X"2F",X"CD",X"74",X"21",X"DD",X"7E",X"05",X"C6",X"03",X"FE",X"07",X"D2",X"C0",
		X"40",X"DD",X"34",X"00",X"DD",X"7E",X"03",X"D6",X"60",X"30",X"01",X"2F",X"87",X"C6",X"10",X"DD",
		X"77",X"0E",X"21",X"00",X"00",X"22",X"C2",X"E2",X"3E",X"FF",X"32",X"71",X"E0",X"C3",X"C0",X"40",
		X"21",X"00",X"02",X"CD",X"81",X"22",X"2A",X"86",X"E2",X"11",X"08",X"00",X"A7",X"ED",X"52",X"38",
		X"03",X"22",X"86",X"E2",X"2A",X"C2",X"E2",X"19",X"7C",X"FE",X"02",X"30",X"03",X"22",X"C2",X"E2",
		X"CD",X"8A",X"23",X"19",X"DD",X"75",X"05",X"DD",X"74",X"06",X"DD",X"4E",X"0E",X"CD",X"99",X"22",
		X"DD",X"7E",X"03",X"C6",X"20",X"CB",X"7F",X"CD",X"A6",X"23",X"21",X"50",X"27",X"19",X"7E",X"DD",
		X"77",X"0D",X"CD",X"C0",X"40",X"DD",X"7E",X"06",X"FE",X"AA",X"38",X"15",X"DD",X"36",X"0F",X"14",
		X"DD",X"34",X"00",X"C9",X"DD",X"36",X"0D",X"4F",X"CD",X"C0",X"40",X"3A",X"2A",X"E7",X"A7",X"28",
		X"28",X"3A",X"2A",X"E7",X"A7",X"C8",X"3A",X"22",X"E0",X"E6",X"03",X"C0",X"21",X"71",X"E0",X"35",
		X"7E",X"FE",X"90",X"CA",X"BD",X"56",X"1E",X"C0",X"CB",X"47",X"20",X"02",X"1E",X"CF",X"FE",X"A6",
		X"30",X"02",X"3E",X"A6",X"C6",X"30",X"C3",X"80",X"40",X"DD",X"35",X"0F",X"CA",X"C8",X"65",X"C9",
		X"22",X"22",X"25",X"26",X"26",X"26",X"26",X"27",X"27",X"27",X"27",X"28",X"28",X"28",X"29",X"29",
		X"29",X"2A",X"2A",X"4F",X"4F",X"4F",X"2A",X"86",X"E2",X"11",X"10",X"00",X"A7",X"ED",X"52",X"38",
		X"28",X"22",X"86",X"E2",X"DD",X"35",X"0F",X"F0",X"DD",X"34",X"0D",X"DD",X"7E",X"0D",X"FE",X"2F",
		X"28",X"04",X"FE",X"33",X"20",X"05",X"D6",X"04",X"DD",X"77",X"0D",X"C3",X"DC",X"25",X"DD",X"7E",
		X"0D",X"FE",X"2E",X"28",X"04",X"FE",X"32",X"20",X"DB",X"DD",X"34",X"00",X"DD",X"36",X"0F",X"08",
		X"C9",X"DD",X"35",X"0F",X"C0",X"C3",X"86",X"57",X"3A",X"87",X"E2",X"2F",X"D6",X"03",X"5F",X"16",
		X"FF",X"CD",X"0D",X"28",X"18",X"1F",X"3A",X"20",X"E0",X"2A",X"08",X"E3",X"A7",X"28",X"E9",X"EE",
		X"05",X"28",X"4A",X"0F",X"30",X"27",X"3A",X"22",X"E0",X"E6",X"07",X"20",X"05",X"3E",X"16",X"CD",
		X"B6",X"5E",X"11",X"E8",X"FF",X"19",X"38",X"02",X"ED",X"52",X"7C",X"32",X"B2",X"E2",X"3D",X"20",
		X"08",X"7D",X"FE",X"A0",X"30",X"03",X"21",X"A0",X"01",X"22",X"08",X"E3",X"C9",X"EB",X"21",X"B2",
		X"E2",X"34",X"7E",X"07",X"07",X"07",X"E6",X"07",X"C6",X"05",X"6F",X"26",X"00",X"19",X"EB",X"2A",
		X"78",X"E0",X"ED",X"52",X"EB",X"30",X"03",X"2A",X"78",X"E0",X"22",X"08",X"E3",X"3A",X"D8",X"E2",
		X"3D",X"C0",X"3A",X"22",X"E0",X"E6",X"0F",X"C0",X"3E",X"17",X"C3",X"B6",X"5E",X"3A",X"05",X"E3",
		X"0E",X"04",X"FE",X"03",X"F0",X"0D",X"FE",X"02",X"F0",X"0D",X"C6",X"01",X"F0",X"0D",X"C6",X"01",
		X"F0",X"0D",X"C9",X"3A",X"0C",X"E0",X"21",X"22",X"E0",X"AE",X"1F",X"D8",X"3A",X"1E",X"E7",X"A7",
		X"28",X"09",X"DD",X"7E",X"04",X"DD",X"86",X"08",X"DD",X"77",X"08",X"5F",X"30",X"03",X"DD",X"34",
		X"09",X"DD",X"56",X"09",X"2A",X"CB",X"E2",X"ED",X"52",X"30",X"04",X"DD",X"36",X"08",X"00",X"DD",
		X"6E",X"0A",X"DD",X"66",X"0B",X"19",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"30",X"03",X"DD",X"34",
		X"0C",X"6C",X"DD",X"66",X"0C",X"ED",X"5B",X"0B",X"E3",X"A7",X"ED",X"52",X"11",X"30",X"00",X"19",
		X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"CB",X"00",X"FE",X"11",X"10",X"00",X"19",X"11",X"20",
		X"01",X"A7",X"ED",X"52",X"D0",X"DD",X"CB",X"00",X"BE",X"01",X"00",X"05",X"FD",X"21",X"50",X"E4",
		X"11",X"10",X"00",X"FD",X"7E",X"00",X"FE",X"17",X"20",X"01",X"0C",X"FD",X"19",X"10",X"F4",X"0D",
		X"28",X"08",X"0E",X"00",X"CD",X"BA",X"22",X"C3",X"C0",X"40",X"DD",X"36",X"0D",X"4E",X"CD",X"C0",
		X"40",X"DD",X"E5",X"E1",X"11",X"10",X"E3",X"01",X"10",X"00",X"ED",X"B0",X"21",X"19",X"04",X"22",
		X"10",X"E3",X"21",X"00",X"00",X"22",X"14",X"E3",X"21",X"50",X"E4",X"11",X"10",X"00",X"06",X"05",
		X"36",X"00",X"19",X"10",X"FB",X"DD",X"6E",X"0E",X"65",X"22",X"11",X"E7",X"2A",X"16",X"E3",X"24",
		X"11",X"30",X"01",X"A7",X"ED",X"52",X"21",X"0D",X"E7",X"7E",X"38",X"03",X"D6",X"01",X"27",X"2B",
		X"77",X"21",X"1D",X"E7",X"34",X"C9",X"DD",X"7E",X"0F",X"E6",X"0F",X"20",X"0F",X"ED",X"5F",X"87",
		X"6F",X"26",X"00",X"29",X"11",X"C0",X"01",X"19",X"29",X"22",X"4F",X"E0",X"DD",X"35",X"0F",X"20",
		X"03",X"DD",X"35",X"00",X"3A",X"22",X"E0",X"DD",X"AE",X"01",X"1F",X"D8",X"3A",X"88",X"E2",X"FE",
		X"03",X"CA",X"E8",X"29",X"CD",X"5D",X"2A",X"38",X"4C",X"DD",X"7E",X"07",X"1F",X"DD",X"7E",X"06",
		X"1F",X"C6",X"04",X"47",X"3A",X"D2",X"E2",X"A7",X"28",X"1A",X"78",X"FE",X"38",X"30",X"15",X"FE",
		X"28",X"30",X"0C",X"CD",X"33",X"2A",X"2A",X"C7",X"E2",X"11",X"00",X"FD",X"19",X"18",X"50",X"CD",
		X"33",X"2A",X"18",X"48",X"DD",X"7E",X"00",X"FE",X"19",X"78",X"28",X"2C",X"30",X"6B",X"FE",X"1A",
		X"30",X"67",X"FE",X"08",X"30",X"19",X"CD",X"33",X"2A",X"30",X"17",X"F5",X"CD",X"80",X"2D",X"2A",
		X"86",X"E2",X"29",X"18",X"2B",X"3C",X"2A",X"C7",X"E2",X"11",X"80",X"FF",X"19",X"18",X"20",X"CD",
		X"33",X"2A",X"F5",X"CD",X"00",X"2B",X"18",X"1B",X"FE",X"1E",X"38",X"40",X"D6",X"2A",X"FE",X"40",
		X"30",X"37",X"3A",X"22",X"E0",X"E6",X"02",X"20",X"30",X"CD",X"47",X"2A",X"2A",X"C7",X"E2",X"F5",
		X"CD",X"BB",X"2A",X"21",X"88",X"E2",X"7E",X"A7",X"20",X"0F",X"DD",X"7E",X"00",X"FE",X"1A",X"20",
		X"08",X"DD",X"36",X"00",X"1A",X"DD",X"36",X"0F",X"5E",X"F1",X"CD",X"85",X"21",X"DD",X"6E",X"0B",
		X"CD",X"E2",X"24",X"CD",X"C4",X"2C",X"38",X"1C",X"C9",X"AF",X"18",X"D0",X"3A",X"22",X"E0",X"E6",
		X"02",X"20",X"F6",X"CD",X"33",X"2A",X"18",X"C4",X"CD",X"5D",X"2A",X"3C",X"38",X"01",X"AF",X"21",
		X"00",X"01",X"18",X"BB",X"DD",X"7E",X"05",X"06",X"40",X"C6",X"08",X"FA",X"04",X"2A",X"FE",X"11",
		X"04",X"38",X"01",X"04",X"DD",X"70",X"0D",X"78",X"D6",X"41",X"28",X"0F",X"3D",X"0E",X"04",X"28",
		X"02",X"0E",X"0C",X"CD",X"BA",X"22",X"38",X"0C",X"79",X"C6",X"04",X"4F",X"CD",X"BA",X"22",X"38",
		X"03",X"C3",X"C0",X"40",X"CB",X"20",X"05",X"DD",X"70",X"05",X"DD",X"36",X"0F",X"01",X"DD",X"36",
		X"00",X"1B",X"C9",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"0E",X"00",X"3F",X"CB",X"11",X"C6",X"1A",
		X"FE",X"35",X"79",X"3C",X"D8",X"AF",X"C9",X"3A",X"C1",X"E2",X"DD",X"96",X"03",X"0E",X"00",X"CB",
		X"11",X"C6",X"40",X"FE",X"81",X"30",X"EE",X"D6",X"44",X"FE",X"F9",X"18",X"E5",X"CD",X"53",X"2C",
		X"D8",X"CD",X"EE",X"23",X"D8",X"CD",X"08",X"2F",X"D8",X"C3",X"33",X"2E",X"3A",X"22",X"E0",X"DD",
		X"AE",X"01",X"1F",X"D8",X"DD",X"35",X"0F",X"20",X"21",X"DD",X"7E",X"0D",X"DD",X"86",X"05",X"E6",
		X"07",X"F6",X"40",X"DD",X"77",X"0D",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"29",X"7C",X"FE",X"08",
		X"38",X"02",X"3E",X"07",X"EE",X"07",X"3C",X"DD",X"77",X"0F",X"DD",X"6E",X"08",X"DD",X"66",X"09",
		X"11",X"14",X"00",X"ED",X"52",X"30",X"03",X"21",X"00",X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",
		X"EB",X"CD",X"C7",X"24",X"CD",X"C4",X"2C",X"DA",X"C0",X"40",X"C9",X"DD",X"7E",X"00",X"FE",X"1A",
		X"20",X"03",X"2A",X"4F",X"E0",X"DD",X"5E",X"08",X"DD",X"56",X"09",X"ED",X"52",X"21",X"F2",X"FF",
		X"38",X"03",X"21",X"0E",X"00",X"19",X"DD",X"75",X"08",X"DD",X"74",X"09",X"EB",X"DD",X"7E",X"00",
		X"2A",X"86",X"E2",X"29",X"ED",X"52",X"38",X"0C",X"FE",X"18",X"C0",X"11",X"80",X"FF",X"19",X"D8",
		X"DD",X"34",X"00",X"C9",X"FE",X"19",X"C0",X"11",X"10",X"00",X"19",X"D8",X"DD",X"35",X"00",X"C9",
		X"DD",X"5E",X"08",X"DD",X"56",X"09",X"21",X"18",X"00",X"18",X"CA",X"21",X"D1",X"E2",X"7E",X"A7",
		X"28",X"01",X"35",X"3A",X"04",X"E7",X"FE",X"02",X"D0",X"2A",X"C9",X"E2",X"ED",X"5B",X"C7",X"E2",
		X"7C",X"A7",X"C8",X"ED",X"52",X"21",X"F2",X"FF",X"38",X"03",X"21",X"0E",X"00",X"19",X"22",X"C7",
		X"E2",X"3A",X"1D",X"E7",X"A7",X"C8",X"3A",X"22",X"E0",X"E6",X"03",X"C0",X"ED",X"5B",X"86",X"E2",
		X"CB",X"3C",X"CB",X"1D",X"AF",X"ED",X"52",X"DE",X"00",X"EB",X"2A",X"27",X"E7",X"19",X"22",X"27",
		X"E7",X"21",X"29",X"E7",X"8E",X"77",X"30",X"16",X"C6",X"04",X"30",X"0A",X"3A",X"0C",X"E7",X"3D",
		X"C8",X"11",X"E0",X"00",X"18",X"0D",X"F0",X"21",X"00",X"FC",X"22",X"28",X"E7",X"C9",X"A7",X"F8",
		X"11",X"C0",X"FF",X"3A",X"60",X"E3",X"A7",X"C0",X"3A",X"88",X"E2",X"FE",X"03",X"C8",X"DD",X"21",
		X"10",X"E3",X"DD",X"7E",X"00",X"A7",X"28",X"09",X"DD",X"21",X"80",X"E3",X"DD",X"7E",X"00",X"A7",
		X"C0",X"2A",X"0B",X"E3",X"19",X"DD",X"75",X"0B",X"DD",X"74",X"0C",X"D5",X"CD",X"60",X"24",X"38",
		X"22",X"DD",X"77",X"03",X"CD",X"71",X"2C",X"38",X"1A",X"2A",X"08",X"E3",X"29",X"DD",X"75",X"08",
		X"DD",X"74",X"09",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"00",X"D1",X"CD",X"C5",X"2B",X"DD",
		X"77",X"0E",X"C9",X"D1",X"C9",X"2A",X"28",X"E7",X"7A",X"ED",X"5B",X"CD",X"E2",X"87",X"38",X"27",
		X"19",X"38",X"03",X"21",X"20",X"00",X"22",X"28",X"E7",X"DD",X"36",X"00",X"19",X"21",X"0C",X"E7",
		X"7E",X"D6",X"01",X"27",X"77",X"21",X"11",X"E7",X"7E",X"D6",X"01",X"30",X"02",X"3E",X"09",X"77",
		X"C6",X"13",X"6F",X"26",X"E7",X"7E",X"C9",X"A7",X"ED",X"52",X"38",X"03",X"21",X"E0",X"FF",X"22",
		X"28",X"E7",X"DD",X"36",X"00",X"18",X"21",X"12",X"E7",X"7E",X"3C",X"FE",X"0A",X"38",X"E0",X"AF",
		X"18",X"DD",X"FE",X"C0",X"38",X"0B",X"21",X"12",X"E7",X"CD",X"36",X"2C",X"21",X"12",X"E7",X"18",
		X"C7",X"21",X"0C",X"E7",X"7E",X"C6",X"01",X"27",X"28",X"01",X"77",X"21",X"11",X"E7",X"CD",X"36",
		X"2C",X"21",X"11",X"E7",X"18",X"D3",X"7E",X"CD",X"F0",X"2B",X"DD",X"BE",X"0E",X"C8",X"4F",X"DD",
		X"7E",X"0E",X"E5",X"21",X"13",X"E7",X"06",X"0A",X"BE",X"28",X"04",X"23",X"10",X"FA",X"76",X"71",
		X"E1",X"77",X"C9",X"3A",X"91",X"E2",X"A7",X"28",X"18",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"C6",
		X"48",X"FE",X"9E",X"30",X"0C",X"21",X"30",X"00",X"DD",X"5E",X"06",X"DD",X"56",X"07",X"ED",X"52",
		X"D0",X"FD",X"21",X"92",X"E2",X"DD",X"5E",X"0B",X"DD",X"56",X"0C",X"DD",X"4E",X"03",X"06",X"04",
		X"FD",X"7E",X"00",X"A7",X"28",X"19",X"FD",X"7E",X"01",X"B9",X"30",X"13",X"FD",X"7E",X"02",X"B9",
		X"38",X"0D",X"FD",X"6E",X"03",X"FD",X"66",X"04",X"ED",X"52",X"30",X"03",X"24",X"28",X"0A",X"EB",
		X"11",X"08",X"00",X"FD",X"19",X"EB",X"10",X"D8",X"C9",X"FD",X"7E",X"05",X"C9",X"DD",X"6E",X"0B",
		X"DD",X"66",X"0C",X"ED",X"5B",X"0B",X"E3",X"ED",X"52",X"09",X"CB",X"2C",X"20",X"04",X"CB",X"1D",
		X"BD",X"C9",X"37",X"C9",X"DD",X"7E",X"07",X"87",X"87",X"4F",X"28",X"05",X"DD",X"7E",X"06",X"C6",
		X"28",X"FE",X"70",X"D8",X"CD",X"12",X"2C",X"AF",X"DD",X"77",X"00",X"C9",X"21",X"C4",X"E2",X"35",
		X"F0",X"23",X"7E",X"2B",X"77",X"3A",X"03",X"E3",X"32",X"C1",X"E2",X"C9",X"21",X"BC",X"E2",X"34",
		X"7E",X"FE",X"12",X"38",X"02",X"36",X"00",X"3A",X"04",X"E7",X"FE",X"02",X"D0",X"CD",X"45",X"2D",
		X"CD",X"8D",X"2D",X"11",X"1D",X"E7",X"1A",X"FE",X"02",X"30",X"0F",X"21",X"89",X"E2",X"3A",X"C6",
		X"E2",X"BE",X"30",X"04",X"EB",X"7E",X"3D",X"C0",X"34",X"C9",X"FD",X"21",X"92",X"E2",X"06",X"04",
		X"FD",X"CB",X"00",X"46",X"28",X"17",X"FD",X"5E",X"03",X"FD",X"56",X"04",X"2A",X"0B",X"E3",X"ED",
		X"52",X"11",X"A0",X"FE",X"19",X"CB",X"7C",X"20",X"04",X"FD",X"36",X"00",X"00",X"11",X"08",X"00",
		X"FD",X"19",X"10",X"DC",X"C9",X"CD",X"6D",X"2D",X"EE",X"1F",X"2A",X"CB",X"E2",X"5C",X"16",X"00",
		X"CB",X"3F",X"30",X"01",X"19",X"28",X"06",X"CB",X"23",X"CB",X"12",X"18",X"F3",X"ED",X"5B",X"7A",
		X"E0",X"ED",X"52",X"38",X"03",X"21",X"00",X"00",X"19",X"22",X"C9",X"E2",X"C9",X"3A",X"0C",X"E7",
		X"FE",X"0A",X"D8",X"D6",X"06",X"FE",X"14",X"D8",X"D6",X"06",X"FE",X"1E",X"D8",X"3E",X"1F",X"C9",
		X"21",X"D1",X"E2",X"7E",X"A7",X"C0",X"36",X"0F",X"3E",X"01",X"C3",X"B6",X"5E",X"21",X"8A",X"E2",
		X"11",X"8E",X"E2",X"01",X"5A",X"1F",X"CD",X"A8",X"2D",X"01",X"2F",X"07",X"CD",X"A8",X"2D",X"01",
		X"2F",X"1F",X"CD",X"A8",X"2D",X"01",X"46",X"0E",X"34",X"7E",X"B9",X"38",X"02",X"36",X"00",X"90",
		X"3E",X"00",X"17",X"12",X"23",X"13",X"C9",X"FD",X"21",X"92",X"E2",X"87",X"87",X"87",X"5F",X"16",
		X"00",X"FD",X"19",X"FD",X"75",X"03",X"FD",X"74",X"04",X"78",X"E6",X"01",X"FD",X"77",X"05",X"78",
		X"E6",X"FE",X"FD",X"77",X"02",X"FD",X"71",X"01",X"FD",X"36",X"00",X"01",X"C9",X"21",X"50",X"E4",
		X"11",X"1F",X"2E",X"06",X"05",X"36",X"17",X"CD",X"1A",X"2E",X"2C",X"CD",X"17",X"2E",X"7D",X"C6",
		X"06",X"6F",X"CD",X"1A",X"2E",X"2C",X"2C",X"36",X"41",X"2C",X"70",X"35",X"2C",X"2C",X"10",X"E5",
		X"21",X"13",X"E7",X"AF",X"77",X"23",X"3C",X"FE",X"0A",X"38",X"F9",X"3E",X"87",X"32",X"0C",X"E7",
		X"21",X"90",X"90",X"22",X"0D",X"E7",X"C9",X"CD",X"1A",X"2E",X"1A",X"23",X"13",X"77",X"C9",X"1C",
		X"67",X"18",X"E0",X"2A",X"3F",X"10",X"80",X"0B",X"8F",X"09",X"80",X"23",X"3F",X"08",X"20",X"04",
		X"8F",X"02",X"20",X"DD",X"E5",X"D1",X"7B",X"EE",X"90",X"5F",X"D5",X"FD",X"E1",X"FD",X"7E",X"00",
		X"D6",X"18",X"FE",X"03",X"30",X"42",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"C6",X"20",X"FE",X"41",
		X"D0",X"D6",X"06",X"47",X"FE",X"35",X"38",X"0E",X"CD",X"BA",X"2E",X"20",X"2B",X"FE",X"69",X"D0",
		X"3E",X"80",X"CB",X"10",X"17",X"C9",X"CD",X"BA",X"2E",X"20",X"1D",X"D6",X"04",X"FE",X"61",X"D0",
		X"11",X"E8",X"FF",X"D6",X"10",X"38",X"13",X"FE",X"41",X"38",X"1E",X"FD",X"6E",X"08",X"FD",X"66",
		X"09",X"19",X"FD",X"75",X"08",X"FD",X"74",X"09",X"AF",X"C9",X"DD",X"6E",X"08",X"DD",X"66",X"09",
		X"19",X"DD",X"75",X"08",X"DD",X"74",X"09",X"AF",X"C9",X"FE",X"1A",X"78",X"38",X"08",X"DD",X"E5",
		X"FD",X"E1",X"EE",X"3F",X"D6",X"0B",X"FE",X"1A",X"3E",X"00",X"17",X"87",X"3D",X"FD",X"77",X"05",
		X"FD",X"36",X"0F",X"01",X"FD",X"36",X"00",X"1B",X"E1",X"C9",X"DD",X"6E",X"0B",X"DD",X"66",X"0C",
		X"FD",X"5E",X"0B",X"FD",X"56",X"0C",X"ED",X"52",X"11",X"34",X"00",X"19",X"24",X"25",X"7D",X"C9",
		X"DD",X"6E",X"0B",X"DD",X"66",X"0C",X"29",X"5C",X"16",X"00",X"7D",X"2A",X"69",X"E0",X"19",X"5E",
		X"53",X"FE",X"70",X"38",X"02",X"23",X"5E",X"7A",X"E6",X"F0",X"67",X"7A",X"E6",X"0F",X"57",X"7B",
		X"E6",X"0F",X"BA",X"38",X"01",X"7A",X"87",X"87",X"87",X"C6",X"24",X"57",X"7B",X"E6",X"F0",X"BC",
		X"30",X"01",X"7C",X"CB",X"3F",X"C6",X"24",X"C9",X"3A",X"04",X"E7",X"A7",X"C8",X"CD",X"D0",X"2E",
		X"DD",X"BE",X"03",X"38",X"03",X"AF",X"37",X"C9",X"7A",X"DD",X"BE",X"03",X"D0",X"3E",X"01",X"C9",
		X"2A",X"86",X"E2",X"11",X"00",X"04",X"CD",X"89",X"23",X"A7",X"ED",X"52",X"30",X"03",X"DD",X"35",
		X"07",X"DD",X"75",X"05",X"DD",X"74",X"06",X"EB",X"29",X"29",X"7C",X"29",X"29",X"84",X"5F",X"6F",
		X"26",X"00",X"54",X"3A",X"C1",X"E2",X"87",X"87",X"DD",X"7E",X"0E",X"3C",X"38",X"30",X"29",X"FE",
		X"02",X"38",X"01",X"19",X"29",X"19",X"CD",X"A2",X"23",X"21",X"F0",X"2F",X"19",X"7E",X"FE",X"38",
		X"38",X"08",X"DD",X"CB",X"0E",X"7E",X"28",X"02",X"C6",X"04",X"DD",X"77",X"0D",X"DD",X"7E",X"06",
		X"DD",X"CB",X"07",X"46",X"28",X"0E",X"FE",X"E8",X"DA",X"B8",X"32",X"C3",X"C0",X"40",X"FE",X"02",
		X"30",X"D2",X"18",X"D2",X"D6",X"28",X"FE",X"1A",X"30",X"5A",X"3A",X"0D",X"E3",X"FE",X"25",X"D0",
		X"6F",X"26",X"00",X"11",X"E4",X"2F",X"19",X"3A",X"03",X"E3",X"86",X"DD",X"96",X"03",X"C6",X"17",
		X"FE",X"2F",X"30",X"49",X"01",X"2F",X"02",X"D6",X"05",X"38",X"16",X"06",X"04",X"FE",X"12",X"38",
		X"05",X"D6",X"12",X"01",X"2B",X"01",X"FE",X"09",X"38",X"07",X"05",X"FE",X"12",X"38",X"02",X"06",
		X"02",X"DD",X"7E",X"0E",X"80",X"F2",X"C9",X"2F",X"AF",X"FE",X"04",X"38",X"02",X"3E",X"03",X"D6",
		X"02",X"DD",X"77",X"0E",X"3A",X"04",X"D0",X"E6",X"40",X"28",X"12",X"79",X"32",X"0D",X"E3",X"3E",
		X"13",X"C3",X"18",X"23",X"D6",X"20",X"30",X"05",X"3E",X"19",X"CD",X"B6",X"5E",X"C3",X"C0",X"40",
		X"3B",X"3A",X"39",X"38",X"38",X"38",X"37",X"37",X"37",X"37",X"36",X"36",X"36",X"35",X"35",X"35",
		X"34",X"34",X"33",X"33",X"F8",X"FC",X"00",X"05",X"09",X"CD",X"62",X"30",X"DD",X"7E",X"07",X"3C",
		X"FE",X"02",X"DA",X"B4",X"32",X"DD",X"7E",X"20",X"DD",X"B6",X"B0",X"C0",X"DD",X"34",X"00",X"3E",
		X"1F",X"32",X"20",X"E3",X"32",X"40",X"E3",X"3E",X"4A",X"32",X"2D",X"E3",X"32",X"4D",X"E3",X"3E",
		X"8E",X"32",X"4E",X"E3",X"AF",X"32",X"2E",X"E3",X"DD",X"7E",X"03",X"D6",X"08",X"32",X"23",X"E3",
		X"C6",X"10",X"32",X"43",X"E3",X"C9",X"CD",X"62",X"30",X"DD",X"36",X"0D",X"49",X"0E",X"14",X"C5",
		X"01",X"50",X"00",X"CD",X"AD",X"2C",X"C1",X"7C",X"A7",X"FA",X"B4",X"32",X"CD",X"BA",X"22",X"C3",
		X"C0",X"40",X"DD",X"7E",X"0E",X"2A",X"86",X"E2",X"5D",X"54",X"29",X"29",X"29",X"A7",X"28",X"04",
		X"19",X"3D",X"20",X"FC",X"29",X"6C",X"26",X"00",X"29",X"29",X"11",X"00",X"01",X"19",X"22",X"52",
		X"E0",X"C3",X"C7",X"24",X"3A",X"60",X"E3",X"A7",X"CA",X"B8",X"32",X"DD",X"7E",X"0E",X"3C",X"FE",
		X"0E",X"28",X"35",X"38",X"35",X"D6",X"02",X"FE",X"80",X"28",X"2D",X"FE",X"8D",X"20",X"2B",X"2A",
		X"66",X"E3",X"7C",X"A7",X"20",X"20",X"7D",X"FE",X"20",X"38",X"1B",X"2A",X"52",X"E0",X"29",X"29",
		X"29",X"29",X"29",X"3A",X"6D",X"E0",X"84",X"30",X"02",X"3E",X"FF",X"DD",X"86",X"0F",X"DD",X"77",
		X"0F",X"30",X"03",X"CD",X"0E",X"31",X"3E",X"0C",X"EE",X"80",X"DD",X"77",X"0E",X"E6",X"0F",X"5F",
		X"16",X"00",X"21",X"F4",X"30",X"19",X"7E",X"A7",X"28",X"08",X"DD",X"7E",X"0D",X"EE",X"01",X"DD",
		X"77",X"0D",X"2A",X"66",X"E3",X"ED",X"52",X"11",X"F3",X"FF",X"19",X"DD",X"75",X"06",X"DD",X"74",
		X"07",X"C3",X"C0",X"40",X"00",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"25",X"FF",X"4A",X"FE",X"6F",X"FD",X"FD",X"21",
		X"E0",X"E3",X"11",X"10",X"00",X"06",X"06",X"FD",X"7E",X"00",X"A7",X"28",X"05",X"FD",X"19",X"10",
		X"F6",X"C9",X"FD",X"36",X"00",X"20",X"FD",X"36",X"0D",X"4C",X"2A",X"52",X"E0",X"FD",X"75",X"08",
		X"FD",X"74",X"09",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"2A",X"66",X"E3",X"11",X"D8",X"FF",X"19",
		X"FD",X"75",X"06",X"FD",X"74",X"07",X"ED",X"5F",X"E6",X"06",X"5F",X"16",X"00",X"21",X"06",X"31",
		X"19",X"5E",X"23",X"56",X"3A",X"63",X"E3",X"DD",X"96",X"03",X"87",X"38",X"08",X"7B",X"ED",X"44",
		X"5F",X"7A",X"ED",X"44",X"57",X"FD",X"72",X"05",X"FD",X"73",X"04",X"FD",X"36",X"0E",X"F0",X"C9",
		X"3A",X"22",X"E0",X"DD",X"AE",X"0D",X"1F",X"D8",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"11",X"C0",
		X"FF",X"19",X"38",X"03",X"21",X"00",X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",X"ED",X"5B",X"86",
		X"E2",X"ED",X"52",X"29",X"EB",X"DD",X"66",X"06",X"DD",X"6E",X"0C",X"19",X"DD",X"74",X"06",X"DD",
		X"75",X"0C",X"DD",X"7E",X"07",X"30",X"01",X"3C",X"CB",X"12",X"30",X"01",X"3D",X"DD",X"77",X"07",
		X"A7",X"28",X"07",X"7C",X"C6",X"10",X"FE",X"20",X"30",X"24",X"DD",X"7E",X"05",X"DD",X"86",X"04",
		X"28",X"03",X"DD",X"77",X"05",X"87",X"6F",X"9F",X"67",X"29",X"DD",X"5E",X"02",X"DD",X"56",X"03",
		X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",X"7C",X"C6",X"08",X"FE",X"D0",X"38",X"05",X"DD",X"36",
		X"00",X"00",X"C9",X"DD",X"7E",X"0B",X"DD",X"46",X"0E",X"CB",X"40",X"20",X"4A",X"C6",X"04",X"DD",
		X"77",X"0B",X"B8",X"38",X"0D",X"67",X"CB",X"38",X"78",X"CB",X"3F",X"80",X"CB",X"C7",X"DD",X"77",
		X"0E",X"7C",X"DD",X"86",X"0A",X"DD",X"77",X"0A",X"30",X"08",X"DD",X"7E",X"0D",X"EE",X"01",X"DD",
		X"77",X"0D",X"CD",X"C0",X"40",X"0E",X"18",X"CD",X"BA",X"22",X"D0",X"DD",X"7E",X"05",X"21",X"FD",
		X"DE",X"87",X"30",X"08",X"7D",X"ED",X"44",X"6F",X"7C",X"ED",X"44",X"67",X"DD",X"74",X"05",X"DD",
		X"75",X"04",X"DD",X"36",X"0E",X"F0",X"C9",X"D6",X"04",X"30",X"04",X"DD",X"35",X"0E",X"AF",X"DD",
		X"77",X"0B",X"18",X"BE",X"DD",X"6E",X"0B",X"CD",X"E2",X"24",X"24",X"28",X"6B",X"25",X"C0",X"DD",
		X"4E",X"0D",X"CD",X"BA",X"22",X"D8",X"DD",X"4E",X"0D",X"79",X"FE",X"2C",X"C8",X"FE",X"40",X"C8",
		X"DD",X"7E",X"07",X"A7",X"C0",X"06",X"00",X"21",X"B8",X"46",X"09",X"EB",X"FD",X"21",X"10",X"E3",
		X"CD",X"77",X"32",X"FD",X"21",X"80",X"E3",X"FD",X"7E",X"00",X"D6",X"18",X"FE",X"03",X"D0",X"FD",
		X"7E",X"07",X"A7",X"C0",X"62",X"6B",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"86",X"23",X"BE",X"D0",
		X"23",X"FD",X"7E",X"06",X"DD",X"96",X"06",X"1F",X"86",X"23",X"BE",X"D0",X"87",X"BE",X"3E",X"FF",
		X"30",X"02",X"3E",X"01",X"FD",X"77",X"05",X"FD",X"36",X"0F",X"01",X"FD",X"36",X"00",X"1B",X"3E",
		X"17",X"C3",X"B6",X"5E",X"AF",X"32",X"88",X"E2",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"6E",X"0B",
		X"CD",X"E2",X"24",X"24",X"20",X"05",X"7D",X"FE",X"D0",X"38",X"ED",X"C3",X"C0",X"40",X"DD",X"6E",
		X"0B",X"CD",X"E2",X"24",X"24",X"28",X"E1",X"25",X"C0",X"3A",X"04",X"D0",X"E6",X"40",X"C8",X"FD",
		X"21",X"00",X"E3",X"FD",X"7E",X"00",X"FE",X"04",X"30",X"4C",X"7D",X"D6",X"08",X"FE",X"40",X"D0",
		X"4F",X"CD",X"29",X"23",X"2A",X"32",X"E3",X"CD",X"42",X"33",X"38",X"0E",X"2A",X"34",X"E3",X"CD",
		X"42",X"33",X"38",X"06",X"2A",X"38",X"E3",X"CD",X"42",X"33",X"47",X"79",X"FE",X"30",X"30",X"19",
		X"78",X"06",X"14",X"D6",X"08",X"30",X"02",X"06",X"10",X"FD",X"70",X"0D",X"FD",X"36",X"00",X"09",
		X"FD",X"36",X"0F",X"0A",X"3E",X"1F",X"C3",X"B6",X"5E",X"FD",X"36",X"00",X"05",X"FD",X"36",X"0F",
		X"0A",X"3E",X"14",X"C3",X"B6",X"5E",X"FE",X"05",X"C0",X"7D",X"D6",X"20",X"D0",X"FD",X"36",X"0F",
		X"01",X"C9",X"FD",X"7E",X"03",X"95",X"38",X"03",X"94",X"38",X"05",X"C6",X"08",X"FE",X"10",X"C9",
		X"7D",X"FE",X"86",X"28",X"04",X"FE",X"26",X"20",X"1B",X"DD",X"7E",X"06",X"D6",X"30",X"30",X"14",
		X"21",X"D8",X"E2",X"CB",X"4E",X"20",X"0D",X"36",X"02",X"23",X"36",X"36",X"3E",X"14",X"CD",X"B6",
		X"5E",X"CD",X"B8",X"32",X"E1",X"C9",X"DD",X"6E",X"0B",X"CD",X"E2",X"24",X"24",X"CA",X"B8",X"32",
		X"25",X"C0",X"3A",X"00",X"E3",X"FE",X"04",X"38",X"03",X"FE",X"0B",X"C0",X"7D",X"D6",X"30",X"FE",
		X"0C",X"D0",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"C6",X"0A",X"FE",X"24",X"D0",X"DD",X"7E",X"0D",
		X"FE",X"06",X"20",X"05",X"3A",X"D8",X"E2",X"A7",X"C8",X"CD",X"B8",X"32",X"DD",X"6E",X"08",X"DD",
		X"66",X"09",X"DD",X"7E",X"0D",X"01",X"80",X"00",X"70",X"09",X"70",X"FE",X"05",X"38",X"08",X"20",
		X"0C",X"23",X"23",X"70",X"ED",X"42",X"70",X"0E",X"01",X"C3",X"73",X"59",X"C9",X"09",X"70",X"18",
		X"F6",X"AF",X"18",X"13",X"DD",X"35",X"0F",X"CA",X"DE",X"57",X"DD",X"7E",X"0F",X"11",X"A4",X"C0",
		X"21",X"9F",X"40",X"E6",X"10",X"20",X"01",X"6F",X"ED",X"53",X"14",X"E2",X"1E",X"94",X"ED",X"53",
		X"18",X"E2",X"1E",X"84",X"ED",X"53",X"1C",X"E2",X"22",X"16",X"E2",X"CD",X"08",X"34",X"22",X"1A",
		X"E2",X"CD",X"08",X"34",X"22",X"1E",X"E2",X"C9",X"7D",X"A7",X"C8",X"2C",X"C9",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"19",X"DD",X"75",X"02",X"DD",X"74",X"03",
		X"DD",X"7E",X"0E",X"FE",X"08",X"30",X"3E",X"4F",X"7C",X"E6",X"FC",X"DD",X"BE",X"0C",X"28",X"72",
		X"79",X"FE",X"06",X"CA",X"B5",X"34",X"30",X"1F",X"CB",X"3F",X"30",X"1B",X"11",X"40",X"00",X"3D",
		X"28",X"08",X"1E",X"A0",X"3D",X"28",X"03",X"11",X"C0",X"FF",X"DD",X"6E",X"0A",X"DD",X"66",X"06",
		X"19",X"DD",X"75",X"0A",X"DD",X"74",X"06",X"DD",X"7E",X"05",X"87",X"3E",X"51",X"CE",X"00",X"DD",
		X"77",X"0D",X"C3",X"C0",X"40",X"21",X"10",X"00",X"20",X"03",X"21",X"F0",X"FF",X"19",X"DD",X"75",
		X"04",X"DD",X"74",X"05",X"11",X"06",X"00",X"CB",X"24",X"30",X"03",X"11",X"FA",X"FF",X"DD",X"6E",
		X"08",X"DD",X"66",X"09",X"19",X"DD",X"75",X"08",X"DD",X"74",X"09",X"EB",X"7B",X"B2",X"20",X"BA",
		X"DD",X"7E",X"0E",X"EE",X"0F",X"DD",X"77",X"0E",X"FE",X"06",X"28",X"BB",X"DD",X"36",X"0C",X"40",
		X"18",X"B5",X"FE",X"E0",X"CA",X"B8",X"32",X"DD",X"36",X"0C",X"E0",X"79",X"FE",X"06",X"DE",X"FE",
		X"DD",X"77",X"0E",X"18",X"A2",X"FD",X"21",X"F0",X"E1",X"11",X"04",X"00",X"06",X"07",X"7C",X"21",
		X"06",X"35",X"BE",X"30",X"07",X"23",X"FD",X"19",X"10",X"F8",X"18",X"8B",X"3E",X"D0",X"32",X"5B",
		X"E0",X"11",X"C0",X"A2",X"DD",X"7E",X"0C",X"FE",X"E0",X"28",X"09",X"7E",X"2F",X"47",X"CD",X"99",
		X"42",X"C3",X"57",X"34",X"78",X"FE",X"07",X"C2",X"57",X"34",X"06",X"C0",X"14",X"CD",X"99",X"42",
		X"78",X"D6",X"10",X"47",X"7A",X"FE",X"A9",X"38",X"F3",X"16",X"00",X"CD",X"99",X"42",X"3E",X"FF",
		X"32",X"D7",X"E2",X"C3",X"57",X"34",X"8C",X"7E",X"68",X"62",X"57",X"48",X"40",X"DD",X"6E",X"0B",
		X"CD",X"E2",X"24",X"24",X"CA",X"B8",X"32",X"25",X"C0",X"3A",X"D8",X"E2",X"A7",X"C0",X"3A",X"00",
		X"E3",X"FE",X"04",X"D0",X"7D",X"D6",X"08",X"FE",X"30",X"D0",X"3A",X"03",X"E3",X"DD",X"96",X"03",
		X"D6",X"03",X"FE",X"12",X"D0",X"21",X"01",X"A4",X"22",X"D8",X"E2",X"C9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"04",X"E7",X"FE",X"02",X"D2",X"BF",X"36",X"21",X"74",X"48",X"CD",X"9C",X"36",X"85",X"6F",
		X"30",X"01",X"24",X"22",X"09",X"E7",X"21",X"A8",X"4C",X"CD",X"9C",X"36",X"22",X"69",X"E0",X"2A",
		X"05",X"E7",X"7C",X"FE",X"02",X"38",X"03",X"3E",X"02",X"67",X"87",X"87",X"84",X"85",X"21",X"E9",
		X"3E",X"CD",X"9F",X"36",X"22",X"CF",X"E2",X"21",X"C0",X"4E",X"CD",X"9C",X"36",X"0F",X"0F",X"0F",
		X"47",X"E6",X"E0",X"57",X"78",X"E6",X"1F",X"28",X"0E",X"47",X"7E",X"F5",X"CD",X"AC",X"36",X"F1",
		X"BE",X"38",X"F7",X"28",X"F5",X"10",X"F3",X"7E",X"BA",X"30",X"0A",X"F5",X"CD",X"AC",X"36",X"F1",
		X"BE",X"38",X"F4",X"28",X"F2",X"22",X"0F",X"E7",X"3E",X"F0",X"32",X"B6",X"E2",X"3E",X"06",X"32",
		X"6C",X"E0",X"11",X"D0",X"FE",X"2A",X"0B",X"E3",X"19",X"22",X"0B",X"E3",X"CD",X"1A",X"38",X"3A",
		X"0B",X"E7",X"A7",X"20",X"F7",X"21",X"6C",X"E0",X"11",X"80",X"00",X"7E",X"FE",X"03",X"20",X"E5",
		X"1E",X"30",X"2A",X"0B",X"E3",X"19",X"22",X"0B",X"E3",X"C3",X"42",X"24",X"3A",X"05",X"E7",X"87",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"3A",X"0C",X"E3",X"C9",X"23",X"7E",X"23",X"23",
		X"FE",X"09",X"28",X"09",X"FE",X"08",X"D0",X"3D",X"2B",X"FE",X"04",X"D0",X"23",X"23",X"C9",X"21",
		X"2A",X"86",X"FD",X"21",X"C4",X"00",X"01",X"15",X"0C",X"C5",X"11",X"00",X"03",X"FD",X"46",X"00",
		X"FD",X"23",X"E5",X"CD",X"8E",X"37",X"2B",X"2B",X"0D",X"10",X"F8",X"15",X"CD",X"8E",X"37",X"2B",
		X"2B",X"0D",X"20",X"F8",X"E1",X"01",X"80",X"00",X"09",X"C1",X"10",X"DD",X"21",X"BE",X"E2",X"36",
		X"00",X"3A",X"0B",X"E3",X"47",X"CD",X"3E",X"37",X"3A",X"05",X"E7",X"87",X"5F",X"16",X"00",X"21",
		X"82",X"03",X"19",X"5E",X"23",X"56",X"21",X"2C",X"80",X"1A",X"4F",X"13",X"1A",X"FE",X"F0",X"38",
		X"08",X"87",X"87",X"87",X"87",X"A9",X"4F",X"18",X"F2",X"77",X"23",X"71",X"23",X"A7",X"20",X"EB",
		X"7D",X"E6",X"1F",X"3E",X"00",X"20",X"F2",X"C5",X"01",X"6C",X"00",X"09",X"C1",X"7C",X"FE",X"8C",
		X"38",X"D9",X"C9",X"3A",X"0B",X"E3",X"21",X"B6",X"E2",X"47",X"96",X"FE",X"05",X"D8",X"70",X"21",
		X"BE",X"E2",X"7E",X"34",X"4F",X"E6",X"07",X"87",X"5F",X"16",X"00",X"21",X"D0",X"00",X"19",X"5E",
		X"23",X"56",X"FD",X"21",X"00",X"00",X"FD",X"19",X"21",X"2A",X"86",X"1E",X"00",X"FD",X"7E",X"00",
		X"A7",X"C8",X"47",X"FD",X"23",X"16",X"CB",X"DD",X"21",X"5D",X"37",X"DD",X"E5",X"17",X"38",X"13",
		X"17",X"38",X"3C",X"17",X"38",X"2C",X"17",X"CD",X"D6",X"37",X"CD",X"F6",X"37",X"D5",X"CD",X"CD",
		X"37",X"D1",X"C9",X"CD",X"D6",X"37",X"CD",X"F6",X"37",X"78",X"E6",X"07",X"83",X"5F",X"CD",X"91",
		X"37",X"73",X"23",X"72",X"7D",X"EE",X"80",X"6F",X"3E",X"0B",X"94",X"67",X"7A",X"EE",X"10",X"57",
		X"2B",X"C9",X"CD",X"D6",X"37",X"CD",X"F6",X"37",X"78",X"E6",X"01",X"C6",X"08",X"18",X"DD",X"CD",
		X"EF",X"37",X"FD",X"7E",X"00",X"CD",X"F6",X"37",X"D5",X"78",X"1F",X"E6",X"0E",X"5F",X"AF",X"57",
		X"ED",X"52",X"78",X"E6",X"03",X"1F",X"57",X"1E",X"00",X"CB",X"1B",X"19",X"D1",X"FD",X"7E",X"00",
		X"FD",X"23",X"E6",X"7F",X"18",X"B7",X"17",X"30",X"0B",X"17",X"30",X"11",X"D5",X"11",X"7E",X"FF",
		X"19",X"D1",X"18",X"0B",X"D5",X"11",X"80",X"00",X"19",X"D1",X"17",X"38",X"02",X"2D",X"2D",X"17",
		X"D0",X"CB",X"E2",X"CB",X"EA",X"C9",X"17",X"30",X"06",X"CB",X"59",X"C0",X"15",X"15",X"C9",X"CB",
		X"59",X"20",X"F9",X"C9",X"FD",X"2A",X"57",X"E0",X"ED",X"4B",X"59",X"E0",X"3A",X"BD",X"E2",X"C3",
		X"D0",X"38",X"3A",X"04",X"E7",X"FE",X"02",X"D2",X"33",X"37",X"3A",X"22",X"E0",X"32",X"5F",X"E0",
		X"3A",X"0B",X"E7",X"3D",X"28",X"DE",X"3D",X"CA",X"B1",X"3C",X"2A",X"0B",X"E3",X"11",X"30",X"01",
		X"19",X"22",X"67",X"E0",X"29",X"7C",X"21",X"B6",X"E2",X"BE",X"C8",X"77",X"87",X"87",X"87",X"87",
		X"32",X"BA",X"E2",X"87",X"4F",X"E6",X"60",X"6F",X"26",X"80",X"22",X"B8",X"E2",X"21",X"00",X"E5",
		X"87",X"6F",X"06",X"10",X"11",X"B7",X"08",X"3A",X"04",X"E7",X"3D",X"28",X"03",X"11",X"BE",X"01",
		X"72",X"23",X"73",X"23",X"72",X"23",X"72",X"23",X"10",X"F6",X"21",X"6C",X"E0",X"7E",X"A7",X"28",
		X"01",X"35",X"2A",X"CF",X"E2",X"3A",X"68",X"E0",X"BE",X"38",X"05",X"23",X"23",X"23",X"18",X"F8",
		X"23",X"7E",X"E6",X"80",X"32",X"D2",X"E2",X"7E",X"E6",X"7F",X"5F",X"16",X"00",X"ED",X"53",X"CD",
		X"E2",X"23",X"6E",X"62",X"29",X"29",X"29",X"29",X"22",X"CB",X"E2",X"21",X"00",X"00",X"22",X"60",
		X"E0",X"21",X"0B",X"E7",X"34",X"2A",X"09",X"E7",X"7E",X"87",X"CB",X"69",X"28",X"05",X"23",X"3C",
		X"22",X"09",X"E7",X"32",X"BD",X"E2",X"6F",X"26",X"00",X"11",X"38",X"4A",X"29",X"29",X"19",X"5E",
		X"23",X"56",X"23",X"ED",X"53",X"BF",X"E2",X"5E",X"23",X"56",X"FD",X"21",X"00",X"00",X"FD",X"19",
		X"0F",X"D6",X"B4",X"FE",X"0C",X"D2",X"93",X"39",X"FD",X"7E",X"00",X"FD",X"23",X"47",X"A7",X"F2",
		X"0D",X"39",X"E6",X"0F",X"87",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",X"21",X"B6",X"47",X"19",
		X"EB",X"2A",X"B8",X"E2",X"78",X"1F",X"1F",X"1F",X"1F",X"E6",X"07",X"C6",X"02",X"47",X"C5",X"CD",
		X"0B",X"3B",X"C1",X"10",X"F9",X"22",X"B8",X"E2",X"FD",X"22",X"57",X"E0",X"C9",X"28",X"4F",X"FE",
		X"40",X"30",X"0F",X"2A",X"B8",X"E2",X"C5",X"11",X"6A",X"48",X"CD",X"0B",X"3B",X"C1",X"10",X"F6",
		X"18",X"E3",X"2A",X"B8",X"E2",X"E6",X"0F",X"57",X"7C",X"E6",X"F0",X"B2",X"67",X"7D",X"E6",X"70",
		X"D6",X"02",X"6F",X"78",X"1F",X"1F",X"E6",X"04",X"FE",X"04",X"DE",X"3F",X"4F",X"E5",X"11",X"7F",
		X"00",X"3E",X"7C",X"06",X"04",X"77",X"2C",X"36",X"09",X"3C",X"19",X"10",X"F8",X"E1",X"11",X"7A",
		X"00",X"CD",X"7C",X"39",X"4F",X"CD",X"83",X"39",X"CD",X"83",X"39",X"CD",X"7C",X"39",X"21",X"39",
		X"E3",X"CD",X"25",X"3B",X"2B",X"2B",X"CD",X"25",X"3B",X"CD",X"25",X"3B",X"2A",X"67",X"E0",X"2E",
		X"90",X"22",X"3B",X"E3",X"3E",X"24",X"32",X"30",X"E3",X"C3",X"61",X"3B",X"06",X"02",X"2C",X"2C",
		X"79",X"18",X"04",X"06",X"03",X"3E",X"80",X"2C",X"2C",X"77",X"3C",X"FE",X"C8",X"28",X"FB",X"10",
		X"F6",X"19",X"C9",X"FD",X"7E",X"00",X"47",X"FD",X"23",X"17",X"30",X"3B",X"17",X"30",X"32",X"17",
		X"D2",X"28",X"3A",X"17",X"30",X"7C",X"17",X"D2",X"66",X"3A",X"17",X"D2",X"D1",X"3A",X"17",X"D2",
		X"00",X"3B",X"17",X"38",X"16",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"FD",X"23",X"FD",X"23",X"FD",
		X"22",X"5D",X"E0",X"FD",X"21",X"00",X"00",X"FD",X"19",X"18",X"C8",X"FD",X"2A",X"5D",X"E0",X"18",
		X"C2",X"78",X"E6",X"3F",X"47",X"18",X"09",X"3A",X"61",X"E0",X"FD",X"AE",X"00",X"4F",X"FD",X"23",
		X"2A",X"B8",X"E2",X"FD",X"5E",X"00",X"FD",X"23",X"3A",X"61",X"E0",X"57",X"CB",X"6A",X"20",X"0E",
		X"73",X"23",X"71",X"23",X"7D",X"E6",X"1F",X"CC",X"4F",X"3B",X"10",X"F4",X"18",X"0C",X"71",X"2B",
		X"73",X"7D",X"2B",X"E6",X"1F",X"CC",X"3C",X"3B",X"10",X"F4",X"22",X"B8",X"E2",X"3A",X"22",X"E0",
		X"21",X"5F",X"E0",X"AE",X"E6",X"FE",X"CA",X"93",X"39",X"FD",X"22",X"57",X"E0",X"ED",X"43",X"59",
		X"E0",X"C9",X"78",X"E6",X"0F",X"47",X"18",X"0D",X"78",X"E6",X"1F",X"47",X"3A",X"61",X"E0",X"FD",
		X"AE",X"00",X"4F",X"FD",X"23",X"2A",X"B8",X"E2",X"3A",X"61",X"E0",X"57",X"CB",X"6A",X"20",X"13",
		X"FD",X"7E",X"00",X"77",X"FD",X"23",X"23",X"71",X"23",X"7D",X"E6",X"1F",X"CC",X"4F",X"3B",X"10",
		X"EF",X"18",X"B7",X"71",X"2B",X"FD",X"7E",X"00",X"77",X"FD",X"23",X"7D",X"2B",X"E6",X"1F",X"CC",
		X"3C",X"3B",X"10",X"EF",X"18",X"A4",X"ED",X"5B",X"60",X"E0",X"3A",X"B8",X"E2",X"E6",X"60",X"87",
		X"6F",X"78",X"E6",X"03",X"B5",X"21",X"00",X"E5",X"CB",X"62",X"28",X"02",X"EE",X"01",X"CB",X"50",
		X"6F",X"20",X"35",X"FD",X"7E",X"00",X"87",X"87",X"FD",X"23",X"CB",X"6A",X"28",X"02",X"EE",X"3C",
		X"85",X"6F",X"FD",X"7E",X"00",X"A7",X"28",X"15",X"83",X"CB",X"62",X"28",X"03",X"D6",X"C0",X"2F",
		X"77",X"FD",X"23",X"CB",X"6A",X"28",X"0B",X"2B",X"2B",X"2B",X"2B",X"18",X"E5",X"FD",X"23",X"C3",
		X"93",X"39",X"23",X"23",X"23",X"23",X"18",X"DA",X"FD",X"7E",X"00",X"83",X"CB",X"62",X"28",X"03",
		X"D6",X"C0",X"2F",X"06",X"10",X"77",X"23",X"23",X"23",X"23",X"10",X"F9",X"FD",X"23",X"C3",X"93",
		X"39",X"2A",X"B8",X"E2",X"57",X"87",X"30",X"06",X"F5",X"7D",X"EE",X"1F",X"6F",X"F1",X"87",X"30",
		X"08",X"7C",X"EE",X"0B",X"67",X"7D",X"EE",X"80",X"6F",X"22",X"B8",X"E2",X"7A",X"0F",X"0F",X"21",
		X"61",X"E0",X"AE",X"E6",X"30",X"77",X"FD",X"7E",X"00",X"2B",X"77",X"FD",X"23",X"C3",X"93",X"39",
		X"17",X"3E",X"10",X"30",X"01",X"87",X"A9",X"4F",X"C3",X"93",X"39",X"01",X"07",X"0A",X"1A",X"77",
		X"23",X"71",X"23",X"13",X"10",X"F8",X"06",X"06",X"3E",X"BC",X"77",X"23",X"71",X"23",X"10",X"FA",
		X"01",X"60",X"00",X"09",X"C9",X"FD",X"7E",X"00",X"FD",X"23",X"47",X"E6",X"07",X"87",X"87",X"87",
		X"C6",X"14",X"77",X"2B",X"78",X"E6",X"F8",X"D6",X"02",X"77",X"2B",X"C9",X"D5",X"CB",X"62",X"11",
		X"A0",X"FF",X"20",X"16",X"11",X"A0",X"00",X"19",X"7C",X"D1",X"FE",X"8C",X"30",X"12",X"C9",X"D5",
		X"CB",X"62",X"11",X"60",X"00",X"28",X"F0",X"11",X"60",X"FF",X"19",X"7C",X"D1",X"FE",X"80",X"D0",
		X"E1",X"21",X"0B",X"E7",X"34",X"ED",X"5B",X"BF",X"E2",X"DD",X"21",X"00",X"00",X"DD",X"19",X"3A",
		X"B8",X"E2",X"87",X"E6",X"C0",X"32",X"B8",X"E2",X"DD",X"7E",X"00",X"47",X"1F",X"1F",X"E6",X"3C",
		X"2A",X"B8",X"E2",X"B5",X"6F",X"DD",X"7E",X"01",X"1F",X"CB",X"1D",X"E6",X"0F",X"F6",X"80",X"67",
		X"22",X"27",X"E0",X"78",X"E6",X"0F",X"C8",X"DD",X"23",X"DD",X"23",X"3D",X"CA",X"42",X"3C",X"3D",
		X"28",X"04",X"FE",X"0A",X"38",X"09",X"21",X"05",X"E7",X"5E",X"1C",X"1D",X"28",X"01",X"3C",X"87",
		X"87",X"5F",X"16",X"00",X"21",X"A9",X"01",X"19",X"5E",X"23",X"56",X"23",X"FD",X"21",X"00",X"00",
		X"FD",X"19",X"7E",X"E6",X"0F",X"47",X"7E",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"4F",X"ED",X"43",
		X"29",X"E0",X"23",X"7E",X"5F",X"E6",X"0F",X"FE",X"0D",X"20",X"0A",X"DD",X"7E",X"FF",X"87",X"30",
		X"04",X"7B",X"EE",X"05",X"5F",X"2A",X"27",X"E0",X"DD",X"7E",X"FF",X"1F",X"E6",X"10",X"AB",X"5F",
		X"FD",X"7E",X"00",X"E6",X"1F",X"47",X"FD",X"7E",X"00",X"FD",X"23",X"87",X"38",X"11",X"87",X"38",
		X"1A",X"87",X"38",X"2C",X"87",X"30",X"35",X"47",X"7B",X"E6",X"0F",X"B0",X"5F",X"18",X"D9",X"FD",
		X"56",X"00",X"FD",X"23",X"CD",X"76",X"3C",X"10",X"F6",X"18",X"D5",X"FD",X"56",X"00",X"FD",X"23",
		X"CD",X"76",X"3C",X"14",X"FD",X"CB",X"FE",X"6E",X"28",X"02",X"15",X"15",X"10",X"F2",X"18",X"C0",
		X"FD",X"56",X"00",X"FD",X"23",X"CD",X"76",X"3C",X"10",X"FB",X"18",X"B4",X"23",X"CD",X"79",X"3C",
		X"18",X"AE",X"DD",X"7E",X"FF",X"07",X"07",X"E6",X"03",X"3C",X"47",X"CB",X"5D",X"28",X"17",X"0E",
		X"5D",X"11",X"48",X"31",X"CD",X"A9",X"3C",X"11",X"19",X"0D",X"CD",X"A3",X"3C",X"11",X"85",X"FF",
		X"19",X"10",X"E8",X"C3",X"78",X"3B",X"0E",X"4D",X"11",X"19",X"0D",X"CD",X"A9",X"3C",X"11",X"48",
		X"31",X"CD",X"A3",X"3C",X"18",X"E7",X"72",X"23",X"73",X"23",X"0D",X"C0",X"21",X"2A",X"E0",X"35",
		X"28",X"1D",X"3A",X"29",X"E0",X"4F",X"2A",X"27",X"E0",X"C5",X"01",X"80",X"00",X"DD",X"CB",X"FF",
		X"6E",X"28",X"01",X"05",X"09",X"22",X"27",X"E0",X"C1",X"7C",X"D6",X"80",X"FE",X"0C",X"D8",X"E1",
		X"C3",X"78",X"3B",X"D5",X"11",X"7D",X"00",X"19",X"D1",X"72",X"23",X"71",X"23",X"73",X"23",X"71",
		X"C9",X"2A",X"0F",X"E7",X"3A",X"BA",X"E2",X"AE",X"E6",X"F0",X"20",X"29",X"7E",X"87",X"87",X"4F",
		X"87",X"5F",X"3A",X"68",X"E0",X"57",X"23",X"7E",X"23",X"22",X"0F",X"E7",X"3D",X"F8",X"FE",X"04",
		X"28",X"0D",X"30",X"16",X"4E",X"23",X"46",X"23",X"22",X"0F",X"E7",X"EB",X"C3",X"B7",X"2D",X"3E",
		X"03",X"32",X"88",X"E2",X"C9",X"AF",X"32",X"0B",X"E7",X"C9",X"D6",X"06",X"38",X"F3",X"20",X"0E",
		X"21",X"60",X"E3",X"7E",X"D6",X"1D",X"28",X"04",X"3D",X"C0",X"3E",X"9E",X"77",X"C9",X"D6",X"03",
		X"30",X"27",X"FD",X"21",X"60",X"E3",X"7E",X"32",X"6D",X"E0",X"E6",X"07",X"FD",X"77",X"0E",X"23",
		X"7E",X"23",X"22",X"0F",X"E7",X"FD",X"77",X"03",X"3A",X"08",X"E7",X"FE",X"02",X"D8",X"FD",X"73",
		X"0B",X"FD",X"72",X"0C",X"FD",X"36",X"00",X"1D",X"C9",X"46",X"23",X"22",X"0F",X"E7",X"FE",X"05",
		X"30",X"3A",X"87",X"21",X"68",X"00",X"85",X"6F",X"30",X"01",X"24",X"7E",X"23",X"66",X"6F",X"78",
		X"CD",X"DD",X"3E",X"4E",X"23",X"EB",X"E5",X"1A",X"13",X"FE",X"10",X"38",X"0C",X"28",X"06",X"77",
		X"23",X"71",X"23",X"18",X"F2",X"A9",X"4F",X"18",X"EE",X"D6",X"02",X"38",X"04",X"85",X"6F",X"18",
		X"E6",X"E1",X"3C",X"C8",X"D5",X"11",X"80",X"00",X"19",X"D1",X"18",X"DA",X"D6",X"16",X"F5",X"21",
		X"6C",X"E0",X"6E",X"2C",X"2D",X"28",X"11",X"E6",X"0F",X"FE",X"08",X"30",X"2B",X"FE",X"05",X"28",
		X"07",X"2D",X"2D",X"2D",X"2D",X"2D",X"28",X"20",X"EB",X"C5",X"FD",X"21",X"F0",X"E3",X"06",X"01",
		X"FE",X"05",X"28",X"0B",X"FD",X"21",X"D0",X"E4",X"11",X"F0",X"FF",X"06",X"0D",X"FD",X"19",X"FD",
		X"7E",X"00",X"A7",X"28",X"05",X"10",X"F6",X"F1",X"F1",X"C9",X"F1",X"FD",X"77",X"03",X"FD",X"75",
		X"0B",X"FD",X"74",X"0C",X"CD",X"DD",X"3E",X"F1",X"FE",X"05",X"CA",X"37",X"3E",X"0E",X"C2",X"FE",
		X"20",X"38",X"02",X"0E",X"D2",X"CB",X"67",X"28",X"01",X"0C",X"E6",X"0F",X"F5",X"F5",X"FD",X"36",
		X"00",X"22",X"21",X"BD",X"05",X"85",X"6F",X"30",X"01",X"24",X"F1",X"87",X"87",X"C6",X"1C",X"CB",
		X"61",X"28",X"02",X"C6",X"14",X"FD",X"77",X"0D",X"6E",X"EB",X"F1",X"51",X"FE",X"08",X"30",X"65",
		X"CB",X"62",X"28",X"04",X"01",X"80",X"01",X"09",X"01",X"04",X"03",X"FE",X"02",X"38",X"14",X"04",
		X"FE",X"03",X"20",X"0F",X"01",X"02",X"03",X"CD",X"13",X"3E",X"1C",X"23",X"23",X"05",X"CD",X"12",
		X"3E",X"1C",X"0C",X"C5",X"7C",X"D6",X"80",X"FE",X"0C",X"30",X"17",X"E5",X"73",X"1C",X"23",X"72",
		X"23",X"10",X"F9",X"E1",X"01",X"80",X"00",X"CB",X"62",X"28",X"01",X"05",X"09",X"C1",X"0D",X"20",
		X"E2",X"C9",X"1C",X"10",X"FD",X"18",X"ED",X"FD",X"36",X"00",X"23",X"FD",X"36",X"0D",X"50",X"01",
		X"03",X"04",X"EB",X"11",X"E4",X"CC",X"CD",X"13",X"3E",X"01",X"80",X"00",X"09",X"01",X"02",X"04",
		X"11",X"E4",X"DC",X"18",X"BE",X"D6",X"08",X"FD",X"77",X"0D",X"FD",X"75",X"08",X"FD",X"74",X"09",
		X"FE",X"05",X"30",X"18",X"C6",X"99",X"77",X"23",X"72",X"FE",X"9D",X"3E",X"00",X"CE",X"9E",X"5F",
		X"3E",X"7F",X"85",X"6F",X"30",X"01",X"24",X"73",X"23",X"72",X"18",X"0A",X"20",X"0D",X"01",X"02",
		X"02",X"1E",X"95",X"CD",X"13",X"3E",X"FD",X"36",X"00",X"25",X"C9",X"FE",X"07",X"20",X"22",X"0E",
		X"09",X"CD",X"CD",X"3E",X"11",X"6F",X"00",X"19",X"06",X"09",X"11",X"C4",X"3E",X"1A",X"77",X"2C",
		X"71",X"2C",X"13",X"10",X"F8",X"11",X"6E",X"00",X"19",X"CD",X"CD",X"3E",X"FD",X"36",X"00",X"28",
		X"C9",X"01",X"02",X"03",X"3E",X"79",X"11",X"7F",X"00",X"77",X"2C",X"36",X"02",X"3E",X"72",X"19",
		X"10",X"F7",X"18",X"C2",X"A5",X"EB",X"ED",X"EC",X"EB",X"EB",X"CC",X"CB",X"A3",X"06",X"08",X"3E",
		X"A5",X"77",X"2C",X"71",X"2C",X"10",X"FA",X"3E",X"A3",X"77",X"2C",X"71",X"C9",X"1F",X"1F",X"1F",
		X"37",X"1F",X"CB",X"19",X"E6",X"8F",X"57",X"59",X"C9",X"07",X"3F",X"4F",X"3F",X"6A",X"3F",X"4F",
		X"3F",X"B2",X"3F",X"1F",X"3F",X"58",X"3F",X"82",X"3F",X"58",X"3F",X"CA",X"3F",X"37",X"3F",X"61",
		X"3F",X"9A",X"3F",X"61",X"3F",X"E2",X"3F",X"0C",X"20",X"90",X"10",X"20",X"65",X"35",X"20",X"90",
		X"39",X"A0",X"98",X"3E",X"A0",X"AC",X"47",X"A0",X"9C",X"4D",X"50",X"A8",X"70",X"72",X"65",X"0C",
		X"20",X"AC",X"10",X"20",X"86",X"35",X"20",X"AC",X"39",X"A0",X"AC",X"3E",X"A0",X"CE",X"47",X"A0",
		X"BB",X"4D",X"50",X"C9",X"70",X"72",X"79",X"0C",X"20",X"D9",X"10",X"20",X"AB",X"35",X"20",X"D9",
		X"39",X"A0",X"D9",X"3E",X"A0",X"F6",X"47",X"A0",X"DF",X"4D",X"50",X"F0",X"70",X"72",X"90",X"30",
		X"24",X"65",X"4C",X"70",X"65",X"70",X"E2",X"80",X"30",X"24",X"8F",X"4C",X"70",X"8F",X"70",X"E2",
		X"A2",X"30",X"24",X"AB",X"4C",X"70",X"AB",X"70",X"E2",X"CE",X"0C",X"20",X"90",X"10",X"20",X"78",
		X"35",X"20",X"90",X"3D",X"A0",X"98",X"40",X"A0",X"AC",X"47",X"A0",X"9C",X"4D",X"50",X"A8",X"70",
		X"72",X"65",X"0C",X"20",X"AC",X"10",X"20",X"8F",X"35",X"20",X"AC",X"3D",X"A0",X"AC",X"40",X"A0",
		X"CE",X"47",X"A0",X"BB",X"4D",X"50",X"C9",X"70",X"72",X"79",X"0C",X"20",X"D9",X"10",X"20",X"C2",
		X"35",X"20",X"D9",X"3D",X"A0",X"D9",X"40",X"A0",X"F6",X"47",X"A0",X"DF",X"4D",X"50",X"F0",X"70",
		X"72",X"90",X"0C",X"20",X"98",X"10",X"20",X"88",X"35",X"20",X"98",X"37",X"A0",X"98",X"3C",X"A0",
		X"AC",X"46",X"A0",X"9C",X"4D",X"50",X"A8",X"70",X"72",X"65",X"0C",X"20",X"BE",X"10",X"20",X"AB",
		X"35",X"20",X"BE",X"37",X"A0",X"AC",X"3C",X"A0",X"CE",X"46",X"A0",X"BB",X"4D",X"50",X"C9",X"70",
		X"72",X"79",X"0C",X"20",X"E4",X"10",X"20",X"CE",X"35",X"20",X"E4",X"37",X"A0",X"D9",X"3C",X"A0",
		X"F6",X"46",X"A0",X"DF",X"4D",X"50",X"F0",X"70",X"72",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"5B",X"E0",X"FD",X"21",X"D0",X"E1",X"01",X"06",X"C2",X"16",X"E0",X"3A",X"04",X"D0",X"E6",
		X"20",X"20",X"04",X"16",X"F0",X"06",X"BA",X"CD",X"A3",X"40",X"CD",X"A3",X"40",X"0E",X"04",X"78",
		X"D6",X"10",X"47",X"D5",X"C5",X"3A",X"5B",X"E0",X"FE",X"60",X"DA",X"B6",X"40",X"CD",X"99",X"42",
		X"CD",X"71",X"44",X"0D",X"20",X"F7",X"CD",X"7E",X"44",X"C1",X"D1",X"7A",X"C6",X"06",X"57",X"C9",
		X"DD",X"7E",X"0D",X"6F",X"26",X"00",X"5F",X"54",X"29",X"29",X"19",X"11",X"F1",X"44",X"19",X"DD",
		X"7E",X"01",X"87",X"16",X"00",X"87",X"30",X"01",X"14",X"5F",X"FD",X"21",X"C0",X"E1",X"FD",X"19",
		X"3A",X"0D",X"E0",X"DD",X"86",X"03",X"86",X"C6",X"0F",X"2F",X"47",X"23",X"5E",X"7B",X"17",X"16",
		X"FF",X"38",X"01",X"14",X"E5",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"19",X"11",X"F9",X"FF",X"19",
		X"22",X"5B",X"E0",X"E1",X"23",X"7E",X"E6",X"0F",X"20",X"24",X"3A",X"06",X"E7",X"FE",X"03",X"38",
		X"02",X"3E",X"02",X"A7",X"28",X"02",X"C6",X"0A",X"86",X"EE",X"C0",X"5F",X"23",X"56",X"23",X"D5",
		X"5E",X"21",X"39",X"41",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"D1",X"AF",X"E9",X"FE",X"07",
		X"3E",X"00",X"20",X"E4",X"DD",X"7E",X"0C",X"18",X"DF",X"E1",X"41",X"FC",X"41",X"81",X"42",X"0C",
		X"42",X"A5",X"41",X"DA",X"41",X"06",X"43",X"1E",X"42",X"18",X"43",X"29",X"43",X"35",X"43",X"8F",
		X"43",X"42",X"43",X"6E",X"43",X"D0",X"41",X"27",X"44",X"32",X"44",X"89",X"42",X"75",X"42",X"38",
		X"44",X"EA",X"41",X"47",X"44",X"34",X"42",X"26",X"42",X"F4",X"41",X"40",X"42",X"63",X"42",X"97",
		X"41",X"5E",X"44",X"FE",X"1A",X"38",X"1C",X"16",X"0C",X"CD",X"C6",X"44",X"38",X"03",X"14",X"14",
		X"14",X"CD",X"EA",X"41",X"CD",X"7D",X"44",X"CD",X"D2",X"42",X"C3",X"89",X"42",X"D6",X"1A",X"FE",
		X"70",X"38",X"E4",X"16",X"06",X"18",X"5D",X"CD",X"D2",X"42",X"CD",X"E4",X"41",X"3E",X"10",X"CD",
		X"74",X"44",X"14",X"18",X"45",X"2A",X"D8",X"E2",X"7C",X"2D",X"28",X"C7",X"2D",X"28",X"DE",X"CD",
		X"C6",X"44",X"38",X"2D",X"21",X"04",X"E7",X"CB",X"46",X"20",X"0B",X"16",X"B0",X"CD",X"CF",X"42",
		X"CD",X"EA",X"41",X"14",X"18",X"21",X"16",X"D9",X"1F",X"38",X"16",X"CB",X"BB",X"05",X"18",X"11",
		X"3A",X"22",X"E0",X"E6",X"02",X"28",X"01",X"14",X"18",X"10",X"CD",X"C6",X"44",X"38",X"02",X"14",
		X"14",X"CD",X"CF",X"42",X"CD",X"EA",X"41",X"CD",X"7D",X"44",X"3A",X"5C",X"E0",X"A7",X"C2",X"D2",
		X"42",X"C3",X"99",X"42",X"CD",X"C6",X"44",X"38",X"03",X"14",X"14",X"14",X"CD",X"D2",X"42",X"CD",
		X"E4",X"41",X"3E",X"09",X"CD",X"80",X"44",X"CD",X"71",X"44",X"18",X"DE",X"48",X"CD",X"6E",X"42",
		X"41",X"EB",X"CD",X"7D",X"44",X"CD",X"C6",X"44",X"38",X"6F",X"14",X"14",X"18",X"6B",X"CD",X"CF",
		X"42",X"CD",X"D2",X"42",X"18",X"C4",X"DD",X"34",X"0F",X"DD",X"7E",X"0F",X"FE",X"10",X"30",X"0A",
		X"FE",X"0A",X"38",X"4D",X"CD",X"CF",X"42",X"C3",X"CF",X"42",X"DD",X"36",X"0F",X"00",X"18",X"41",
		X"CD",X"C6",X"44",X"38",X"3C",X"3A",X"04",X"E7",X"3D",X"28",X"14",X"48",X"CD",X"EA",X"41",X"CD",
		X"71",X"44",X"6A",X"16",X"BA",X"CD",X"EA",X"41",X"41",X"55",X"CD",X"7D",X"44",X"18",X"2A",X"16",
		X"DB",X"18",X"1E",X"CD",X"C6",X"44",X"38",X"19",X"14",X"14",X"14",X"14",X"18",X"13",X"62",X"7B",
		X"C6",X"80",X"6F",X"18",X"17",X"48",X"CD",X"6E",X"42",X"EB",X"CD",X"85",X"42",X"41",X"CD",X"7D",
		X"44",X"48",X"CD",X"89",X"42",X"CD",X"7D",X"44",X"41",X"62",X"6B",X"24",X"3A",X"5C",X"E0",X"A7",
		X"20",X"39",X"CD",X"99",X"42",X"CD",X"72",X"44",X"EB",X"FD",X"70",X"60",X"FD",X"73",X"61",X"FD",
		X"72",X"62",X"3A",X"5B",X"E0",X"D6",X"08",X"FD",X"77",X"63",X"FD",X"70",X"00",X"FD",X"73",X"01",
		X"FD",X"72",X"02",X"FD",X"77",X"03",X"FD",X"70",X"A0",X"FD",X"73",X"A1",X"FD",X"72",X"A2",X"FD",
		X"77",X"A3",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"C9",X"CD",X"72",X"44",X"EB",X"CD",
		X"D2",X"42",X"FD",X"36",X"62",X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"A2",X"00",X"FD",X"23",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"C9",X"78",X"FE",X"A0",X"30",X"0D",X"3A",X"5C",X"E0",X"A7",
		X"20",X"E8",X"3A",X"5B",X"E0",X"D6",X"08",X"18",X"BD",X"3A",X"5C",X"E0",X"A7",X"20",X"D7",X"3A",
		X"5B",X"E0",X"D6",X"08",X"18",X"A4",X"CD",X"D2",X"42",X"CD",X"6E",X"42",X"EB",X"CD",X"7D",X"44",
		X"3E",X"08",X"CD",X"74",X"44",X"C3",X"EA",X"41",X"CD",X"89",X"42",X"14",X"3E",X"F8",X"CD",X"80",
		X"44",X"3E",X"18",X"CD",X"74",X"44",X"C3",X"89",X"42",X"CD",X"D2",X"42",X"CD",X"89",X"42",X"CD",
		X"71",X"44",X"C3",X"EA",X"41",X"CD",X"EA",X"41",X"3E",X"10",X"CD",X"74",X"44",X"CD",X"7D",X"44",
		X"18",X"EA",X"3E",X"F9",X"CD",X"99",X"44",X"CD",X"EA",X"41",X"3E",X"F9",X"CD",X"80",X"44",X"CD",
		X"71",X"44",X"CD",X"EA",X"41",X"14",X"3E",X"FD",X"CD",X"80",X"44",X"3E",X"15",X"CD",X"74",X"44",
		X"CD",X"89",X"42",X"CD",X"7D",X"44",X"3E",X"13",X"CD",X"74",X"44",X"C3",X"89",X"42",X"3E",X"F8",
		X"CD",X"80",X"44",X"3E",X"03",X"CD",X"B9",X"44",X"3E",X"08",X"CD",X"80",X"44",X"CD",X"2C",X"43",
		X"15",X"15",X"CD",X"7E",X"44",X"3E",X"20",X"CD",X"74",X"44",X"CB",X"B3",X"C3",X"2C",X"43",X"3E",
		X"F8",X"CD",X"99",X"44",X"DD",X"CB",X"0B",X"66",X"20",X"02",X"16",X"01",X"3A",X"1D",X"E7",X"A7",
		X"28",X"0E",X"CD",X"81",X"42",X"41",X"CD",X"7D",X"44",X"7A",X"EE",X"00",X"67",X"C3",X"6F",X"42",
		X"78",X"FE",X"A0",X"38",X"3F",X"D6",X"10",X"47",X"CD",X"22",X"44",X"CD",X"22",X"44",X"7A",X"EE",
		X"00",X"67",X"6B",X"CB",X"BD",X"EB",X"3A",X"5C",X"E0",X"A7",X"20",X"17",X"78",X"C6",X"10",X"FD",
		X"77",X"00",X"FD",X"75",X"01",X"FD",X"74",X"02",X"3A",X"5B",X"E0",X"D6",X"08",X"FD",X"77",X"03",
		X"C3",X"B6",X"42",X"FD",X"36",X"02",X"00",X"C3",X"DA",X"42",X"62",X"6B",X"24",X"18",X"D6",X"62",
		X"6B",X"24",X"18",X"0F",X"48",X"CD",X"1C",X"44",X"CD",X"1C",X"44",X"7A",X"EE",X"00",X"67",X"7B",
		X"C6",X"80",X"6F",X"3A",X"5C",X"E0",X"A7",X"20",X"0C",X"CD",X"F2",X"42",X"CD",X"72",X"44",X"EB",
		X"CD",X"F2",X"42",X"18",X"5D",X"CD",X"DA",X"42",X"EB",X"C3",X"DA",X"42",X"CD",X"EF",X"43",X"41",
		X"18",X"03",X"CD",X"EA",X"43",X"18",X"56",X"48",X"CD",X"2C",X"43",X"41",X"CD",X"7D",X"44",X"C3",
		X"2C",X"43",X"48",X"CD",X"89",X"42",X"18",X"F3",X"CD",X"EA",X"41",X"3E",X"F6",X"CD",X"80",X"44",
		X"7A",X"EE",X"0F",X"57",X"C3",X"EA",X"41",X"78",X"06",X"07",X"FE",X"A0",X"38",X"0A",X"CD",X"56",
		X"44",X"11",X"50",X"00",X"FD",X"19",X"06",X"04",X"CD",X"DA",X"42",X"10",X"FB",X"C9",X"CD",X"81",
		X"42",X"CD",X"C6",X"44",X"D8",X"3E",X"24",X"FD",X"77",X"5A",X"FD",X"77",X"FA",X"FD",X"77",X"9A",
		X"C9",X"14",X"3E",X"F0",X"CB",X"7B",X"20",X"02",X"ED",X"44",X"80",X"47",X"C9",X"14",X"3E",X"F0",
		X"CB",X"73",X"20",X"02",X"ED",X"44",X"E5",X"2A",X"5B",X"E0",X"CB",X"7F",X"28",X"01",X"25",X"85",
		X"6F",X"30",X"01",X"24",X"22",X"5B",X"E0",X"E1",X"C9",X"CD",X"DD",X"44",X"C6",X"78",X"D5",X"57",
		X"CB",X"73",X"1E",X"C1",X"20",X"02",X"1E",X"01",X"3A",X"1D",X"E7",X"A7",X"28",X"06",X"CD",X"EA",
		X"41",X"D1",X"41",X"C9",X"CD",X"E7",X"42",X"18",X"F8",X"CD",X"DD",X"44",X"C6",X"82",X"D5",X"57",
		X"CD",X"EA",X"41",X"D1",X"41",X"C9",X"3A",X"1E",X"E7",X"A7",X"C8",X"21",X"D4",X"E2",X"35",X"F2",
		X"D9",X"44",X"2B",X"7E",X"23",X"77",X"23",X"34",X"2B",X"23",X"7E",X"1F",X"C9",X"48",X"CD",X"74",
		X"44",X"DD",X"7E",X"0E",X"D6",X"05",X"38",X"02",X"D6",X"05",X"3C",X"83",X"5F",X"DD",X"7E",X"0E",
		X"C9",X"FE",X"0F",X"80",X"B6",X"32",X"F8",X"0F",X"80",X"B3",X"02",X"F9",X"0F",X"00",X"B1",X"08",
		X"F9",X"0F",X"00",X"B3",X"02",X"F3",X"0F",X"00",X"B6",X"32",X"FB",X"0F",X"80",X"C2",X"34",X"F1",
		X"0F",X"80",X"BF",X"36",X"F9",X"0F",X"00",X"BB",X"0A",X"00",X"0F",X"00",X"BF",X"36",X"F6",X"0F",
		X"00",X"C2",X"34",X"F2",X"0F",X"80",X"D3",X"30",X"F4",X"0F",X"80",X"D0",X"02",X"F7",X"0F",X"00",
		X"CA",X"30",X"FD",X"0F",X"00",X"D0",X"02",X"FF",X"0F",X"00",X"D3",X"30",X"F9",X"0F",X"00",X"19",
		X"00",X"F7",X"0F",X"00",X"32",X"04",X"F0",X"0B",X"00",X"36",X"10",X"F6",X"0D",X"00",X"3A",X"12",
		X"F9",X"FE",X"C0",X"2E",X"04",X"FA",X"00",X"C0",X"32",X"04",X"01",X"FC",X"C0",X"36",X"10",X"FB",
		X"02",X"C0",X"3A",X"12",X"F8",X"12",X"00",X"2E",X"04",X"FA",X"0F",X"80",X"32",X"04",X"01",X"0B",
		X"80",X"36",X"10",X"FB",X"0D",X"80",X"3A",X"12",X"F8",X"FE",X"40",X"2E",X"04",X"F7",X"00",X"40",
		X"32",X"04",X"F0",X"FC",X"40",X"36",X"10",X"F6",X"02",X"40",X"3A",X"12",X"E9",X"12",X"80",X"2E",
		X"04",X"F8",X"0F",X"80",X"20",X"38",X"F1",X"0F",X"00",X"1B",X"06",X"F1",X"0F",X"00",X"1B",X"06",
		X"F1",X"0F",X"00",X"1B",X"06",X"F9",X"0F",X"00",X"20",X"38",X"F1",X"12",X"00",X"25",X"0C",X"F9",
		X"14",X"00",X"2C",X"00",X"F9",X"16",X"00",X"27",X"00",X"F9",X"08",X"00",X"29",X"0E",X"F9",X"0A",
		X"00",X"2A",X"0E",X"F9",X"0D",X"00",X"2B",X"0E",X"04",X"0F",X"00",X"3D",X"14",X"F8",X"0B",X"00",
		X"41",X"04",X"07",X"0B",X"00",X"45",X"14",X"F9",X"0D",X"00",X"49",X"04",X"ED",X"0F",X"80",X"3D",
		X"14",X"F9",X"0B",X"80",X"41",X"04",X"EA",X"0B",X"80",X"45",X"14",X"F8",X"0D",X"80",X"49",X"04",
		X"F9",X"0F",X"07",X"70",X"28",X"F9",X"0D",X"07",X"6F",X"28",X"F9",X"0C",X"07",X"6E",X"28",X"F9",
		X"0B",X"07",X"6D",X"28",X"F9",X"0A",X"07",X"6C",X"28",X"F5",X"08",X"07",X"6A",X"22",X"F1",X"15",
		X"07",X"66",X"04",X"EF",X"14",X"07",X"61",X"20",X"E9",X"0F",X"07",X"5B",X"1E",X"FC",X"08",X"87",
		X"6A",X"22",X"00",X"15",X"87",X"66",X"04",X"02",X"14",X"87",X"61",X"20",X"08",X"0F",X"87",X"5B",
		X"1E",X"FB",X"15",X"8A",X"52",X"18",X"F1",X"17",X"0A",X"4D",X"16",X"F5",X"15",X"0A",X"52",X"18",
		X"08",X"0F",X"8A",X"58",X"1A",X"F5",X"06",X"4A",X"52",X"18",X"F1",X"08",X"4A",X"4D",X"16",X"FB",
		X"06",X"CA",X"52",X"18",X"E9",X"0F",X"0A",X"58",X"1A",X"00",X"00",X"00",X"00",X"00",X"F1",X"1B",
		X"05",X"71",X"24",X"F9",X"07",X"0A",X"17",X"26",X"F9",X"07",X"0A",X"18",X"26",X"F9",X"07",X"0A",
		X"17",X"28",X"F9",X"07",X"0A",X"18",X"28",X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"2C",X"09",X"1F",X"00",X"97",X"2E",X"F8",X"0B",X"00",X"19",X"1C",X"F8",X"0B",X"80",X"19",X"1C",
		X"10",X"21",X"19",X"25",X"0D",X"1F",X"0C",X"18",X"11",X"1D",X"19",X"18",X"10",X"1F",X"0C",X"18",
		X"0C",X"1D",X"19",X"18",X"11",X"23",X"28",X"43",X"09",X"13",X"0F",X"11",X"FA",X"18",X"05",X"18",
		X"FB",X"18",X"08",X"1B",X"00",X"1D",X"04",X"1B",X"FF",X"19",X"04",X"13",X"02",X"1E",X"04",X"20",
		X"01",X"18",X"05",X"18",X"01",X"18",X"08",X"1B",X"02",X"1D",X"04",X"1B",X"FE",X"19",X"04",X"13",
		X"F9",X"1E",X"04",X"20",X"00",X"24",X"03",X"14",X"01",X"24",X"05",X"16",X"06",X"29",X"03",X"16",
		X"05",X"25",X"03",X"12",X"08",X"28",X"03",X"18",X"07",X"24",X"03",X"14",X"07",X"24",X"05",X"16",
		X"08",X"29",X"03",X"16",X"04",X"25",X"03",X"12",X"FF",X"2A",X"03",X"18",X"18",X"31",X"0D",X"1B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"65",X"19",X"23",X"F0",X"00",X"84",X"67",X"F8",X"AE",X"05",X"A0",X"02",X"B6",X"02",X"8D",X"00",
		X"23",X"68",X"A0",X"E2",X"02",X"CC",X"04",X"A0",X"00",X"00",X"40",X"82",X"86",X"02",X"EA",X"08",
		X"A0",X"00",X"00",X"10",X"66",X"AE",X"04",X"B0",X"B5",X"02",X"AC",X"00",X"00",X"22",X"90",X"B8",
		X"BD",X"08",X"C0",X"42",X"00",X"28",X"56",X"A4",X"02",X"EA",X"04",X"C0",X"00",X"00",X"20",X"72",
		X"9A",X"02",X"9F",X"08",X"E0",X"00",X"00",X"18",X"46",X"CC",X"05",X"E0",X"B8",X"00",X"00",X"00",
		X"33",X"CC",X"09",X"90",X"02",X"A5",X"00",X"00",X"37",X"90",X"AE",X"06",X"A0",X"04",X"C8",X"00",
		X"00",X"24",X"72",X"A9",X"02",X"9F",X"06",X"F0",X"58",X"20",X"4C",X"88",X"AE",X"06",X"B0",X"B5",
		X"02",X"8D",X"00",X"00",X"24",X"A0",X"9B",X"98",X"96",X"BB",X"97",X"96",X"BB",X"95",X"94",X"B6",
		X"9C",X"A8",X"84",X"8F",X"BB",X"BB",X"8C",X"B8",X"B1",X"B7",X"9D",X"A9",X"85",X"BB",X"8C",X"BB",
		X"8D",X"BB",X"AC",X"B2",X"9E",X"AA",X"89",X"86",X"8D",X"BB",X"8E",X"8F",X"AD",X"B3",X"9F",X"AB",
		X"8A",X"87",X"8E",X"BB",X"BB",X"BB",X"AE",X"B4",X"9A",X"A6",X"8B",X"88",X"BB",X"8C",X"BB",X"84",
		X"AC",X"B2",X"9B",X"A7",X"BB",X"BD",X"BB",X"8D",X"BB",X"85",X"AD",X"B3",X"9C",X"A8",X"8C",X"BB",
		X"BB",X"BB",X"BB",X"BD",X"AE",X"B4",X"9A",X"A6",X"BD",X"BB",X"BB",X"BB",X"8C",X"BA",X"AF",X"B5",
		X"9B",X"A7",X"BB",X"BB",X"8C",X"BB",X"8D",X"B9",X"B0",X"B6",X"9C",X"A8",X"BB",X"BB",X"8D",X"BB",
		X"BB",X"B8",X"B1",X"B7",X"9A",X"A6",X"BB",X"BB",X"BB",X"BB",X"BB",X"8C",X"AC",X"B2",X"9B",X"A7",
		X"89",X"86",X"BB",X"8C",X"BB",X"8D",X"AD",X"B3",X"9C",X"A8",X"8A",X"87",X"BB",X"8D",X"BB",X"BD",
		X"AE",X"B4",X"9D",X"A9",X"8B",X"88",X"BB",X"8E",X"BB",X"BA",X"AF",X"B5",X"9E",X"AA",X"BD",X"BB",
		X"8C",X"BB",X"84",X"B9",X"B0",X"B6",X"9F",X"AB",X"BB",X"BB",X"8D",X"BB",X"85",X"B8",X"B1",X"B7",
		X"9D",X"93",X"92",X"8F",X"91",X"92",X"BB",X"91",X"90",X"B2",X"80",X"81",X"82",X"80",X"81",X"82",
		X"80",X"81",X"82",X"83",X"7E",X"48",X"D6",X"48",X"2E",X"49",X"86",X"49",X"DE",X"49",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"04",X"05",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"07",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",
		X"0A",X"0A",X"0A",X"0B",X"0C",X"40",X"0D",X"0E",X"0F",X"45",X"47",X"42",X"12",X"40",X"49",X"0A",
		X"4B",X"4C",X"4D",X"0B",X"0D",X"0E",X"44",X"17",X"18",X"17",X"18",X"46",X"10",X"45",X"46",X"46",
		X"46",X"46",X"46",X"46",X"46",X"46",X"2E",X"25",X"24",X"29",X"26",X"2C",X"3C",X"30",X"20",X"2B",
		X"2F",X"30",X"29",X"2B",X"27",X"3E",X"25",X"29",X"24",X"26",X"2A",X"3C",X"23",X"20",X"21",X"2B",
		X"27",X"24",X"38",X"2C",X"31",X"32",X"22",X"3E",X"28",X"3C",X"32",X"2C",X"29",X"2E",X"27",X"2B",
		X"2B",X"21",X"2F",X"3D",X"30",X"21",X"2B",X"27",X"21",X"2B",X"2B",X"27",X"2B",X"2B",X"26",X"2C",
		X"36",X"33",X"27",X"2B",X"2B",X"26",X"2C",X"38",X"31",X"3B",X"28",X"35",X"33",X"34",X"2C",X"39",
		X"20",X"26",X"19",X"1A",X"1D",X"1C",X"1B",X"1C",X"1B",X"1A",X"1B",X"1A",X"1B",X"1A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"04",X"05",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"07",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"0A",
		X"0A",X"0A",X"0A",X"4B",X"4C",X"4C",X"4D",X"0B",X"0C",X"0D",X"0E",X"0F",X"45",X"47",X"12",X"40",
		X"13",X"14",X"15",X"40",X"0D",X"0E",X"44",X"17",X"18",X"17",X"18",X"46",X"10",X"45",X"46",X"46",
		X"46",X"46",X"46",X"46",X"46",X"46",X"2A",X"2C",X"31",X"30",X"2C",X"33",X"3A",X"22",X"31",X"38",
		X"2A",X"32",X"33",X"23",X"28",X"3D",X"28",X"33",X"31",X"32",X"28",X"3E",X"31",X"22",X"23",X"2A",
		X"23",X"3C",X"2A",X"32",X"3D",X"2C",X"32",X"33",X"3C",X"31",X"3A",X"23",X"2C",X"38",X"22",X"28",
		X"32",X"28",X"33",X"3E",X"23",X"2A",X"2C",X"28",X"33",X"31",X"28",X"28",X"33",X"33",X"31",X"28",
		X"39",X"22",X"33",X"2C",X"31",X"32",X"23",X"3D",X"22",X"36",X"28",X"39",X"31",X"3D",X"33",X"3B",
		X"2C",X"37",X"19",X"1C",X"1D",X"1C",X"1D",X"1C",X"1B",X"1A",X"1B",X"1A",X"1B",X"1A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"04",X"04",X"05",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"07",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"45",X"47",X"12",X"40",X"49",X"4B",X"4C",X"4D",
		X"0B",X"13",X"15",X"0D",X"43",X"17",X"18",X"17",X"18",X"17",X"18",X"46",X"10",X"45",X"46",X"46",
		X"46",X"46",X"46",X"46",X"46",X"46",X"E6",X"00",X"00",X"11",X"17",X"13",X"00",X"11",X"17",X"13",
		X"07",X"11",X"33",X"13",X"0E",X"11",X"E2",X"13",X"0E",X"11",X"E2",X"13",X"0E",X"11",X"E2",X"13",
		X"13",X"11",X"F7",X"13",X"18",X"11",X"59",X"14",X"18",X"11",X"59",X"14",X"18",X"11",X"59",X"14",
		X"18",X"11",X"59",X"14",X"06",X"11",X"70",X"14",X"06",X"11",X"D2",X"14",X"06",X"11",X"D2",X"14",
		X"06",X"11",X"E2",X"14",X"06",X"11",X"1E",X"15",X"21",X"11",X"97",X"15",X"21",X"11",X"97",X"15",
		X"21",X"11",X"AB",X"15",X"21",X"11",X"BE",X"15",X"1D",X"11",X"E9",X"15",X"1D",X"11",X"E9",X"15",
		X"26",X"11",X"35",X"16",X"2D",X"11",X"26",X"17",X"30",X"11",X"09",X"18",X"2B",X"11",X"09",X"18",
		X"35",X"11",X"28",X"18",X"3A",X"11",X"42",X"18",X"48",X"11",X"66",X"18",X"4F",X"11",X"66",X"18",
		X"66",X"11",X"87",X"18",X"6D",X"11",X"7D",X"18",X"8A",X"11",X"61",X"18",X"91",X"11",X"61",X"18",
		X"AC",X"11",X"82",X"18",X"B3",X"11",X"78",X"18",X"C4",X"11",X"44",X"18",X"D2",X"11",X"23",X"18",
		X"06",X"11",X"8F",X"19",X"06",X"11",X"43",X"19",X"D5",X"11",X"EC",X"17",X"D5",X"11",X"EC",X"17",
		X"DA",X"11",X"45",X"19",X"DD",X"11",X"8A",X"19",X"06",X"11",X"1C",X"15",X"06",X"11",X"E0",X"14",
		X"E0",X"11",X"02",X"1B",X"E7",X"11",X"CE",X"1A",X"EC",X"11",X"D3",X"1A",X"F3",X"11",X"04",X"1B",
		X"06",X"11",X"D7",X"1B",X"00",X"13",X"25",X"1C",X"F7",X"12",X"27",X"1C",X"06",X"11",X"33",X"1D",
		X"06",X"11",X"31",X"1D",X"00",X"13",X"25",X"1C",X"F7",X"12",X"E9",X"1D",X"06",X"11",X"A2",X"1D",
		X"06",X"11",X"A0",X"1D",X"00",X"13",X"E7",X"1D",X"09",X"13",X"61",X"1E",X"0E",X"13",X"61",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"12",X"77",X"1E",X"2F",X"12",X"EC",X"1E",
		X"14",X"12",X"98",X"1E",X"C9",X"12",X"7B",X"20",X"1D",X"12",X"B1",X"1E",X"56",X"12",X"57",X"1F",
		X"26",X"12",X"D0",X"1E",X"C4",X"12",X"63",X"20",X"2F",X"12",X"EC",X"1E",X"D4",X"12",X"97",X"20",
		X"3C",X"12",X"11",X"1F",X"0B",X"12",X"77",X"1E",X"3C",X"12",X"11",X"1F",X"D4",X"12",X"97",X"20",
		X"63",X"12",X"76",X"1F",X"14",X"12",X"98",X"1E",X"85",X"12",X"C3",X"1F",X"49",X"12",X"32",X"1F",
		X"B2",X"12",X"2C",X"20",X"A7",X"12",X"10",X"20",X"BD",X"12",X"4C",X"20",X"EC",X"12",X"D9",X"20",
		X"C9",X"12",X"7B",X"20",X"74",X"12",X"9C",X"1F",X"E1",X"12",X"B7",X"20",X"96",X"12",X"E9",X"1F",
		X"E1",X"12",X"B7",X"20",X"3C",X"12",X"11",X"1F",X"3C",X"12",X"11",X"1F",X"3C",X"12",X"11",X"1F",
		X"2F",X"12",X"EC",X"1E",X"1D",X"12",X"B1",X"1E",X"49",X"12",X"32",X"1F",X"D4",X"12",X"97",X"20",
		X"85",X"12",X"C3",X"1F",X"EC",X"12",X"D9",X"20",X"49",X"12",X"32",X"1F",X"56",X"12",X"57",X"1F",
		X"96",X"12",X"E9",X"1F",X"85",X"12",X"C3",X"1F",X"E1",X"12",X"B7",X"20",X"06",X"11",X"48",X"47",
		X"85",X"12",X"C3",X"1F",X"06",X"11",X"53",X"47",X"26",X"12",X"D0",X"1E",X"06",X"11",X"5C",X"47",
		X"26",X"12",X"D0",X"1E",X"06",X"11",X"65",X"47",X"1D",X"12",X"B1",X"1E",X"06",X"11",X"6F",X"47",
		X"96",X"12",X"E9",X"1F",X"06",X"11",X"77",X"47",X"C4",X"12",X"63",X"20",X"06",X"11",X"80",X"47",
		X"EC",X"12",X"D9",X"20",X"06",X"11",X"89",X"47",X"BD",X"12",X"4C",X"20",X"06",X"11",X"91",X"47",
		X"56",X"12",X"57",X"1F",X"06",X"11",X"9A",X"47",X"E1",X"12",X"B7",X"20",X"06",X"11",X"A3",X"47",
		X"49",X"12",X"32",X"1F",X"06",X"11",X"AC",X"47",X"2B",X"11",X"09",X"18",X"2B",X"11",X"09",X"18",
		X"35",X"11",X"28",X"18",X"41",X"11",X"42",X"18",X"58",X"11",X"66",X"18",X"5F",X"11",X"66",X"18",
		X"72",X"11",X"87",X"18",X"79",X"11",X"7D",X"18",X"80",X"11",X"87",X"18",X"85",X"11",X"7D",X"18",
		X"98",X"11",X"61",X"18",X"9D",X"11",X"61",X"18",X"A0",X"11",X"61",X"18",X"A5",X"11",X"61",X"18",
		X"BA",X"11",X"82",X"18",X"BF",X"11",X"78",X"18",X"CB",X"11",X"44",X"18",X"D2",X"11",X"23",X"18",
		X"05",X"12",X"24",X"17",X"08",X"12",X"33",X"16",X"21",X"11",X"BC",X"15",X"21",X"11",X"A9",X"15",
		X"26",X"11",X"13",X"16",X"FC",X"11",X"EC",X"16",X"FA",X"11",X"FC",X"17",X"FA",X"11",X"FC",X"17",
		X"FF",X"11",X"EA",X"16",X"02",X"12",X"11",X"16",X"00",X"00",X"B2",X"4C",X"00",X"00",X"62",X"4D",
		X"00",X"00",X"0F",X"1F",X"3F",X"5E",X"2F",X"0C",X"0A",X"0E",X"0F",X"0E",X"2E",X"1D",X"1B",X"39",
		X"4F",X"6E",X"0D",X"2B",X"09",X"2D",X"2F",X"1F",X"3F",X"5E",X"0F",X"0E",X"0F",X"2D",X"1F",X"2B",
		X"4B",X"69",X"0F",X"0E",X"2F",X"4E",X"2E",X"0B",X"09",X"0E",X"1D",X"2B",X"1B",X"39",X"1F",X"3F",
		X"5E",X"2B",X"09",X"07",X"0F",X"2D",X"1F",X"3E",X"2A",X"3E",X"5E",X"7C",X"2E",X"1D",X"2D",X"2C",
		X"1F",X"3D",X"5F",X"5D",X"3B",X"59",X"2D",X"1F",X"1F",X"39",X"19",X"07",X"2E",X"1D",X"0F",X"1E",
		X"3F",X"5F",X"2F",X"4E",X"2E",X"2B",X"09",X"2D",X"3E",X"5E",X"2C",X"8A",X"9A",X"BC",X"9F",X"9E",
		X"3E",X"5C",X"0A",X"28",X"4F",X"5E",X"3D",X"5B",X"69",X"8A",X"6F",X"8D",X"8F",X"5E",X"8F",X"AD",
		X"CF",X"CD",X"9F",X"9E",X"BE",X"CD",X"9D",X"9E",X"CD",X"7D",X"6A",X"08",X"04",X"24",X"03",X"2D",
		X"7F",X"BE",X"5E",X"7D",X"9F",X"7C",X"BD",X"6C",X"3C",X"35",X"27",X"6C",X"DD",X"DE",X"1D",X"2A",
		X"26",X"13",X"2E",X"5D",X"8D",X"BC",X"CE",X"9F",X"0F",X"02",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"1F",X"2C",X"29",X"1D",X"2D",X"4C",X"1C",X"5D",X"2C",X"1A",X"18",X"2D",X"4C",X"5A",
		X"5F",X"0D",X"2D",X"4C",X"6E",X"7C",X"1C",X"2C",X"1C",X"5D",X"1D",X"2D",X"3C",X"2A",X"2A",X"1A",
		X"07",X"24",X"4D",X"6F",X"1D",X"2C",X"2A",X"2C",X"4E",X"6D",X"2C",X"2A",X"4A",X"69",X"2D",X"2C",
		X"0A",X"0D",X"2F",X"4F",X"1E",X"2C",X"1C",X"2A",X"1B",X"39",X"1F",X"2C",X"1A",X"08",X"06",X"14",
		X"2E",X"1D",X"3F",X"5D",X"1B",X"2B",X"19",X"39",X"2D",X"2C",X"4C",X"5A",X"1C",X"2F",X"2E",X"3D",
		X"5F",X"7C",X"0F",X"0D",X"2D",X"1B",X"19",X"17",X"3D",X"5F",X"7D",X"2B",X"49",X"69",X"1A",X"2A",
		X"1A",X"3B",X"49",X"6D",X"3D",X"5D",X"7A",X"29",X"47",X"66",X"8D",X"7F",X"9D",X"6C",X"8D",X"7D",
		X"9D",X"8D",X"AD",X"8C",X"9D",X"7E",X"9C",X"BC",X"5C",X"5A",X"18",X"28",X"27",X"15",X"24",X"23",
		X"4A",X"8B",X"69",X"5B",X"2D",X"3C",X"5F",X"7D",X"9D",X"9E",X"BD",X"AF",X"BD",X"BC",X"8D",X"8C",
		X"AD",X"AC",X"9D",X"8B",X"49",X"35",X"59",X"7B",X"28",X"12",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CA",X"4E",X"8A",X"4F",X"5B",X"51",X"55",X"52",X"D5",X"54",X"FF",X"00",X"6C",X"24",X"58",X"78",
		X"0B",X"58",X"80",X"0B",X"58",X"D2",X"24",X"28",X"4A",X"24",X"70",X"AA",X"24",X"30",X"3A",X"24",
		X"28",X"DC",X"24",X"38",X"E0",X"24",X"38",X"30",X"24",X"68",X"5A",X"24",X"90",X"A7",X"24",X"38",
		X"4C",X"24",X"38",X"64",X"2F",X"10",X"6D",X"2E",X"10",X"A2",X"24",X"28",X"22",X"24",X"28",X"25",
		X"24",X"08",X"90",X"24",X"68",X"90",X"01",X"60",X"FF",X"98",X"0B",X"60",X"A0",X"0B",X"60",X"B0",
		X"2D",X"88",X"CA",X"25",X"60",X"DA",X"24",X"20",X"E8",X"0D",X"10",X"F0",X"0D",X"10",X"F8",X"0D",
		X"10",X"00",X"0D",X"10",X"24",X"24",X"90",X"28",X"0A",X"90",X"30",X"0A",X"90",X"38",X"0A",X"90",
		X"40",X"0A",X"90",X"68",X"0D",X"10",X"6C",X"24",X"08",X"70",X"0D",X"10",X"78",X"0D",X"10",X"80",
		X"0D",X"10",X"A8",X"0C",X"90",X"B0",X"0C",X"90",X"B4",X"24",X"90",X"B8",X"0C",X"90",X"C0",X"0C",
		X"90",X"EC",X"24",X"08",X"30",X"01",X"00",X"60",X"32",X"24",X"38",X"38",X"0B",X"40",X"40",X"0B",
		X"40",X"6C",X"24",X"68",X"90",X"01",X"60",X"FF",X"98",X"0B",X"60",X"A0",X"0B",X"60",X"B0",X"2D",
		X"88",X"B8",X"0D",X"10",X"C0",X"0D",X"10",X"E8",X"0A",X"90",X"F0",X"0A",X"90",X"F6",X"24",X"60",
		X"F8",X"0A",X"90",X"00",X"0A",X"90",X"FF",X"00",X"E0",X"00",X"30",X"50",X"20",X"32",X"39",X"10",
		X"60",X"31",X"80",X"62",X"3A",X"A0",X"DA",X"39",X"90",X"FB",X"50",X"28",X"FD",X"39",X"18",X"1C",
		X"34",X"80",X"28",X"31",X"78",X"2A",X"3A",X"98",X"60",X"3D",X"60",X"7C",X"33",X"20",X"7E",X"3A",
		X"10",X"AB",X"34",X"10",X"D8",X"32",X"88",X"FA",X"3B",X"98",X"FA",X"3A",X"20",X"12",X"34",X"80",
		X"31",X"33",X"80",X"33",X"3A",X"A0",X"3C",X"32",X"18",X"40",X"34",X"58",X"6B",X"30",X"78",X"6D",
		X"39",X"98",X"91",X"32",X"88",X"BA",X"38",X"90",X"E2",X"33",X"20",X"E4",X"3D",X"10",X"14",X"31",
		X"68",X"18",X"33",X"68",X"48",X"34",X"18",X"55",X"33",X"10",X"60",X"33",X"80",X"62",X"3A",X"A0",
		X"9A",X"3B",X"28",X"C0",X"34",X"30",X"0A",X"3D",X"70",X"0C",X"32",X"20",X"0E",X"39",X"10",X"12",
		X"32",X"20",X"14",X"39",X"10",X"3A",X"39",X"20",X"3A",X"3B",X"88",X"7A",X"38",X"90",X"94",X"32",
		X"68",X"96",X"38",X"88",X"CC",X"34",X"88",X"F0",X"50",X"20",X"F2",X"3A",X"10",X"16",X"50",X"18",
		X"48",X"31",X"78",X"4A",X"3D",X"98",X"60",X"34",X"40",X"78",X"33",X"20",X"7A",X"39",X"10",X"9A",
		X"30",X"90",X"A0",X"32",X"80",X"DC",X"51",X"40",X"F9",X"33",X"20",X"FB",X"38",X"10",X"1C",X"30",
		X"70",X"1C",X"3D",X"90",X"1E",X"3D",X"90",X"24",X"34",X"88",X"30",X"05",X"38",X"33",X"20",X"3C",
		X"33",X"20",X"50",X"05",X"58",X"51",X"20",X"5A",X"39",X"10",X"60",X"33",X"78",X"62",X"39",X"98",
		X"76",X"50",X"38",X"78",X"38",X"28",X"80",X"09",X"23",X"88",X"98",X"33",X"38",X"9A",X"39",X"28",
		X"A0",X"33",X"38",X"B0",X"30",X"18",X"BC",X"31",X"58",X"CA",X"34",X"18",X"D6",X"33",X"40",X"DA",
		X"33",X"38",X"DC",X"3A",X"28",X"E6",X"30",X"58",X"F0",X"33",X"18",X"F4",X"30",X"58",X"04",X"31",
		X"40",X"08",X"32",X"28",X"0A",X"39",X"18",X"18",X"32",X"40",X"28",X"31",X"50",X"38",X"32",X"58",
		X"3C",X"32",X"58",X"5A",X"3A",X"10",X"60",X"34",X"38",X"6C",X"32",X"58",X"6E",X"39",X"48",X"70",
		X"32",X"28",X"7C",X"32",X"30",X"80",X"51",X"28",X"90",X"33",X"70",X"94",X"33",X"70",X"96",X"39",
		X"90",X"AB",X"33",X"50",X"B0",X"33",X"50",X"B4",X"33",X"50",X"B8",X"33",X"50",X"BC",X"34",X"68",
		X"C7",X"31",X"78",X"C9",X"3D",X"98",X"CA",X"50",X"48",X"CB",X"3A",X"68",X"D8",X"3D",X"60",X"F2",
		X"32",X"18",X"F4",X"38",X"38",X"F4",X"51",X"48",X"FA",X"31",X"50",X"FC",X"50",X"20",X"FC",X"39",
		X"40",X"14",X"32",X"30",X"16",X"39",X"20",X"27",X"32",X"40",X"3A",X"3B",X"28",X"48",X"32",X"50",
		X"4C",X"32",X"50",X"5C",X"32",X"38",X"5C",X"3D",X"18",X"5E",X"3D",X"18",X"60",X"3D",X"18",X"84",
		X"32",X"60",X"8A",X"32",X"60",X"8B",X"38",X"80",X"90",X"34",X"78",X"9C",X"32",X"30",X"9C",X"32",
		X"90",X"9E",X"3A",X"20",X"BA",X"38",X"40",X"DC",X"32",X"80",X"EC",X"32",X"78",X"FA",X"38",X"68",
		X"FA",X"3C",X"A0",X"1C",X"32",X"20",X"1E",X"3D",X"10",X"3A",X"39",X"20",X"40",X"30",X"58",X"44",
		X"51",X"20",X"46",X"3A",X"10",X"50",X"33",X"40",X"62",X"34",X"70",X"70",X"30",X"70",X"72",X"3D",
		X"90",X"74",X"3D",X"90",X"78",X"51",X"40",X"00",X"00",X"FF",X"00",X"FF",X"00",X"72",X"24",X"58",
		X"78",X"0B",X"58",X"80",X"0B",X"58",X"CA",X"24",X"18",X"42",X"24",X"20",X"92",X"24",X"68",X"DA",
		X"24",X"08",X"2A",X"24",X"40",X"DA",X"24",X"88",X"40",X"24",X"38",X"44",X"24",X"38",X"62",X"24",
		X"90",X"BA",X"24",X"38",X"22",X"24",X"18",X"30",X"2F",X"68",X"39",X"2E",X"68",X"D2",X"24",X"38",
		X"02",X"24",X"28",X"05",X"24",X"08",X"30",X"24",X"38",X"90",X"01",X"00",X"60",X"94",X"24",X"68",
		X"98",X"0B",X"40",X"A0",X"0B",X"40",X"B0",X"2D",X"30",X"C2",X"24",X"80",X"02",X"24",X"68",X"10",
		X"01",X"60",X"FF",X"18",X"0B",X"60",X"20",X"0B",X"60",X"30",X"2D",X"88",X"48",X"0D",X"10",X"4A",
		X"25",X"60",X"50",X"0D",X"10",X"54",X"24",X"08",X"58",X"0D",X"10",X"60",X"0D",X"10",X"88",X"0A",
		X"90",X"90",X"0A",X"90",X"98",X"0A",X"90",X"9A",X"24",X"68",X"A0",X"0A",X"90",X"C8",X"0D",X"10",
		X"D0",X"0D",X"10",X"D8",X"0D",X"10",X"DC",X"24",X"08",X"E0",X"0D",X"10",X"F8",X"0C",X"90",X"00",
		X"0C",X"90",X"28",X"0D",X"10",X"28",X"0A",X"90",X"30",X"0D",X"10",X"30",X"0A",X"90",X"34",X"24",
		X"08",X"38",X"01",X"00",X"60",X"38",X"0D",X"10",X"38",X"0A",X"90",X"40",X"0D",X"10",X"40",X"0A",
		X"90",X"42",X"25",X"60",X"56",X"2D",X"20",X"68",X"0D",X"10",X"68",X"0A",X"90",X"70",X"0D",X"10",
		X"70",X"0A",X"90",X"78",X"01",X"60",X"FF",X"78",X"0D",X"10",X"78",X"0A",X"90",X"7A",X"24",X"70",
		X"80",X"0D",X"10",X"80",X"0A",X"90",X"A8",X"0D",X"10",X"B0",X"0D",X"10",X"B8",X"0D",X"10",X"BC",
		X"24",X"08",X"C0",X"0D",X"10",X"E8",X"0A",X"90",X"F0",X"0A",X"90",X"F8",X"0A",X"90",X"00",X"0A",
		X"90",X"FF",X"00",X"E0",X"00",X"2C",X"31",X"78",X"2E",X"39",X"98",X"5B",X"50",X"18",X"6A",X"32",
		X"90",X"75",X"32",X"20",X"76",X"39",X"10",X"A0",X"31",X"70",X"A2",X"3A",X"90",X"B4",X"34",X"50",
		X"DA",X"38",X"18",X"EB",X"32",X"20",X"ED",X"39",X"10",X"20",X"32",X"28",X"22",X"39",X"18",X"3A",
		X"3B",X"28",X"4A",X"32",X"90",X"60",X"3D",X"50",X"64",X"34",X"50",X"6C",X"31",X"90",X"7C",X"50",
		X"20",X"7E",X"39",X"10",X"83",X"32",X"98",X"A4",X"52",X"10",X"B4",X"30",X"80",X"B6",X"39",X"A0",
		X"BB",X"52",X"08",X"CC",X"34",X"80",X"D7",X"31",X"80",X"1C",X"51",X"28",X"1C",X"51",X"28",X"1E",
		X"39",X"18",X"28",X"34",X"40",X"40",X"31",X"80",X"58",X"34",X"30",X"74",X"32",X"28",X"76",X"38",
		X"18",X"98",X"30",X"80",X"9A",X"3A",X"A0",X"BA",X"39",X"20",X"BA",X"3B",X"88",X"C6",X"34",X"68",
		X"DC",X"34",X"30",X"FC",X"52",X"78",X"FE",X"3A",X"98",X"1A",X"32",X"18",X"1C",X"3A",X"08",X"24",
		X"34",X"68",X"56",X"52",X"80",X"58",X"3D",X"A0",X"5B",X"32",X"08",X"7A",X"38",X"90",X"A8",X"31",
		X"80",X"AA",X"3A",X"A0",X"F4",X"34",X"50",X"18",X"50",X"20",X"18",X"50",X"20",X"1A",X"39",X"10",
		X"2C",X"31",X"88",X"45",X"52",X"78",X"47",X"39",X"98",X"5A",X"39",X"90",X"68",X"34",X"78",X"88",
		X"52",X"00",X"9A",X"3A",X"18",X"AA",X"3D",X"60",X"AC",X"32",X"90",X"BB",X"52",X"08",X"D8",X"34",
		X"48",X"FA",X"3B",X"28",X"30",X"05",X"33",X"34",X"48",X"3B",X"30",X"88",X"50",X"05",X"55",X"31",
		X"68",X"57",X"38",X"88",X"80",X"09",X"43",X"60",X"8A",X"51",X"30",X"8C",X"38",X"20",X"BA",X"39",
		X"20",X"BA",X"3B",X"88",X"D8",X"34",X"58",X"DC",X"52",X"08",X"EB",X"3D",X"A0",X"FC",X"52",X"10",
		X"0C",X"31",X"78",X"0E",X"39",X"98",X"14",X"34",X"70",X"1A",X"32",X"28",X"1A",X"3D",X"18",X"1C",
		X"3D",X"18",X"30",X"05",X"3B",X"32",X"98",X"41",X"32",X"30",X"45",X"32",X"30",X"4A",X"32",X"28",
		X"4C",X"3A",X"18",X"4C",X"30",X"80",X"50",X"05",X"53",X"31",X"78",X"6A",X"30",X"68",X"6C",X"39",
		X"88",X"70",X"31",X"60",X"7C",X"51",X"28",X"7E",X"3C",X"18",X"80",X"09",X"63",X"80",X"85",X"50",
		X"38",X"87",X"39",X"28",X"91",X"51",X"20",X"A2",X"50",X"40",X"A4",X"38",X"30",X"B0",X"34",X"60",
		X"B2",X"50",X"28",X"B6",X"52",X"20",X"CC",X"51",X"38",X"CE",X"39",X"28",X"DA",X"50",X"20",X"E1",
		X"34",X"58",X"EB",X"52",X"10",X"EC",X"32",X"40",X"ED",X"39",X"30",X"F8",X"51",X"38",X"FA",X"38",
		X"28",X"0C",X"51",X"48",X"10",X"50",X"38",X"12",X"38",X"28",X"1B",X"34",X"80",X"1C",X"32",X"30",
		X"1E",X"3A",X"20",X"2C",X"50",X"40",X"34",X"51",X"30",X"36",X"38",X"20",X"3C",X"50",X"28",X"3E",
		X"39",X"18",X"42",X"32",X"90",X"48",X"52",X"40",X"48",X"3D",X"30",X"5A",X"39",X"20",X"69",X"32",
		X"20",X"6B",X"38",X"10",X"75",X"50",X"20",X"77",X"39",X"10",X"80",X"50",X"70",X"81",X"3A",X"90",
		X"82",X"34",X"90",X"A8",X"52",X"70",X"AC",X"31",X"70",X"AE",X"39",X"90",X"B1",X"52",X"68",X"B6",
		X"52",X"60",X"BB",X"52",X"58",X"C0",X"52",X"50",X"D0",X"50",X"48",X"E0",X"34",X"88",X"EA",X"51",
		X"80",X"EC",X"3C",X"A0",X"F0",X"05",X"F1",X"32",X"30",X"F5",X"50",X"38",X"F9",X"51",X"38",X"FB",
		X"3D",X"28",X"FC",X"52",X"08",X"0B",X"50",X"28",X"0C",X"52",X"78",X"0D",X"38",X"18",X"0D",X"39",
		X"98",X"10",X"05",X"18",X"32",X"20",X"1C",X"32",X"20",X"1C",X"34",X"90",X"1D",X"38",X"10",X"2B",
		X"52",X"08",X"40",X"09",X"70",X"80",X"54",X"50",X"30",X"56",X"34",X"58",X"5A",X"3D",X"18",X"5B",
		X"51",X"28",X"5C",X"3D",X"18",X"5E",X"3D",X"18",X"68",X"32",X"40",X"6C",X"32",X"30",X"7A",X"3C",
		X"10",X"8C",X"51",X"20",X"8C",X"30",X"50",X"95",X"50",X"48",X"99",X"34",X"18",X"A0",X"50",X"50",
		X"A9",X"32",X"30",X"BA",X"3A",X"20",X"C4",X"50",X"38",X"C6",X"39",X"28",X"CC",X"51",X"30",X"CE",
		X"38",X"20",X"D2",X"34",X"50",X"DC",X"32",X"30",X"DE",X"3D",X"20",X"E9",X"51",X"10",X"EB",X"32",
		X"48",X"00",X"32",X"40",X"05",X"34",X"40",X"10",X"51",X"38",X"14",X"50",X"38",X"16",X"38",X"28",
		X"1B",X"51",X"30",X"1D",X"39",X"20",X"47",X"52",X"78",X"50",X"34",X"18",X"53",X"30",X"88",X"54",
		X"51",X"30",X"54",X"3D",X"20",X"56",X"3D",X"20",X"64",X"32",X"08",X"64",X"52",X"70",X"7A",X"3A",
		X"90",X"60",X"00",X"50",X"00",X"FF",X"00",X"72",X"24",X"58",X"78",X"0B",X"58",X"80",X"0B",X"58",
		X"80",X"24",X"88",X"0C",X"24",X"98",X"22",X"24",X"20",X"72",X"24",X"68",X"BA",X"24",X"08",X"EC",
		X"24",X"40",X"52",X"24",X"68",X"DA",X"24",X"98",X"02",X"24",X"90",X"02",X"24",X"90",X"1C",X"24",
		X"38",X"23",X"24",X"38",X"42",X"24",X"90",X"9A",X"24",X"38",X"E2",X"24",X"18",X"45",X"24",X"40",
		X"46",X"2F",X"68",X"4F",X"2E",X"68",X"E2",X"24",X"28",X"E5",X"24",X"08",X"1A",X"24",X"38",X"5A",
		X"24",X"68",X"90",X"01",X"60",X"FF",X"95",X"24",X"38",X"98",X"0B",X"60",X"A0",X"0B",X"60",X"AE",
		X"2D",X"80",X"C8",X"0D",X"10",X"CA",X"25",X"60",X"D0",X"0D",X"10",X"D8",X"0D",X"10",X"E0",X"0D",
		X"10",X"E0",X"24",X"38",X"08",X"0A",X"90",X"10",X"0A",X"90",X"18",X"0A",X"90",X"1C",X"24",X"90",
		X"20",X"0A",X"90",X"48",X"0D",X"10",X"50",X"0D",X"10",X"58",X"0D",X"10",X"5C",X"24",X"08",X"60",
		X"0D",X"10",X"78",X"24",X"60",X"78",X"0C",X"90",X"80",X"0C",X"90",X"B2",X"24",X"20",X"C0",X"24",
		X"38",X"D0",X"01",X"00",X"60",X"D8",X"0B",X"40",X"E0",X"0B",X"40",X"E0",X"24",X"68",X"EE",X"2D",
		X"30",X"F4",X"24",X"68",X"1A",X"24",X"98",X"30",X"01",X"60",X"FF",X"38",X"0B",X"60",X"40",X"0B",
		X"60",X"40",X"24",X"38",X"50",X"02",X"00",X"60",X"58",X"0D",X"10",X"5C",X"24",X"08",X"60",X"0D",
		X"10",X"62",X"25",X"60",X"76",X"2D",X"20",X"76",X"01",X"60",X"FF",X"78",X"0A",X"90",X"7C",X"24",
		X"60",X"80",X"0A",X"90",X"98",X"0D",X"10",X"9C",X"24",X"08",X"A0",X"0D",X"10",X"A0",X"24",X"38",
		X"B8",X"0A",X"90",X"BC",X"24",X"90",X"C0",X"0A",X"90",X"B0",X"00",X"A0",X"00",X"06",X"DF",X"70",
		X"DE",X"84",X"DF",X"A2",X"DD",X"B8",X"DF",X"28",X"DD",X"40",X"DF",X"50",X"DE",X"80",X"DF",X"10",
		X"DD",X"20",X"DF",X"70",X"DE",X"84",X"DF",X"A0",X"DD",X"B0",X"DF",X"C0",X"DD",X"D6",X"DF",X"F0",
		X"DE",X"10",X"DF",X"98",X"DD",X"B0",X"DF",X"A0",X"DF",X"90",X"DF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"81",X"00",X"41",X"20",X"2D",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",
		X"20",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"21",X"1C",X"E0",X"36",X"04",X"FB",
		X"CD",X"77",X"5E",X"C3",X"C3",X"56",X"0A",X"0A",X"0E",X"0E",X"14",X"0B",X"0B",X"10",X"10",X"18",
		X"0D",X"0D",X"13",X"13",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"D9",X"CD",X"8A",X"5B",X"3A",X"FF",X"E0",X"A7",X"F2",X"D9",X"56",X"CD",X"5E",X"57",X"01",
		X"03",X"00",X"10",X"FE",X"0D",X"20",X"FB",X"D9",X"08",X"FB",X"C9",X"CD",X"03",X"5C",X"CD",X"EA",
		X"5C",X"CD",X"77",X"5E",X"CD",X"D7",X"5E",X"3E",X"68",X"32",X"26",X"E7",X"3E",X"04",X"32",X"05",
		X"E7",X"32",X"2A",X"E7",X"32",X"1D",X"E7",X"32",X"1E",X"E7",X"C3",X"17",X"5F",X"AF",X"21",X"1C",
		X"E0",X"77",X"FB",X"CD",X"54",X"5D",X"CD",X"5C",X"6C",X"CD",X"02",X"5B",X"CD",X"F7",X"5B",X"CD",
		X"D7",X"5E",X"C3",X"17",X"5F",X"00",X"00",X"00",X"00",X"CD",X"DA",X"5B",X"3A",X"00",X"D0",X"2F",
		X"32",X"26",X"E0",X"CB",X"4F",X"28",X"15",X"3A",X"04",X"D0",X"CB",X"67",X"20",X"0E",X"21",X"1C",
		X"E0",X"CB",X"4E",X"20",X"07",X"3A",X"00",X"D0",X"E6",X"01",X"20",X"F9",X"CD",X"5E",X"57",X"FD",
		X"E5",X"DD",X"E5",X"CD",X"2C",X"5A",X"CD",X"E7",X"6C",X"CD",X"B9",X"5A",X"3A",X"12",X"E0",X"A7",
		X"20",X"05",X"3E",X"02",X"32",X"1E",X"E0",X"21",X"1C",X"E0",X"46",X"CB",X"78",X"20",X"15",X"CB",
		X"48",X"20",X"1F",X"3A",X"1E",X"E0",X"A7",X"20",X"21",X"CB",X"50",X"20",X"15",X"3A",X"1D",X"E0",
		X"A7",X"C2",X"5A",X"56",X"CB",X"40",X"28",X"0A",X"CD",X"00",X"21",X"CD",X"0F",X"62",X"21",X"B5",
		X"E2",X"34",X"DD",X"E1",X"FD",X"E1",X"D9",X"08",X"FB",X"C9",X"36",X"02",X"31",X"00",X"E8",X"FB",
		X"CD",X"77",X"5E",X"CD",X"1C",X"5B",X"28",X"FB",X"CD",X"CE",X"5E",X"C3",X"17",X"5F",X"21",X"22",
		X"E0",X"34",X"20",X"16",X"E5",X"2A",X"76",X"E0",X"23",X"22",X"76",X"E0",X"3A",X"1C",X"E0",X"87",
		X"30",X"07",X"2A",X"74",X"E0",X"23",X"22",X"74",X"E0",X"E1",X"7E",X"23",X"E6",X"0F",X"20",X"01",
		X"34",X"23",X"35",X"23",X"35",X"C9",X"3A",X"F0",X"E3",X"FE",X"26",X"C8",X"ED",X"5B",X"17",X"E0",
		X"2A",X"05",X"E7",X"7D",X"B4",X"20",X"07",X"CB",X"72",X"28",X"03",X"11",X"80",X"02",X"CB",X"B2",
		X"CD",X"AD",X"61",X"3A",X"F0",X"E3",X"FE",X"26",X"C8",X"31",X"00",X"E8",X"21",X"1C",X"E0",X"35",
		X"FB",X"F2",X"A4",X"56",X"CD",X"D9",X"63",X"21",X"1C",X"E0",X"CB",X"66",X"28",X"0C",X"CD",X"27",
		X"5C",X"3A",X"03",X"E7",X"A7",X"28",X"06",X"CD",X"27",X"5C",X"C3",X"17",X"5F",X"3A",X"04",X"D0",
		X"CB",X"4F",X"3E",X"C0",X"28",X"02",X"3E",X"78",X"CD",X"F9",X"5B",X"C3",X"17",X"5F",X"31",X"00",
		X"E8",X"21",X"1C",X"E0",X"35",X"FB",X"CD",X"D9",X"63",X"CD",X"F3",X"5B",X"01",X"00",X"0C",X"CD",
		X"7A",X"5E",X"3E",X"01",X"32",X"03",X"E7",X"3E",X"1B",X"CD",X"B6",X"5E",X"21",X"1C",X"E0",X"CB",
		X"66",X"28",X"28",X"21",X"AD",X"58",X"CD",X"92",X"59",X"3A",X"1C",X"E0",X"1F",X"1F",X"1F",X"E6",
		X"01",X"3C",X"11",X"80",X"FF",X"FD",X"19",X"CD",X"0C",X"5A",X"CD",X"F3",X"5B",X"CD",X"C5",X"6A",
		X"CD",X"27",X"5C",X"3A",X"03",X"E7",X"A7",X"28",X"A4",X"18",X"0C",X"21",X"C3",X"58",X"CD",X"92",
		X"59",X"CD",X"F3",X"5B",X"CD",X"C5",X"6A",X"3A",X"1B",X"E0",X"1F",X"30",X"55",X"CD",X"42",X"5C",
		X"28",X"03",X"CD",X"27",X"5C",X"CD",X"F3",X"5B",X"CD",X"77",X"5E",X"21",X"D0",X"58",X"CD",X"8A",
		X"59",X"3E",X"11",X"A7",X"28",X"3C",X"3D",X"27",X"32",X"27",X"E0",X"FD",X"21",X"24",X"89",X"CD",
		X"00",X"5A",X"3E",X"40",X"32",X"24",X"E0",X"3A",X"24",X"E0",X"A7",X"3A",X"27",X"E0",X"28",X"E3",
		X"3A",X"1E",X"E0",X"A7",X"20",X"0B",X"21",X"F1",X"58",X"CD",X"A5",X"59",X"CD",X"02",X"5B",X"18",
		X"E6",X"CD",X"1C",X"5B",X"28",X"E1",X"CD",X"9A",X"58",X"CD",X"9A",X"58",X"CD",X"77",X"5E",X"C3",
		X"17",X"5F",X"F3",X"AF",X"32",X"1C",X"E0",X"C3",X"A4",X"56",X"21",X"00",X"00",X"22",X"00",X"E7",
		X"22",X"02",X"E7",X"7C",X"32",X"2B",X"E7",X"CD",X"F5",X"5E",X"C3",X"27",X"5C",X"A4",X"81",X"00",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"20",X"21",X"A4",X"83",X"00",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"21",
		X"32",X"84",X"00",X"54",X"4F",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"45",X"20",X"47",
		X"41",X"4D",X"45",X"20",X"22",X"A4",X"86",X"00",X"54",X"49",X"4D",X"45",X"20",X"20",X"20",X"20",
		X"21",X"A8",X"84",X"00",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",X"4F",X"49",X"4E",X"20",
		X"20",X"21",X"CD",X"12",X"38",X"CD",X"BD",X"60",X"21",X"51",X"E0",X"3A",X"22",X"E0",X"46",X"77",
		X"A8",X"28",X"1F",X"CB",X"67",X"20",X"0F",X"CB",X"5F",X"20",X"11",X"CD",X"DC",X"2C",X"CD",X"FD",
		X"60",X"CD",X"36",X"61",X"18",X"0C",X"CD",X"DB",X"63",X"CD",X"96",X"61",X"CD",X"EC",X"2C",X"CD",
		X"FF",X"63",X"3A",X"82",X"E2",X"21",X"83",X"E2",X"BE",X"28",X"C7",X"5F",X"16",X"E6",X"DD",X"21",
		X"00",X"00",X"DD",X"19",X"DD",X"4E",X"00",X"CB",X"21",X"20",X"13",X"21",X"82",X"E2",X"BE",X"20",
		X"05",X"C6",X"04",X"E6",X"7F",X"77",X"DD",X"E5",X"C1",X"79",X"C6",X"04",X"18",X"D7",X"06",X"00",
		X"DD",X"70",X"00",X"DD",X"7E",X"01",X"21",X"56",X"59",X"E5",X"21",X"86",X"59",X"09",X"4E",X"23",
		X"66",X"69",X"E9",X"21",X"83",X"E2",X"6E",X"26",X"E6",X"71",X"23",X"77",X"23",X"73",X"23",X"72",
		X"2C",X"7D",X"E6",X"7F",X"32",X"83",X"E2",X"C9",X"48",X"5C",X"CD",X"DC",X"59",X"CD",X"CA",X"59",
		X"18",X"FB",X"CD",X"DC",X"59",X"CD",X"CA",X"59",X"3E",X"05",X"32",X"24",X"E0",X"3A",X"24",X"E0",
		X"A7",X"20",X"FA",X"18",X"F0",X"3A",X"22",X"E0",X"CB",X"67",X"20",X"DE",X"CD",X"DC",X"59",X"7E",
		X"23",X"FE",X"21",X"C8",X"FE",X"23",X"28",X"0F",X"FE",X"22",X"28",X"F0",X"FD",X"36",X"00",X"00",
		X"11",X"80",X"00",X"FD",X"19",X"18",X"E8",X"23",X"18",X"E5",X"7E",X"23",X"FE",X"21",X"28",X"19",
		X"FE",X"23",X"28",X"12",X"FE",X"25",X"28",X"13",X"FE",X"22",X"20",X"17",X"5E",X"23",X"56",X"23",
		X"FD",X"21",X"00",X"00",X"FD",X"19",X"4E",X"23",X"C9",X"E1",X"C9",X"46",X"23",X"CD",X"F3",X"59",
		X"10",X"FB",X"C9",X"FD",X"77",X"00",X"FD",X"71",X"01",X"11",X"80",X"00",X"FD",X"19",X"C9",X"7E",
		X"F5",X"11",X"80",X"00",X"1F",X"1F",X"1F",X"1F",X"CD",X"0C",X"5A",X"F1",X"E6",X"0F",X"C6",X"30",
		X"FD",X"77",X"00",X"FD",X"19",X"C9",X"7E",X"F5",X"1F",X"1F",X"1F",X"1F",X"CD",X"20",X"5A",X"F1",
		X"11",X"80",X"00",X"10",X"E7",X"E6",X"0F",X"20",X"E3",X"04",X"18",X"E4",X"21",X"10",X"E0",X"11",
		X"12",X"E0",X"3A",X"00",X"D0",X"CD",X"5C",X"5A",X"21",X"11",X"E0",X"13",X"3A",X"02",X"D0",X"1F",
		X"F6",X"04",X"CD",X"5C",X"5A",X"21",X"0E",X"E0",X"01",X"02",X"00",X"CD",X"B1",X"5A",X"23",X"0E",
		X"20",X"CD",X"B1",X"5A",X"3A",X"21",X"E0",X"B0",X"32",X"01",X"D0",X"C9",X"1F",X"1F",X"1F",X"CB",
		X"16",X"1F",X"CB",X"16",X"7E",X"E6",X"55",X"FE",X"50",X"28",X"0E",X"7E",X"E6",X"AA",X"C0",X"21",
		X"56",X"E0",X"34",X"7E",X"E6",X"0F",X"C0",X"18",X"28",X"2B",X"2B",X"36",X"0C",X"3E",X"13",X"CD",
		X"BE",X"5E",X"21",X"72",X"E0",X"7E",X"C6",X"01",X"27",X"77",X"23",X"7E",X"CE",X"00",X"27",X"77",
		X"1A",X"FE",X"01",X"28",X"11",X"FE",X"08",X"30",X"0B",X"21",X"1D",X"E0",X"34",X"BE",X"C0",X"AF",
		X"77",X"3C",X"18",X"02",X"D6",X"08",X"21",X"1E",X"E0",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",
		X"C9",X"7E",X"A7",X"C8",X"35",X"78",X"B1",X"47",X"C9",X"3A",X"1C",X"E0",X"07",X"30",X"20",X"11",
		X"01",X"D0",X"CB",X"67",X"28",X"07",X"3A",X"14",X"E0",X"3D",X"28",X"01",X"13",X"21",X"1F",X"E0",
		X"1A",X"2F",X"47",X"E6",X"03",X"77",X"78",X"07",X"07",X"07",X"E6",X"05",X"23",X"77",X"C9",X"11",
		X"70",X"E0",X"3A",X"2A",X"E7",X"A7",X"3E",X"DF",X"20",X"15",X"2A",X"0B",X"E3",X"29",X"29",X"29",
		X"29",X"29",X"7C",X"2A",X"6E",X"E0",X"BE",X"20",X"D4",X"23",X"7E",X"23",X"22",X"6E",X"E0",X"12",
		X"18",X"CB",X"21",X"12",X"5B",X"CD",X"8A",X"59",X"FD",X"21",X"82",X"8D",X"3A",X"1E",X"E0",X"C3",
		X"00",X"5A",X"02",X"8A",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"21",X"21",X"56",X"5B",X"CD",
		X"A5",X"59",X"CD",X"02",X"5B",X"21",X"67",X"5B",X"3A",X"1E",X"E0",X"3D",X"28",X"03",X"21",X"78",
		X"5B",X"CD",X"8A",X"59",X"3A",X"26",X"E0",X"E6",X"03",X"C8",X"1F",X"3A",X"1E",X"E0",X"06",X"80",
		X"38",X"06",X"D6",X"01",X"27",X"C8",X"06",X"90",X"D6",X"01",X"27",X"F3",X"32",X"1E",X"E0",X"78",
		X"32",X"1C",X"E0",X"3C",X"FB",X"C9",X"A8",X"84",X"00",X"20",X"50",X"55",X"53",X"48",X"20",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"20",X"21",X"A0",X"84",X"00",X"4F",X"4E",X"4C",X"59",X"20",X"31",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"21",X"A0",X"84",X"00",X"31",X"20",X"4F",X"52",X"20",
		X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"21",X"21",X"6B",X"E0",X"7E",X"FE",X"04",
		X"30",X"0D",X"34",X"21",X"00",X"E1",X"11",X"A0",X"C9",X"01",X"60",X"00",X"ED",X"B0",X"C9",X"21",
		X"60",X"E1",X"11",X"C0",X"C8",X"01",X"40",X"00",X"ED",X"B0",X"0E",X"20",X"11",X"A0",X"C8",X"ED",
		X"B0",X"11",X"40",X"C9",X"01",X"40",X"00",X"ED",X"B0",X"0E",X"20",X"1E",X"20",X"ED",X"B0",X"11",
		X"40",X"C8",X"0E",X"40",X"ED",X"B0",X"0E",X"20",X"1E",X"20",X"ED",X"B0",X"2A",X"80",X"E2",X"7D",
		X"32",X"00",X"90",X"7C",X"32",X"00",X"A0",X"C9",X"18",X"C5",X"2A",X"84",X"E2",X"7D",X"BC",X"C8",
		X"26",X"E0",X"7E",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"7D",X"3C",X"E6",X"07",X"32",
		X"84",X"E2",X"C9",X"3E",X"40",X"18",X"02",X"3E",X"C0",X"32",X"24",X"E0",X"3A",X"24",X"E0",X"A7",
		X"20",X"FA",X"C9",X"21",X"00",X"E0",X"01",X"80",X"07",X"CD",X"1E",X"5C",X"21",X"65",X"03",X"22",
		X"09",X"E0",X"21",X"9C",X"6C",X"11",X"7C",X"E0",X"01",X"4B",X"00",X"ED",X"B0",X"C9",X"36",X"00",
		X"23",X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"21",X"1C",X"E0",X"7E",X"EE",X"08",X"77",X"21",X"00",
		X"E7",X"11",X"2C",X"E7",X"01",X"2C",X"00",X"41",X"1A",X"4F",X"7E",X"12",X"71",X"23",X"13",X"10",
		X"F7",X"C9",X"3A",X"1C",X"E0",X"CB",X"5F",X"C9",X"4F",X"87",X"87",X"81",X"4F",X"06",X"00",X"3A",
		X"F0",X"E3",X"FE",X"26",X"C8",X"21",X"C2",X"5C",X"09",X"5E",X"23",X"56",X"23",X"E5",X"2A",X"07",
		X"E7",X"19",X"22",X"07",X"E7",X"E1",X"3A",X"1C",X"E0",X"A7",X"F0",X"11",X"00",X"E7",X"06",X"03",
		X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"ED",X"5B",X"01",X"E7",X"2A",X"09",X"E0",X"A7",
		X"ED",X"52",X"38",X"0B",X"20",X"16",X"21",X"08",X"E0",X"3A",X"00",X"E7",X"96",X"38",X"0D",X"3A",
		X"00",X"E7",X"32",X"08",X"E0",X"ED",X"53",X"09",X"E0",X"CD",X"B9",X"5C",X"FD",X"21",X"B6",X"8C",
		X"CD",X"42",X"5C",X"28",X"04",X"FD",X"21",X"B2",X"8C",X"21",X"02",X"E7",X"06",X"01",X"CD",X"16",
		X"5A",X"2B",X"CD",X"16",X"5A",X"2B",X"C3",X"FF",X"59",X"21",X"0A",X"E0",X"FD",X"21",X"BA",X"8C",
		X"18",X"EA",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"02",X"00",X"05",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"01",X"00",X"01",X"00",X"3A",X"03",X"D0",X"2F",X"47",X"E6",
		X"03",X"6F",X"87",X"85",X"C6",X"0A",X"2E",X"00",X"CB",X"3F",X"CB",X"1D",X"CB",X"3F",X"CB",X"1D",
		X"00",X"00",X"00",X"67",X"22",X"17",X"E0",X"78",X"1F",X"1F",X"21",X"A1",X"64",X"CB",X"47",X"28",
		X"03",X"21",X"66",X"56",X"22",X"19",X"E0",X"1F",X"32",X"1B",X"E0",X"1F",X"21",X"04",X"D0",X"CB",
		X"56",X"21",X"12",X"E0",X"28",X"1E",X"3C",X"E6",X"0F",X"CB",X"5F",X"28",X"01",X"3C",X"77",X"23",
		X"77",X"3A",X"04",X"D0",X"2F",X"47",X"CD",X"3C",X"5D",X"CD",X"3C",X"5D",X"78",X"1F",X"47",X"E6",
		X"01",X"23",X"77",X"C9",X"47",X"3C",X"E6",X"03",X"77",X"78",X"1F",X"1F",X"E6",X"03",X"FE",X"02",
		X"DE",X"F5",X"18",X"DB",X"CD",X"98",X"5F",X"21",X"00",X"80",X"01",X"00",X"0C",X"CD",X"1E",X"5C",
		X"21",X"24",X"5E",X"CD",X"8A",X"59",X"CD",X"02",X"5B",X"21",X"15",X"5E",X"CD",X"92",X"59",X"11",
		X"27",X"E0",X"01",X"20",X"00",X"3A",X"15",X"E0",X"A7",X"20",X"34",X"CD",X"B7",X"5D",X"CD",X"00",
		X"5E",X"7E",X"FE",X"32",X"20",X"20",X"3E",X"53",X"32",X"32",X"E0",X"32",X"3B",X"E0",X"21",X"35",
		X"E0",X"7E",X"87",X"D6",X"30",X"FE",X"3A",X"38",X"06",X"D6",X"0A",X"77",X"2B",X"3E",X"31",X"77",
		X"21",X"27",X"E0",X"CD",X"92",X"59",X"3A",X"1D",X"E0",X"A7",X"20",X"FA",X"C3",X"F7",X"5B",X"CD",
		X"EB",X"5D",X"CD",X"F5",X"5D",X"18",X"E9",X"21",X"38",X"5E",X"ED",X"B0",X"21",X"2A",X"E0",X"3A",
		X"12",X"E0",X"11",X"08",X"00",X"FE",X"08",X"38",X"12",X"C6",X"28",X"77",X"19",X"36",X"53",X"23",
		X"23",X"23",X"36",X"31",X"11",X"06",X"00",X"19",X"36",X"00",X"C9",X"3D",X"C8",X"11",X"0B",X"00",
		X"19",X"C6",X"31",X"77",X"11",X"06",X"00",X"19",X"36",X"53",X"C9",X"21",X"40",X"56",X"ED",X"B0",
		X"21",X"2E",X"E0",X"18",X"CA",X"CD",X"00",X"5E",X"21",X"2E",X"E0",X"3A",X"13",X"E0",X"18",X"C2",
		X"21",X"27",X"E0",X"CD",X"92",X"59",X"2A",X"27",X"E0",X"11",X"FC",X"FF",X"19",X"22",X"27",X"E0",
		X"21",X"2A",X"E0",X"34",X"C9",X"A8",X"83",X"00",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",
		X"4F",X"49",X"4E",X"21",X"1A",X"83",X"01",X"5D",X"31",X"39",X"38",X"33",X"20",X"49",X"52",X"45",
		X"4D",X"20",X"43",X"4F",X"52",X"50",X"2E",X"21",X"22",X"82",X"00",X"31",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"20",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0C",X"21",X"00",X"80",X"7D",X"E6",X"01",X"77",X"2C",
		X"20",X"F9",X"24",X"10",X"F6",X"18",X"09",X"01",X"00",X"10",X"21",X"00",X"80",X"CD",X"1E",X"5C",
		X"21",X"00",X"E1",X"01",X"82",X"01",X"CD",X"1E",X"5C",X"3A",X"14",X"E0",X"3D",X"28",X"09",X"21",
		X"1C",X"E0",X"AF",X"CB",X"5E",X"28",X"01",X"3C",X"32",X"21",X"E0",X"21",X"04",X"D0",X"AE",X"21",
		X"0D",X"E0",X"36",X"00",X"1F",X"30",X"02",X"36",X"00",X"F3",X"AF",X"CD",X"BE",X"5E",X"FB",X"C9",
		X"F3",X"CD",X"B6",X"5E",X"FB",X"C9",X"E5",X"21",X"1C",X"E0",X"CB",X"7E",X"E1",X"F0",X"E5",X"2A",
		X"85",X"E2",X"26",X"E0",X"77",X"7D",X"3C",X"E6",X"07",X"32",X"85",X"E2",X"E1",X"C9",X"CD",X"E3",
		X"5E",X"CD",X"77",X"5E",X"C3",X"55",X"6A",X"CD",X"FC",X"5E",X"21",X"CD",X"55",X"22",X"6E",X"E0",
		X"C3",X"77",X"5E",X"CD",X"E6",X"5E",X"CD",X"27",X"5C",X"21",X"00",X"E7",X"01",X"2C",X"00",X"CD",
		X"1E",X"5C",X"CD",X"00",X"2E",X"21",X"00",X"1E",X"22",X"07",X"E7",X"C9",X"21",X"03",X"E7",X"01",
		X"29",X"00",X"18",X"EB",X"CD",X"89",X"5E",X"CD",X"36",X"5F",X"AF",X"CD",X"B0",X"5E",X"CD",X"18",
		X"64",X"CD",X"00",X"36",X"C3",X"98",X"5F",X"CD",X"04",X"5F",X"21",X"1C",X"E0",X"34",X"CD",X"C1",
		X"64",X"3E",X"0F",X"00",X"00",X"00",X"3A",X"04",X"E7",X"A7",X"28",X"02",X"C6",X"07",X"C6",X"18",
		X"CD",X"B0",X"5E",X"C3",X"02",X"59",X"21",X"00",X"E1",X"01",X"00",X"06",X"CD",X"1E",X"5C",X"DD",
		X"21",X"00",X"E3",X"DD",X"36",X"03",X"60",X"DD",X"36",X"06",X"30",X"11",X"10",X"00",X"3E",X"04",
		X"DD",X"19",X"DD",X"77",X"01",X"3C",X"FE",X"18",X"38",X"F6",X"21",X"05",X"E7",X"7E",X"E6",X"01",
		X"2B",X"77",X"3A",X"1D",X"E7",X"A7",X"28",X"29",X"3A",X"12",X"E7",X"32",X"11",X"E7",X"3A",X"0D",
		X"E7",X"32",X"0C",X"E7",X"2A",X"25",X"E7",X"2E",X"30",X"22",X"0B",X"E3",X"7C",X"32",X"25",X"E7",
		X"FE",X"54",X"3E",X"02",X"38",X"07",X"3E",X"02",X"32",X"04",X"E7",X"3E",X"0E",X"32",X"00",X"E3",
		X"C9",X"CD",X"DD",X"2D",X"26",X"00",X"18",X"DF",X"21",X"06",X"60",X"CD",X"8A",X"59",X"3A",X"16",
		X"E0",X"A7",X"20",X"06",X"21",X"9D",X"60",X"CD",X"8A",X"59",X"CD",X"36",X"61",X"CD",X"E4",X"61",
		X"06",X"00",X"CD",X"CD",X"60",X"CD",X"FD",X"60",X"CD",X"99",X"5C",X"3A",X"1C",X"E0",X"CB",X"67",
		X"28",X"0F",X"CD",X"27",X"5C",X"CD",X"9C",X"5C",X"CD",X"27",X"5C",X"21",X"A3",X"60",X"CD",X"8A",
		X"59",X"21",X"93",X"8C",X"01",X"06",X"0F",X"CD",X"00",X"60",X"21",X"13",X"8D",X"06",X"08",X"CD",
		X"00",X"60",X"21",X"26",X"8D",X"01",X"01",X"04",X"11",X"AA",X"60",X"CD",X"F7",X"5F",X"01",X"0B",
		X"0F",X"21",X"12",X"8E",X"11",X"AE",X"60",X"1A",X"77",X"2C",X"71",X"2C",X"13",X"10",X"F8",X"C9",
		X"71",X"2C",X"2C",X"10",X"FB",X"C9",X"3C",X"8C",X"01",X"48",X"49",X"2D",X"53",X"43",X"4F",X"52",
		X"45",X"22",X"BA",X"8C",X"04",X"20",X"20",X"20",X"20",X"30",X"30",X"22",X"38",X"8C",X"01",X"31",
		X"55",X"50",X"22",X"B6",X"8C",X"06",X"20",X"20",X"20",X"20",X"30",X"30",X"22",X"B2",X"8C",X"06",
		X"20",X"20",X"20",X"20",X"20",X"20",X"22",X"0E",X"8C",X"01",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0C",X"22",X"0C",X"8C",X"01",X"0D",X"52",X"41",X"4E",X"4B",X"20",X"16",X"22",X"0A",X"8C",X"04",
		X"0D",X"20",X"20",X"20",X"20",X"20",X"16",X"22",X"08",X"8C",X"01",X"17",X"18",X"18",X"18",X"18",
		X"18",X"19",X"22",X"86",X"8C",X"01",X"53",X"50",X"45",X"45",X"44",X"22",X"84",X"8C",X"00",X"20",
		X"20",X"20",X"22",X"04",X"8E",X"01",X"5B",X"5C",X"22",X"12",X"8F",X"01",X"60",X"61",X"22",X"18",
		X"8F",X"01",X"62",X"63",X"22",X"1E",X"8F",X"01",X"64",X"65",X"22",X"24",X"8F",X"01",X"66",X"67",
		X"22",X"2A",X"8F",X"01",X"68",X"69",X"22",X"2E",X"8F",X"01",X"6A",X"6B",X"21",X"04",X"8E",X"01",
		X"5E",X"5F",X"21",X"34",X"8C",X"01",X"32",X"55",X"50",X"21",X"4C",X"45",X"55",X"46",X"71",X"6D",
		X"6D",X"70",X"6F",X"6F",X"6E",X"6D",X"6D",X"70",X"6F",X"6F",X"6E",X"6D",X"6C",X"21",X"B5",X"E2",
		X"7E",X"FE",X"1D",X"D8",X"36",X"00",X"2A",X"21",X"E7",X"23",X"22",X"21",X"E7",X"3A",X"05",X"E7",
		X"87",X"87",X"87",X"4F",X"87",X"81",X"11",X"8A",X"04",X"2A",X"0B",X"E3",X"0E",X"FF",X"0C",X"ED",
		X"52",X"30",X"FB",X"81",X"21",X"92",X"8D",X"06",X"0F",X"D6",X"08",X"38",X"07",X"36",X"28",X"2C",
		X"2C",X"10",X"F6",X"C9",X"C6",X"28",X"77",X"AF",X"2C",X"2C",X"10",X"FA",X"C9",X"FD",X"21",X"84",
		X"8C",X"2A",X"08",X"E3",X"06",X"00",X"3A",X"16",X"E0",X"A7",X"28",X"19",X"11",X"BC",X"02",X"CD",
		X"1A",X"61",X"11",X"46",X"00",X"CD",X"1A",X"61",X"1E",X"07",X"AF",X"ED",X"52",X"3C",X"30",X"FB",
		X"19",X"3D",X"C3",X"20",X"5A",X"11",X"D4",X"03",X"CD",X"1A",X"61",X"11",X"62",X"00",X"CD",X"1A",
		X"61",X"11",X"0A",X"00",X"18",X"E4",X"01",X"00",X"05",X"3A",X"04",X"E7",X"FE",X"02",X"28",X"30",
		X"11",X"10",X"00",X"FD",X"21",X"50",X"E4",X"3A",X"1D",X"E7",X"A7",X"28",X"09",X"11",X"70",X"00",
		X"06",X"02",X"FD",X"21",X"10",X"E3",X"D5",X"FD",X"7E",X"00",X"A7",X"28",X"0E",X"FD",X"5E",X"0B",
		X"FD",X"56",X"0C",X"2A",X"0B",X"E3",X"ED",X"52",X"30",X"01",X"0C",X"D1",X"FD",X"19",X"10",X"E6",
		X"21",X"0C",X"E7",X"7E",X"81",X"27",X"30",X"02",X"3E",X"99",X"23",X"77",X"FD",X"21",X"0A",X"8D",
		X"CD",X"27",X"6C",X"7E",X"23",X"BE",X"D0",X"7E",X"D6",X"01",X"27",X"77",X"3E",X"02",X"CD",X"48",
		X"5C",X"3E",X"11",X"C3",X"B0",X"5E",X"3A",X"22",X"E0",X"E6",X"10",X"28",X"0C",X"3A",X"08",X"E7",
		X"FE",X"02",X"30",X"05",X"3E",X"12",X"CD",X"B0",X"5E",X"ED",X"5B",X"62",X"E0",X"2A",X"07",X"E7",
		X"A7",X"ED",X"52",X"30",X"32",X"21",X"00",X"00",X"22",X"07",X"E7",X"CD",X"E4",X"61",X"3A",X"04",
		X"D0",X"CB",X"77",X"C8",X"21",X"F0",X"E3",X"7E",X"FE",X"26",X"28",X"07",X"3E",X"C0",X"32",X"FF",
		X"E3",X"36",X"26",X"21",X"00",X"E3",X"7E",X"FE",X"03",X"28",X"03",X"FE",X"0F",X"C0",X"C6",X"07",
		X"77",X"C3",X"29",X"23",X"2A",X"07",X"E7",X"7C",X"FE",X"1E",X"38",X"03",X"21",X"00",X"1E",X"22",
		X"07",X"E7",X"29",X"29",X"7C",X"21",X"92",X"8C",X"06",X"0F",X"D6",X"08",X"38",X"07",X"36",X"09",
		X"2C",X"2C",X"10",X"F6",X"C9",X"C6",X"09",X"77",X"2C",X"2C",X"3E",X"01",X"10",X"F9",X"C9",X"3A",
		X"04",X"E7",X"FE",X"02",X"30",X"39",X"2A",X"0B",X"E3",X"01",X"D0",X"FF",X"09",X"22",X"80",X"E2",
		X"3A",X"0C",X"E3",X"FE",X"54",X"D8",X"3A",X"00",X"E3",X"FE",X"04",X"D0",X"3E",X"54",X"32",X"26",
		X"E7",X"21",X"1C",X"E0",X"35",X"31",X"00",X"E8",X"FB",X"2A",X"04",X"E3",X"E5",X"2A",X"08",X"E3",
		X"E5",X"CD",X"04",X"5F",X"E1",X"22",X"08",X"E3",X"E1",X"22",X"04",X"E3",X"C3",X"1A",X"5F",X"3A",
		X"00",X"E3",X"FE",X"0F",X"C0",X"CD",X"72",X"63",X"3A",X"0C",X"E3",X"D6",X"6D",X"30",X"2E",X"C6",
		X"02",X"38",X"30",X"3A",X"08",X"E7",X"A7",X"C8",X"21",X"22",X"E0",X"CB",X"46",X"C8",X"21",X"64",
		X"E0",X"35",X"F0",X"3A",X"2A",X"E7",X"A7",X"C0",X"FD",X"21",X"10",X"E3",X"FD",X"7E",X"00",X"A7",
		X"28",X"76",X"FD",X"21",X"C0",X"E3",X"FD",X"7E",X"00",X"A7",X"28",X"6C",X"C9",X"3E",X"10",X"32",
		X"00",X"E3",X"C9",X"3D",X"C0",X"3A",X"2A",X"E7",X"A7",X"C0",X"FD",X"21",X"70",X"E3",X"FD",X"7E",
		X"00",X"A7",X"C0",X"3A",X"05",X"E7",X"87",X"D6",X"02",X"D8",X"6F",X"26",X"00",X"11",X"51",X"63",
		X"19",X"5E",X"23",X"56",X"EB",X"FD",X"E5",X"D1",X"13",X"13",X"AF",X"06",X"0E",X"12",X"13",X"10",
		X"FC",X"7E",X"FD",X"77",X"03",X"23",X"11",X"00",X"02",X"C6",X"20",X"87",X"30",X"03",X"11",X"00",
		X"FE",X"FD",X"73",X"04",X"FD",X"72",X"05",X"7E",X"FD",X"77",X"06",X"23",X"7E",X"FD",X"77",X"0C",
		X"3A",X"05",X"E7",X"87",X"D6",X"02",X"FD",X"77",X"0E",X"FD",X"36",X"00",X"27",X"11",X"10",X"00",
		X"FD",X"19",X"23",X"7E",X"A7",X"20",X"BE",X"C9",X"FD",X"36",X"03",X"60",X"FD",X"36",X"06",X"A8",
		X"FD",X"36",X"07",X"00",X"3A",X"03",X"E3",X"06",X"03",X"D6",X"30",X"38",X"02",X"10",X"FA",X"ED",
		X"5F",X"4F",X"E6",X"03",X"23",X"23",X"BE",X"C8",X"77",X"0F",X"38",X"0C",X"87",X"80",X"3D",X"FE",
		X"04",X"38",X"04",X"EE",X"02",X"E6",X"03",X"47",X"78",X"EE",X"03",X"D6",X"02",X"FD",X"77",X"0E",
		X"2B",X"79",X"E6",X"0F",X"4F",X"E5",X"2A",X"08",X"E3",X"29",X"7C",X"29",X"84",X"D6",X"40",X"2F",
		X"81",X"E1",X"86",X"2B",X"77",X"FD",X"36",X"00",X"1C",X"ED",X"5F",X"E6",X"03",X"FD",X"77",X"0C",
		X"C9",X"59",X"63",X"63",X"63",X"6A",X"63",X"6E",X"63",X"EF",X"F0",X"80",X"F7",X"E0",X"88",X"FF",
		X"D0",X"90",X"00",X"C8",X"E0",X"40",X"D0",X"D0",X"48",X"00",X"FF",X"D8",X"70",X"00",X"FF",X"D0",
		X"90",X"00",X"3A",X"0C",X"E3",X"FE",X"54",X"28",X"09",X"FE",X"56",X"C0",X"21",X"9E",X"63",X"C3",
		X"AC",X"59",X"3A",X"05",X"E7",X"87",X"21",X"94",X"63",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"C3",X"8A",X"59",X"9E",X"63",X"AB",X"63",X"B6",X"63",X"C2",X"63",X"CD",X"63",X"04",X"84",
		X"02",X"4C",X"41",X"53",X"20",X"56",X"45",X"47",X"41",X"53",X"21",X"84",X"84",X"02",X"48",X"4F",
		X"55",X"53",X"54",X"4F",X"4E",X"21",X"04",X"84",X"02",X"53",X"54",X"2E",X"4C",X"4F",X"55",X"49",
		X"53",X"21",X"84",X"84",X"02",X"43",X"48",X"49",X"43",X"41",X"47",X"4F",X"21",X"04",X"84",X"02",
		X"4E",X"45",X"57",X"20",X"59",X"4F",X"52",X"4B",X"21",X"3E",X"FF",X"47",X"3A",X"1C",X"E0",X"21",
		X"F1",X"63",X"CB",X"5F",X"28",X"03",X"21",X"F8",X"63",X"CB",X"68",X"CA",X"AC",X"59",X"C3",X"8A",
		X"59",X"38",X"8C",X"01",X"31",X"55",X"50",X"21",X"34",X"8C",X"01",X"32",X"55",X"50",X"21",X"2A",
		X"08",X"E3",X"11",X"72",X"00",X"06",X"0C",X"ED",X"52",X"38",X"02",X"10",X"FA",X"78",X"C6",X"04",
		X"32",X"D3",X"E2",X"C6",X"1F",X"C9",X"00",X"00",X"2A",X"05",X"E7",X"7D",X"24",X"25",X"28",X"07",
		X"C6",X"05",X"25",X"28",X"02",X"C6",X"05",X"5F",X"16",X"00",X"2A",X"19",X"E0",X"19",X"4E",X"06",
		X"00",X"ED",X"43",X"62",X"E0",X"21",X"74",X"64",X"19",X"19",X"56",X"1E",X"50",X"ED",X"53",X"64",
		X"E0",X"23",X"7E",X"32",X"C5",X"E2",X"3E",X"28",X"32",X"C6",X"E2",X"3A",X"06",X"E7",X"FE",X"03",
		X"38",X"02",X"3E",X"02",X"21",X"04",X"E7",X"46",X"10",X"02",X"C6",X"03",X"87",X"5F",X"16",X"00",
		X"21",X"B0",X"64",X"19",X"5E",X"23",X"56",X"EB",X"22",X"78",X"E0",X"29",X"11",X"C0",X"FF",X"19",
		X"22",X"7A",X"E0",X"C9",X"12",X"18",X"11",X"16",X"10",X"15",X"0F",X"13",X"0E",X"12",X"0D",X"10",
		X"0C",X"10",X"0B",X"0E",X"0A",X"0D",X"09",X"0C",X"08",X"0A",X"07",X"0A",X"06",X"08",X"06",X"07",
		X"06",X"06",X"07",X"07",X"0B",X"0B",X"0F",X"08",X"08",X"0C",X"0C",X"11",X"09",X"09",X"0D",X"0D",
		X"13",X"08",X"08",X"0B",X"0B",X"10",X"09",X"09",X"0D",X"0D",X"13",X"0A",X"0A",X"0F",X"0F",X"15",
		X"C0",X"05",X"D8",X"06",X"37",X"08",X"10",X"05",X"06",X"06",X"42",X"07",X"3E",X"10",X"C3",X"B0",
		X"5E",X"3A",X"1E",X"E7",X"A7",X"20",X"F5",X"21",X"54",X"65",X"3A",X"06",X"E7",X"FE",X"03",X"38",
		X"02",X"3E",X"02",X"87",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"5E",X"23",X"56",X"EB",X"CD",X"8A",
		X"59",X"21",X"7D",X"65",X"CD",X"8A",X"59",X"21",X"8F",X"65",X"CD",X"8A",X"59",X"3A",X"06",X"E7",
		X"A7",X"20",X"13",X"3A",X"1C",X"E0",X"87",X"30",X"0D",X"3E",X"1C",X"CD",X"B0",X"5E",X"CD",X"F7",
		X"5B",X"3E",X"58",X"CD",X"F9",X"5B",X"3E",X"28",X"CD",X"F9",X"5B",X"3E",X"10",X"CD",X"B0",X"5E",
		X"3E",X"15",X"CD",X"B0",X"5E",X"06",X"03",X"21",X"90",X"C0",X"22",X"18",X"E2",X"78",X"C6",X"9B",
		X"6F",X"26",X"88",X"22",X"1A",X"E2",X"3E",X"28",X"CD",X"F9",X"5B",X"3E",X"10",X"CD",X"B0",X"5E",
		X"10",X"E5",X"21",X"86",X"65",X"CD",X"8A",X"59",X"3E",X"9B",X"32",X"1A",X"E2",X"3E",X"28",X"CD",
		X"F9",X"5B",X"21",X"6C",X"65",X"CD",X"AC",X"59",X"21",X"8F",X"65",X"CD",X"AC",X"59",X"3E",X"01",
		X"32",X"1E",X"E7",X"C9",X"5A",X"65",X"63",X"65",X"6C",X"65",X"2A",X"83",X"02",X"77",X"72",X"72",
		X"43",X"43",X"21",X"2A",X"83",X"02",X"79",X"77",X"72",X"43",X"43",X"21",X"2A",X"83",X"02",X"73",
		X"74",X"72",X"72",X"43",X"43",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"21",X"2A",X"87",X"02",
		X"52",X"45",X"41",X"44",X"59",X"21",X"2A",X"87",X"02",X"53",X"54",X"41",X"52",X"54",X"21",X"18",
		X"84",X"02",X"4C",X"4F",X"53",X"20",X"41",X"4E",X"47",X"45",X"4C",X"45",X"53",X"21",X"3E",X"00",
		X"32",X"26",X"E7",X"21",X"05",X"E7",X"34",X"7E",X"FE",X"05",X"38",X"15",X"AF",X"77",X"23",X"34",
		X"FD",X"21",X"14",X"89",X"47",X"21",X"1D",X"E7",X"01",X"08",X"00",X"CD",X"1E",X"5C",X"C3",X"F5",
		X"5E",X"21",X"02",X"01",X"22",X"1D",X"E7",X"C9",X"21",X"1C",X"E0",X"35",X"31",X"00",X"E8",X"FB",
		X"CD",X"D9",X"63",X"AF",X"CD",X"B0",X"5E",X"3A",X"05",X"E7",X"FE",X"04",X"28",X"0F",X"3E",X"1D",
		X"CD",X"B0",X"5E",X"CD",X"47",X"66",X"3E",X"1A",X"CD",X"B0",X"5E",X"18",X"08",X"3E",X"1E",X"CD",
		X"B0",X"5E",X"CD",X"47",X"66",X"06",X"00",X"3E",X"04",X"CD",X"F9",X"5B",X"3A",X"05",X"E7",X"FE",
		X"04",X"20",X"1F",X"FD",X"21",X"F0",X"E1",X"C5",X"06",X"06",X"FD",X"7E",X"03",X"3D",X"FD",X"77",
		X"A3",X"FD",X"77",X"03",X"FD",X"77",X"63",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",
		X"E9",X"C1",X"78",X"32",X"80",X"E2",X"04",X"FE",X"18",X"38",X"CC",X"CD",X"72",X"66",X"CD",X"1E",
		X"67",X"CD",X"EA",X"68",X"3A",X"05",X"E7",X"FE",X"04",X"20",X"03",X"CD",X"E1",X"69",X"CD",X"9E",
		X"65",X"CD",X"F7",X"5B",X"C3",X"17",X"5F",X"3E",X"80",X"CD",X"F9",X"5B",X"CD",X"D1",X"33",X"21",
		X"00",X"80",X"CD",X"6A",X"66",X"0E",X"16",X"06",X"2B",X"CD",X"6C",X"66",X"36",X"03",X"11",X"11",
		X"00",X"19",X"06",X"44",X"CD",X"6C",X"66",X"0D",X"20",X"ED",X"06",X"80",X"36",X"00",X"23",X"10",
		X"FB",X"C9",X"3A",X"05",X"E7",X"FE",X"04",X"30",X"25",X"21",X"A4",X"66",X"CD",X"8A",X"59",X"3A",
		X"05",X"E7",X"C6",X"73",X"FD",X"77",X"00",X"FD",X"36",X"01",X"04",X"3A",X"05",X"E7",X"87",X"4F",
		X"06",X"00",X"21",X"16",X"67",X"09",X"5E",X"23",X"56",X"23",X"EB",X"C3",X"8A",X"59",X"21",X"F4",
		X"66",X"C3",X"8A",X"59",X"40",X"83",X"04",X"43",X"48",X"45",X"43",X"4B",X"50",X"4F",X"49",X"4E",
		X"54",X"20",X"2F",X"20",X"21",X"3E",X"83",X"05",X"40",X"20",X"4C",X"41",X"53",X"20",X"56",X"45",
		X"47",X"41",X"53",X"20",X"40",X"21",X"3E",X"83",X"05",X"40",X"20",X"48",X"4F",X"55",X"53",X"54",
		X"4F",X"4E",X"20",X"40",X"21",X"3E",X"83",X"05",X"40",X"20",X"53",X"54",X"2E",X"4C",X"4F",X"55",
		X"49",X"53",X"20",X"40",X"21",X"3E",X"83",X"05",X"40",X"20",X"43",X"48",X"49",X"43",X"41",X"47",
		X"4F",X"20",X"40",X"21",X"C0",X"82",X"04",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",
		X"41",X"54",X"49",X"4F",X"4E",X"22",X"3E",X"83",X"05",X"40",X"20",X"4E",X"45",X"57",X"20",X"59",
		X"4F",X"52",X"4B",X"20",X"40",X"21",X"B5",X"66",X"C6",X"66",X"D5",X"66",X"E5",X"66",X"21",X"8F",
		X"67",X"CD",X"8A",X"59",X"FD",X"21",X"A3",X"67",X"CD",X"DD",X"67",X"3E",X"20",X"CD",X"F9",X"5B",
		X"3A",X"0D",X"E7",X"FD",X"BE",X"09",X"38",X"05",X"CD",X"DD",X"67",X"18",X"F3",X"21",X"A2",X"81",
		X"11",X"FC",X"FF",X"FD",X"BE",X"03",X"38",X"09",X"19",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"18",
		X"F2",X"01",X"01",X"09",X"79",X"EE",X"05",X"4F",X"C5",X"CD",X"46",X"68",X"3E",X"10",X"CD",X"F9",
		X"5B",X"C1",X"10",X"F0",X"EB",X"FD",X"66",X"02",X"FD",X"6E",X"01",X"22",X"27",X"E0",X"21",X"80",
		X"05",X"19",X"CD",X"9B",X"68",X"3E",X"10",X"CD",X"F9",X"5B",X"21",X"96",X"81",X"06",X"04",X"C5",
		X"CD",X"53",X"68",X"2B",X"2B",X"2B",X"2B",X"C1",X"10",X"F5",X"3E",X"10",X"C3",X"F9",X"5B",X"A6",
		X"81",X"05",X"52",X"41",X"4E",X"4B",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",
		X"4F",X"49",X"4E",X"54",X"53",X"21",X"01",X"00",X"02",X"02",X"40",X"01",X"03",X"20",X"01",X"04",
		X"00",X"01",X"05",X"80",X"00",X"06",X"60",X"00",X"07",X"30",X"00",X"11",X"24",X"00",X"16",X"22",
		X"00",X"21",X"20",X"00",X"31",X"18",X"00",X"41",X"16",X"00",X"51",X"14",X"00",X"61",X"12",X"00",
		X"71",X"10",X"00",X"81",X"08",X"00",X"91",X"06",X"00",X"99",X"00",X"00",X"A0",X"FD",X"23",X"FD",
		X"23",X"FD",X"23",X"FD",X"E5",X"21",X"A2",X"81",X"CD",X"FB",X"67",X"2B",X"2B",X"2B",X"2B",X"7D",
		X"FE",X"88",X"30",X"F4",X"FD",X"E1",X"3E",X"15",X"C3",X"F9",X"5B",X"11",X"80",X"00",X"FD",X"7E",
		X"00",X"FE",X"A0",X"30",X"4E",X"E5",X"CD",X"65",X"68",X"FD",X"7E",X"03",X"FE",X"A0",X"30",X"47",
		X"D6",X"01",X"27",X"FD",X"BE",X"00",X"28",X"09",X"36",X"1A",X"19",X"36",X"1B",X"19",X"CD",X"65",
		X"68",X"36",X"2D",X"19",X"7C",X"FE",X"87",X"38",X"F8",X"0E",X"2D",X"CD",X"7D",X"68",X"DD",X"21",
		X"5F",X"68",X"06",X"06",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"19",X"10",X"F7",X"E1",X"FD",X"23",
		X"FD",X"23",X"FD",X"23",X"3E",X"01",X"E5",X"23",X"06",X"14",X"11",X"80",X"00",X"77",X"19",X"10",
		X"FC",X"E1",X"C9",X"E5",X"AF",X"18",X"F1",X"36",X"1A",X"19",X"36",X"1B",X"19",X"18",X"C2",X"30",
		X"30",X"20",X"50",X"54",X"53",X"F5",X"1F",X"1F",X"1F",X"1F",X"E6",X"0F",X"28",X"03",X"CD",X"74",
		X"68",X"F1",X"E6",X"0F",X"F6",X"30",X"77",X"19",X"C9",X"FD",X"21",X"26",X"E0",X"06",X"00",X"FD",
		X"7E",X"02",X"CD",X"91",X"68",X"FD",X"7E",X"01",X"F5",X"1F",X"1F",X"1F",X"1F",X"CD",X"91",X"68",
		X"F1",X"04",X"E6",X"0F",X"20",X"DE",X"10",X"DC",X"71",X"19",X"C9",X"E5",X"2A",X"27",X"E0",X"7D",
		X"D6",X"01",X"27",X"6F",X"7C",X"DE",X"00",X"27",X"67",X"22",X"27",X"E0",X"E1",X"D8",X"E5",X"0E",
		X"2D",X"11",X"80",X"00",X"CD",X"79",X"68",X"AF",X"32",X"F0",X"E3",X"3A",X"05",X"E7",X"D6",X"04",
		X"28",X"02",X"3E",X"07",X"CD",X"48",X"5C",X"CD",X"E4",X"61",X"3E",X"04",X"CD",X"F9",X"5B",X"3A",
		X"27",X"E0",X"E6",X"03",X"20",X"C6",X"3E",X"13",X"CD",X"B0",X"5E",X"18",X"BF",X"ED",X"5B",X"23",
		X"E7",X"22",X"23",X"E7",X"ED",X"52",X"C6",X"02",X"18",X"21",X"21",X"C1",X"69",X"11",X"27",X"E0",
		X"01",X"20",X"00",X"ED",X"B0",X"2A",X"21",X"E7",X"3A",X"05",X"E7",X"FE",X"04",X"3A",X"16",X"E0",
		X"DA",X"DD",X"68",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"E5",X"87",X"5F",X"16",X"00",
		X"21",X"D9",X"69",X"19",X"5E",X"23",X"56",X"E1",X"EB",X"AF",X"47",X"C6",X"01",X"27",X"30",X"01",
		X"04",X"ED",X"52",X"30",X"F6",X"21",X"39",X"E0",X"CD",X"AF",X"69",X"3A",X"16",X"E0",X"A7",X"20",
		X"06",X"21",X"5E",X"5F",X"22",X"3C",X"E0",X"21",X"27",X"E0",X"CD",X"8A",X"59",X"CD",X"F3",X"5B",
		X"3A",X"05",X"E7",X"5F",X"16",X"00",X"FE",X"04",X"20",X"0E",X"21",X"2B",X"E7",X"7E",X"A7",X"3A",
		X"0D",X"E7",X"28",X"03",X"BE",X"30",X"01",X"77",X"21",X"C2",X"E0",X"19",X"FD",X"21",X"90",X"88",
		X"3A",X"0D",X"E7",X"BE",X"30",X"12",X"77",X"CD",X"78",X"69",X"21",X"97",X"69",X"CD",X"8A",X"59",
		X"3E",X"11",X"CD",X"B0",X"5E",X"C3",X"F3",X"5B",X"E5",X"21",X"86",X"69",X"CD",X"8A",X"59",X"E1",
		X"CD",X"27",X"6C",X"C3",X"F7",X"5B",X"10",X"82",X"01",X"54",X"4F",X"44",X"41",X"59",X"3F",X"53",
		X"20",X"42",X"45",X"53",X"54",X"20",X"21",X"0C",X"81",X"05",X"59",X"4F",X"55",X"20",X"53",X"45",
		X"54",X"20",X"41",X"20",X"4E",X"45",X"57",X"20",X"52",X"45",X"43",X"4F",X"52",X"44",X"21",X"11",
		X"01",X"00",X"F5",X"78",X"A7",X"28",X"03",X"C6",X"30",X"77",X"19",X"F1",X"06",X"02",X"C3",X"88",
		X"68",X"96",X"81",X"01",X"41",X"56",X"45",X"52",X"41",X"47",X"45",X"20",X"53",X"50",X"45",X"45",
		X"44",X"20",X"20",X"20",X"20",X"20",X"5B",X"5C",X"21",X"7D",X"83",X"18",X"B8",X"32",X"69",X"47",
		X"93",X"CD",X"F7",X"5B",X"21",X"97",X"69",X"CD",X"AC",X"59",X"21",X"32",X"6A",X"CD",X"8A",X"59",
		X"21",X"00",X"00",X"22",X"27",X"E0",X"AF",X"CD",X"48",X"5C",X"2A",X"27",X"E0",X"7D",X"C6",X"01",
		X"27",X"6F",X"7C",X"CE",X"00",X"27",X"67",X"22",X"27",X"E0",X"21",X"8C",X"84",X"0E",X"00",X"CD",
		X"79",X"68",X"2A",X"07",X"E7",X"25",X"FA",X"26",X"6A",X"22",X"07",X"E7",X"CD",X"E4",X"61",X"3E",
		X"06",X"CD",X"F9",X"5B",X"18",X"D0",X"21",X"00",X"00",X"22",X"07",X"E7",X"CD",X"E4",X"61",X"C3",
		X"F3",X"5B",X"10",X"82",X"04",X"20",X"20",X"20",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"20",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",X"22",X"8C",X"84",X"04",X"20",X"20",X"20",X"30",X"30",
		X"20",X"50",X"54",X"53",X"21",X"C9",X"3A",X"04",X"D0",X"CB",X"6F",X"C0",X"21",X"8C",X"6A",X"CD",
		X"8A",X"59",X"AF",X"F5",X"FD",X"21",X"20",X"89",X"CD",X"00",X"5A",X"3E",X"50",X"32",X"25",X"E0",
		X"21",X"26",X"E0",X"7E",X"4E",X"A9",X"A1",X"1F",X"38",X"09",X"3A",X"25",X"E0",X"47",X"79",X"10",
		X"F3",X"F1",X"C9",X"CD",X"9E",X"65",X"F1",X"C6",X"01",X"27",X"18",X"D7",X"30",X"82",X"00",X"50",
		X"49",X"43",X"54",X"55",X"52",X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"53",X"45",
		X"54",X"22",X"28",X"84",X"00",X"4E",X"45",X"58",X"54",X"20",X"31",X"50",X"20",X"42",X"55",X"54",
		X"54",X"4F",X"4E",X"22",X"20",X"84",X"00",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"20",X"3D",
		X"20",X"20",X"20",X"20",X"21",X"21",X"BB",X"E0",X"11",X"00",X"E7",X"CD",X"A0",X"6B",X"D8",X"0E",
		X"03",X"EB",X"ED",X"B0",X"EB",X"3A",X"2B",X"E7",X"77",X"06",X"03",X"23",X"36",X"00",X"10",X"FB",
		X"0E",X"09",X"21",X"B4",X"E0",X"CD",X"9A",X"6B",X"38",X"14",X"06",X"07",X"C5",X"4E",X"1A",X"77",
		X"79",X"12",X"23",X"13",X"10",X"F7",X"C1",X"11",X"F2",X"FF",X"19",X"0D",X"20",X"E7",X"C5",X"CD",
		X"5C",X"6C",X"C1",X"21",X"FF",X"FF",X"22",X"29",X"E0",X"AF",X"32",X"28",X"E0",X"3E",X"20",X"CD",
		X"F9",X"5B",X"AF",X"32",X"23",X"E0",X"CD",X"11",X"6C",X"3E",X"41",X"77",X"CD",X"F4",X"6B",X"21",
		X"22",X"E0",X"3A",X"27",X"E0",X"AE",X"28",X"F7",X"7E",X"32",X"27",X"E0",X"E6",X"1F",X"28",X"28",
		X"E6",X"0F",X"CC",X"C8",X"6B",X"2A",X"1F",X"E0",X"ED",X"5B",X"29",X"E0",X"22",X"29",X"E0",X"7A",
		X"AC",X"A4",X"E6",X"01",X"28",X"17",X"CD",X"D9",X"6B",X"21",X"28",X"E0",X"34",X"7E",X"FE",X"03",
		X"38",X"BB",X"CD",X"11",X"6C",X"C3",X"F3",X"5B",X"CD",X"D9",X"6B",X"18",X"D8",X"3A",X"23",X"E0",
		X"FE",X"32",X"30",X"30",X"7D",X"57",X"21",X"2B",X"E0",X"A7",X"28",X"B3",X"AB",X"A2",X"06",X"1C",
		X"20",X"06",X"35",X"20",X"AA",X"06",X"0B",X"7A",X"70",X"1F",X"38",X"0D",X"CD",X"11",X"6C",X"7E",
		X"3D",X"FE",X"41",X"30",X"96",X"3E",X"5A",X"18",X"92",X"CD",X"11",X"6C",X"7E",X"3C",X"FE",X"5B",
		X"30",X"87",X"18",X"87",X"CD",X"11",X"6C",X"36",X"00",X"C9",X"11",X"07",X"00",X"EB",X"19",X"EB",
		X"E5",X"D5",X"06",X"03",X"A7",X"1A",X"9E",X"23",X"13",X"10",X"FA",X"D1",X"E1",X"C9",X"79",X"87",
		X"87",X"5F",X"87",X"91",X"6F",X"26",X"00",X"3E",X"2C",X"93",X"5F",X"16",X"81",X"FD",X"21",X"00",
		X"00",X"FD",X"19",X"11",X"7E",X"E0",X"19",X"C9",X"CD",X"AE",X"6B",X"11",X"80",X"00",X"06",X"11",
		X"FD",X"36",X"00",X"00",X"FD",X"19",X"10",X"F8",X"C9",X"CD",X"AE",X"6B",X"79",X"C6",X"01",X"27",
		X"06",X"01",X"CD",X"17",X"5A",X"FD",X"19",X"CD",X"AC",X"5C",X"FD",X"19",X"FD",X"19",X"23",X"23",
		X"23",X"CD",X"27",X"6C",X"CD",X"03",X"6C",X"06",X"03",X"7E",X"FD",X"77",X"00",X"23",X"FD",X"19",
		X"10",X"F7",X"C9",X"CD",X"AE",X"6B",X"11",X"80",X"08",X"FD",X"19",X"11",X"80",X"00",X"23",X"23",
		X"C9",X"CD",X"03",X"6C",X"3A",X"28",X"E0",X"3C",X"FD",X"36",X"01",X"05",X"3D",X"C8",X"FD",X"36",
		X"01",X"01",X"FD",X"19",X"2C",X"18",X"F1",X"7E",X"A7",X"28",X"20",X"06",X"01",X"CD",X"16",X"5A",
		X"7E",X"FE",X"20",X"38",X"02",X"E6",X"0F",X"3D",X"FE",X"03",X"38",X"02",X"3E",X"03",X"87",X"C6",
		X"0E",X"CD",X"45",X"6C",X"3C",X"FD",X"77",X"00",X"FD",X"19",X"C9",X"3E",X"A2",X"06",X"06",X"FD",
		X"77",X"00",X"FD",X"36",X"01",X"41",X"3C",X"FD",X"19",X"10",X"F4",X"C9",X"CD",X"66",X"5E",X"21",
		X"71",X"6C",X"CD",X"8A",X"59",X"0E",X"00",X"CD",X"D9",X"6B",X"0C",X"79",X"FE",X"0A",X"38",X"F7",
		X"C9",X"B6",X"82",X"01",X"42",X"45",X"53",X"54",X"20",X"31",X"30",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"53",X"22",X"30",X"81",X"01",X"4E",X"4F",X"2E",X"20",X"53",X"43",X"4F",X"52",X"45",
		X"20",X"20",X"52",X"41",X"4E",X"4B",X"20",X"4E",X"41",X"4D",X"45",X"21",X"00",X"65",X"03",X"01",
		X"49",X"45",X"4F",X"00",X"27",X"03",X"03",X"52",X"52",X"54",X"00",X"94",X"02",X"02",X"45",X"53",
		X"45",X"00",X"48",X"02",X"10",X"4D",X"45",X"4D",X"00",X"19",X"02",X"00",X"4E",X"55",X"4F",X"00",
		X"61",X"01",X"11",X"4F",X"53",X"49",X"00",X"33",X"01",X"00",X"54",X"41",X"49",X"00",X"96",X"00",
		X"00",X"52",X"57",X"49",X"00",X"72",X"00",X"00",X"41",X"41",X"57",X"00",X"50",X"00",X"00",X"56",
		X"54",X"41",X"75",X"60",X"45",X"30",X"15",X"2A",X"04",X"E7",X"2D",X"2D",X"C0",X"3A",X"22",X"E0",
		X"87",X"0E",X"85",X"FD",X"21",X"61",X"6D",X"24",X"25",X"28",X"0D",X"21",X"D7",X"E2",X"CB",X"4E",
		X"C8",X"1F",X"0E",X"80",X"FD",X"21",X"59",X"6D",X"06",X"01",X"E6",X"3F",X"28",X"04",X"05",X"E6",
		X"1F",X"C0",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"FD",X"23",X"FD",X"23",X"FD",X"7E",X"00",X"FD",
		X"23",X"FE",X"FE",X"30",X"25",X"D6",X"50",X"38",X"0C",X"11",X"7E",X"00",X"D6",X"50",X"38",X"04",
		X"D6",X"50",X"1D",X"1D",X"19",X"C6",X"50",X"28",X"02",X"C6",X"60",X"10",X"10",X"BE",X"C0",X"71",
		X"3E",X"C0",X"23",X"B6",X"77",X"23",X"0C",X"04",X"18",X"D2",X"28",X"C6",X"C9",X"5F",X"79",X"BE",
		X"C0",X"73",X"23",X"7E",X"E6",X"8F",X"77",X"18",X"EC",X"34",X"8A",X"01",X"02",X"03",X"A8",X"00",
		X"FF",X"B0",X"81",X"0D",X"61",X"63",X"64",X"FE",X"AE",X"83",X"16",X"68",X"6A",X"6E",X"FE",X"32",
		X"87",X"2C",X"FE",X"B0",X"89",X"39",X"3A",X"8D",X"91",X"E4",X"45",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
