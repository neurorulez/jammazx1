library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity colony7_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of colony7_prog is
	type rom is array(0 to  22527) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7E",X"D7",X"D4",X"7E",X"D7",X"AA",X"7E",X"D7",X"B6",X"7E",X"D7",X"BC",X"7E",X"D7",X"C2",
		X"7E",X"D7",X"C8",X"7E",X"D7",X"CE",X"7E",X"D7",X"B0",X"A7",X"A0",X"5A",X"26",X"FB",X"39",X"A7",
		X"A4",X"31",X"A9",X"01",X"00",X"5A",X"26",X"F7",X"39",X"5F",X"D7",X"00",X"F7",X"D0",X"00",X"B6",
		X"CC",X"00",X"C6",X"02",X"D7",X"00",X"F7",X"D0",X"00",X"39",X"D6",X"04",X"56",X"56",X"56",X"D8",
		X"04",X"56",X"06",X"03",X"06",X"04",X"39",X"34",X"02",X"A6",X"80",X"BD",X"EF",X"3E",X"A6",X"80",
		X"26",X"F9",X"35",X"02",X"39",X"7E",X"F9",X"01",X"7E",X"EB",X"A2",X"7E",X"F6",X"75",X"7E",X"E4",
		X"0F",X"7E",X"DE",X"32",X"7E",X"FE",X"E5",X"7E",X"EB",X"17",X"02",X"04",X"03",X"05",X"03",X"05",
		X"04",X"07",X"86",X"03",X"97",X"00",X"B7",X"D0",X"00",X"7E",X"C0",X"00",X"1A",X"10",X"7F",X"D0",
		X"00",X"86",X"38",X"B7",X"C3",X"FC",X"8E",X"CC",X"00",X"6F",X"01",X"6F",X"03",X"6F",X"05",X"6F",
		X"07",X"86",X"C0",X"A7",X"84",X"86",X"FF",X"A7",X"02",X"6F",X"04",X"6F",X"06",X"CC",X"34",X"3C",
		X"A7",X"01",X"E7",X"03",X"A7",X"05",X"E7",X"07",X"6C",X"01",X"6F",X"84",X"6F",X"02",X"10",X"CE",
		X"C0",X"00",X"CC",X"38",X"3F",X"B7",X"C3",X"FC",X"F7",X"CC",X"02",X"8E",X"C0",X"10",X"CC",X"00",
		X"00",X"ED",X"83",X"8C",X"A0",X"00",X"26",X"F9",X"1C",X"EF",X"CC",X"A5",X"A0",X"1F",X"9B",X"DD",
		X"03",X"BD",X"F9",X"01",X"96",X"07",X"26",X"FC",X"C6",X"10",X"D7",X"07",X"8E",X"A1",X"76",X"9F",
		X"A4",X"BD",X"E8",X"91",X"BD",X"FE",X"C1",X"BD",X"FE",X"C9",X"BD",X"D3",X"0C",X"BD",X"D7",X"1D",
		X"BD",X"EC",X"CE",X"BD",X"F5",X"AE",X"BD",X"EA",X"D0",X"BD",X"DD",X"47",X"BD",X"EE",X"B9",X"BD",
		X"EB",X"88",X"96",X"0B",X"2A",X"09",X"BD",X"FD",X"20",X"BD",X"EF",X"A1",X"BD",X"F0",X"51",X"9E",
		X"A4",X"9F",X"A0",X"8E",X"A1",X"3E",X"9F",X"A6",X"BD",X"F6",X"04",X"BD",X"D1",X"9D",X"BD",X"F3",
		X"AA",X"BD",X"E2",X"79",X"BD",X"E3",X"32",X"BD",X"E0",X"44",X"BD",X"E0",X"97",X"BD",X"E1",X"5D",
		X"9E",X"A4",X"9F",X"A2",X"BD",X"FA",X"A0",X"BD",X"F2",X"0B",X"BD",X"F2",X"88",X"BD",X"F2",X"C6",
		X"BD",X"E8",X"85",X"BD",X"F3",X"4A",X"BD",X"E8",X"E1",X"BD",X"EE",X"FF",X"BD",X"F0",X"91",X"BD",
		X"E9",X"CD",X"BD",X"F9",X"E5",X"96",X"93",X"27",X"11",X"91",X"95",X"27",X"0D",X"81",X"0E",X"22",
		X"04",X"D6",X"0B",X"2A",X"05",X"B7",X"CC",X"02",X"97",X"95",X"BD",X"ED",X"A2",X"86",X"3F",X"B7",
		X"CC",X"02",X"96",X"7D",X"27",X"02",X"0A",X"7D",X"96",X"80",X"27",X"02",X"0A",X"80",X"96",X"94",
		X"27",X"08",X"0A",X"94",X"26",X"04",X"0F",X"93",X"0F",X"95",X"96",X"07",X"27",X"0C",X"96",X"6C",
		X"27",X"08",X"0F",X"6C",X"BD",X"EB",X"17",X"BD",X"D6",X"F9",X"7E",X"D0",X"D4",X"96",X"63",X"10",
		X"26",X"00",X"E8",X"96",X"7E",X"27",X"03",X"0A",X"7E",X"39",X"96",X"7A",X"91",X"21",X"10",X"24",
		X"00",X"D9",X"96",X"20",X"10",X"27",X"00",X"D3",X"96",X"7B",X"27",X"16",X"0A",X"7B",X"96",X"88",
		X"10",X"27",X"00",X"C7",X"D6",X"89",X"27",X"01",X"5A",X"8E",X"FE",X"91",X"BD",X"FB",X"41",X"7E",
		X"D2",X"8B",X"96",X"8E",X"27",X"36",X"86",X"20",X"97",X"7B",X"CC",X"00",X"D6",X"97",X"88",X"97",
		X"8E",X"10",X"8E",X"20",X"18",X"BD",X"D0",X"19",X"10",X"8E",X"21",X"00",X"BD",X"D0",X"19",X"BD",
		X"D0",X"19",X"8E",X"FE",X"7D",X"10",X"8E",X"84",X"14",X"BD",X"D0",X"47",X"BD",X"F8",X"EA",X"8E",
		X"D5",X"A7",X"10",X"8E",X"78",X"20",X"BD",X"D0",X"47",X"7E",X"D2",X"8B",X"0A",X"20",X"BD",X"D0",
		X"3A",X"96",X"1F",X"4A",X"81",X"0F",X"23",X"02",X"86",X"0F",X"48",X"48",X"48",X"8E",X"D2",X"8C",
		X"31",X"86",X"8E",X"B7",X"DC",X"CE",X"AA",X"10",X"A6",X"46",X"27",X"07",X"30",X"88",X"10",X"33",
		X"48",X"20",X"F5",X"0C",X"7A",X"EC",X"A1",X"ED",X"46",X"DC",X"03",X"85",X"24",X"26",X"0E",X"5D",
		X"2B",X"06",X"0D",X"77",X"26",X"06",X"20",X"05",X"0D",X"76",X"27",X"01",X"50",X"E7",X"41",X"C4",
		X"1F",X"CB",X"10",X"D7",X"7B",X"E6",X"A0",X"3D",X"AB",X"A0",X"A7",X"C4",X"CC",X"00",X"00",X"ED",
		X"44",X"A7",X"08",X"BD",X"D0",X"3A",X"C4",X"1F",X"CB",X"10",X"E7",X"84",X"DC",X"03",X"E6",X"A0",
		X"3D",X"AB",X"A0",X"A7",X"06",X"BD",X"D0",X"3A",X"C4",X"78",X"26",X"02",X"CB",X"08",X"E7",X"02",
		X"96",X"03",X"E6",X"A0",X"3D",X"AB",X"A0",X"8B",X"C0",X"A7",X"0A",X"39",X"EB",X"A2",X"40",X"B0",
		X"28",X"60",X"02",X"01",X"EB",X"A2",X"40",X"B0",X"28",X"60",X"02",X"01",X"EB",X"A2",X"40",X"B0",
		X"30",X"60",X"02",X"01",X"EB",X"A2",X"40",X"B0",X"28",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",
		X"28",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",X"2C",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",
		X"2C",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",X"30",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",
		X"30",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",X"30",X"60",X"03",X"01",X"EB",X"A2",X"40",X"B0",
		X"30",X"60",X"03",X"01",X"EB",X"A2",X"34",X"B8",X"28",X"60",X"04",X"01",X"EB",X"A2",X"34",X"B8",
		X"28",X"60",X"04",X"01",X"EB",X"A2",X"34",X"B8",X"2C",X"60",X"04",X"01",X"EB",X"A2",X"34",X"B8",
		X"2C",X"60",X"04",X"01",X"EB",X"A2",X"34",X"B8",X"30",X"60",X"04",X"01",X"96",X"11",X"10",X"26",
		X"02",X"E5",X"96",X"58",X"10",X"27",X"02",X"C7",X"96",X"12",X"10",X"27",X"02",X"D9",X"8B",X"99",
		X"19",X"97",X"12",X"0F",X"0E",X"4F",X"5F",X"DD",X"19",X"DD",X"1B",X"DD",X"1D",X"DD",X"58",X"97",
		X"0C",X"97",X"0D",X"8E",X"A0",X"1F",X"ED",X"81",X"8C",X"A0",X"3F",X"26",X"F9",X"86",X"1E",X"97",
		X"20",X"BD",X"F9",X"01",X"96",X"0E",X"27",X"09",X"97",X"0D",X"86",X"33",X"97",X"0F",X"BD",X"EB",
		X"17",X"0F",X"0D",X"CC",X"99",X"14",X"97",X"0F",X"D7",X"6F",X"BD",X"EB",X"17",X"96",X"0B",X"8A",
		X"80",X"97",X"0B",X"0C",X"11",X"8E",X"FE",X"A5",X"B6",X"CC",X"00",X"44",X"24",X"03",X"8E",X"FE",
		X"B1",X"9F",X"13",X"CC",X"1C",X"00",X"D7",X"20",X"DD",X"2F",X"DD",X"49",X"4C",X"DD",X"33",X"DD",
		X"4D",X"CC",X"06",X"00",X"DD",X"31",X"DD",X"4B",X"4C",X"DD",X"35",X"DD",X"4F",X"F6",X"CC",X"00",
		X"C4",X"03",X"58",X"8E",X"D0",X"6A",X"3A",X"EC",X"84",X"97",X"38",X"97",X"52",X"D7",X"9E",X"0F",
		X"37",X"0F",X"51",X"CC",X"FF",X"88",X"97",X"6E",X"8E",X"D6",X"9C",X"10",X"8E",X"78",X"40",X"BD",
		X"D0",X"47",X"C6",X"11",X"10",X"8E",X"6E",X"60",X"BD",X"D0",X"47",X"C6",X"88",X"8E",X"D6",X"CF",
		X"10",X"8E",X"55",X"48",X"BD",X"D0",X"47",X"86",X"31",X"BD",X"EF",X"3E",X"C6",X"AA",X"8E",X"D6",
		X"E0",X"10",X"8E",X"28",X"20",X"BD",X"D0",X"47",X"96",X"0E",X"26",X"12",X"96",X"12",X"26",X"53",
		X"C6",X"88",X"8E",X"D6",X"C2",X"10",X"8E",X"5F",X"50",X"BD",X"D0",X"47",X"20",X"45",X"C6",X"11",
		X"8E",X"D6",X"B7",X"10",X"8E",X"69",X"58",X"BD",X"D0",X"47",X"C6",X"88",X"8E",X"D6",X"CF",X"10",
		X"8E",X"37",X"48",X"BD",X"D0",X"47",X"86",X"32",X"BD",X"EF",X"3E",X"96",X"12",X"26",X"1D",X"10",
		X"8E",X"4B",X"78",X"BD",X"D0",X"47",X"8E",X"D6",X"C2",X"10",X"8E",X"5F",X"50",X"BD",X"D0",X"47",
		X"8E",X"D6",X"C2",X"10",X"8E",X"41",X"50",X"BD",X"D0",X"47",X"20",X"07",X"10",X"8E",X"46",X"78",
		X"BD",X"D0",X"47",X"96",X"07",X"26",X"FC",X"86",X"10",X"96",X"92",X"81",X"03",X"10",X"27",X"01",
		X"81",X"97",X"07",X"BD",X"E8",X"91",X"BD",X"FE",X"C1",X"BD",X"FE",X"C9",X"27",X"41",X"96",X"93",
		X"B7",X"CC",X"02",X"8E",X"D5",X"A7",X"10",X"8E",X"5F",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",
		X"10",X"8E",X"4B",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",X"10",X"8E",X"41",X"20",X"BD",X"D0",
		X"47",X"96",X"0E",X"27",X"1A",X"96",X"92",X"26",X"16",X"C6",X"88",X"8E",X"D6",X"DD",X"10",X"8E",
		X"46",X"78",X"BD",X"D0",X"47",X"CC",X"3F",X"00",X"B7",X"CC",X"02",X"D7",X"93",X"D7",X"94",X"96",
		X"59",X"10",X"26",X"01",X"2D",X"96",X"58",X"10",X"27",X"00",X"91",X"0F",X"58",X"96",X"0E",X"26",
		X"23",X"96",X"12",X"27",X"8E",X"8B",X"99",X"19",X"97",X"12",X"BD",X"FE",X"E5",X"CC",X"24",X"00",
		X"DD",X"2F",X"4C",X"DD",X"33",X"CC",X"09",X"00",X"DD",X"31",X"4C",X"DD",X"35",X"96",X"9E",X"97",
		X"38",X"7E",X"D5",X"C2",X"96",X"92",X"44",X"10",X"25",X"FF",X"68",X"96",X"12",X"10",X"27",X"FF",
		X"62",X"8B",X"99",X"19",X"97",X"12",X"26",X"10",X"96",X"92",X"26",X"0C",X"C6",X"88",X"8E",X"D6",
		X"C2",X"10",X"8E",X"41",X"50",X"BD",X"D0",X"47",X"BD",X"FE",X"E5",X"0C",X"92",X"CC",X"24",X"00",
		X"DD",X"2F",X"4C",X"DD",X"33",X"CC",X"09",X"00",X"DD",X"31",X"4C",X"DD",X"35",X"96",X"9E",X"97",
		X"38",X"8E",X"D5",X"A7",X"10",X"8E",X"5F",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",X"10",X"8E",
		X"55",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",X"10",X"8E",X"4B",X"20",X"BD",X"D0",X"47",X"8E",
		X"D5",X"A7",X"10",X"8E",X"46",X"20",X"BD",X"D0",X"47",X"7E",X"D4",X"33",X"96",X"57",X"10",X"27",
		X"FF",X"01",X"0F",X"57",X"96",X"0E",X"10",X"27",X"FE",X"F9",X"96",X"92",X"44",X"44",X"10",X"25",
		X"FE",X"F1",X"96",X"12",X"10",X"27",X"FE",X"EB",X"8B",X"99",X"19",X"97",X"12",X"26",X"10",X"96",
		X"92",X"26",X"0C",X"C6",X"88",X"8E",X"D6",X"C2",X"10",X"8E",X"5F",X"50",X"BD",X"D0",X"47",X"BD",
		X"FE",X"E5",X"96",X"92",X"8A",X"02",X"97",X"92",X"CC",X"24",X"00",X"DD",X"49",X"4C",X"DD",X"4D",
		X"CC",X"09",X"00",X"DD",X"4B",X"4C",X"DD",X"4F",X"96",X"9E",X"97",X"52",X"8E",X"D5",X"A7",X"10",
		X"8E",X"4B",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",X"10",X"8E",X"46",X"20",X"BD",X"D0",X"47",
		X"8E",X"D5",X"A7",X"10",X"8E",X"41",X"20",X"BD",X"D0",X"47",X"8E",X"D5",X"A7",X"10",X"8E",X"37",
		X"20",X"BD",X"D0",X"47",X"7E",X"D4",X"33",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"00",X"8E",X"80",X"00",X"CC",X"00",X"00",X"ED",X"83",X"8C",X"28",X"00",X"26",X"F9",X"9E",
		X"13",X"EC",X"84",X"10",X"AE",X"02",X"BD",X"D0",X"19",X"0F",X"92",X"BD",X"F9",X"BD",X"39",X"96",
		X"57",X"27",X"FB",X"96",X"12",X"81",X"02",X"25",X"0E",X"8B",X"98",X"19",X"97",X"12",X"4F",X"97",
		X"57",X"4C",X"97",X"0E",X"7E",X"D3",X"25",X"0F",X"57",X"0F",X"58",X"39",X"0C",X"0C",X"86",X"02",
		X"F6",X"CC",X"00",X"54",X"24",X"01",X"4C",X"91",X"0C",X"27",X"2C",X"0F",X"0D",X"BD",X"F9",X"01",
		X"9E",X"13",X"30",X"04",X"9F",X"13",X"EC",X"84",X"10",X"AE",X"02",X"BD",X"D0",X"19",X"96",X"0E",
		X"27",X"09",X"0C",X"0D",X"86",X"33",X"97",X"0F",X"BD",X"EB",X"17",X"0F",X"0D",X"CC",X"99",X"14",
		X"97",X"0F",X"D7",X"6F",X"7E",X"EB",X"17",X"4F",X"97",X"0B",X"97",X"11",X"97",X"0D",X"97",X"6F",
		X"9E",X"13",X"EC",X"04",X"10",X"AE",X"06",X"BD",X"D0",X"19",X"96",X"19",X"91",X"1C",X"22",X"1C",
		X"26",X"0E",X"96",X"1A",X"91",X"1D",X"22",X"14",X"26",X"06",X"96",X"1B",X"91",X"1E",X"24",X"0C",
		X"CC",X"33",X"88",X"DD",X"9C",X"BD",X"FB",X"DD",X"0C",X"0D",X"20",X"03",X"BD",X"FB",X"D8",X"CC",
		X"80",X"88",X"97",X"6B",X"8E",X"FA",X"7C",X"10",X"8E",X"8A",X"14",X"BD",X"D0",X"47",X"10",X"8E",
		X"84",X"14",X"BD",X"D0",X"47",X"96",X"9C",X"97",X"0F",X"0F",X"0D",X"BD",X"EB",X"17",X"96",X"0E",
		X"27",X"09",X"96",X"9D",X"97",X"0F",X"0C",X"0D",X"BD",X"EB",X"17",X"39",X"45",X"58",X"54",X"45",
		X"4E",X"44",X"45",X"44",X"40",X"57",X"45",X"41",X"50",X"4F",X"4E",X"52",X"59",X"00",X"31",X"40",
		X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"50",X"45",X"52",X"40",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"00",X"44",X"45",X"50",X"4F",X"53",X"49",X"54",X"40",X"43",X"4F",X"49",X"4E",X"00",X"50",
		X"52",X"45",X"53",X"53",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"00",X"4F",X"52",X"00",
		X"50",X"52",X"45",X"53",X"53",X"40",X"46",X"49",X"52",X"45",X"40",X"54",X"4F",X"40",X"53",X"54",
		X"41",X"52",X"54",X"40",X"47",X"41",X"4D",X"45",X"00",X"96",X"37",X"26",X"1F",X"8E",X"A0",X"19",
		X"96",X"0D",X"27",X"03",X"8E",X"A0",X"1C",X"A6",X"84",X"91",X"38",X"2D",X"0F",X"0C",X"37",X"86",
		X"AA",X"97",X"0F",X"7E",X"EB",X"17",X"91",X"93",X"25",X"02",X"DD",X"93",X"39",X"96",X"6B",X"27",
		X"09",X"96",X"70",X"26",X"02",X"0A",X"6B",X"0F",X"63",X"39",X"96",X"0B",X"9A",X"11",X"9A",X"74",
		X"26",X"F5",X"96",X"77",X"94",X"76",X"27",X"EF",X"86",X"02",X"97",X"00",X"B7",X"D0",X"00",X"BD",
		X"C0",X"00",X"4F",X"97",X"00",X"B7",X"D0",X"00",X"39",X"34",X"36",X"8E",X"CE",X"AE",X"10",X"AE",
		X"81",X"27",X"07",X"EC",X"81",X"BD",X"D0",X"19",X"20",X"F4",X"10",X"8E",X"0B",X"5C",X"86",X"B0",
		X"A7",X"A4",X"BD",X"D8",X"06",X"BD",X"D8",X"3C",X"BD",X"C7",X"F0",X"BD",X"D8",X"72",X"CC",X"BD",
		X"EC",X"8E",X"BF",X"BE",X"10",X"8E",X"B1",X"BC",X"CE",X"0C",X"98",X"BD",X"D8",X"C6",X"CC",X"BD",
		X"EC",X"8E",X"BF",X"BE",X"10",X"8E",X"B1",X"BC",X"CE",X"0F",X"70",X"BD",X"D8",X"C6",X"CC",X"5D",
		X"EC",X"8E",X"5F",X"5E",X"10",X"8E",X"51",X"5C",X"CE",X"12",X"E3",X"BD",X"D8",X"C6",X"BD",X"C8",
		X"70",X"BD",X"D8",X"D6",X"BD",X"D9",X"3D",X"35",X"36",X"39",X"34",X"10",X"C6",X"33",X"20",X"28",
		X"34",X"10",X"C6",X"22",X"20",X"22",X"34",X"10",X"C6",X"AA",X"20",X"1C",X"34",X"10",X"C6",X"44",
		X"20",X"16",X"34",X"10",X"C6",X"88",X"20",X"10",X"34",X"10",X"C6",X"55",X"20",X"0A",X"34",X"10",
		X"C6",X"BB",X"20",X"04",X"34",X"10",X"C6",X"11",X"E7",X"E2",X"EC",X"A4",X"44",X"1F",X"01",X"86",
		X"F0",X"25",X"02",X"86",X"0F",X"A4",X"84",X"A7",X"84",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",
		X"A6",X"E0",X"25",X"09",X"84",X"F0",X"AA",X"84",X"A7",X"84",X"35",X"10",X"39",X"84",X"0F",X"AA",
		X"84",X"A7",X"84",X"35",X"10",X"39",X"34",X"26",X"10",X"8E",X"1D",X"0D",X"CC",X"52",X"52",X"ED",
		X"A1",X"ED",X"A4",X"10",X"8E",X"1E",X"0D",X"CC",X"20",X"20",X"ED",X"A1",X"ED",X"A4",X"31",X"A9",
		X"01",X"01",X"A7",X"A4",X"31",X"A9",X"00",X"FE",X"A7",X"A4",X"CC",X"22",X"2C",X"31",X"A9",X"FE",
		X"00",X"A7",X"A4",X"31",X"A9",X"01",X"00",X"ED",X"A4",X"35",X"26",X"39",X"34",X"26",X"10",X"8E",
		X"1D",X"EE",X"CC",X"52",X"52",X"ED",X"A1",X"ED",X"A4",X"10",X"8E",X"1E",X"EE",X"CC",X"20",X"20",
		X"ED",X"A1",X"ED",X"A4",X"31",X"A9",X"00",X"FE",X"A7",X"A4",X"31",X"A9",X"01",X"02",X"A7",X"A4",
		X"CC",X"2C",X"22",X"31",X"A9",X"FE",X"00",X"E7",X"A4",X"31",X"A9",X"00",X"FF",X"ED",X"A4",X"35",
		X"26",X"39",X"CC",X"33",X"33",X"8E",X"33",X"33",X"10",X"8E",X"33",X"33",X"CE",X"12",X"81",X"36",
		X"32",X"CC",X"03",X"30",X"8E",X"33",X"30",X"10",X"8E",X"33",X"30",X"CE",X"13",X"83",X"36",X"02",
		X"36",X"02",X"36",X"36",X"36",X"02",X"CC",X"11",X"11",X"8E",X"11",X"11",X"10",X"8E",X"11",X"11",
		X"CE",X"14",X"84",X"36",X"36",X"36",X"32",X"86",X"AA",X"8E",X"8A",X"AA",X"10",X"8E",X"8A",X"AA",
		X"CE",X"15",X"83",X"36",X"30",X"36",X"32",X"86",X"80",X"8E",X"80",X"80",X"10",X"8E",X"80",X"80",
		X"CE",X"16",X"81",X"36",X"32",X"39",X"36",X"32",X"8E",X"1E",X"CF",X"10",X"8E",X"FD",X"DF",X"33",
		X"C9",X"01",X"05",X"7E",X"CF",X"E4",X"CC",X"22",X"22",X"8E",X"22",X"22",X"10",X"8E",X"22",X"22",
		X"CE",X"0F",X"C8",X"36",X"36",X"36",X"36",X"CE",X"12",X"C8",X"36",X"36",X"36",X"36",X"CE",X"15",
		X"C8",X"36",X"36",X"36",X"36",X"CE",X"0C",X"C8",X"36",X"36",X"36",X"36",X"CC",X"33",X"33",X"8E",
		X"33",X"43",X"10",X"8E",X"43",X"33",X"CE",X"0E",X"C6",X"36",X"36",X"36",X"06",X"CE",X"11",X"C6",
		X"36",X"36",X"36",X"06",X"CE",X"14",X"C6",X"36",X"36",X"36",X"06",X"CE",X"0B",X"C3",X"36",X"06",
		X"36",X"06",X"36",X"02",X"8E",X"34",X"34",X"CE",X"0D",X"C4",X"36",X"12",X"36",X"02",X"CE",X"10",
		X"C4",X"36",X"12",X"36",X"02",X"CE",X"13",X"C4",X"36",X"12",X"36",X"02",X"39",X"86",X"0C",X"10",
		X"8E",X"03",X"3C",X"CE",X"0E",X"CF",X"36",X"22",X"C6",X"03",X"8E",X"33",X"3C",X"CE",X"12",X"D5",
		X"36",X"02",X"36",X"04",X"36",X"10",X"36",X"10",X"36",X"22",X"CC",X"33",X"33",X"8E",X"33",X"33",
		X"10",X"8E",X"33",X"33",X"CE",X"11",X"D3",X"36",X"32",X"CC",X"11",X"11",X"8E",X"11",X"11",X"10",
		X"8E",X"11",X"11",X"CE",X"0F",X"D6",X"36",X"36",X"36",X"32",X"CE",X"13",X"D6",X"36",X"36",X"36",
		X"32",X"CC",X"8A",X"AA",X"8E",X"8A",X"AA",X"10",X"8E",X"8A",X"AA",X"CE",X"10",X"D5",X"36",X"36",
		X"36",X"24",X"CE",X"14",X"D5",X"36",X"36",X"36",X"24",X"CC",X"80",X"80",X"8E",X"80",X"80",X"10",
		X"8E",X"80",X"80",X"CE",X"15",X"D3",X"36",X"32",X"39",X"34",X"72",X"86",X"01",X"97",X"00",X"B7",
		X"D0",X"00",X"0C",X"75",X"C1",X"24",X"10",X"25",X"02",X"F7",X"C1",X"2F",X"22",X"59",X"96",X"7C",
		X"85",X"80",X"10",X"26",X"02",X"EB",X"8A",X"80",X"97",X"7C",X"CC",X"0A",X"20",X"BD",X"D7",X"16",
		X"96",X"82",X"26",X"0B",X"0C",X"82",X"CE",X"CE",X"36",X"BD",X"DC",X"D9",X"BD",X"DD",X"FA",X"CE",
		X"CD",X"DA",X"BD",X"DC",X"D9",X"CC",X"50",X"00",X"8E",X"00",X"00",X"10",X"8E",X"50",X"50",X"CE",
		X"0D",X"2D",X"36",X"36",X"4F",X"5F",X"10",X"8E",X"00",X"00",X"CE",X"0E",X"30",X"36",X"36",X"36",
		X"36",X"C6",X"07",X"CE",X"0F",X"27",X"36",X"12",X"33",X"C9",X"01",X"03",X"5A",X"26",X"F7",X"CE",
		X"13",X"2A",X"36",X"12",X"7E",X"DC",X"CE",X"C1",X"43",X"10",X"25",X"02",X"94",X"C1",X"53",X"22",
		X"61",X"96",X"7C",X"85",X"40",X"10",X"26",X"02",X"88",X"8A",X"40",X"97",X"7C",X"CC",X"08",X"20",
		X"BD",X"D7",X"16",X"CE",X"CB",X"6A",X"BD",X"DC",X"D9",X"CC",X"50",X"50",X"8E",X"50",X"50",X"10",
		X"8E",X"50",X"50",X"CE",X"0B",X"51",X"36",X"36",X"36",X"32",X"4F",X"5F",X"8E",X"00",X"00",X"10",
		X"8E",X"00",X"00",X"CE",X"0C",X"4E",X"36",X"36",X"CE",X"0D",X"4F",X"36",X"36",X"36",X"10",X"CE",
		X"0E",X"54",X"36",X"36",X"36",X"36",X"36",X"36",X"CE",X"0F",X"54",X"36",X"36",X"36",X"36",X"36",
		X"36",X"CE",X"10",X"52",X"36",X"36",X"36",X"36",X"36",X"10",X"CE",X"11",X"4E",X"36",X"36",X"7E",
		X"DC",X"CE",X"C1",X"6B",X"10",X"25",X"02",X"29",X"C1",X"6F",X"22",X"49",X"96",X"7C",X"85",X"20",
		X"10",X"26",X"02",X"1D",X"8A",X"20",X"97",X"7C",X"CC",X"09",X"20",X"BD",X"D7",X"16",X"96",X"87",
		X"85",X"04",X"26",X"06",X"8A",X"04",X"97",X"87",X"0C",X"7F",X"CE",X"CC",X"9C",X"BD",X"DC",X"D9",
		X"10",X"8E",X"B0",X"B0",X"8E",X"00",X"00",X"86",X"B0",X"CE",X"0F",X"70",X"36",X"32",X"4F",X"10",
		X"8E",X"00",X"00",X"CE",X"10",X"70",X"36",X"32",X"CE",X"11",X"70",X"36",X"32",X"CE",X"12",X"6F",
		X"36",X"12",X"7E",X"DC",X"CE",X"C1",X"79",X"10",X"25",X"01",X"D6",X"C1",X"83",X"22",X"4E",X"96",
		X"7C",X"85",X"10",X"10",X"26",X"01",X"CA",X"8A",X"10",X"97",X"7C",X"CC",X"08",X"20",X"BD",X"D7",
		X"16",X"CE",X"CB",X"08",X"BD",X"DC",X"D9",X"CC",X"B0",X"B0",X"8E",X"00",X"00",X"10",X"8E",X"00",
		X"00",X"CE",X"11",X"81",X"36",X"02",X"36",X"16",X"CC",X"00",X"00",X"CE",X"12",X"81",X"36",X"32",
		X"CE",X"13",X"83",X"36",X"36",X"36",X"12",X"CE",X"14",X"84",X"36",X"36",X"36",X"32",X"CE",X"15",
		X"83",X"36",X"36",X"36",X"12",X"CE",X"16",X"81",X"36",X"32",X"7E",X"DC",X"CE",X"C1",X"93",X"10",
		X"25",X"01",X"7E",X"C1",X"97",X"22",X"49",X"96",X"7C",X"85",X"08",X"10",X"26",X"01",X"72",X"8A",
		X"08",X"97",X"7C",X"CC",X"09",X"20",X"BD",X"D7",X"16",X"96",X"87",X"85",X"02",X"26",X"06",X"8A",
		X"02",X"97",X"87",X"0C",X"7F",X"CE",X"CC",X"08",X"BD",X"DC",X"D9",X"86",X"B0",X"8E",X"00",X"00",
		X"10",X"8E",X"B0",X"B0",X"CE",X"0C",X"98",X"36",X"32",X"4F",X"10",X"8E",X"00",X"00",X"CE",X"0D",
		X"98",X"36",X"32",X"CE",X"0E",X"98",X"36",X"32",X"CE",X"0F",X"97",X"36",X"12",X"7E",X"DC",X"CE",
		X"C1",X"BB",X"10",X"25",X"01",X"2B",X"C1",X"C7",X"22",X"75",X"96",X"7C",X"85",X"04",X"10",X"26",
		X"01",X"1F",X"8A",X"04",X"97",X"7C",X"CC",X"08",X"20",X"BD",X"D7",X"16",X"CE",X"CD",X"48",X"BD",
		X"DC",X"D9",X"4F",X"5F",X"8E",X"00",X"00",X"10",X"8E",X"00",X"00",X"CE",X"0C",X"C8",X"36",X"36",
		X"36",X"36",X"CE",X"0D",X"C4",X"36",X"32",X"CE",X"0E",X"C6",X"36",X"36",X"36",X"10",X"CE",X"0F",
		X"C8",X"36",X"36",X"36",X"36",X"CE",X"10",X"C4",X"36",X"32",X"CE",X"11",X"C6",X"36",X"36",X"36",
		X"10",X"CE",X"12",X"C8",X"36",X"36",X"36",X"36",X"CE",X"13",X"C4",X"36",X"32",X"CE",X"14",X"C6",
		X"36",X"36",X"36",X"10",X"CE",X"15",X"C8",X"36",X"36",X"36",X"36",X"CE",X"0B",X"C3",X"CC",X"BB",
		X"BB",X"8E",X"BB",X"BB",X"10",X"8E",X"BB",X"BB",X"36",X"10",X"36",X"36",X"7E",X"DC",X"CE",X"C1",
		X"CB",X"10",X"25",X"00",X"AC",X"C1",X"D5",X"22",X"56",X"96",X"7C",X"85",X"02",X"10",X"26",X"00",
		X"A0",X"8A",X"02",X"97",X"7C",X"CC",X"08",X"20",X"BD",X"D7",X"16",X"CE",X"CC",X"E6",X"BD",X"DC",
		X"D9",X"4F",X"5F",X"8E",X"00",X"00",X"10",X"8E",X"00",X"00",X"CE",X"0E",X"CF",X"36",X"12",X"CE",
		X"0F",X"D6",X"36",X"36",X"36",X"32",X"CE",X"10",X"D5",X"36",X"36",X"36",X"12",X"CE",X"11",X"D3",
		X"36",X"32",X"CE",X"12",X"D5",X"36",X"36",X"36",X"12",X"CE",X"13",X"D6",X"36",X"36",X"36",X"32",
		X"CE",X"14",X"D5",X"36",X"36",X"36",X"12",X"CE",X"15",X"D3",X"36",X"32",X"7E",X"DC",X"CE",X"C1",
		X"DD",X"25",X"4E",X"C1",X"E2",X"22",X"4A",X"96",X"7C",X"85",X"01",X"26",X"44",X"8A",X"01",X"97",
		X"7C",X"CC",X"09",X"20",X"BD",X"D7",X"16",X"96",X"87",X"85",X"01",X"26",X"06",X"8A",X"01",X"97",
		X"87",X"0C",X"7F",X"CE",X"CC",X"52",X"BD",X"DC",X"D9",X"86",X"50",X"8E",X"50",X"00",X"10",X"8E",
		X"00",X"50",X"CE",X"12",X"E3",X"36",X"32",X"4F",X"10",X"8E",X"00",X"00",X"8E",X"00",X"00",X"CE",
		X"13",X"E3",X"36",X"32",X"CE",X"14",X"E3",X"36",X"32",X"CE",X"15",X"E2",X"36",X"12",X"7E",X"DC",
		X"CE",X"A6",X"E4",X"34",X"04",X"1F",X"02",X"E6",X"A4",X"27",X"05",X"4C",X"E6",X"E4",X"20",X"F5",
		X"35",X"04",X"48",X"1F",X"02",X"BD",X"DD",X"04",X"CC",X"01",X"01",X"BD",X"D7",X"16",X"4F",X"97",
		X"00",X"B7",X"D0",X"00",X"35",X"72",X"7E",X"E9",X"02",X"34",X"16",X"8E",X"AF",X"C8",X"A6",X"06",
		X"27",X"04",X"30",X"08",X"20",X"F8",X"EC",X"C1",X"27",X"17",X"ED",X"84",X"EC",X"C1",X"ED",X"04",
		X"EC",X"C1",X"ED",X"06",X"AF",X"9F",X"A0",X"9A",X"DC",X"9A",X"C3",X"00",X"02",X"DD",X"9A",X"20",
		X"DD",X"35",X"16",X"39",X"34",X"56",X"8E",X"AF",X"C8",X"CE",X"DD",X"31",X"A6",X"06",X"27",X"04",
		X"30",X"08",X"20",X"F8",X"EC",X"C1",X"27",X"16",X"10",X"AF",X"84",X"ED",X"04",X"EC",X"C1",X"ED",
		X"06",X"AF",X"9F",X"A0",X"9A",X"DC",X"9A",X"C3",X"00",X"02",X"DD",X"9A",X"20",X"DE",X"35",X"56",
		X"39",X"01",X"FF",X"D0",X"10",X"02",X"FF",X"D0",X"13",X"02",X"00",X"D0",X"13",X"01",X"01",X"D0",
		X"10",X"02",X"01",X"D0",X"13",X"00",X"00",X"10",X"8E",X"A7",X"B8",X"CE",X"A7",X"B8",X"AE",X"A1",
		X"26",X"03",X"0F",X"75",X"39",X"96",X"09",X"26",X"02",X"6A",X"04",X"34",X"20",X"EC",X"84",X"AB",
		X"04",X"EB",X"05",X"C1",X"08",X"23",X"08",X"C1",X"F8",X"24",X"04",X"81",X"0C",X"22",X"17",X"EC",
		X"06",X"2A",X"0F",X"EC",X"84",X"44",X"1F",X"02",X"86",X"F0",X"25",X"02",X"86",X"0F",X"A4",X"A4",
		X"A7",X"A4",X"6F",X"06",X"20",X"57",X"ED",X"02",X"44",X"10",X"AE",X"06",X"2B",X"1C",X"1F",X"02",
		X"86",X"0F",X"25",X"02",X"86",X"F0",X"A4",X"A4",X"27",X"06",X"EC",X"02",X"ED",X"84",X"20",X"3B",
		X"EC",X"02",X"ED",X"84",X"86",X"D0",X"A7",X"06",X"20",X"25",X"1F",X"02",X"86",X"0F",X"25",X"02",
		X"86",X"F0",X"A4",X"A4",X"27",X"19",X"EC",X"84",X"44",X"1F",X"02",X"86",X"F0",X"25",X"02",X"86",
		X"0F",X"A4",X"A4",X"A7",X"A4",X"EC",X"02",X"ED",X"84",X"86",X"01",X"A7",X"06",X"20",X"0C",X"AF",
		X"9F",X"A0",X"A4",X"10",X"9E",X"A4",X"31",X"22",X"10",X"9F",X"A4",X"AF",X"C1",X"35",X"20",X"AE",
		X"A1",X"10",X"26",X"FF",X"70",X"CC",X"00",X"00",X"DF",X"9A",X"10",X"9F",X"9C",X"11",X"93",X"9C",
		X"27",X"07",X"ED",X"C1",X"11",X"93",X"9C",X"26",X"F9",X"39",X"34",X"36",X"4F",X"5F",X"8E",X"00",
		X"00",X"10",X"8E",X"00",X"00",X"CE",X"0F",X"2F",X"36",X"36",X"36",X"06",X"CE",X"10",X"2F",X"36",
		X"36",X"36",X"06",X"CE",X"11",X"2E",X"36",X"32",X"CE",X"12",X"2D",X"36",X"12",X"CE",X"13",X"2D",
		X"36",X"12",X"CE",X"14",X"2D",X"36",X"12",X"CE",X"15",X"2B",X"6F",X"C4",X"35",X"36",X"39",X"7E",
		X"DF",X"71",X"34",X"70",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"ED",X"02",
		X"ED",X"04",X"ED",X"06",X"ED",X"08",X"ED",X"0A",X"ED",X"0C",X"30",X"89",X"01",X"00",X"ED",X"84",
		X"ED",X"02",X"ED",X"04",X"ED",X"06",X"ED",X"08",X"ED",X"0A",X"30",X"89",X"01",X"00",X"ED",X"02",
		X"ED",X"04",X"ED",X"06",X"ED",X"08",X"30",X"89",X"01",X"00",X"ED",X"04",X"ED",X"06",X"EC",X"22",
		X"ED",X"A4",X"44",X"1F",X"01",X"E6",X"24",X"CE",X"DE",X"A3",X"EE",X"C5",X"EC",X"C1",X"2B",X"20",
		X"ED",X"84",X"EC",X"C1",X"ED",X"02",X"EC",X"C1",X"ED",X"04",X"EC",X"C1",X"ED",X"06",X"EC",X"C1",
		X"ED",X"08",X"EC",X"C1",X"ED",X"0A",X"EC",X"C1",X"ED",X"0C",X"30",X"89",X"01",X"00",X"20",X"DC",
		X"35",X"70",X"39",X"DE",X"AF",X"DE",X"BF",X"DE",X"CF",X"DE",X"ED",X"DF",X"0B",X"DF",X"37",X"30",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"30",
		X"33",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"33",
		X"03",X"03",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"10",X"13",X"00",
		X"00",X"00",X"13",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"33",X"33",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"10",X"13",X"10",X"00",X"00",
		X"00",X"10",X"13",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"33",X"30",X"30",X"30",X"33",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"10",X"10",X"13",X"10",X"00",X"00",X"00",X"00",X"00",
		X"10",X"13",X"10",X"10",X"00",X"00",X"00",X"33",X"03",X"03",X"C3",X"D3",X"E3",X"03",X"03",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"03",X"03",X"03",X"03",X"03",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"D0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"0F",X"8D",X"CC",X"07",X"18",X"DD",X"93",X"BD",X"F9",X"D6",X"0C",X"7A",X"34",X"10",X"CE",
		X"DF",X"37",X"EC",X"A4",X"44",X"1F",X"01",X"EC",X"C1",X"85",X"01",X"26",X"20",X"ED",X"84",X"EC",
		X"C1",X"ED",X"02",X"EC",X"C1",X"ED",X"04",X"EC",X"C1",X"ED",X"06",X"EC",X"C1",X"ED",X"08",X"EC",
		X"C1",X"ED",X"0A",X"EC",X"C1",X"ED",X"0C",X"30",X"89",X"01",X"00",X"20",X"DA",X"8E",X"AA",X"50",
		X"CE",X"E0",X"04",X"A6",X"06",X"27",X"04",X"30",X"08",X"20",X"F8",X"EC",X"A4",X"E3",X"C1",X"ED",
		X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EC",X"E9",X"ED",X"06",X"AF",X"9F",X"A0",X"A8",X"DC",X"A8",
		X"C3",X"00",X"02",X"DD",X"A8",X"11",X"83",X"E0",X"44",X"26",X"D8",X"EC",X"A4",X"44",X"1F",X"01",
		X"0C",X"6C",X"8E",X"A0",X"19",X"96",X"0D",X"27",X"03",X"8E",X"A0",X"1C",X"A6",X"02",X"9B",X"29",
		X"19",X"A7",X"02",X"A6",X"01",X"99",X"28",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",X"19",X"A7",
		X"84",X"35",X"10",X"39",X"00",X"00",X"FC",X"FA",X"00",X"02",X"FC",X"FC",X"00",X"08",X"FC",X"03",
		X"00",X"0A",X"FC",X"05",X"00",X"0C",X"FC",X"07",X"02",X"02",X"FF",X"FC",X"02",X"04",X"FD",X"FE",
		X"02",X"06",X"FD",X"02",X"02",X"08",X"FF",X"03",X"02",X"0A",X"FF",X"05",X"04",X"02",X"00",X"FC",
		X"04",X"04",X"01",X"FE",X"04",X"06",X"01",X"01",X"04",X"08",X"00",X"03",X"06",X"04",X"03",X"FE",
		X"06",X"06",X"03",X"01",X"96",X"0B",X"2A",X"0F",X"96",X"7A",X"27",X"0B",X"96",X"6F",X"9A",X"7E",
		X"9A",X"8D",X"BA",X"BF",X"AA",X"27",X"01",X"39",X"96",X"1F",X"4A",X"26",X"06",X"96",X"20",X"81",
		X"0A",X"22",X"F4",X"0C",X"8D",X"CC",X"0B",X"FF",X"BD",X"D7",X"16",X"10",X"8E",X"A1",X"1C",X"CC",
		X"DE",X"32",X"ED",X"26",X"6F",X"24",X"BD",X"D0",X"3A",X"C4",X"01",X"27",X"0E",X"96",X"77",X"26",
		X"0E",X"C6",X"01",X"E7",X"25",X"CC",X"E8",X"08",X"ED",X"A4",X"39",X"96",X"76",X"26",X"F2",X"6F",
		X"25",X"CC",X"E8",X"F8",X"ED",X"A4",X"39",X"96",X"8D",X"26",X"01",X"39",X"10",X"8E",X"A1",X"1C",
		X"C6",X"80",X"A6",X"25",X"26",X"01",X"5F",X"96",X"2A",X"DB",X"09",X"1F",X"01",X"86",X"01",X"97",
		X"00",X"B7",X"D0",X"00",X"AE",X"84",X"4F",X"97",X"00",X"B7",X"D0",X"00",X"1F",X"10",X"AB",X"A4",
		X"EB",X"21",X"ED",X"22",X"C1",X"08",X"10",X"23",X"00",X"81",X"C1",X"F8",X"24",X"7D",X"9E",X"A4",
		X"10",X"AF",X"81",X"9F",X"A4",X"4F",X"C1",X"10",X"25",X"2E",X"C1",X"F0",X"22",X"2A",X"86",X"02",
		X"C1",X"18",X"25",X"24",X"C1",X"E8",X"22",X"20",X"86",X"04",X"C1",X"20",X"25",X"1A",X"C1",X"E0",
		X"22",X"16",X"86",X"06",X"C1",X"28",X"25",X"10",X"C1",X"D8",X"22",X"0C",X"86",X"08",X"C1",X"30",
		X"25",X"06",X"C1",X"D0",X"22",X"02",X"86",X"0A",X"A7",X"24",X"96",X"8D",X"2B",X"8D",X"A6",X"25",
		X"27",X"28",X"EC",X"22",X"D1",X"2C",X"25",X"83",X"86",X"E6",X"CB",X"05",X"8E",X"C0",X"01",X"10",
		X"8E",X"A1",X"14",X"ED",X"A4",X"AF",X"24",X"8E",X"F1",X"48",X"AF",X"26",X"0C",X"8C",X"00",X"8D",
		X"86",X"10",X"97",X"91",X"CC",X"0C",X"30",X"7E",X"D7",X"16",X"EC",X"22",X"D1",X"2B",X"10",X"22",
		X"FF",X"59",X"86",X"E6",X"CB",X"05",X"8E",X"C0",X"FF",X"20",X"D4",X"0F",X"8D",X"EC",X"A4",X"44",
		X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"86",X"08",X"B7",X"BF",X"AA",X"39",X"96",X"8C",X"26",
		X"01",X"39",X"10",X"8E",X"A1",X"14",X"0A",X"91",X"26",X"0F",X"86",X"10",X"97",X"91",X"A6",X"24",
		X"4C",X"81",X"C6",X"23",X"02",X"86",X"C6",X"A7",X"24",X"A6",X"24",X"C6",X"40",X"DB",X"09",X"1F",
		X"01",X"86",X"01",X"97",X"00",X"B7",X"D0",X"00",X"AE",X"84",X"4F",X"97",X"00",X"B7",X"D0",X"00",
		X"1F",X"10",X"AB",X"A4",X"EB",X"25",X"EB",X"21",X"ED",X"22",X"81",X"40",X"22",X"2E",X"0F",X"8C",
		X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"ED",X"02",X"ED",X"89",X"01",X"00",
		X"ED",X"89",X"01",X"02",X"86",X"47",X"A7",X"A4",X"E6",X"25",X"2B",X"08",X"0D",X"77",X"26",X"42",
		X"BD",X"EA",X"68",X"39",X"0D",X"76",X"26",X"3A",X"BD",X"EA",X"38",X"39",X"9E",X"A4",X"10",X"AF",
		X"81",X"9F",X"A4",X"39",X"0F",X"8C",X"CC",X"07",X"10",X"DD",X"93",X"0C",X"6C",X"34",X"10",X"8E",
		X"A0",X"19",X"96",X"0D",X"27",X"03",X"8E",X"A0",X"1C",X"A6",X"02",X"9B",X"29",X"19",X"A7",X"02",
		X"A6",X"01",X"99",X"28",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",X"19",X"A7",X"84",X"35",X"10",
		X"0C",X"7A",X"34",X"30",X"8E",X"AA",X"50",X"10",X"8E",X"A1",X"14",X"CE",X"E2",X"39",X"A6",X"06",
		X"27",X"04",X"30",X"08",X"20",X"F8",X"EC",X"A4",X"E3",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"04",
		X"CC",X"ED",X"80",X"ED",X"06",X"AF",X"9F",X"A0",X"A8",X"DC",X"A8",X"C3",X"00",X"02",X"DD",X"A8",
		X"11",X"83",X"E2",X"79",X"26",X"D8",X"35",X"30",X"39",X"00",X"00",X"FE",X"FE",X"00",X"01",X"FD",
		X"00",X"00",X"02",X"FE",X"02",X"01",X"00",X"FF",X"FD",X"01",X"01",X"FC",X"FE",X"01",X"01",X"FC",
		X"02",X"01",X"01",X"00",X"04",X"01",X"02",X"FF",X"03",X"02",X"00",X"01",X"FD",X"02",X"01",X"00",
		X"FC",X"02",X"01",X"04",X"FE",X"02",X"01",X"04",X"02",X"02",X"02",X"01",X"03",X"03",X"00",X"02",
		X"FE",X"03",X"01",X"03",X"00",X"03",X"02",X"02",X"02",X"96",X"0B",X"2A",X"18",X"96",X"6F",X"26",
		X"14",X"96",X"7E",X"26",X"10",X"96",X"7A",X"27",X"0C",X"96",X"84",X"26",X"08",X"96",X"8F",X"2B",
		X"04",X"DC",X"24",X"26",X"01",X"39",X"4D",X"27",X"0C",X"0D",X"8F",X"26",X"08",X"91",X"20",X"25",
		X"F4",X"0C",X"8F",X"20",X"06",X"D1",X"20",X"25",X"EC",X"03",X"8F",X"0C",X"84",X"10",X"8E",X"A1",
		X"26",X"8E",X"E6",X"82",X"D6",X"03",X"86",X"13",X"3D",X"48",X"48",X"30",X"86",X"30",X"86",X"AF",
		X"28",X"EC",X"81",X"ED",X"A4",X"CC",X"03",X"03",X"ED",X"24",X"CC",X"E4",X"0F",X"ED",X"26",X"31",
		X"2A",X"EC",X"81",X"ED",X"A1",X"EC",X"81",X"ED",X"A1",X"EC",X"81",X"ED",X"A1",X"6F",X"A0",X"BD",
		X"D0",X"3A",X"C4",X"07",X"CB",X"08",X"E7",X"A4",X"D6",X"03",X"C4",X"03",X"58",X"8E",X"E7",X"1C",
		X"3A",X"AE",X"84",X"A6",X"80",X"A7",X"23",X"AF",X"21",X"8E",X"E3",X"25",X"10",X"8E",X"8A",X"AC",
		X"C6",X"88",X"BD",X"D0",X"47",X"8E",X"E3",X"2E",X"10",X"8E",X"84",X"AC",X"BD",X"D0",X"47",X"8E",
		X"00",X"02",X"10",X"8E",X"84",X"AC",X"CE",X"A0",X"26",X"0F",X"6D",X"BD",X"EB",X"32",X"8E",X"FE",
		X"78",X"BD",X"D0",X"47",X"39",X"41",X"44",X"56",X"49",X"53",X"4F",X"52",X"53",X"00",X"40",X"40",
		X"40",X"00",X"96",X"84",X"26",X"01",X"39",X"10",X"8E",X"A1",X"26",X"EC",X"2A",X"1F",X"01",X"E6",
		X"A8",X"10",X"3A",X"86",X"01",X"97",X"00",X"B7",X"D0",X"00",X"AE",X"84",X"4F",X"97",X"00",X"B7",
		X"D0",X"00",X"1F",X"10",X"AB",X"A4",X"EB",X"21",X"ED",X"22",X"9E",X"A4",X"10",X"AF",X"81",X"9F",
		X"A4",X"A6",X"A8",X"10",X"8B",X"02",X"84",X"07",X"A7",X"A8",X"10",X"6A",X"A8",X"11",X"26",X"62",
		X"BD",X"D0",X"3A",X"C4",X"07",X"CB",X"08",X"E7",X"A8",X"11",X"AE",X"A8",X"12",X"A6",X"80",X"2B",
		X"11",X"A7",X"A8",X"14",X"AF",X"A8",X"12",X"8E",X"E7",X"8B",X"30",X"86",X"EC",X"84",X"ED",X"24",
		X"20",X"40",X"0F",X"84",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"9E",X"A4",
		X"30",X"1E",X"9F",X"A4",X"ED",X"84",X"8E",X"E3",X"2E",X"10",X"8E",X"84",X"D4",X"BD",X"D0",X"47",
		X"96",X"8B",X"27",X"18",X"8E",X"F6",X"57",X"10",X"8E",X"8A",X"AC",X"C6",X"44",X"BD",X"D0",X"47",
		X"C6",X"CC",X"10",X"8E",X"84",X"AC",X"BD",X"D0",X"47",X"7E",X"E3",X"36",X"BD",X"FB",X"D8",X"7E",
		X"E3",X"36",X"6A",X"2D",X"10",X"26",X"FF",X"5E",X"A6",X"2F",X"27",X"0F",X"6A",X"2E",X"27",X"0B",
		X"A7",X"2D",X"A6",X"2C",X"AB",X"2B",X"A7",X"2B",X"7E",X"E3",X"36",X"AE",X"28",X"30",X"08",X"AF",
		X"28",X"EC",X"81",X"26",X"05",X"8E",X"E6",X"82",X"20",X"F5",X"ED",X"22",X"EC",X"81",X"ED",X"2A",
		X"EC",X"81",X"ED",X"2C",X"EC",X"81",X"ED",X"2E",X"6F",X"A8",X"10",X"39",X"7E",X"E5",X"A7",X"34",
		X"70",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"ED",X"02",X"ED",X"04",X"ED",
		X"06",X"30",X"89",X"01",X"00",X"ED",X"84",X"ED",X"02",X"ED",X"04",X"ED",X"06",X"30",X"89",X"01",
		X"00",X"ED",X"84",X"ED",X"02",X"ED",X"04",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"E6",X"A8",
		X"14",X"CE",X"E4",X"6F",X"24",X"03",X"CE",X"E4",X"7B",X"EE",X"C5",X"C6",X"03",X"10",X"AE",X"C1",
		X"10",X"AF",X"84",X"10",X"AE",X"C1",X"10",X"AF",X"02",X"10",X"AE",X"C1",X"10",X"AF",X"04",X"10",
		X"AE",X"C1",X"10",X"AF",X"06",X"30",X"89",X"01",X"00",X"5A",X"26",X"E1",X"35",X"70",X"39",X"E4",
		X"87",X"E4",X"9F",X"E4",X"B7",X"E4",X"CF",X"E4",X"E7",X"E4",X"FF",X"E5",X"17",X"E5",X"2F",X"E5",
		X"47",X"E5",X"47",X"E5",X"77",X"E5",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"8A",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"8A",X"8A",X"80",X"00",X"00",X"00",X"80",
		X"80",X"84",X"84",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"8A",X"4A",X"8A",X"80",X"00",X"00",X"80",X"8A",X"8A",X"8A",X"8A",X"8A",X"80",X"00",X"00",
		X"00",X"40",X"40",X"40",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"A8",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"08",
		X"08",X"A8",X"A8",X"08",X"08",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"08",X"08",X"04",X"08",X"08",X"00",X"00",X"08",X"08",X"A8",X"A8",X"A8",X"08",X"08",X"00",X"00",
		X"A0",X"A4",X"A4",X"A4",X"A0",X"00",X"00",X"0F",X"84",X"CC",X"07",X"18",X"BD",X"D7",X"16",X"0C",
		X"7A",X"34",X"30",X"CE",X"E4",X"FF",X"EC",X"A4",X"44",X"24",X"03",X"CE",X"E5",X"8F",X"1F",X"01",
		X"C6",X"03",X"10",X"AE",X"C1",X"10",X"AF",X"84",X"10",X"AE",X"C1",X"10",X"AF",X"02",X"10",X"AE",
		X"C1",X"10",X"AF",X"04",X"10",X"AE",X"C1",X"10",X"AF",X"06",X"30",X"89",X"01",X"00",X"5A",X"26",
		X"E1",X"10",X"AE",X"62",X"8E",X"AA",X"50",X"CE",X"E6",X"5E",X"A6",X"06",X"27",X"04",X"30",X"08",
		X"20",X"F8",X"EC",X"A4",X"E3",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EC",X"E9",X"ED",
		X"06",X"AF",X"9F",X"A0",X"A8",X"DC",X"A8",X"C3",X"00",X"02",X"DD",X"A8",X"11",X"83",X"E6",X"82",
		X"26",X"D8",X"0C",X"6C",X"8E",X"A0",X"19",X"96",X"0D",X"27",X"03",X"8E",X"A0",X"1C",X"A6",X"02",
		X"9B",X"27",X"19",X"A7",X"02",X"A6",X"01",X"99",X"26",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",
		X"19",X"A7",X"84",X"8E",X"E3",X"2E",X"10",X"8E",X"84",X"D4",X"BD",X"D0",X"47",X"96",X"8B",X"27",
		X"17",X"8E",X"F6",X"57",X"10",X"8E",X"8A",X"AC",X"C6",X"44",X"BD",X"D0",X"47",X"C6",X"CC",X"10",
		X"8E",X"84",X"AC",X"BD",X"D0",X"47",X"20",X"03",X"BD",X"FB",X"D8",X"35",X"30",X"39",X"00",X"00",
		X"00",X"FB",X"00",X"02",X"FD",X"FD",X"00",X"04",X"FB",X"00",X"02",X"00",X"FD",X"03",X"02",X"02",
		X"00",X"05",X"02",X"04",X"03",X"03",X"02",X"06",X"04",X"02",X"04",X"02",X"05",X"00",X"04",X"04",
		X"03",X"FD",X"C0",X"28",X"C2",X"90",X"00",X"24",X"00",X"00",X"D2",X"5E",X"C3",X"90",X"08",X"01",
		X"0A",X"01",X"E2",X"64",X"C3",X"E0",X"F8",X"01",X"0A",X"01",X"F1",X"65",X"C3",X"90",X"F8",X"02",
		X"02",X"02",X"F3",X"6C",X"C3",X"80",X"00",X"30",X"00",X"00",X"F3",X"C0",X"C3",X"80",X"F8",X"02",
		X"06",X"02",X"EA",X"D2",X"C3",X"50",X"00",X"20",X"00",X"00",X"B2",X"EA",X"C3",X"50",X"F8",X"02",
		X"0C",X"02",X"98",X"D4",X"C3",X"F0",X"00",X"40",X"00",X"00",X"C8",X"64",X"C3",X"F0",X"08",X"02",
		X"18",X"02",X"AF",X"6B",X"C3",X"B0",X"00",X"20",X"00",X"00",X"E7",X"83",X"C3",X"B0",X"F8",X"02",
		X"0E",X"02",X"E3",X"A6",X"C3",X"40",X"00",X"18",X"00",X"00",X"B9",X"A6",X"C3",X"40",X"08",X"02",
		X"0C",X"02",X"A9",X"C4",X"C3",X"A0",X"00",X"18",X"00",X"00",X"C7",X"E2",X"C3",X"A0",X"08",X"02",
		X"0E",X"02",X"E6",X"D0",X"C3",X"10",X"00",X"5E",X"00",X"00",X"A0",X"2C",X"C3",X"10",X"F8",X"02",
		X"10",X"02",X"C0",X"1A",X"C3",X"80",X"00",X"08",X"00",X"00",X"00",X"00",X"E7",X"24",X"E7",X"41",
		X"E7",X"5E",X"E7",X"78",X"00",X"02",X"04",X"06",X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"06",
		X"04",X"02",X"00",X"02",X"04",X"06",X"08",X"0A",X"0A",X"0A",X"0A",X"08",X"06",X"04",X"02",X"00",
		X"FF",X"00",X"02",X"04",X"06",X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"06",X"04",
		X"02",X"04",X"06",X"08",X"0A",X"0A",X"0A",X"0A",X"08",X"06",X"04",X"02",X"00",X"FF",X"00",X"02",
		X"04",X"06",X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"06",X"04",X"02",X"04",X"06",X"08",X"0A",
		X"0A",X"0A",X"08",X"06",X"04",X"02",X"00",X"FF",X"00",X"02",X"04",X"06",X"08",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"08",X"06",X"04",X"02",X"00",X"FF",X"03",X"03",X"03",X"03",X"03",
		X"03",X"04",X"04",X"05",X"07",X"06",X"08",X"BD",X"DD",X"FA",X"CC",X"FE",X"DC",X"8E",X"FE",X"CF",
		X"10",X"8E",X"FD",X"4C",X"CE",X"0F",X"2F",X"36",X"36",X"CC",X"CD",X"E4",X"36",X"02",X"8E",X"FC",
		X"DF",X"10",X"8E",X"ED",X"F0",X"CE",X"10",X"2F",X"36",X"36",X"CC",X"E0",X"F0",X"36",X"02",X"8E",
		X"CF",X"DE",X"10",X"8E",X"EC",X"C0",X"CE",X"11",X"2E",X"36",X"34",X"CC",X"CE",X"FD",X"8E",X"D4",
		X"FD",X"10",X"8E",X"CF",X"EC",X"CE",X"12",X"2D",X"36",X"12",X"CE",X"13",X"2D",X"36",X"24",X"CC",
		X"CE",X"C0",X"8E",X"E4",X"DF",X"CE",X"14",X"2D",X"36",X"12",X"CE",X"15",X"2B",X"E7",X"C4",X"86",
		X"7F",X"97",X"8A",X"39",X"34",X"76",X"C6",X"11",X"8E",X"11",X"11",X"10",X"8E",X"11",X"11",X"96",
		X"87",X"85",X"04",X"26",X"28",X"8A",X"04",X"97",X"87",X"CE",X"10",X"70",X"36",X"34",X"C6",X"13",
		X"8E",X"13",X"13",X"10",X"8E",X"13",X"13",X"CE",X"11",X"70",X"36",X"34",X"C6",X"B1",X"8E",X"B1",
		X"B1",X"10",X"8E",X"B1",X"B1",X"CE",X"0F",X"70",X"36",X"34",X"35",X"76",X"39",X"85",X"02",X"26",
		X"28",X"8A",X"02",X"97",X"87",X"CE",X"0D",X"98",X"36",X"34",X"C6",X"13",X"8E",X"13",X"13",X"10",
		X"8E",X"13",X"13",X"CE",X"0E",X"98",X"36",X"34",X"C6",X"B1",X"8E",X"B1",X"B1",X"10",X"8E",X"B1",
		X"B1",X"CE",X"0C",X"98",X"36",X"34",X"35",X"76",X"39",X"85",X"01",X"26",X"25",X"8A",X"01",X"97",
		X"87",X"CE",X"13",X"E3",X"36",X"34",X"C6",X"13",X"8E",X"13",X"13",X"10",X"8E",X"13",X"13",X"CE",
		X"14",X"E3",X"36",X"34",X"C6",X"51",X"8E",X"51",X"51",X"10",X"8E",X"51",X"51",X"CE",X"12",X"E3",
		X"36",X"34",X"35",X"76",X"39",X"0D",X"8A",X"27",X"07",X"0A",X"8A",X"26",X"03",X"BD",X"DD",X"FA",
		X"39",X"B6",X"CC",X"04",X"26",X"04",X"97",X"15",X"20",X"1D",X"F6",X"CC",X"04",X"94",X"15",X"D7",
		X"15",X"1F",X"89",X"43",X"9A",X"16",X"D7",X"16",X"43",X"27",X"0C",X"8E",X"A0",X"52",X"30",X"01",
		X"44",X"24",X"02",X"6C",X"84",X"26",X"F7",X"B6",X"CC",X"00",X"48",X"BA",X"CC",X"06",X"26",X"04",
		X"97",X"17",X"20",X"1C",X"1F",X"89",X"94",X"17",X"D7",X"17",X"1F",X"89",X"43",X"9A",X"18",X"D7",
		X"18",X"43",X"27",X"0C",X"8E",X"A0",X"5A",X"30",X"01",X"44",X"24",X"02",X"6C",X"84",X"26",X"F7",
		X"39",X"10",X"8E",X"A5",X"76",X"CE",X"A5",X"76",X"AE",X"A1",X"27",X"45",X"EC",X"84",X"AB",X"04",
		X"EB",X"05",X"ED",X"02",X"C1",X"03",X"25",X"0A",X"C1",X"FC",X"22",X"06",X"81",X"43",X"22",X"0D",
		X"20",X"30",X"6F",X"06",X"EC",X"84",X"44",X"1F",X"01",X"6F",X"84",X"20",X"0C",X"AF",X"9F",X"A0",
		X"A4",X"AF",X"C1",X"9E",X"A4",X"30",X"02",X"9F",X"A4",X"AE",X"A1",X"26",X"CF",X"CC",X"00",X"00",
		X"DF",X"AA",X"10",X"9F",X"9C",X"11",X"93",X"9C",X"27",X"07",X"ED",X"C1",X"11",X"93",X"9C",X"26",
		X"F9",X"39",X"C1",X"14",X"10",X"25",X"00",X"BC",X"C1",X"ED",X"10",X"22",X"00",X"B6",X"44",X"10",
		X"AF",X"E3",X"1F",X"02",X"6D",X"A4",X"26",X"09",X"10",X"AE",X"E1",X"81",X"06",X"23",X"B3",X"20",
		X"BC",X"81",X"19",X"24",X"06",X"10",X"AE",X"E1",X"7E",X"D9",X"A9",X"34",X"16",X"6F",X"06",X"EC",
		X"84",X"44",X"1F",X"01",X"6F",X"84",X"35",X"16",X"C1",X"14",X"25",X"E9",X"C1",X"EB",X"22",X"E5",
		X"C1",X"E5",X"25",X"02",X"C6",X"E4",X"81",X"1C",X"22",X"07",X"4C",X"1F",X"02",X"6D",X"A4",X"26",
		X"F5",X"4C",X"1F",X"02",X"CC",X"00",X"00",X"ED",X"A4",X"ED",X"22",X"ED",X"24",X"ED",X"26",X"31",
		X"A9",X"FF",X"00",X"ED",X"A4",X"ED",X"22",X"ED",X"24",X"ED",X"26",X"31",X"A9",X"FF",X"00",X"ED",
		X"A4",X"ED",X"22",X"ED",X"24",X"ED",X"A9",X"FF",X"02",X"EC",X"26",X"84",X"F0",X"C4",X"F0",X"ED",
		X"26",X"31",X"A9",X"FF",X"00",X"A6",X"21",X"84",X"F0",X"A7",X"21",X"A6",X"24",X"84",X"F0",X"A7",
		X"24",X"10",X"AE",X"E1",X"CC",X"03",X"08",X"BD",X"D7",X"16",X"7E",X"E9",X"19",X"96",X"73",X"26",
		X"09",X"96",X"0B",X"2A",X"1E",X"86",X"40",X"97",X"0B",X"39",X"96",X"7C",X"43",X"26",X"14",X"96",
		X"0B",X"2A",X"10",X"96",X"76",X"26",X"02",X"8D",X"4F",X"96",X"77",X"26",X"02",X"8D",X"79",X"86",
		X"20",X"97",X"0B",X"39",X"44",X"10",X"AF",X"E3",X"1F",X"02",X"6D",X"A4",X"26",X"06",X"10",X"AE",
		X"E1",X"7E",X"E9",X"0D",X"10",X"AE",X"E1",X"5D",X"2B",X"17",X"0D",X"76",X"10",X"26",X"EF",X"99",
		X"C1",X"09",X"10",X"25",X"EF",X"93",X"C1",X"13",X"10",X"22",X"EF",X"8D",X"8D",X"1A",X"7E",X"E9",
		X"02",X"0D",X"77",X"10",X"26",X"EF",X"82",X"C1",X"EB",X"10",X"25",X"EF",X"7C",X"C1",X"F6",X"10",
		X"22",X"EF",X"76",X"8D",X"33",X"7E",X"E9",X"02",X"34",X"50",X"0C",X"76",X"0C",X"74",X"0A",X"73",
		X"96",X"0B",X"2A",X"06",X"CC",X"0F",X"40",X"BD",X"D7",X"16",X"8E",X"B7",X"6C",X"CE",X"EA",X"98",
		X"EC",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EB",X"6D",X"ED",X"06",X"30",X"08",X"11",
		X"83",X"EA",X"B4",X"26",X"EB",X"35",X"50",X"39",X"34",X"50",X"0C",X"77",X"0C",X"74",X"0A",X"73",
		X"96",X"0B",X"2A",X"06",X"CC",X"0F",X"40",X"BD",X"D7",X"16",X"8E",X"B7",X"A4",X"CE",X"EA",X"B4",
		X"EC",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EB",X"6D",X"ED",X"06",X"30",X"08",X"11",
		X"83",X"EA",X"D0",X"26",X"EB",X"35",X"50",X"39",X"3A",X"0D",X"03",X"03",X"3A",X"0F",X"04",X"03",
		X"3C",X"0D",X"04",X"02",X"3C",X"0F",X"05",X"02",X"3E",X"0D",X"05",X"01",X"3E",X"0F",X"06",X"01",
		X"40",X"0D",X"06",X"00",X"3A",X"EE",X"03",X"FD",X"3A",X"F0",X"04",X"FD",X"3C",X"EE",X"04",X"FE",
		X"3C",X"F0",X"05",X"FE",X"3E",X"EE",X"05",X"FF",X"3E",X"F0",X"06",X"FF",X"40",X"F0",X"06",X"00",
		X"96",X"74",X"26",X"01",X"39",X"8E",X"B7",X"6C",X"10",X"9E",X"A4",X"A6",X"06",X"27",X"25",X"96",
		X"70",X"26",X"05",X"A6",X"04",X"4A",X"A7",X"04",X"EC",X"04",X"AB",X"84",X"EB",X"01",X"ED",X"02",
		X"81",X"3A",X"24",X"0E",X"6F",X"06",X"EC",X"84",X"44",X"1F",X"03",X"CC",X"00",X"00",X"ED",X"C4",
		X"20",X"02",X"AF",X"A1",X"30",X"08",X"8C",X"B7",X"DC",X"25",X"D0",X"10",X"9C",X"A4",X"26",X"03",
		X"0F",X"74",X"39",X"10",X"9F",X"A4",X"39",X"96",X"0D",X"27",X"09",X"CE",X"A0",X"1C",X"10",X"8E",
		X"84",X"70",X"20",X"07",X"CE",X"A0",X"19",X"10",X"8E",X"8A",X"70",X"D6",X"0F",X"8E",X"00",X"03",
		X"0F",X"6D",X"A6",X"C4",X"44",X"44",X"44",X"44",X"26",X"09",X"8C",X"00",X"01",X"27",X"04",X"0D",
		X"6D",X"27",X"09",X"8A",X"30",X"BD",X"EF",X"3E",X"0C",X"6D",X"20",X"02",X"31",X"28",X"A6",X"C0",
		X"84",X"0F",X"26",X"09",X"8C",X"00",X"01",X"27",X"04",X"0D",X"6D",X"27",X"09",X"8A",X"30",X"BD",
		X"EF",X"3E",X"0C",X"6D",X"20",X"02",X"31",X"28",X"30",X"1F",X"26",X"C6",X"39",X"34",X"10",X"EC",
		X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",
		X"CC",X"88",X"88",X"ED",X"84",X"35",X"10",X"39",X"96",X"6F",X"27",X"12",X"0A",X"6F",X"26",X"0E",
		X"86",X"14",X"97",X"6F",X"96",X"6E",X"27",X"03",X"4F",X"20",X"01",X"4A",X"97",X"6E",X"39",X"7E",
		X"ED",X"03",X"34",X"50",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"ED",X"02",
		X"ED",X"04",X"ED",X"06",X"30",X"89",X"01",X"00",X"ED",X"84",X"ED",X"02",X"ED",X"04",X"ED",X"06",
		X"8E",X"EB",X"FE",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"03",X"25",X"03",X"8E",X"EC",X"5E",X"EC",
		X"24",X"C1",X"0C",X"27",X"0E",X"4D",X"26",X"09",X"CC",X"09",X"02",X"A7",X"24",X"EB",X"25",X"E7",
		X"25",X"6A",X"24",X"58",X"58",X"58",X"3A",X"EC",X"81",X"ED",X"C4",X"EC",X"81",X"ED",X"42",X"EC",
		X"81",X"ED",X"44",X"EC",X"81",X"ED",X"46",X"33",X"C9",X"01",X"00",X"EC",X"81",X"ED",X"C4",X"EC",
		X"81",X"ED",X"42",X"EC",X"81",X"ED",X"44",X"EC",X"84",X"ED",X"46",X"35",X"50",X"39",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"00",X"00",X"00",X"00",X"00",X"20",X"C2",X"D2",X"20",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"02",X"00",X"00",X"00",X"00",X"20",X"C2",X"D2",X"E2",X"20",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"00",X"00",X"00",X"20",X"20",X"C2",X"D2",X"E2",X"20",X"20",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"00",X"00",X"20",X"20",X"C2",X"D2",X"E2",X"F2",X"20",X"20",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"2C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"2C",
		X"2D",X"02",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"02",X"2C",
		X"2D",X"2E",X"02",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"02",X"02",
		X"2C",X"2D",X"2E",X"02",X"02",X"00",X"00",X"00",X"20",X"20",X"20",X"00",X"00",X"00",X"02",X"02",
		X"2C",X"2D",X"2E",X"2F",X"02",X"02",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"8E",X"A1",
		X"3E",X"10",X"AE",X"84",X"27",X"12",X"CC",X"00",X"00",X"ED",X"81",X"EE",X"26",X"ED",X"26",X"0A",
		X"7A",X"AD",X"5D",X"10",X"AE",X"84",X"26",X"EE",X"39",X"34",X"50",X"EC",X"A4",X"44",X"1F",X"01",
		X"CC",X"00",X"00",X"EE",X"84",X"ED",X"84",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"EF",X"84",
		X"35",X"50",X"39",X"34",X"10",X"CC",X"04",X"0C",X"BD",X"D7",X"16",X"BD",X"F8",X"EA",X"8E",X"AA",
		X"50",X"CE",X"ED",X"60",X"A6",X"06",X"27",X"04",X"30",X"08",X"20",X"F8",X"EC",X"A4",X"E3",X"C1",
		X"ED",X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EC",X"E9",X"ED",X"06",X"AF",X"9F",X"A0",X"A8",X"DC",
		X"A8",X"C3",X"00",X"02",X"DD",X"A8",X"11",X"83",X"ED",X"80",X"26",X"D8",X"0C",X"6C",X"8E",X"A0",
		X"19",X"96",X"0D",X"27",X"03",X"8E",X"A0",X"1C",X"A6",X"02",X"9B",X"23",X"19",X"A7",X"02",X"A6",
		X"01",X"99",X"22",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",X"19",X"A7",X"84",X"35",X"10",X"39",
		X"00",X"00",X"FC",X"FC",X"00",X"02",X"FB",X"00",X"00",X"04",X"FC",X"04",X"00",X"06",X"00",X"05",
		X"02",X"00",X"00",X"FB",X"02",X"02",X"04",X"FC",X"02",X"04",X"05",X"00",X"02",X"06",X"04",X"04",
		X"34",X"10",X"EC",X"A4",X"44",X"1F",X"01",X"86",X"00",X"A7",X"84",X"EC",X"22",X"ED",X"A4",X"44",
		X"1F",X"01",X"25",X"07",X"86",X"80",X"A7",X"84",X"35",X"10",X"39",X"86",X"08",X"A7",X"84",X"35",
		X"10",X"39",X"0F",X"08",X"8E",X"A1",X"76",X"CE",X"A1",X"76",X"10",X"AE",X"84",X"27",X"2C",X"CC",
		X"00",X"00",X"ED",X"81",X"96",X"07",X"27",X"17",X"AB",X"21",X"B1",X"C8",X"00",X"22",X"09",X"96",
		X"07",X"AB",X"23",X"B1",X"C8",X"00",X"25",X"07",X"0C",X"08",X"10",X"AF",X"C1",X"20",X"03",X"AD",
		X"B8",X"06",X"10",X"AE",X"84",X"26",X"D8",X"96",X"08",X"26",X"C7",X"39",X"34",X"10",X"EC",X"A4",
		X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"A7",X"02",X"ED",X"89",X"01",X"00",X"A7",X"89",
		X"01",X"02",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"25",X"11",X"CC",X"0D",X"C2",X"ED",X"84",
		X"CC",X"0F",X"E0",X"A7",X"02",X"E7",X"89",X"01",X"01",X"35",X"10",X"39",X"CC",X"0C",X"D0",X"A7",
		X"01",X"E7",X"89",X"01",X"00",X"CC",X"2E",X"F0",X"ED",X"89",X"01",X"01",X"35",X"10",X"39",X"34",
		X"10",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"A7",X"02",X"ED",X"89",X"01",
		X"00",X"A7",X"89",X"01",X"02",X"35",X"10",X"39",X"34",X"10",X"EC",X"A4",X"44",X"1F",X"01",X"CC",
		X"00",X"00",X"A7",X"03",X"A7",X"89",X"01",X"03",X"ED",X"89",X"02",X"00",X"ED",X"89",X"02",X"02",
		X"ED",X"89",X"02",X"04",X"A7",X"89",X"02",X"06",X"A7",X"89",X"03",X"03",X"A7",X"89",X"04",X"03",
		X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"25",X"27",X"CC",X"01",X"1D",X"A7",X"03",X"E7",X"89",
		X"01",X"03",X"CC",X"10",X"10",X"ED",X"89",X"02",X"00",X"ED",X"89",X"02",X"05",X"4C",X"A7",X"89",
		X"03",X"03",X"CC",X"D0",X"0D",X"ED",X"89",X"02",X"02",X"A7",X"89",X"02",X"04",X"35",X"10",X"39",
		X"CC",X"01",X"01",X"ED",X"89",X"02",X"00",X"ED",X"89",X"02",X"05",X"CC",X"0D",X"D0",X"ED",X"89",
		X"02",X"02",X"A7",X"89",X"02",X"04",X"5C",X"E7",X"89",X"03",X"03",X"CC",X"11",X"10",X"A7",X"89",
		X"01",X"03",X"E7",X"89",X"04",X"03",X"35",X"10",X"39",X"96",X"63",X"26",X"41",X"CE",X"A9",X"B8",
		X"9E",X"A4",X"EF",X"81",X"9F",X"A4",X"8E",X"F8",X"B5",X"5F",X"96",X"0B",X"2A",X"03",X"F6",X"CC",
		X"04",X"C4",X"0F",X"58",X"3A",X"EC",X"C4",X"AB",X"84",X"EB",X"01",X"81",X"50",X"24",X"04",X"86",
		X"50",X"20",X"06",X"81",X"F6",X"23",X"02",X"86",X"F6",X"C1",X"0E",X"24",X"04",X"C6",X"0E",X"20",
		X"06",X"C1",X"E9",X"23",X"02",X"C6",X"E9",X"ED",X"42",X"8E",X"EE",X"38",X"AF",X"46",X"39",X"96",
		X"02",X"27",X"03",X"0A",X"02",X"39",X"96",X"63",X"26",X"F4",X"BD",X"D0",X"3A",X"C4",X"1E",X"D7",
		X"02",X"8E",X"A1",X"56",X"3A",X"10",X"AE",X"84",X"27",X"04",X"4F",X"BD",X"EF",X"2E",X"96",X"03",
		X"C6",X"B0",X"3D",X"8B",X"50",X"D6",X"04",X"ED",X"84",X"10",X"9E",X"03",X"20",X"02",X"1E",X"02",
		X"44",X"1E",X"02",X"25",X"04",X"84",X"70",X"20",X"02",X"84",X"07",X"A7",X"A4",X"39",X"34",X"14",
		X"80",X"30",X"2A",X"0B",X"1F",X"20",X"80",X"06",X"C6",X"08",X"1F",X"02",X"35",X"14",X"39",X"C6",
		X"18",X"3D",X"8E",X"C7",X"00",X"30",X"8B",X"86",X"01",X"D6",X"00",X"97",X"00",X"B7",X"D0",X"00",
		X"D7",X"01",X"C6",X"04",X"6F",X"A0",X"A6",X"80",X"A4",X"E4",X"A7",X"A0",X"A6",X"80",X"A4",X"E4",
		X"A7",X"A0",X"A6",X"80",X"A4",X"E4",X"A7",X"A0",X"A6",X"80",X"A4",X"E4",X"A7",X"A0",X"A6",X"80",
		X"A4",X"E4",X"A7",X"A0",X"A6",X"80",X"A4",X"E4",X"A7",X"A0",X"6F",X"A4",X"31",X"A9",X"00",X"F9",
		X"5A",X"26",X"D1",X"31",X"A9",X"FC",X"08",X"D6",X"01",X"D7",X"00",X"F7",X"D0",X"00",X"35",X"14",
		X"39",X"96",X"59",X"27",X"4D",X"0F",X"59",X"96",X"88",X"26",X"47",X"96",X"6F",X"27",X"15",X"0F",
		X"6F",X"CC",X"FF",X"99",X"97",X"6E",X"D7",X"0F",X"0C",X"6C",X"8E",X"D5",X"A7",X"10",X"8E",X"60",
		X"20",X"BD",X"D0",X"47",X"8E",X"A0",X"B0",X"CE",X"A9",X"C0",X"CC",X"02",X"02",X"BD",X"D7",X"16",
		X"EC",X"84",X"27",X"1F",X"8E",X"A0",X"C4",X"CE",X"A9",X"C8",X"EC",X"84",X"27",X"15",X"8E",X"A0",
		X"D8",X"CE",X"A9",X"D0",X"EC",X"84",X"27",X"0B",X"8E",X"A0",X"EC",X"CE",X"A9",X"D8",X"EC",X"84",
		X"27",X"01",X"39",X"FC",X"A9",X"B8",X"C3",X"04",X"03",X"ED",X"84",X"80",X"40",X"C0",X"10",X"44",
		X"54",X"ED",X"02",X"44",X"54",X"ED",X"04",X"44",X"54",X"ED",X"06",X"44",X"54",X"ED",X"08",X"44",
		X"54",X"ED",X"0A",X"6F",X"0C",X"C6",X"ED",X"F0",X"A9",X"B9",X"C0",X"03",X"54",X"E7",X"0E",X"54",
		X"E7",X"0F",X"54",X"E7",X"88",X"10",X"54",X"E7",X"88",X"11",X"54",X"E7",X"88",X"12",X"CC",X"80",
		X"80",X"ED",X"C4",X"ED",X"C8",X"28",X"CC",X"ED",X"DC",X"ED",X"46",X"ED",X"C8",X"2E",X"A7",X"44",
		X"A7",X"C8",X"2C",X"96",X"76",X"26",X"02",X"6F",X"44",X"96",X"77",X"26",X"03",X"6F",X"C8",X"2C",
		X"39",X"96",X"5A",X"27",X"3B",X"0F",X"5A",X"96",X"7D",X"9A",X"7E",X"9A",X"88",X"26",X"31",X"0C",
		X"7F",X"96",X"7F",X"81",X"03",X"23",X"03",X"0A",X"7F",X"39",X"86",X"30",X"97",X"7D",X"8E",X"A1",
		X"00",X"CE",X"A9",X"E0",X"CC",X"05",X"0C",X"DD",X"93",X"EC",X"84",X"26",X"13",X"BD",X"EF",X"F3",
		X"CC",X"F1",X"48",X"ED",X"46",X"ED",X"C8",X"2E",X"FC",X"A9",X"B8",X"DD",X"96",X"BD",X"E7",X"F4",
		X"39",X"8E",X"A0",X"B0",X"10",X"8E",X"A9",X"C0",X"EC",X"84",X"26",X"0C",X"30",X"88",X"14",X"31",
		X"28",X"10",X"8C",X"A9",X"E8",X"2D",X"F1",X"39",X"6C",X"0C",X"A6",X"0C",X"85",X"F8",X"27",X"3C",
		X"CC",X"EE",X"1F",X"ED",X"26",X"ED",X"A8",X"2E",X"10",X"8C",X"A9",X"E0",X"27",X"26",X"DE",X"A4",
		X"A6",X"24",X"26",X"03",X"10",X"AF",X"C1",X"A6",X"A8",X"2C",X"26",X"07",X"1F",X"20",X"C3",X"00",
		X"28",X"ED",X"C1",X"DF",X"A4",X"CC",X"00",X"00",X"ED",X"84",X"34",X"10",X"BD",X"F1",X"C1",X"35",
		X"10",X"7E",X"F0",X"98",X"CC",X"00",X"00",X"ED",X"84",X"7E",X"F1",X"89",X"A7",X"0D",X"EC",X"84",
		X"EB",X"88",X"10",X"1F",X"03",X"CC",X"40",X"10",X"64",X"0D",X"24",X"04",X"E3",X"06",X"20",X"07",
		X"1E",X"03",X"EB",X"88",X"10",X"1E",X"03",X"64",X"0D",X"24",X"04",X"E3",X"04",X"20",X"06",X"1E",
		X"03",X"EB",X"0F",X"1E",X"03",X"64",X"0D",X"24",X"04",X"E3",X"02",X"20",X"06",X"1E",X"03",X"EB",
		X"0E",X"1E",X"03",X"ED",X"22",X"EF",X"A8",X"2A",X"A7",X"A8",X"2A",X"DE",X"A4",X"A6",X"24",X"26",
		X"03",X"10",X"AF",X"C1",X"A6",X"A8",X"2C",X"26",X"07",X"1F",X"20",X"C3",X"00",X"28",X"ED",X"C1",
		X"DF",X"A4",X"7E",X"F0",X"9C",X"7E",X"E1",X"D4",X"34",X"10",X"EC",X"A4",X"44",X"1F",X"01",X"CC",
		X"00",X"00",X"ED",X"84",X"A7",X"02",X"ED",X"89",X"01",X"00",X"A7",X"89",X"01",X"02",X"EC",X"22",
		X"ED",X"A4",X"44",X"1F",X"01",X"25",X"10",X"CC",X"08",X"88",X"ED",X"84",X"A7",X"02",X"C6",X"80",
		X"E7",X"89",X"01",X"01",X"35",X"10",X"39",X"CC",X"08",X"80",X"A7",X"01",X"E7",X"89",X"01",X"00",
		X"86",X"88",X"ED",X"89",X"01",X"01",X"35",X"10",X"39",X"FD",X"A9",X"E2",X"FF",X"AA",X"0A",X"B7",
		X"AA",X"0A",X"8E",X"A9",X"E0",X"10",X"8E",X"AA",X"08",X"DE",X"A4",X"B6",X"A9",X"E4",X"26",X"02",
		X"AF",X"C1",X"B6",X"AA",X"0C",X"26",X"03",X"10",X"AF",X"C1",X"DF",X"A4",X"8E",X"B8",X"5C",X"10",
		X"9E",X"AC",X"86",X"08",X"97",X"83",X"CC",X"ED",X"80",X"DE",X"33",X"DF",X"9C",X"DE",X"2F",X"20",
		X"1D",X"8E",X"B8",X"5C",X"10",X"9E",X"AC",X"86",X"10",X"97",X"83",X"CC",X"D0",X"0A",X"DE",X"35",
		X"DF",X"9C",X"DE",X"31",X"0D",X"77",X"26",X"04",X"0D",X"76",X"27",X"02",X"08",X"83",X"DD",X"9E",
		X"FC",X"A9",X"B8",X"C3",X"04",X"03",X"DD",X"98",X"A6",X"06",X"27",X"04",X"30",X"08",X"20",X"F8",
		X"AF",X"A1",X"DC",X"98",X"ED",X"84",X"30",X"04",X"EF",X"81",X"DC",X"9E",X"ED",X"81",X"96",X"83",
		X"33",X"C6",X"11",X"93",X"9C",X"26",X"E1",X"10",X"9F",X"AC",X"39",X"10",X"8E",X"BE",X"38",X"CE",
		X"BE",X"38",X"AE",X"A1",X"27",X"F4",X"6A",X"04",X"27",X"2F",X"86",X"01",X"97",X"00",X"B7",X"D0",
		X"00",X"86",X"C6",X"E6",X"05",X"DB",X"09",X"AF",X"E3",X"1F",X"01",X"EC",X"84",X"AE",X"E1",X"0F",
		X"00",X"7F",X"D0",X"00",X"AB",X"84",X"EB",X"01",X"ED",X"02",X"81",X"48",X"22",X"19",X"34",X"16",
		X"44",X"1F",X"01",X"A6",X"84",X"35",X"16",X"27",X"0E",X"6F",X"06",X"EC",X"84",X"44",X"1F",X"01",
		X"CC",X"00",X"00",X"ED",X"84",X"20",X"18",X"81",X"FB",X"22",X"EE",X"C1",X"05",X"25",X"EA",X"C1",
		X"FB",X"22",X"E6",X"AF",X"9F",X"A0",X"A4",X"AF",X"C1",X"9E",X"A4",X"30",X"02",X"9F",X"A4",X"AE",
		X"A1",X"26",X"A3",X"CC",X"00",X"00",X"DF",X"AC",X"10",X"9F",X"9C",X"11",X"93",X"9C",X"27",X"07",
		X"ED",X"C1",X"11",X"93",X"9C",X"26",X"F9",X"39",X"DE",X"A0",X"96",X"5B",X"26",X"05",X"11",X"93",
		X"A2",X"26",X"01",X"39",X"AE",X"C1",X"EC",X"02",X"8E",X"BE",X"38",X"10",X"AE",X"81",X"27",X"EE",
		X"A1",X"22",X"22",X"F7",X"8B",X"08",X"A1",X"22",X"23",X"18",X"E1",X"23",X"22",X"14",X"CB",X"08",
		X"E1",X"23",X"23",X"0C",X"AE",X"5E",X"10",X"9E",X"A6",X"AF",X"A1",X"10",X"9F",X"A6",X"20",X"CE",
		X"C0",X"08",X"80",X"08",X"20",X"D5",X"96",X"5B",X"27",X"7F",X"0F",X"5B",X"96",X"0B",X"2A",X"79",
		X"96",X"88",X"9A",X"7E",X"9A",X"82",X"26",X"71",X"97",X"8B",X"97",X"84",X"0C",X"82",X"BD",X"E7",
		X"97",X"CC",X"0D",X"04",X"BD",X"D7",X"16",X"DE",X"A6",X"10",X"9E",X"A0",X"10",X"9C",X"A2",X"27",
		X"06",X"AE",X"A1",X"AF",X"C1",X"20",X"F5",X"DF",X"A6",X"CE",X"FE",X"00",X"8E",X"B8",X"5C",X"10",
		X"9E",X"AC",X"A6",X"06",X"27",X"04",X"30",X"08",X"20",X"F8",X"AF",X"A1",X"CC",X"A0",X"80",X"ED",
		X"84",X"30",X"04",X"EF",X"81",X"CC",X"F3",X"88",X"ED",X"81",X"33",X"C8",X"10",X"11",X"83",X"FF",
		X"00",X"26",X"DF",X"10",X"9F",X"AC",X"CC",X"40",X"0C",X"97",X"7E",X"D7",X"80",X"0C",X"81",X"8E",
		X"A5",X"76",X"9F",X"AA",X"10",X"AE",X"84",X"27",X"10",X"EC",X"A4",X"44",X"1F",X"03",X"CC",X"00",
		X"00",X"A7",X"C4",X"A7",X"26",X"ED",X"81",X"20",X"EB",X"39",X"96",X"81",X"26",X"01",X"39",X"96",
		X"80",X"26",X"FB",X"0F",X"81",X"CC",X"0E",X"04",X"BD",X"D7",X"16",X"CE",X"FE",X"00",X"8E",X"B8",
		X"5C",X"10",X"9E",X"AC",X"A6",X"06",X"27",X"04",X"30",X"08",X"20",X"F8",X"AF",X"A1",X"CC",X"A0",
		X"80",X"ED",X"84",X"30",X"04",X"EF",X"81",X"CC",X"ED",X"80",X"ED",X"81",X"33",X"48",X"11",X"83",
		X"FF",X"00",X"26",X"E0",X"10",X"9F",X"AC",X"39",X"34",X"10",X"EC",X"A4",X"44",X"1F",X"01",X"86",
		X"00",X"A7",X"84",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"25",X"07",X"86",X"40",X"A7",X"84",
		X"35",X"10",X"39",X"86",X"04",X"A7",X"84",X"35",X"10",X"39",X"10",X"8E",X"AA",X"10",X"CE",X"B7",
		X"DC",X"A6",X"26",X"26",X"0C",X"31",X"28",X"33",X"C8",X"10",X"10",X"8C",X"AA",X"50",X"26",X"F1",
		X"39",X"6A",X"C4",X"26",X"66",X"A6",X"41",X"26",X"2D",X"BD",X"D0",X"3A",X"A6",X"47",X"27",X"10",
		X"6F",X"48",X"A6",X"42",X"8B",X"40",X"2B",X"04",X"86",X"F8",X"20",X"0A",X"86",X"08",X"20",X"06",
		X"86",X"08",X"54",X"24",X"01",X"40",X"A7",X"43",X"C4",X"03",X"CB",X"02",X"E7",X"44",X"86",X"01",
		X"94",X"04",X"8B",X"02",X"A7",X"41",X"E6",X"44",X"27",X"0C",X"6A",X"44",X"A7",X"C4",X"A6",X"42",
		X"AB",X"43",X"A7",X"42",X"20",X"25",X"BD",X"D0",X"3A",X"A6",X"47",X"27",X"16",X"C4",X"1F",X"CB",
		X"30",X"A6",X"4A",X"84",X"07",X"40",X"8B",X"07",X"48",X"48",X"48",X"A7",X"E2",X"EB",X"E0",X"E7",
		X"47",X"20",X"04",X"C4",X"1F",X"CB",X"30",X"E7",X"C4",X"6F",X"41",X"86",X"01",X"97",X"00",X"B7",
		X"D0",X"00",X"A6",X"4A",X"E6",X"42",X"1F",X"01",X"AE",X"84",X"9F",X"9E",X"DB",X"09",X"1F",X"01",
		X"AE",X"84",X"4F",X"97",X"00",X"B7",X"D0",X"00",X"1F",X"10",X"AB",X"A4",X"EB",X"21",X"ED",X"22",
		X"A1",X"46",X"22",X"5D",X"A6",X"47",X"26",X"55",X"C1",X"A5",X"22",X"2C",X"C1",X"55",X"23",X"04",
		X"D6",X"04",X"2B",X"24",X"CC",X"08",X"80",X"E7",X"47",X"E0",X"42",X"54",X"54",X"54",X"ED",X"43",
		X"E7",X"48",X"E7",X"49",X"C5",X"08",X"26",X"08",X"CC",X"02",X"02",X"ED",X"C4",X"7E",X"F5",X"53",
		X"CC",X"01",X"01",X"ED",X"C4",X"7E",X"F5",X"53",X"86",X"F8",X"A7",X"47",X"E6",X"42",X"54",X"54",
		X"54",X"ED",X"43",X"E7",X"48",X"E7",X"49",X"C5",X"08",X"26",X"0A",X"CC",X"02",X"02",X"ED",X"C4",
		X"6C",X"47",X"7E",X"F5",X"53",X"CC",X"01",X"01",X"ED",X"C4",X"7E",X"F5",X"53",X"A6",X"A4",X"20",
		X"02",X"6F",X"47",X"81",X"E8",X"23",X"3A",X"C1",X"F0",X"24",X"4A",X"C1",X"08",X"23",X"6D",X"E6",
		X"47",X"10",X"2B",X"00",X"8E",X"E6",X"42",X"2E",X"26",X"81",X"F4",X"25",X"0C",X"CC",X"40",X"00",
		X"ED",X"42",X"86",X"08",X"ED",X"C4",X"7E",X"F5",X"53",X"A6",X"45",X"26",X"72",X"6F",X"43",X"CB",
		X"40",X"2A",X"66",X"86",X"F8",X"A7",X"45",X"AB",X"42",X"A7",X"42",X"6F",X"43",X"20",X"64",X"E6",
		X"21",X"C1",X"1C",X"23",X"2F",X"C1",X"D8",X"22",X"04",X"6F",X"45",X"20",X"56",X"A6",X"47",X"2B",
		X"52",X"C1",X"F0",X"25",X"0B",X"CC",X"00",X"00",X"ED",X"42",X"86",X"08",X"ED",X"C4",X"20",X"43",
		X"E6",X"42",X"6F",X"48",X"CB",X"40",X"1C",X"FD",X"2E",X"DF",X"A6",X"45",X"26",X"31",X"A6",X"42",
		X"2E",X"C1",X"20",X"25",X"A6",X"47",X"2B",X"2B",X"C1",X"08",X"22",X"0B",X"CC",X"80",X"00",X"ED",
		X"42",X"86",X"08",X"ED",X"C4",X"20",X"1C",X"E6",X"42",X"6F",X"48",X"CB",X"C0",X"1C",X"FD",X"2E",
		X"B8",X"A6",X"45",X"26",X"0A",X"A6",X"42",X"2F",X"9A",X"86",X"08",X"A7",X"45",X"6F",X"43",X"AB",
		X"42",X"A7",X"42",X"9E",X"A4",X"10",X"AF",X"81",X"9F",X"A4",X"A6",X"48",X"10",X"27",X"FE",X"55",
		X"EC",X"26",X"10",X"83",X"EB",X"A2",X"10",X"26",X"FE",X"4B",X"A6",X"49",X"27",X"05",X"6A",X"49",
		X"7E",X"F3",X"B5",X"86",X"0E",X"A7",X"49",X"8E",X"B6",X"6C",X"A6",X"06",X"27",X"0A",X"30",X"08",
		X"8C",X"B7",X"6C",X"26",X"F5",X"7E",X"F3",X"B5",X"CC",X"ED",X"80",X"ED",X"06",X"EC",X"A4",X"CB",
		X"03",X"ED",X"84",X"86",X"FE",X"D6",X"9F",X"2B",X"04",X"C6",X"02",X"20",X"02",X"C6",X"FE",X"ED",
		X"04",X"AF",X"9F",X"A0",X"AA",X"9E",X"AA",X"30",X"02",X"9F",X"AA",X"7E",X"F3",X"B5",X"10",X"8E",
		X"A5",X"B8",X"CE",X"A5",X"B8",X"AE",X"A1",X"27",X"4A",X"EC",X"84",X"AB",X"04",X"EB",X"05",X"ED",
		X"02",X"81",X"45",X"23",X"0C",X"81",X"F8",X"24",X"08",X"C1",X"08",X"23",X"04",X"C1",X"F8",X"25",
		X"0E",X"6F",X"06",X"EC",X"84",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",X"84",X"20",X"0C",X"AF",
		X"9F",X"A0",X"A4",X"AF",X"C1",X"9E",X"A4",X"30",X"02",X"9F",X"A4",X"AE",X"A1",X"26",X"CA",X"CC",
		X"00",X"00",X"DF",X"A8",X"10",X"9F",X"9C",X"11",X"93",X"9C",X"27",X"07",X"ED",X"C1",X"11",X"93",
		X"9C",X"26",X"F9",X"39",X"96",X"63",X"26",X"04",X"96",X"78",X"27",X"01",X"39",X"96",X"7A",X"9B",
		X"7E",X"91",X"21",X"24",X"F7",X"96",X"6F",X"26",X"F3",X"96",X"84",X"26",X"15",X"C6",X"44",X"8E",
		X"F6",X"57",X"10",X"8E",X"8A",X"AC",X"BD",X"D0",X"47",X"C6",X"CC",X"10",X"8E",X"84",X"AC",X"BD",
		X"D0",X"47",X"86",X"70",X"97",X"8B",X"97",X"86",X"CC",X"00",X"10",X"DD",X"AE",X"8E",X"B7",X"DC",
		X"10",X"8E",X"F6",X"6A",X"CE",X"AA",X"10",X"A6",X"46",X"27",X"07",X"30",X"88",X"10",X"33",X"48",
		X"20",X"F5",X"0A",X"78",X"7E",X"D2",X"33",X"43",X"41",X"55",X"54",X"49",X"4F",X"4E",X"40",X"40",
		X"00",X"53",X"43",X"4F",X"55",X"54",X"40",X"40",X"40",X"00",X"F6",X"75",X"1F",X"D0",X"00",X"B0",
		X"00",X"02",X"7E",X"F7",X"F6",X"34",X"70",X"EC",X"A4",X"44",X"1F",X"01",X"CC",X"00",X"00",X"ED",
		X"84",X"ED",X"02",X"ED",X"04",X"ED",X"06",X"A7",X"08",X"30",X"89",X"01",X"00",X"ED",X"84",X"ED",
		X"02",X"ED",X"04",X"ED",X"06",X"A7",X"08",X"30",X"89",X"01",X"00",X"ED",X"84",X"ED",X"02",X"ED",
		X"04",X"ED",X"06",X"A7",X"08",X"30",X"89",X"01",X"00",X"ED",X"84",X"ED",X"02",X"ED",X"04",X"ED",
		X"06",X"A7",X"08",X"CE",X"F6",X"F6",X"EC",X"22",X"ED",X"A4",X"44",X"1F",X"01",X"25",X"03",X"CE",
		X"F7",X"00",X"96",X"AE",X"81",X"08",X"27",X"0A",X"0A",X"AF",X"26",X"06",X"C6",X"10",X"8B",X"02",
		X"DD",X"AE",X"EE",X"C6",X"10",X"AE",X"C1",X"EC",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"02",X"EC",
		X"C1",X"ED",X"04",X"EC",X"C1",X"ED",X"06",X"A6",X"C0",X"A7",X"08",X"30",X"89",X"01",X"00",X"31",
		X"3F",X"26",X"E4",X"35",X"70",X"39",X"F7",X"0A",X"F7",X"15",X"F7",X"29",X"F7",X"46",X"F7",X"63",
		X"F7",X"89",X"F7",X"94",X"F7",X"9F",X"F7",X"B3",X"F7",X"D0",X"00",X"01",X"04",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"0D",X"0E",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"40",X"44",X"40",X"44",X"40",X"00",X"00",X"00",X"00",X"C0",X"40",X"00",
		X"40",X"D0",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"0D",X"0E",X"0D",X"00",X"00",X"00",
		X"00",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"00",X"00",X"0C",X"44",X"0E",X"C0",X"0F",X"44",
		X"0D",X"00",X"00",X"00",X"04",X"00",X"00",X"0D",X"0E",X"0F",X"0E",X"0D",X"00",X"00",X"A4",X"A4",
		X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"00",X"44",X"00",X"40",X"4C",X"40",X"00",X"44",X"00",
		X"0C",X"44",X"0E",X"00",X"00",X"00",X"0F",X"44",X"0D",X"00",X"01",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"44",X"40",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"D4",X"E4",X"D4",X"04",X"00",X"00",X"00",X"00",X"0C",X"44",X"00",X"44",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0A",X"0A",X"DA",X"EA",X"DA",X"0A",X"0A",X"00",X"00",X"40",X"44",
		X"40",X"4C",X"40",X"44",X"40",X"00",X"00",X"C0",X"40",X"E0",X"00",X"F0",X"40",X"D0",X"00",X"00",
		X"00",X"04",X"0A",X"0A",X"DA",X"EA",X"FA",X"EA",X"DA",X"0A",X"0A",X"40",X"44",X"40",X"44",X"44",
		X"44",X"40",X"44",X"40",X"00",X"44",X"00",X"00",X"C0",X"00",X"00",X"44",X"00",X"C0",X"40",X"E0",
		X"00",X"00",X"00",X"F0",X"40",X"D0",X"34",X"10",X"96",X"84",X"26",X"07",X"34",X"20",X"BD",X"FB",
		X"D8",X"35",X"20",X"CC",X"3F",X"00",X"D7",X"86",X"D7",X"8B",X"94",X"04",X"8B",X"30",X"97",X"78",
		X"CC",X"06",X"18",X"BD",X"D7",X"16",X"8E",X"AA",X"50",X"CE",X"F8",X"75",X"A6",X"06",X"27",X"04",
		X"30",X"08",X"20",X"F8",X"EC",X"A4",X"E3",X"C1",X"ED",X"84",X"EC",X"C1",X"ED",X"04",X"CC",X"EC",
		X"E9",X"ED",X"06",X"AF",X"9F",X"A0",X"A8",X"DC",X"A8",X"C3",X"00",X"02",X"DD",X"A8",X"11",X"83",
		X"F8",X"B5",X"26",X"D8",X"EC",X"A4",X"44",X"1F",X"01",X"4F",X"A7",X"08",X"A7",X"89",X"01",X"08",
		X"A7",X"89",X"02",X"08",X"A7",X"89",X"03",X"08",X"0C",X"6C",X"8E",X"A0",X"19",X"96",X"0D",X"27",
		X"03",X"8E",X"A0",X"1C",X"A6",X"01",X"8B",X"01",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",X"19",
		X"A7",X"84",X"35",X"10",X"39",X"00",X"00",X"00",X"FB",X"00",X"02",X"FE",X"FC",X"00",X"04",X"FD",
		X"FD",X"00",X"06",X"FC",X"FE",X"02",X"00",X"FB",X"00",X"02",X"02",X"FC",X"02",X"02",X"04",X"FD",
		X"03",X"02",X"06",X"FE",X"04",X"04",X"00",X"00",X"05",X"04",X"02",X"02",X"04",X"04",X"04",X"03",
		X"03",X"04",X"06",X"04",X"02",X"06",X"00",X"05",X"00",X"06",X"02",X"04",X"FE",X"06",X"04",X"03",
		X"FD",X"06",X"06",X"02",X"FC",X"00",X"00",X"FD",X"00",X"00",X"03",X"FE",X"02",X"00",X"FD",X"FE",
		X"FE",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"02",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"00",X"46",X"49",X"47",X"48",X"54",X"45",X"52",X"53",X"00",X"C6",X"AA",
		X"8E",X"F8",X"D5",X"10",X"8E",X"8A",X"14",X"BD",X"D0",X"47",X"34",X"20",X"C6",X"AA",X"10",X"8E",
		X"84",X"2C",X"96",X"20",X"9B",X"7A",X"0D",X"8B",X"27",X"01",X"4A",X"BD",X"FD",X"38",X"35",X"20",
		X"39",X"0C",X"0A",X"8E",X"C0",X"00",X"CC",X"00",X"00",X"ED",X"81",X"8C",X"C0",X"10",X"26",X"F9",
		X"1F",X"40",X"C4",X"FE",X"1F",X"01",X"CC",X"00",X"00",X"A7",X"82",X"8C",X"A0",X"6C",X"26",X"F9",
		X"8E",X"A0",X"00",X"ED",X"83",X"8C",X"00",X"00",X"26",X"F9",X"10",X"8E",X"80",X"00",X"CC",X"01",
		X"00",X"BD",X"D0",X"19",X"10",X"8E",X"81",X"58",X"CC",X"11",X"1E",X"BD",X"D0",X"1F",X"10",X"8E",
		X"81",X"A8",X"CC",X"11",X"1E",X"BD",X"D0",X"1F",X"CC",X"80",X"80",X"FD",X"A9",X"B8",X"10",X"8E",
		X"1C",X"14",X"CC",X"22",X"D8",X"BD",X"D0",X"19",X"10",X"8E",X"1B",X"14",X"CC",X"44",X"D8",X"BD",
		X"D0",X"19",X"10",X"8E",X"1A",X"14",X"CC",X"84",X"D8",X"BD",X"D0",X"19",X"86",X"01",X"D6",X"00",
		X"97",X"00",X"B7",X"D0",X"00",X"D7",X"01",X"BD",X"D7",X"49",X"96",X"01",X"97",X"00",X"B7",X"D0",
		X"00",X"BD",X"FE",X"E5",X"0F",X"64",X"00",X"0A",X"96",X"0A",X"26",X"FC",X"8E",X"A5",X"B8",X"9F",
		X"A8",X"8E",X"A5",X"76",X"9F",X"AA",X"8E",X"BE",X"38",X"9F",X"AC",X"8E",X"A7",X"B8",X"9F",X"9A",
		X"CC",X"02",X"C0",X"97",X"73",X"D7",X"7B",X"BD",X"FB",X"D8",X"BD",X"F8",X"DE",X"BD",X"FD",X"5F",
		X"BD",X"D0",X"3A",X"C4",X"3F",X"CB",X"30",X"D7",X"78",X"96",X"11",X"27",X"13",X"C6",X"88",X"8E",
		X"D6",X"D5",X"10",X"8E",X"78",X"60",X"BD",X"D0",X"47",X"96",X"0D",X"8B",X"31",X"BD",X"EF",X"3E",
		X"4F",X"5F",X"DD",X"59",X"97",X"5B",X"D6",X"03",X"86",X"40",X"3D",X"8B",X"40",X"90",X"1F",X"90",
		X"1F",X"B7",X"BF",X"AA",X"39",X"96",X"0B",X"2B",X"0C",X"85",X"40",X"26",X"0D",X"85",X"20",X"26",
		X"05",X"85",X"10",X"26",X"11",X"39",X"96",X"75",X"26",X"FB",X"96",X"74",X"26",X"F7",X"CC",X"C0",
		X"10",X"D7",X"0B",X"97",X"10",X"39",X"96",X"10",X"27",X"03",X"0A",X"10",X"39",X"86",X"80",X"97",
		X"0B",X"0A",X"1F",X"0F",X"20",X"96",X"37",X"2F",X"17",X"00",X"37",X"BD",X"F9",X"01",X"C6",X"99",
		X"8E",X"FE",X"86",X"10",X"8E",X"60",X"58",X"BD",X"D0",X"47",X"96",X"0E",X"27",X"44",X"20",X"2F",
		X"96",X"0E",X"27",X"14",X"8E",X"A0",X"1F",X"10",X"8E",X"A0",X"39",X"EC",X"84",X"EE",X"A4",X"ED",
		X"A1",X"EF",X"81",X"8C",X"A0",X"39",X"26",X"F3",X"96",X"0D",X"91",X"0E",X"10",X"27",X"DB",X"AC",
		X"0C",X"0D",X"BD",X"F9",X"01",X"9E",X"13",X"EC",X"84",X"10",X"AE",X"02",X"BD",X"D0",X"19",X"96",
		X"0D",X"88",X"01",X"97",X"0D",X"86",X"33",X"97",X"0F",X"BD",X"EB",X"17",X"96",X"0D",X"88",X"01",
		X"97",X"0D",X"CC",X"99",X"14",X"97",X"0F",X"D7",X"6F",X"7E",X"EB",X"17",X"40",X"40",X"47",X"41",
		X"4D",X"45",X"40",X"40",X"00",X"40",X"40",X"4F",X"56",X"45",X"52",X"40",X"40",X"00",X"53",X"51",
		X"55",X"41",X"44",X"52",X"4F",X"4E",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"96",X"20",X"9A",X"84",X"9A",X"8D",X"9A",X"8C",X"9A",X"7A",X"9A",X"63",X"27",X"01",X"39",X"0F",
		X"85",X"0F",X"8F",X"0F",X"90",X"BD",X"F9",X"D6",X"96",X"11",X"26",X"04",X"C6",X"02",X"20",X"09",
		X"D6",X"1F",X"5C",X"C1",X"63",X"23",X"02",X"C6",X"63",X"D7",X"1F",X"5A",X"C1",X"0F",X"23",X"02",
		X"C6",X"0F",X"58",X"58",X"58",X"8E",X"FD",X"78",X"10",X"8E",X"A0",X"20",X"3A",X"3A",X"86",X"07",
		X"EE",X"81",X"EF",X"A1",X"4A",X"26",X"F9",X"A6",X"84",X"A7",X"A4",X"8E",X"A5",X"76",X"9F",X"AA",
		X"10",X"AE",X"84",X"27",X"10",X"EC",X"A4",X"44",X"1F",X"03",X"CC",X"00",X"00",X"A7",X"C4",X"A7",
		X"26",X"ED",X"81",X"20",X"EB",X"96",X"03",X"84",X"3F",X"8B",X"30",X"97",X"78",X"BD",X"FB",X"D8",
		X"C6",X"22",X"8E",X"00",X"02",X"10",X"8E",X"84",X"14",X"CE",X"A0",X"22",X"0F",X"6D",X"BD",X"EB",
		X"32",X"8E",X"FE",X"78",X"BD",X"D0",X"47",X"0C",X"8E",X"D6",X"11",X"26",X"01",X"39",X"D6",X"6F",
		X"26",X"FB",X"86",X"80",X"97",X"7B",X"8E",X"FE",X"91",X"D6",X"89",X"C1",X"09",X"22",X"02",X"0C",
		X"89",X"58",X"3A",X"D6",X"7C",X"C5",X"80",X"26",X"11",X"96",X"82",X"27",X"04",X"A6",X"84",X"20",
		X"02",X"A6",X"01",X"10",X"8E",X"20",X"21",X"BD",X"FC",X"37",X"C5",X"40",X"26",X"09",X"A6",X"01",
		X"10",X"8E",X"20",X"43",X"BD",X"FC",X"37",X"C5",X"20",X"26",X"13",X"96",X"87",X"85",X"04",X"27",
		X"04",X"A6",X"84",X"20",X"02",X"A6",X"01",X"10",X"8E",X"20",X"62",X"BD",X"FC",X"37",X"C5",X"10",
		X"26",X"09",X"A6",X"01",X"10",X"8E",X"20",X"78",X"BD",X"FC",X"37",X"C5",X"08",X"26",X"13",X"96",
		X"87",X"85",X"02",X"27",X"04",X"A6",X"84",X"20",X"02",X"A6",X"01",X"10",X"8E",X"20",X"8E",X"BD",
		X"FC",X"37",X"C5",X"04",X"26",X"09",X"A6",X"01",X"10",X"8E",X"20",X"AF",X"BD",X"FC",X"37",X"C5",
		X"02",X"26",X"09",X"A6",X"01",X"10",X"8E",X"20",X"C5",X"BD",X"FC",X"37",X"C5",X"01",X"26",X"13",
		X"96",X"87",X"85",X"01",X"27",X"04",X"A6",X"84",X"20",X"02",X"A6",X"01",X"10",X"8E",X"20",X"DB",
		X"BD",X"FC",X"37",X"86",X"01",X"97",X"88",X"39",X"CC",X"88",X"33",X"DD",X"9C",X"C6",X"66",X"8E",
		X"FA",X"8E",X"10",X"8E",X"8A",X"AC",X"BD",X"D0",X"47",X"10",X"8E",X"84",X"AC",X"BD",X"D0",X"47",
		X"DC",X"9C",X"0D",X"0D",X"27",X"02",X"1E",X"89",X"DD",X"9C",X"96",X"1F",X"26",X"01",X"4C",X"D6",
		X"9C",X"0D",X"0E",X"27",X"2A",X"10",X"8E",X"84",X"B4",X"0D",X"0D",X"27",X"06",X"D6",X"9D",X"10",
		X"8E",X"84",X"D4",X"BD",X"FD",X"38",X"96",X"39",X"26",X"01",X"4C",X"D6",X"9D",X"10",X"8E",X"84",
		X"D4",X"0D",X"0D",X"27",X"06",X"D6",X"9C",X"10",X"8E",X"84",X"B4",X"BD",X"FD",X"38",X"39",X"10",
		X"8E",X"84",X"C4",X"BD",X"FD",X"38",X"39",X"34",X"06",X"0D",X"7B",X"2A",X"17",X"0C",X"6C",X"CE",
		X"A0",X"19",X"D6",X"0D",X"27",X"03",X"CE",X"A0",X"1C",X"AB",X"41",X"19",X"A7",X"41",X"A6",X"C4",
		X"89",X"00",X"A7",X"C4",X"A6",X"E4",X"44",X"44",X"84",X"3C",X"27",X"0C",X"31",X"3B",X"CE",X"FC",
		X"A8",X"33",X"C6",X"48",X"33",X"C6",X"8D",X"1D",X"A6",X"E0",X"84",X"0F",X"CE",X"FC",X"A8",X"48",
		X"48",X"33",X"C6",X"48",X"33",X"C6",X"8D",X"0D",X"CE",X"FC",X"A8",X"8D",X"08",X"CE",X"FC",X"A8",
		X"8D",X"03",X"35",X"04",X"39",X"EC",X"C1",X"ED",X"A4",X"EC",X"C1",X"ED",X"22",X"EC",X"C1",X"ED",
		X"A9",X"01",X"00",X"EC",X"C1",X"ED",X"A9",X"01",X"02",X"EC",X"C1",X"ED",X"A9",X"02",X"00",X"EC",
		X"C1",X"ED",X"A9",X"02",X"02",X"31",X"25",X"39",X"88",X"80",X"80",X"88",X"88",X"00",X"00",X"88",
		X"80",X"80",X"80",X"80",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"80",X"00",
		X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"88",
		X"00",X"80",X"80",X"88",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"88",X"88",X"80",X"80",X"88",
		X"80",X"00",X"00",X"80",X"80",X"80",X"80",X"88",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"88",X"80",X"80",X"88",X"88",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"08",X"00",X"00",
		X"00",X"00",X"80",X"08",X"80",X"80",X"80",X"80",X"88",X"80",X"80",X"88",X"88",X"80",X"80",X"88",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"88",X"88",X"80",X"80",X"88",X"80",X"80",X"80",X"80",
		X"96",X"86",X"26",X"01",X"39",X"0A",X"86",X"26",X"FB",X"86",X"32",X"97",X"86",X"96",X"20",X"81",
		X"62",X"24",X"F1",X"0C",X"20",X"7E",X"F8",X"EA",X"34",X"02",X"81",X"09",X"22",X"0F",X"86",X"40",
		X"BD",X"EF",X"3E",X"A6",X"E4",X"8A",X"30",X"BD",X"EF",X"3E",X"35",X"02",X"39",X"6F",X"E2",X"6C",
		X"E4",X"80",X"0A",X"81",X"09",X"22",X"F8",X"A7",X"61",X"A6",X"E0",X"8A",X"30",X"20",X"E1",X"CC",
		X"31",X"88",X"10",X"8E",X"8A",X"60",X"BD",X"EF",X"3E",X"96",X"0E",X"27",X"0A",X"CC",X"32",X"88",
		X"10",X"8E",X"84",X"60",X"BD",X"EF",X"3E",X"39",X"1E",X"02",X"00",X"25",X"00",X"15",X"05",X"00",
		X"01",X"00",X"C0",X"6E",X"86",X"00",X"10",X"00",X"1E",X"03",X"00",X"50",X"00",X"11",X"07",X"50",
		X"01",X"00",X"C0",X"6E",X"86",X"00",X"10",X"00",X"1E",X"03",X"00",X"75",X"00",X"11",X"10",X"00",
		X"02",X"50",X"C0",X"6E",X"86",X"00",X"10",X"00",X"1E",X"03",X"01",X"00",X"00",X"11",X"10",X"00",
		X"02",X"50",X"C0",X"6E",X"86",X"00",X"14",X"00",X"1E",X"03",X"01",X"00",X"00",X"0E",X"20",X"00",
		X"05",X"00",X"C1",X"6E",X"86",X"00",X"0C",X"00",X"1E",X"03",X"01",X"25",X"00",X"07",X"20",X"00",
		X"05",X"00",X"C2",X"6E",X"86",X"00",X"1A",X"00",X"1E",X"03",X"01",X"25",X"15",X"07",X"20",X"00",
		X"05",X"00",X"C1",X"6E",X"86",X"14",X"08",X"00",X"1E",X"03",X"01",X"50",X"15",X"07",X"25",X"00",
		X"07",X"50",X"C1",X"6E",X"86",X"00",X"08",X"00",X"1E",X"03",X"01",X"50",X"15",X"07",X"25",X"00",
		X"07",X"50",X"C2",X"6E",X"86",X"00",X"0F",X"00",X"1E",X"03",X"01",X"75",X"15",X"07",X"30",X"00",
		X"07",X"50",X"C1",X"6E",X"86",X"1C",X"12",X"00",X"1E",X"03",X"01",X"75",X"15",X"07",X"30",X"00",
		X"07",X"50",X"C2",X"6E",X"86",X"13",X"07",X"00",X"1E",X"03",X"02",X"00",X"15",X"07",X"40",X"00",
		X"10",X"00",X"C2",X"6E",X"86",X"00",X"18",X"00",X"1E",X"03",X"02",X"00",X"15",X"07",X"40",X"00",
		X"10",X"00",X"C2",X"6E",X"86",X"16",X"0B",X"00",X"1E",X"03",X"02",X"25",X"15",X"07",X"40",X"00",
		X"10",X"00",X"C2",X"6E",X"86",X"16",X"0B",X"00",X"1E",X"03",X"02",X"25",X"15",X"07",X"40",X"00",
		X"10",X"00",X"C2",X"6E",X"86",X"16",X"0B",X"00",X"1E",X"03",X"02",X"50",X"15",X"07",X"50",X"00",
		X"10",X"00",X"C3",X"6E",X"86",X"16",X"0B",X"00",X"40",X"50",X"54",X"53",X"00",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"00",X"42",X"4F",X"4E",X"55",X"53",X"40",X"54",X"55",X"52",X"4E",
		X"00",X"01",X"02",X"02",X"05",X"05",X"10",X"08",X"15",X"10",X"20",X"15",X"30",X"20",X"50",X"50",
		X"50",X"50",X"50",X"50",X"50",X"11",X"28",X"81",X"58",X"11",X"50",X"81",X"58",X"11",X"50",X"81",
		X"58",X"11",X"1B",X"81",X"58",X"11",X"36",X"81",X"58",X"11",X"50",X"81",X"58",X"11",X"50",X"81",
		X"58",X"96",X"61",X"27",X"03",X"7E",X"D0",X"7C",X"39",X"96",X"60",X"27",X"FB",X"0F",X"60",X"96",
		X"12",X"81",X"99",X"27",X"F3",X"8B",X"01",X"19",X"97",X"12",X"BD",X"FE",X"E5",X"CC",X"10",X"04",
		X"BD",X"D7",X"16",X"4C",X"39",X"10",X"8E",X"0C",X"DE",X"96",X"12",X"44",X"44",X"44",X"44",X"8D",
		X"04",X"96",X"12",X"84",X"0F",X"CE",X"C7",X"00",X"C6",X"18",X"3D",X"33",X"CB",X"86",X"01",X"D6",
		X"00",X"97",X"00",X"B7",X"D0",X"00",X"D7",X"01",X"C6",X"04",X"86",X"55",X"A7",X"A0",X"8E",X"00",
		X"06",X"A6",X"C4",X"84",X"BB",X"A7",X"A4",X"A6",X"C0",X"43",X"84",X"55",X"AA",X"A4",X"A7",X"A0",
		X"30",X"1F",X"26",X"ED",X"86",X"55",X"A7",X"A4",X"31",X"A9",X"00",X"F9",X"5A",X"26",X"DB",X"31",
		X"A9",X"FC",X"08",X"96",X"01",X"97",X"00",X"B7",X"D0",X"00",X"39",X"7F",X"D0",X"00",X"96",X"63",
		X"26",X"05",X"96",X"6E",X"B7",X"C0",X"09",X"96",X"0A",X"2A",X"18",X"8E",X"FF",X"B7",X"96",X"64",
		X"AE",X"86",X"CE",X"C0",X"00",X"EC",X"81",X"ED",X"C1",X"11",X"83",X"C0",X"10",X"26",X"F6",X"0F",
		X"0A",X"20",X"22",X"26",X"20",X"0A",X"05",X"2A",X"1C",X"C6",X"07",X"D7",X"05",X"0C",X"06",X"D6",
		X"06",X"C4",X"03",X"8E",X"FF",X"BB",X"96",X"64",X"AE",X"86",X"3A",X"EC",X"84",X"FD",X"C0",X"0C",
		X"EC",X"02",X"FD",X"C0",X"0E",X"B6",X"CC",X"00",X"0F",X"07",X"CC",X"38",X"02",X"B7",X"C3",X"FC",
		X"DB",X"09",X"C4",X"07",X"D7",X"09",X"D6",X"70",X"5C",X"C4",X"07",X"D7",X"70",X"26",X"12",X"96",
		X"6F",X"26",X"0E",X"96",X"78",X"2F",X"02",X"0A",X"78",X"B6",X"BF",X"AA",X"27",X"03",X"7A",X"BF",
		X"AA",X"96",X"00",X"B7",X"D0",X"00",X"3B",X"FF",X"C7",X"FF",X"DF",X"FF",X"BF",X"FF",X"D7",X"E0",
		X"3F",X"38",X"00",X"E0",X"3F",X"38",X"00",X"00",X"E0",X"07",X"A4",X"3F",X"65",X"87",X"27",X"FF",
		X"FF",X"3A",X"13",X"E0",X"3F",X"38",X"00",X"07",X"FF",X"C0",X"3F",X"07",X"FF",X"C0",X"3F",X"00",
		X"3F",X"17",X"07",X"38",X"00",X"00",X"00",X"00",X"FF",X"C0",X"38",X"07",X"FF",X"C0",X"3F",X"84",
		X"D0",X"7C",X"D0",X"7C",X"D0",X"7C",X"D0",X"7C",X"FF",X"3B",X"D0",X"7C",X"D0",X"7C",X"D0",X"7C",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",
		X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"00",
		X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"00",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"00",
		X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",
		X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FE",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FE",X"FF",
		X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FE",X"01",
		X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",
		X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",
		X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"02",
		X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"02",
		X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",
		X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"02",X"01",
		X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"FF",X"01",X"00",X"02",X"FF",
		X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",
		X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FE",
		X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FF",X"FF",X"FE",X"00",X"FF",X"00",X"FE",
		X"00",X"FF",X"FF",X"FE",X"00",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",
		X"FF",X"00",X"FE",X"FF",X"FF",X"00",X"FE",X"FF",X"FF",X"00",X"FE",X"FF",X"FF",X"00",X"FE",X"00",
		X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"01",X"FF",X"00",X"FE",X"00",
		X"FF",X"00",X"FE",X"01",X"FF",X"00",X"FE",X"01",X"FE",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",
		X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"02",X"FF",X"01",X"00",X"01",X"FF",X"01",
		X"00",X"01",X"FF",X"02",X"00",X"01",X"FF",X"02",X"00",X"01",X"FF",X"02",X"00",X"01",X"00",X"02",
		X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"01",X"01",X"02",X"00",X"01",X"00",X"02",
		X"00",X"01",X"01",X"02",X"00",X"01",X"01",X"02",X"01",X"02",X"01",X"01",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"00",X"01",X"01",
		X"01",X"00",X"02",X"01",X"01",X"00",X"02",X"01",X"01",X"00",X"02",X"01",X"01",X"00",X"02",X"00",
		X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"01",X"00",X"02",X"FF",X"01",X"00",X"02",X"00",
		X"01",X"00",X"02",X"FF",X"01",X"00",X"02",X"FF",X"02",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",
		X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FE",X"01",X"FF",X"00",X"FF",X"01",X"FF",
		X"00",X"FF",X"01",X"FE",X"00",X"FF",X"01",X"FE",X"00",X"FF",X"01",X"FE",X"00",X"FF",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"FF",X"FE",X"00",X"FF",X"FF",X"FE",X"00",X"FE",
		X"FF",X"FE",X"00",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"FE",X"FF",X"FF",X"00",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"00",X"FE",X"FF",X"FE",X"00",
		X"FE",X"00",X"FE",X"00",X"FF",X"00",X"FE",X"00",X"FE",X"01",X"FF",X"00",X"FE",X"01",X"FE",X"00",
		X"FE",X"01",X"FF",X"00",X"FE",X"01",X"FE",X"01",X"FF",X"01",X"FE",X"01",X"FF",X"01",X"FE",X"01",
		X"FF",X"01",X"FF",X"01",X"FE",X"02",X"FF",X"01",X"FF",X"01",X"FF",X"02",X"FF",X"01",X"FF",X"02",
		X"FF",X"02",X"00",X"01",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"00",X"01",X"FF",X"02",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"01",X"02",X"00",X"01",X"01",X"02",X"00",X"02",
		X"01",X"02",X"00",X"01",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"02",X"01",
		X"02",X"01",X"01",X"00",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"00",X"02",X"01",X"02",X"00",
		X"02",X"00",X"02",X"00",X"01",X"00",X"02",X"00",X"02",X"FF",X"01",X"00",X"02",X"FF",X"02",X"00",
		X"02",X"FF",X"01",X"00",X"02",X"FF",X"02",X"FF",X"01",X"FF",X"02",X"FF",X"01",X"FF",X"02",X"FF",
		X"01",X"FF",X"01",X"FF",X"02",X"FE",X"01",X"FF",X"01",X"FF",X"01",X"FE",X"01",X"FF",X"01",X"FE",
		X"01",X"FE",X"00",X"FF",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"00",X"FF",X"01",X"FE",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"FF",X"FE",X"00",X"FE",X"FF",X"FE",X"00",X"FE",
		X"FF",X"FE",X"00",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"FE",X"FF",X"FE",X"00",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"00",X"FE",X"FF",X"FE",X"00",
		X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FE",X"00",
		X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FF",X"01",X"FE",X"01",
		X"FF",X"01",X"FE",X"02",X"FF",X"01",X"FE",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"01",X"FF",X"02",
		X"FF",X"02",X"00",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"00",X"02",X"FF",X"02",X"00",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"00",X"02",
		X"01",X"02",X"00",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"01",X"01",X"02",
		X"01",X"01",X"02",X"02",X"01",X"01",X"02",X"02",X"02",X"01",X"02",X"01",X"01",X"01",X"02",X"01",
		X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"00",
		X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"FF",X"02",X"00",X"02",X"FF",X"02",X"00",
		X"02",X"FF",X"02",X"00",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"01",X"FF",X"02",X"FF",
		X"01",X"FF",X"02",X"FE",X"01",X"FF",X"02",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FF",X"01",X"FE",
		X"01",X"FE",X"00",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FE",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"00",X"FD",X"00",X"FE",X"FF",X"FE",X"00",X"FE",X"FF",X"FE",X"00",X"FD",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FF",X"FF",
		X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"00",X"FE",X"FF",X"FD",X"00",
		X"FE",X"00",X"FE",X"00",X"FD",X"00",X"FE",X"00",X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FD",X"00",
		X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"02",X"FE",X"01",X"FE",X"02",X"FF",X"01",
		X"FE",X"02",X"FF",X"01",X"FE",X"02",X"FF",X"01",X"FE",X"02",X"FF",X"02",X"FE",X"02",X"FF",X"01",
		X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"00",X"02",X"FF",X"02",X"00",X"03",
		X"00",X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"01",X"02",X"00",X"02",X"01",X"02",X"00",X"03",
		X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"01",X"01",
		X"02",X"02",X"01",X"01",X"02",X"02",X"01",X"01",X"02",X"02",X"02",X"01",X"02",X"02",X"01",X"01",
		X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"01",X"02",X"00",X"02",X"01",X"03",X"00",
		X"02",X"00",X"02",X"00",X"03",X"00",X"02",X"00",X"02",X"FF",X"02",X"00",X"02",X"FF",X"03",X"00",
		X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FE",X"02",X"FF",X"02",X"FE",X"01",X"FF",
		X"02",X"FE",X"01",X"FF",X"02",X"FE",X"01",X"FF",X"02",X"FE",X"01",X"FE",X"02",X"FE",X"01",X"FF",
		X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"00",X"FE",X"01",X"FE",X"00",X"FD",
		X"00",X"FD",X"00",X"FD",X"00",X"FE",X"00",X"FD",X"FF",X"FD",X"00",X"FD",X"FF",X"FD",X"00",X"FE",
		X"FF",X"FD",X"FF",X"FE",X"FF",X"FD",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FD",X"FF",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FD",X"FE",X"FE",X"FF",
		X"FD",X"FF",X"FE",X"FF",X"FD",X"FF",X"FE",X"FF",X"FD",X"FF",X"FD",X"00",X"FD",X"FF",X"FE",X"00",
		X"FD",X"00",X"FD",X"00",X"FE",X"00",X"FD",X"00",X"FD",X"01",X"FD",X"00",X"FD",X"01",X"FE",X"01",
		X"FD",X"01",X"FE",X"02",X"FD",X"01",X"FE",X"02",X"FE",X"02",X"FE",X"01",X"FD",X"02",X"FE",X"01",
		X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FF",X"02",X"FE",X"03",X"FF",X"02",
		X"FF",X"03",X"FF",X"02",X"FF",X"03",X"FF",X"02",X"FF",X"03",X"00",X"03",X"FF",X"03",X"00",X"02",
		X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"01",X"03",X"00",X"03",X"01",X"03",X"00",X"02",
		X"01",X"03",X"01",X"02",X"01",X"03",X"01",X"02",X"02",X"02",X"01",X"02",X"02",X"03",X"01",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"03",X"02",X"02",X"01",
		X"03",X"01",X"02",X"01",X"03",X"01",X"02",X"01",X"03",X"01",X"03",X"00",X"03",X"01",X"02",X"00",
		X"03",X"00",X"03",X"00",X"02",X"00",X"03",X"00",X"03",X"FF",X"03",X"00",X"03",X"FF",X"02",X"00",
		X"03",X"FF",X"02",X"FF",X"03",X"FF",X"02",X"FF",X"02",X"FE",X"02",X"FF",X"03",X"FE",X"02",X"FF",
		X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"01",X"FE",X"02",X"FD",X"01",X"FE",
		X"01",X"FD",X"01",X"FE",X"01",X"FD",X"01",X"FE",X"01",X"FD",X"00",X"FD",X"01",X"FD",X"00",X"FE",
		X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"F0",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"FF",X"0F",X"00",X"F0",X"0F",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"00",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",
		X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"0F",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"FF",X"0F",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"8E",X"C8",X"16",X"10",X"AE",X"81",X"2B",X"07",X"EC",X"81",X"BD",X"D0",X"1F",X"20",X"F4",X"10",
		X"AE",X"81",X"EC",X"81",X"BD",X"D0",X"19",X"EC",X"81",X"27",X"0A",X"10",X"AE",X"81",X"A7",X"A4",
		X"5A",X"26",X"F8",X"20",X"F2",X"39",X"0E",X"24",X"33",X"08",X"0E",X"26",X"33",X"08",X"0F",X"2A",
		X"88",X"05",X"0F",X"2B",X"88",X"05",X"0F",X"2C",X"88",X"05",X"FF",X"FF",X"0E",X"27",X"22",X"09",
		X"03",X"06",X"15",X"25",X"12",X"25",X"0F",X"25",X"13",X"27",X"13",X"28",X"13",X"29",X"30",X"02",
		X"14",X"25",X"11",X"25",X"11",X"0A",X"0F",X"27",X"0F",X"28",X"0F",X"29",X"0F",X"2D",X"0F",X"2E",
		X"10",X"29",X"10",X"2D",X"14",X"2A",X"14",X"2B",X"14",X"2C",X"10",X"06",X"10",X"27",X"10",X"28",
		X"10",X"2E",X"11",X"29",X"11",X"2D",X"15",X"2B",X"18",X"02",X"13",X"2B",X"12",X"2B",X"00",X"00",
		X"8E",X"CE",X"68",X"10",X"AE",X"81",X"27",X"07",X"EC",X"81",X"BD",X"D0",X"19",X"20",X"F4",X"39",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",
		X"00",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0F",X"FF",X"0F",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0F",X"0F",X"FF",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"F0",X"00",X"FF",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"F0",X"0F",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"FF",X"F0",X"00",X"00",X"F0",X"FF",
		X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"0F",X"F0",
		X"00",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"FF",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"FF",X"00",
		X"00",X"0F",X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"FF",X"0F",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"0F",X"0F",X"0F",X"0F",X"F0",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"0F",X"FF",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"F0",X"F0",X"0F",X"00",X"0F",X"F0",X"00",X"00",
		X"F0",X"0F",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"00",X"00",X"0F",X"00",X"FF",X"00",
		X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"0F",X"00",X"00",X"00",X"00",X"0F",X"F0",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"0F",X"F0",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"7E",X"01",X"FB",X"D0",X"07",X"24",X"7E",
		X"02",X"05",X"D0",X"0D",X"24",X"7E",X"02",X"FC",X"D0",X"07",X"24",X"7E",X"01",X"FD",X"D0",X"0D",
		X"24",X"7E",X"03",X"01",X"D0",X"01",X"24",X"7E",X"01",X"05",X"D0",X"04",X"24",X"7E",X"02",X"FE",
		X"D0",X"07",X"24",X"7E",X"01",X"03",X"D0",X"04",X"24",X"7E",X"01",X"01",X"D0",X"07",X"24",X"7E",
		X"01",X"FF",X"D0",X"04",X"24",X"7E",X"03",X"FF",X"D0",X"01",X"24",X"7E",X"02",X"00",X"D0",X"04",
		X"24",X"7E",X"03",X"03",X"D0",X"01",X"24",X"7E",X"03",X"FD",X"D0",X"04",X"24",X"7E",X"04",X"00",
		X"D0",X"01",X"24",X"7E",X"02",X"02",X"D0",X"04",X"00",X"00",X"1C",X"4A",X"01",X"FD",X"D0",X"01",
		X"1C",X"4A",X"01",X"FE",X"D0",X"0A",X"1C",X"4A",X"02",X"FE",X"D0",X"01",X"1C",X"4A",X"03",X"FE",
		X"D0",X"01",X"1C",X"4A",X"01",X"FF",X"D0",X"01",X"1C",X"4A",X"02",X"FF",X"D0",X"0A",X"1C",X"4A",
		X"03",X"FF",X"D0",X"01",X"1C",X"4A",X"02",X"00",X"D0",X"0A",X"1C",X"4A",X"04",X"00",X"D0",X"01",
		X"1C",X"4A",X"01",X"01",X"D0",X"01",X"1C",X"4A",X"02",X"01",X"D0",X"01",X"1C",X"4A",X"03",X"01",
		X"D0",X"0A",X"1C",X"4A",X"01",X"02",X"D0",X"0A",X"1C",X"4A",X"02",X"02",X"D0",X"01",X"1C",X"4A",
		X"03",X"02",X"D0",X"01",X"1C",X"4A",X"01",X"03",X"D0",X"01",X"1C",X"4A",X"02",X"03",X"D0",X"0A",
		X"1C",X"4A",X"03",X"03",X"D0",X"01",X"1C",X"4A",X"04",X"01",X"D0",X"01",X"1C",X"4A",X"04",X"02",
		X"D0",X"16",X"1C",X"4A",X"05",X"01",X"D0",X"16",X"1C",X"4A",X"05",X"FF",X"D0",X"0A",X"1C",X"4A",
		X"04",X"FF",X"D0",X"01",X"1C",X"4A",X"04",X"FE",X"D0",X"16",X"1C",X"4A",X"03",X"FD",X"D0",X"01",
		X"1C",X"4A",X"02",X"FD",X"D0",X"16",X"00",X"00",X"18",X"96",X"03",X"FE",X"D0",X"01",X"18",X"96",
		X"02",X"FF",X"D0",X"04",X"18",X"96",X"03",X"FF",X"D0",X"01",X"18",X"96",X"04",X"FF",X"D0",X"04",
		X"18",X"96",X"02",X"00",X"D0",X"01",X"18",X"96",X"04",X"00",X"D0",X"04",X"18",X"96",X"01",X"01",
		X"D0",X"01",X"18",X"96",X"02",X"01",X"D0",X"01",X"18",X"96",X"03",X"01",X"D0",X"04",X"18",X"96",
		X"04",X"01",X"D0",X"01",X"18",X"96",X"02",X"02",X"D0",X"01",X"18",X"96",X"03",X"02",X"D0",X"01",
		X"00",X"00",X"24",X"E0",X"03",X"FE",X"D0",X"01",X"24",X"E0",X"02",X"FF",X"D0",X"04",X"24",X"E0",
		X"03",X"FF",X"D0",X"01",X"24",X"E0",X"04",X"FF",X"D0",X"04",X"24",X"E0",X"02",X"00",X"D0",X"01",
		X"24",X"E0",X"04",X"00",X"D0",X"04",X"24",X"E0",X"01",X"01",X"D0",X"01",X"24",X"E0",X"02",X"01",
		X"D0",X"01",X"24",X"E0",X"03",X"01",X"D0",X"04",X"24",X"E0",X"04",X"01",X"D0",X"01",X"24",X"E0",
		X"02",X"02",X"D0",X"01",X"24",X"E0",X"03",X"02",X"D0",X"01",X"00",X"00",X"1E",X"6D",X"03",X"FE",
		X"D0",X"01",X"1E",X"6D",X"02",X"FF",X"D0",X"04",X"1E",X"6D",X"03",X"FF",X"D0",X"01",X"1E",X"6D",
		X"04",X"FF",X"D0",X"04",X"1E",X"6D",X"02",X"00",X"D0",X"01",X"1E",X"6D",X"04",X"00",X"D0",X"04",
		X"1E",X"6D",X"01",X"01",X"D0",X"01",X"1E",X"6D",X"02",X"01",X"D0",X"01",X"1E",X"6D",X"03",X"01",
		X"D0",X"04",X"1E",X"6D",X"04",X"01",X"D0",X"01",X"1E",X"6D",X"02",X"02",X"D0",X"01",X"1E",X"6D",
		X"03",X"02",X"D0",X"01",X"00",X"00",X"20",X"D1",X"03",X"FE",X"D0",X"04",X"20",X"D1",X"04",X"FE",
		X"D0",X"04",X"20",X"D1",X"05",X"FE",X"D0",X"0A",X"20",X"D1",X"02",X"FF",X"D0",X"04",X"20",X"D1",
		X"03",X"FF",X"D0",X"04",X"20",X"D1",X"04",X"FF",X"D0",X"01",X"20",X"D1",X"03",X"00",X"D0",X"07",
		X"20",X"D1",X"05",X"00",X"D0",X"07",X"20",X"D1",X"02",X"01",X"D0",X"0A",X"20",X"D1",X"03",X"01",
		X"D0",X"07",X"20",X"D1",X"04",X"01",X"D0",X"07",X"20",X"D1",X"05",X"01",X"D0",X"0A",X"20",X"D1",
		X"03",X"02",X"D0",X"01",X"20",X"D1",X"04",X"02",X"D0",X"01",X"20",X"D1",X"05",X"02",X"D0",X"0A",
		X"20",X"D1",X"05",X"FF",X"D0",X"01",X"00",X"00",X"20",X"C1",X"03",X"FD",X"D0",X"04",X"20",X"C1",
		X"04",X"FD",X"D0",X"0A",X"20",X"C1",X"02",X"FE",X"D0",X"04",X"20",X"C1",X"03",X"FE",X"D0",X"04",
		X"20",X"C1",X"04",X"FE",X"D0",X"04",X"20",X"C1",X"05",X"FE",X"D0",X"0A",X"20",X"C1",X"01",X"FF",
		X"D0",X"04",X"20",X"C1",X"02",X"FF",X"D0",X"0A",X"20",X"C1",X"03",X"FF",X"D0",X"04",X"20",X"C1",
		X"04",X"FF",X"D0",X"04",X"20",X"C1",X"05",X"FF",X"D0",X"04",X"20",X"C1",X"02",X"00",X"D0",X"0A",
		X"20",X"C1",X"05",X"00",X"D0",X"0A",X"20",X"C1",X"01",X"01",X"D0",X"16",X"20",X"C1",X"02",X"01",
		X"D0",X"04",X"20",X"C1",X"03",X"01",X"D0",X"16",X"20",X"C1",X"04",X"01",X"D0",X"0A",X"20",X"C1",
		X"05",X"01",X"D0",X"16",X"20",X"C1",X"02",X"02",X"D0",X"16",X"20",X"C1",X"03",X"02",X"D0",X"16",
		X"20",X"C1",X"04",X"02",X"D0",X"16",X"20",X"C1",X"05",X"02",X"D0",X"0A",X"20",X"C1",X"03",X"03",
		X"D0",X"16",X"20",X"C1",X"04",X"03",X"D0",X"16",X"00",X"00",X"1E",X"27",X"03",X"FF",X"D0",X"04",
		X"1E",X"27",X"04",X"FF",X"D0",X"04",X"1E",X"27",X"03",X"00",X"D0",X"04",X"1E",X"27",X"04",X"00",
		X"D0",X"04",X"1E",X"27",X"02",X"01",X"D0",X"04",X"1E",X"27",X"03",X"01",X"D0",X"04",X"1E",X"27",
		X"01",X"02",X"D0",X"04",X"1E",X"27",X"02",X"02",X"D0",X"04",X"1E",X"27",X"01",X"03",X"D0",X"16",
		X"1E",X"27",X"02",X"03",X"D0",X"16",X"1E",X"27",X"03",X"03",X"D0",X"16",X"1E",X"27",X"03",X"02",
		X"D0",X"16",X"1E",X"27",X"04",X"01",X"D0",X"04",X"1E",X"27",X"04",X"02",X"D0",X"04",X"1E",X"27",
		X"04",X"03",X"D0",X"04",X"00",X"00",X"24",X"2B",X"03",X"FF",X"D0",X"01",X"24",X"2B",X"04",X"FF",
		X"D0",X"0D",X"24",X"2B",X"03",X"00",X"D0",X"0D",X"24",X"2B",X"04",X"00",X"D0",X"01",X"24",X"2B",
		X"02",X"01",X"D0",X"0D",X"24",X"2B",X"03",X"01",X"D0",X"0D",X"24",X"2B",X"01",X"02",X"D0",X"01",
		X"24",X"2B",X"02",X"02",X"D0",X"0D",X"00",X"00",X"0B",X"45",X"50",X"10",X"0B",X"46",X"51",X"0B",
		X"0C",X"48",X"11",X"06",X"0D",X"47",X"11",X"08",X"0E",X"42",X"02",X"02",X"0E",X"44",X"12",X"0E",
		X"0E",X"52",X"02",X"02",X"0F",X"42",X"22",X"12",X"10",X"44",X"10",X"04",X"10",X"48",X"11",X"06",
		X"10",X"4E",X"10",X"04",X"11",X"48",X"10",X"06",X"10",X"49",X"14",X"04",X"0F",X"43",X"42",X"04",
		X"0F",X"49",X"42",X"04",X"0F",X"4F",X"42",X"04",X"0E",X"49",X"42",X"04",X"00",X"00",X"07",X"00",
		X"55",X"FF",X"08",X"00",X"55",X"FF",X"09",X"00",X"55",X"71",X"09",X"71",X"5B",X"2D",X"09",X"9E",
		X"55",X"14",X"09",X"B2",X"5B",X"07",X"09",X"B9",X"55",X"46",X"0A",X"00",X"55",X"5D",X"0A",X"5D",
		X"BB",X"63",X"0A",X"C0",X"55",X"3F",X"0B",X"00",X"55",X"45",X"0B",X"5D",X"BB",X"4E",X"0B",X"B6",
		X"B0",X"04",X"0B",X"BA",X"BB",X"04",X"0B",X"C3",X"55",X"3C",X"0C",X"00",X"55",X"39",X"0C",X"39",
		X"50",X"04",X"0C",X"5E",X"B0",X"03",X"0C",X"61",X"BB",X"3C",X"0C",X"9D",X"B0",X"0B",X"0C",X"C8",
		X"55",X"37",X"0D",X"00",X"55",X"33",X"0D",X"33",X"50",X"04",X"0D",X"64",X"BB",X"2E",X"0D",X"CB",
		X"55",X"34",X"0E",X"00",X"55",X"21",X"0E",X"21",X"50",X"11",X"0E",X"65",X"B0",X"03",X"0E",X"68",
		X"BB",X"27",X"0E",X"8D",X"B0",X"02",X"0E",X"CF",X"55",X"30",X"0F",X"00",X"55",X"21",X"0F",X"69",
		X"BB",X"23",X"0F",X"D7",X"55",X"28",X"10",X"00",X"55",X"1E",X"10",X"70",X"B0",X"04",X"10",X"74",
		X"BB",X"18",X"10",X"DB",X"55",X"24",X"11",X"00",X"55",X"1D",X"11",X"76",X"BB",X"14",X"11",X"DC",
		X"55",X"23",X"12",X"00",X"55",X"1D",X"12",X"DD",X"55",X"22",X"13",X"00",X"55",X"1B",X"13",X"E4",
		X"55",X"1B",X"14",X"00",X"55",X"19",X"14",X"E6",X"55",X"19",X"15",X"00",X"55",X"19",X"15",X"E8",
		X"55",X"17",X"16",X"00",X"55",X"16",X"16",X"16",X"50",X"02",X"16",X"E9",X"55",X"16",X"17",X"00",
		X"55",X"16",X"17",X"E9",X"55",X"16",X"18",X"00",X"55",X"15",X"18",X"15",X"50",X"01",X"18",X"EB",
		X"55",X"14",X"19",X"00",X"55",X"14",X"19",X"EC",X"55",X"13",X"1A",X"00",X"55",X"14",X"1A",X"EC",
		X"55",X"13",X"1B",X"00",X"55",X"14",X"1B",X"EC",X"55",X"13",X"1C",X"00",X"55",X"14",X"1C",X"EC",
		X"55",X"13",X"1D",X"00",X"55",X"0B",X"1D",X"0B",X"50",X"09",X"1D",X"EB",X"50",X"08",X"1D",X"F3",
		X"55",X"0B",X"1E",X"00",X"55",X"08",X"1E",X"08",X"50",X"03",X"1E",X"F5",X"50",X"02",X"1E",X"F7",
		X"55",X"08",X"1F",X"00",X"50",X"08",X"1F",X"F7",X"55",X"08",X"20",X"F7",X"55",X"08",X"21",X"F8",
		X"55",X"07",X"00",X"00",X"36",X"34",X"CC",X"13",X"30",X"8E",X"D3",X"C3",X"10",X"8E",X"E3",X"13",
		X"33",X"C9",X"01",X"05",X"36",X"32",X"8E",X"30",X"30",X"33",X"C9",X"01",X"04",X"36",X"14",X"39",
		X"96",X"63",X"30",X"8D",X"00",X"02",X"6E",X"96",X"C0",X"1A",X"C0",X"27",X"C1",X"C5",X"C2",X"9C",
		X"C2",X"B2",X"C3",X"37",X"C3",X"A9",X"D0",X"72",X"C4",X"3B",X"BD",X"C4",X"4D",X"CC",X"02",X"FF",
		X"97",X"64",X"97",X"63",X"D7",X"0A",X"39",X"BD",X"D0",X"64",X"C6",X"04",X"D7",X"63",X"CC",X"00",
		X"A0",X"DD",X"69",X"8E",X"5D",X"7E",X"CC",X"0A",X"0A",X"ED",X"81",X"ED",X"84",X"30",X"89",X"00",
		X"FE",X"CC",X"A0",X"A0",X"ED",X"81",X"ED",X"84",X"30",X"1A",X"CC",X"AA",X"AA",X"ED",X"81",X"ED",
		X"84",X"30",X"1A",X"8C",X"63",X"00",X"25",X"DE",X"8E",X"5D",X"7E",X"CC",X"0A",X"0A",X"ED",X"81",
		X"ED",X"84",X"30",X"89",X"00",X"FE",X"CC",X"A0",X"A0",X"ED",X"81",X"ED",X"81",X"CC",X"AA",X"AA",
		X"ED",X"81",X"ED",X"81",X"8C",X"63",X"00",X"25",X"E2",X"8E",X"6B",X"7D",X"CC",X"AA",X"AA",X"ED",
		X"81",X"ED",X"81",X"ED",X"84",X"30",X"17",X"CC",X"0A",X"0A",X"ED",X"81",X"ED",X"81",X"A7",X"84",
		X"30",X"89",X"00",X"FC",X"CC",X"A0",X"A0",X"ED",X"81",X"ED",X"81",X"A7",X"84",X"30",X"16",X"8C",
		X"70",X"46",X"25",X"D8",X"8E",X"6B",X"7D",X"CC",X"AA",X"AA",X"ED",X"81",X"ED",X"81",X"ED",X"81",
		X"CC",X"0A",X"0A",X"ED",X"81",X"ED",X"81",X"A7",X"84",X"30",X"89",X"00",X"FC",X"CC",X"A0",X"A0",
		X"ED",X"81",X"ED",X"81",X"A7",X"80",X"8C",X"70",X"B4",X"25",X"DC",X"10",X"8E",X"70",X"4A",X"C6",
		X"6C",X"86",X"AA",X"BD",X"D0",X"19",X"8E",X"63",X"52",X"CC",X"AA",X"AA",X"ED",X"84",X"30",X"89",
		X"00",X"FF",X"86",X"0A",X"ED",X"81",X"86",X"A0",X"A7",X"84",X"30",X"89",X"00",X"FE",X"86",X"AA",
		X"ED",X"84",X"30",X"89",X"00",X"FF",X"ED",X"84",X"30",X"89",X"00",X"FF",X"8C",X"70",X"46",X"25",
		X"E1",X"8E",X"63",X"AC",X"CC",X"AA",X"AA",X"ED",X"84",X"30",X"89",X"01",X"00",X"86",X"A0",X"ED",
		X"81",X"86",X"0A",X"A7",X"84",X"30",X"89",X"00",X"FF",X"86",X"AA",X"ED",X"84",X"30",X"89",X"01",
		X"01",X"ED",X"84",X"30",X"89",X"01",X"00",X"8C",X"70",X"B4",X"25",X"E1",X"8E",X"6C",X"5E",X"9F",
		X"67",X"8E",X"64",X"5E",X"CE",X"C5",X"11",X"86",X"07",X"BD",X"C4",X"BB",X"8E",X"6A",X"6C",X"9F",
		X"67",X"8E",X"61",X"6C",X"CE",X"C5",X"81",X"86",X"07",X"BD",X"C4",X"BB",X"10",X"8E",X"61",X"7E",
		X"CC",X"CC",X"08",X"BD",X"D0",X"1F",X"10",X"8E",X"61",X"7F",X"CC",X"DD",X"08",X"BD",X"D0",X"1F",
		X"10",X"8E",X"61",X"80",X"CC",X"EE",X"08",X"BD",X"D0",X"1F",X"10",X"8E",X"61",X"81",X"CC",X"FF",
		X"08",X"BD",X"D0",X"1F",X"8E",X"6B",X"86",X"9F",X"67",X"8E",X"62",X"86",X"CE",X"C5",X"FF",X"86",
		X"07",X"BD",X"C4",X"BB",X"8E",X"6C",X"96",X"9F",X"67",X"8E",X"64",X"96",X"CE",X"C6",X"7D",X"86",
		X"08",X"BD",X"C4",X"BB",X"8E",X"61",X"A2",X"9F",X"67",X"8E",X"5D",X"A2",X"CE",X"C6",X"FD",X"86",
		X"04",X"7E",X"C4",X"BB",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"00",X"31",X"39",X"38",
		X"31",X"40",X"54",X"41",X"49",X"54",X"4F",X"40",X"41",X"4D",X"45",X"52",X"49",X"43",X"41",X"40",
		X"43",X"4F",X"52",X"50",X"00",X"BD",X"C4",X"44",X"26",X"E4",X"C6",X"06",X"D7",X"63",X"CC",X"01",
		X"80",X"DD",X"69",X"C6",X"22",X"8E",X"C1",X"A4",X"10",X"8E",X"48",X"60",X"BD",X"D0",X"47",X"8E",
		X"34",X"55",X"86",X"0A",X"A7",X"84",X"8E",X"35",X"55",X"86",X"AA",X"A7",X"84",X"8E",X"36",X"55",
		X"A7",X"84",X"8E",X"3F",X"56",X"9F",X"67",X"8E",X"31",X"56",X"CE",X"C7",X"1D",X"86",X"10",X"BD",
		X"C4",X"BB",X"8E",X"3C",X"75",X"9F",X"67",X"8E",X"31",X"75",X"CE",X"C8",X"DD",X"86",X"10",X"BD",
		X"C4",X"BB",X"8E",X"3E",X"92",X"CC",X"A0",X"A0",X"A7",X"80",X"ED",X"84",X"8E",X"3D",X"93",X"CC",
		X"AA",X"AA",X"ED",X"84",X"8E",X"3C",X"94",X"A7",X"84",X"8E",X"3F",X"95",X"9F",X"67",X"8E",X"31",
		X"95",X"CE",X"CA",X"3D",X"86",X"07",X"BD",X"C4",X"BB",X"8E",X"3F",X"A3",X"9F",X"67",X"8E",X"3A",
		X"A3",X"CE",X"CB",X"01",X"86",X"04",X"BD",X"C4",X"BB",X"8E",X"30",X"8A",X"86",X"0A",X"A7",X"84",
		X"8E",X"31",X"72",X"9F",X"67",X"8E",X"25",X"72",X"CE",X"CB",X"29",X"86",X"0C",X"BD",X"C4",X"BB",
		X"8E",X"1C",X"18",X"9F",X"67",X"CE",X"CC",X"6D",X"8E",X"18",X"18",X"86",X"04",X"BD",X"C4",X"BB",
		X"8E",X"1C",X"21",X"9F",X"67",X"CE",X"CC",X"8D",X"8E",X"18",X"21",X"86",X"04",X"BD",X"C4",X"BB",
		X"C6",X"22",X"8E",X"C1",X"AD",X"10",X"8E",X"18",X"30",X"BD",X"D0",X"47",X"8E",X"2D",X"91",X"9F",
		X"67",X"8E",X"2A",X"91",X"CE",X"CC",X"49",X"86",X"06",X"7E",X"C4",X"BB",X"BD",X"C4",X"44",X"26",
		X"10",X"BD",X"C4",X"FC",X"0C",X"77",X"0C",X"76",X"CC",X"F7",X"08",X"97",X"66",X"D7",X"65",X"D7",
		X"63",X"39",X"0A",X"65",X"2A",X"FB",X"D6",X"66",X"CB",X"09",X"C1",X"6C",X"24",X"42",X"D7",X"66",
		X"8E",X"CC",X"AD",X"3A",X"A6",X"07",X"27",X"24",X"34",X"10",X"10",X"8E",X"CE",X"CD",X"10",X"AE",
		X"A6",X"CE",X"BF",X"96",X"9E",X"A4",X"EF",X"81",X"9F",X"A4",X"AE",X"A4",X"AF",X"46",X"AE",X"22",
		X"AF",X"C4",X"AF",X"42",X"AE",X"24",X"A6",X"26",X"A7",X"84",X"35",X"10",X"EE",X"84",X"10",X"AE",
		X"02",X"EC",X"04",X"DD",X"67",X"A6",X"08",X"BD",X"C4",X"DB",X"A6",X"06",X"97",X"65",X"20",X"36",
		X"86",X"1E",X"CE",X"CE",X"F3",X"33",X"C6",X"AE",X"C4",X"10",X"AE",X"42",X"E6",X"44",X"BD",X"C4",
		X"70",X"80",X"05",X"2A",X"ED",X"CC",X"30",X"30",X"8E",X"44",X"29",X"ED",X"81",X"ED",X"84",X"8E",
		X"44",X"89",X"ED",X"81",X"ED",X"84",X"8E",X"44",X"CA",X"ED",X"81",X"ED",X"84",X"C6",X"0A",X"D7",
		X"63",X"CC",X"00",X"C0",X"DD",X"69",X"39",X"BD",X"C4",X"44",X"26",X"11",X"8E",X"80",X"00",X"CC",
		X"00",X"00",X"ED",X"83",X"8C",X"24",X"00",X"26",X"F9",X"C6",X"0C",X"D7",X"63",X"39",X"31",X"40",
		X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"40",X"50",X"4C",
		X"41",X"59",X"00",X"32",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"40",X"45",X"58",X"54",
		X"45",X"4E",X"44",X"45",X"44",X"40",X"57",X"45",X"41",X"50",X"4F",X"4E",X"52",X"59",X"00",X"49",
		X"4E",X"49",X"54",X"49",X"41",X"4C",X"40",X"43",X"4F",X"4C",X"4F",X"4E",X"49",X"45",X"53",X"00",
		X"42",X"4F",X"4E",X"55",X"53",X"40",X"43",X"4F",X"4C",X"4F",X"4E",X"59",X"40",X"41",X"54",X"00",
		X"32",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"FF",X"BD",X"C4",X"44",X"26",X"9F",X"10",X"8E",
		X"68",X"2C",X"8E",X"C3",X"4E",X"C6",X"22",X"8D",X"3B",X"10",X"8E",X"40",X"11",X"8D",X"35",X"10",
		X"8E",X"60",X"44",X"8E",X"C3",X"7F",X"8D",X"2C",X"10",X"8E",X"58",X"2D",X"8D",X"26",X"10",X"8E",
		X"38",X"44",X"8E",X"C3",X"7F",X"8D",X"1D",X"10",X"8E",X"30",X"2D",X"8D",X"17",X"BD",X"D0",X"29",
		X"C6",X"44",X"10",X"8E",X"60",X"34",X"85",X"01",X"27",X"0D",X"8E",X"C3",X"A2",X"8D",X"05",X"8E",
		X"C3",X"A2",X"20",X"0B",X"7E",X"D0",X"47",X"8E",X"C3",X"A0",X"8D",X"F8",X"8E",X"C3",X"A0",X"10",
		X"8E",X"38",X"34",X"8D",X"EF",X"84",X"03",X"48",X"8E",X"D0",X"6A",X"30",X"86",X"C6",X"55",X"A6",
		X"84",X"10",X"8E",X"59",X"A9",X"8D",X"66",X"A6",X"01",X"10",X"8E",X"31",X"A9",X"8D",X"5E",X"8E",
		X"C3",X"A4",X"10",X"8E",X"59",X"AF",X"8D",X"48",X"8E",X"C3",X"A4",X"10",X"8E",X"31",X"AF",X"8D",
		X"3F",X"C6",X"0E",X"D7",X"63",X"CC",X"01",X"C0",X"DD",X"69",X"39",X"8D",X"07",X"26",X"FB",X"0F",
		X"63",X"7E",X"C4",X"FC",X"9E",X"69",X"30",X"1F",X"27",X"02",X"9F",X"69",X"39",X"1F",X"40",X"C4",
		X"FE",X"1F",X"01",X"CC",X"00",X"00",X"A7",X"82",X"8C",X"A0",X"64",X"26",X"F9",X"0C",X"77",X"0C",
		X"76",X"CE",X"A0",X"00",X"8E",X"00",X"00",X"36",X"16",X"11",X"83",X"00",X"00",X"26",X"F8",X"39",
		X"34",X"02",X"A6",X"80",X"8D",X"07",X"A6",X"80",X"2A",X"FA",X"35",X"02",X"39",X"34",X"04",X"CE",
		X"CF",X"33",X"C6",X"12",X"3D",X"33",X"CB",X"C6",X"03",X"37",X"02",X"A4",X"E4",X"A7",X"A0",X"37",
		X"02",X"A4",X"E4",X"A7",X"A0",X"37",X"02",X"A4",X"E4",X"A7",X"A0",X"37",X"02",X"A4",X"E4",X"A7",
		X"A0",X"37",X"02",X"A4",X"E4",X"A7",X"A0",X"37",X"02",X"A4",X"E4",X"A7",X"A4",X"31",X"A9",X"00",
		X"FB",X"5A",X"26",X"D5",X"31",X"A9",X"FD",X"06",X"35",X"04",X"39",X"34",X"02",X"A6",X"E4",X"97",
		X"65",X"37",X"06",X"ED",X"81",X"0A",X"65",X"26",X"F8",X"CC",X"00",X"FF",X"E0",X"E4",X"E0",X"E4",
		X"CB",X"01",X"30",X"8B",X"9C",X"67",X"25",X"E5",X"35",X"02",X"39",X"34",X"02",X"A6",X"E4",X"97",
		X"65",X"37",X"06",X"ED",X"A1",X"0A",X"65",X"26",X"F8",X"CC",X"00",X"FF",X"E0",X"E4",X"E0",X"E4",
		X"CB",X"01",X"31",X"AB",X"10",X"9C",X"67",X"25",X"E4",X"35",X"02",X"39",X"BD",X"D0",X"55",X"86",
		X"88",X"97",X"0F",X"0F",X"0D",X"BD",X"D0",X"67",X"96",X"0E",X"27",X"EF",X"0C",X"0D",X"7E",X"D0",
		X"67",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"CD",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"DE",X"DE",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FC",X"FC",X"CD",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"DE",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",
		X"CD",X"CD",X"00",X"00",X"00",X"0D",X"0E",X"00",X"00",X"00",X"00",X"0F",X"DE",X"DD",X"EC",X"DD",
		X"EE",X"FF",X"CC",X"DD",X"EE",X"FF",X"EE",X"DD",X"CC",X"FF",X"EE",X"DD",X"CC",X"DD",X"EE",X"FF",
		X"CC",X"D0",X"E0",X"FF",X"EE",X"DD",X"CC",X"F0",X"E0",X"D0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0E",X"0F",X"00",
		X"0D",X"0C",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"CC",X"DD",X"EE",X"FF",X"EE",X"DD",X"CC",
		X"FF",X"0E",X"0D",X"0C",X"0D",X"EF",X"FC",X"CD",X"DE",X"EF",X"F0",X"00",X"EE",X"DD",X"CC",X"FF",
		X"EE",X"DD",X"EE",X"FF",X"CC",X"DD",X"EE",X"FF",X"00",X"00",X"00",X"EE",X"DD",X"CC",X"FF",X"E0",
		X"E0",X"FC",X"CD",X"DE",X"EF",X"F0",X"00",X"00",X"00",X"E0",X"DE",X"CD",X"FC",X"0F",X"FF",X"CC",
		X"DD",X"EE",X"FF",X"00",X"00",X"00",X"00",X"00",X"E0",X"DE",X"CD",X"CC",X"FC",X"CD",X"DE",X"EF",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"CC",X"CC",X"DD",X"EE",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"CC",X"D0",X"E0",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FE",X"FE",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"DC",X"ED",X"ED",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"CF",X"CF",X"CF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",
		X"ED",X"ED",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"CF",X"CF",
		X"CF",X"00",X"00",X"00",X"00",X"FF",X"CC",X"0D",X"0E",X"0F",X"DC",X"DC",X"ED",X"ED",X"ED",X"00",
		X"00",X"00",X"00",X"FF",X"CC",X"DD",X"EE",X"FF",X"CC",X"DD",X"EE",X"DD",X"CC",X"0F",X"0E",X"0D",
		X"0C",X"00",X"00",X"D0",X"E0",X"F0",X"C0",X"DD",X"EE",X"DD",X"CC",X"FF",X"EE",X"DD",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"D0",X"C0",X"00",X"00",X"00",
		X"0C",X"0C",X"CD",X"CD",X"CD",X"CD",X"CD",X"CD",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0C",X"CD",
		X"DD",X"DE",X"DE",X"EF",X"EF",X"EF",X"EF",X"DE",X"DE",X"DD",X"CD",X"0C",X"00",X"0C",X"CD",X"DD",
		X"EE",X"EF",X"F0",X"00",X"00",X"00",X"00",X"F0",X"EF",X"EE",X"DD",X"CD",X"0C",X"CC",X"DD",X"EE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"DD",X"CC",X"CC",X"DD",X"EE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"EE",X"DD",X"CC",X"C0",X"DC",X"DD",
		X"EE",X"FE",X"0F",X"00",X"00",X"00",X"00",X"0F",X"FE",X"EE",X"DD",X"DC",X"C0",X"00",X"C0",X"DC",
		X"DD",X"ED",X"ED",X"FE",X"FE",X"FE",X"FE",X"ED",X"ED",X"DD",X"DC",X"C0",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"0A",X"0A",X"00",X"00",X"00",X"0A",X"A0",X"33",X"00",X"33",X"A0",X"0A",X"00",X"AA",X"00",X"33",
		X"30",X"03",X"00",X"AA",X"00",X"00",X"A0",X"3A",X"3A",X"3A",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"22",X"00",X"00",X"0A",X"AA",
		X"A2",X"A2",X"21",X"21",X"21",X"21",X"21",X"21",X"21",X"A2",X"A2",X"AA",X"AA",X"0A",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"22",X"00",X"0A",X"AA",X"A2",
		X"21",X"19",X"11",X"11",X"11",X"12",X"12",X"12",X"1A",X"1A",X"1A",X"1A",X"A1",X"A1",X"AA",X"AA",
		X"0A",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"A0",X"AA",X"2A",X"00",X"AA",X"22",X"11",
		X"11",X"99",X"11",X"11",X"12",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"1A",X"A1",
		X"A1",X"AA",X"0A",X"AA",X"A2",X"A2",X"A2",X"A2",X"A2",X"AA",X"0A",X"00",X"00",X"AA",X"22",X"11",
		X"11",X"99",X"11",X"11",X"22",X"2A",X"AA",X"AA",X"A0",X"00",X"00",X"A0",X"A0",X"A0",X"AA",X"AA",
		X"AA",X"1A",X"A1",X"21",X"11",X"11",X"11",X"11",X"21",X"21",X"A2",X"AA",X"00",X"AA",X"22",X"11",
		X"11",X"99",X"11",X"11",X"22",X"A2",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"22",X"11",X"12",X"2A",X"AA",X"AA",X"1A",X"11",X"21",X"AA",X"00",X"AA",X"2A",X"12",
		X"11",X"91",X"99",X"11",X"21",X"22",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"11",X"11",X"22",X"AA",X"00",X"00",X"AA",X"AA",X"11",X"22",X"00",X"A0",X"AA",X"2A",
		X"12",X"11",X"91",X"19",X"11",X"22",X"22",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"AA",X"1A",X"11",X"21",X"A2",X"AA",X"AA",X"A1",X"21",X"11",X"22",X"00",X"00",X"00",X"A0",
		X"AA",X"2A",X"12",X"11",X"99",X"11",X"21",X"22",X"A2",X"AA",X"AA",X"0A",X"00",X"00",X"0A",X"0A",
		X"0A",X"0A",X"AA",X"AA",X"1A",X"11",X"11",X"11",X"12",X"12",X"2A",X"AA",X"00",X"00",X"00",X"00",
		X"A0",X"AA",X"2A",X"22",X"11",X"91",X"19",X"19",X"21",X"A2",X"A2",X"AA",X"AA",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"2A",X"2A",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"AA",X"2A",X"2A",X"11",X"11",X"91",X"21",X"21",X"A2",X"A2",X"A2",X"A2",X"A2",
		X"A2",X"22",X"21",X"22",X"A2",X"AA",X"AA",X"AA",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"AA",X"1A",X"1A",X"11",X"11",X"11",X"11",X"21",X"11",
		X"11",X"11",X"11",X"21",X"22",X"22",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"AA",X"AA",X"1A",X"1A",X"1A",
		X"1A",X"1A",X"1A",X"12",X"22",X"22",X"22",X"AA",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"99",X"29",X"21",
		X"A2",X"A2",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"1A",X"99",X"19",X"11",X"11",X"21",
		X"22",X"A2",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"11",
		X"11",X"11",X"21",X"21",X"21",X"21",X"22",X"A2",X"A2",X"A2",X"A2",X"22",X"99",X"11",X"11",X"11",
		X"21",X"22",X"A2",X"AA",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"92",X"92",
		X"92",X"19",X"19",X"11",X"11",X"11",X"11",X"11",X"11",X"21",X"21",X"21",X"11",X"11",X"11",X"11",
		X"11",X"12",X"22",X"22",X"A2",X"AA",X"AA",X"AA",X"0A",X"00",X"00",X"0A",X"00",X"AA",X"AA",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"12",X"12",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"2A",X"2A",X"2A",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A2",X"A1",X"A9",
		X"A1",X"A1",X"A1",X"A2",X"A2",X"A2",X"AA",X"A0",X"AA",X"A1",X"A1",X"A1",X"A1",X"A1",X"AA",X"AA",
		X"0A",X"AA",X"A2",X"A2",X"A2",X"00",X"0A",X"AA",X"21",X"11",X"21",X"22",X"AA",X"AA",X"22",X"99",
		X"11",X"11",X"11",X"12",X"22",X"22",X"AA",X"AA",X"A2",X"11",X"12",X"12",X"12",X"12",X"11",X"21",
		X"A2",X"AA",X"12",X"99",X"22",X"AA",X"AA",X"A2",X"11",X"11",X"11",X"22",X"AA",X"AA",X"22",X"99",
		X"11",X"22",X"AA",X"AA",X"AA",X"AA",X"AA",X"22",X"11",X"11",X"22",X"AA",X"A0",X"A0",X"AA",X"11",
		X"22",X"AA",X"22",X"99",X"21",X"A2",X"22",X"21",X"11",X"11",X"11",X"11",X"22",X"AA",X"AA",X"11",
		X"99",X"11",X"A2",X"AA",X"AA",X"A0",X"AA",X"2A",X"12",X"11",X"22",X"AA",X"0A",X"0A",X"AA",X"11",
		X"22",X"AA",X"AA",X"22",X"99",X"11",X"11",X"11",X"12",X"22",X"22",X"19",X"11",X"AA",X"AA",X"2A",
		X"91",X"11",X"22",X"AA",X"AA",X"00",X"00",X"AA",X"2A",X"12",X"12",X"21",X"21",X"21",X"11",X"12",
		X"22",X"AA",X"AA",X"22",X"91",X"11",X"11",X"12",X"2A",X"AA",X"22",X"91",X"12",X"00",X"AA",X"AA",
		X"2A",X"2A",X"2A",X"AA",X"AA",X"AA",X"00",X"00",X"A0",X"AA",X"AA",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"A0",X"00",X"A0",X"AA",X"2A",X"2A",X"2A",X"2A",X"A0",X"A0",X"AA",X"1A",X"2A",X"00",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",
		X"00",X"00",X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"A0",X"A0",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"A2",X"A2",X"22",
		X"22",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"22",X"29",X"21",X"21",X"22",X"AA",
		X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"22",X"99",X"11",X"11",X"22",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"AA",X"22",X"91",X"11",X"11",X"22",X"A2",X"AA",X"0A",X"00",X"00",
		X"00",X"AA",X"AA",X"AA",X"22",X"11",X"11",X"11",X"11",X"22",X"A2",X"AA",X"0A",X"00",X"00",X"AA",
		X"AA",X"AA",X"22",X"11",X"11",X"11",X"11",X"11",X"22",X"22",X"AA",X"AA",X"00",X"22",X"AA",X"A2",
		X"11",X"99",X"11",X"22",X"12",X"11",X"11",X"21",X"22",X"AA",X"AA",X"2A",X"AA",X"22",X"11",X"11",
		X"22",X"2A",X"2A",X"12",X"11",X"19",X"21",X"22",X"A2",X"AA",X"22",X"11",X"19",X"11",X"2A",X"AA",
		X"AA",X"2A",X"12",X"91",X"19",X"11",X"22",X"22",X"11",X"19",X"12",X"22",X"AA",X"AA",X"A0",X"AA",
		X"AA",X"2A",X"12",X"12",X"12",X"2A",X"2A",X"2A",X"2A",X"2A",X"AA",X"A0",X"00",X"00",X"A0",X"AA",
		X"AA",X"2A",X"2A",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",
		X"A0",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"A2",X"AA",X"AA",X"0A",X"00",X"00",X"00",
		X"00",X"22",X"22",X"AA",X"AA",X"0A",X"00",X"00",X"00",X"2A",X"2A",X"2A",X"AA",X"AA",X"AA",X"0A",
		X"00",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"01",X"11",X"00",X"00",X"11",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"01",X"11",X"11",X"11",X"1F",X"11",X"11",
		X"11",X"11",X"11",X"10",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"11",X"1F",
		X"11",X"11",X"F1",X"11",X"1F",X"1F",X"11",X"11",X"11",X"1F",X"11",X"11",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"11",X"1F",X"11",X"11",X"11",X"F1",X"11",X"1F",X"11",X"11",
		X"11",X"11",X"F1",X"11",X"11",X"11",X"01",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"11",
		X"11",X"1A",X"1A",X"11",X"11",X"11",X"12",X"02",X"02",X"10",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"00",X"AA",X"AA",X"12",X"11",X"19",X"11",X"22",
		X"0A",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"AA",X"AA",X"11",X"99",X"19",X"21",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"AA",X"2A",X"11",X"99",X"11",
		X"21",X"22",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"12",X"91",X"99",X"11",X"11",X"22",X"AA",X"0A",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"AA",X"AA",X"11",X"91",
		X"19",X"11",X"21",X"22",X"AA",X"AA",X"0A",X"00",X"00",X"AA",X"AA",X"AA",X"0A",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"11",X"99",X"91",X"11",X"21",X"22",X"AA",X"AA",X"0A",
		X"00",X"AA",X"AA",X"22",X"A2",X"A2",X"AA",X"AA",X"0A",X"0A",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"12",X"99",X"19",X"11",X"21",X"22",X"A2",X"AA",X"AA",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"02",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"22",X"00",X"22",
		X"00",X"20",X"20",X"20",X"20",X"20",X"00",X"20",X"20",X"00",X"20",X"20",X"00",X"00",X"0A",X"A2",
		X"A0",X"A0",X"A0",X"0A",X"00",X"AA",X"00",X"22",X"02",X"02",X"00",X"00",X"AA",X"AA",X"00",X"22",
		X"00",X"00",X"22",X"00",X"AA",X"00",X"A0",X"2A",X"2A",X"2A",X"0A",X"A0",X"00",X"00",X"0A",X"A0",
		X"A2",X"A2",X"A0",X"0A",X"00",X"AA",X"00",X"22",X"00",X"00",X"20",X"00",X"AA",X"AA",X"00",X"22",
		X"00",X"00",X"02",X"00",X"AA",X"00",X"A0",X"0A",X"2A",X"2A",X"0A",X"A0",X"00",X"CE",X"A7",X"50",
		X"1B",X"51",X"1B",X"08",X"02",X"14",X"CE",X"7F",X"50",X"1B",X"52",X"1B",X"08",X"00",X"14",X"CE",
		X"57",X"50",X"1B",X"53",X"1B",X"64",X"00",X"14",X"CD",X"55",X"50",X"50",X"51",X"50",X"08",X"04",
		X"0F",X"CD",X"37",X"50",X"50",X"52",X"50",X"08",X"00",X"0F",X"CD",X"19",X"50",X"50",X"53",X"50",
		X"64",X"00",X"0F",X"CD",X"BB",X"50",X"7C",X"51",X"7C",X"08",X"06",X"12",X"CD",X"97",X"50",X"7C",
		X"52",X"7C",X"08",X"00",X"12",X"CD",X"73",X"50",X"7C",X"53",X"7C",X"64",X"00",X"12",X"CE",X"2F",
		X"50",X"BC",X"51",X"BC",X"08",X"08",X"14",X"CE",X"07",X"50",X"BC",X"52",X"BC",X"08",X"00",X"14",
		X"CD",X"DF",X"50",X"BC",X"53",X"BC",X"64",X"00",X"14",X"04",X"40",X"40",X"40",X"04",X"00",X"44",
		X"40",X"40",X"40",X"44",X"00",X"44",X"40",X"40",X"40",X"44",X"00",X"44",X"40",X"40",X"40",X"44",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"40",X"00",X"44",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"40",X"04",X"04",X"04",X"00",X"00",X"44",X"04",X"04",X"04",X"44",
		X"00",X"44",X"04",X"04",X"04",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"04",X"44",
		X"04",X"04",X"00",X"44",X"40",X"40",X"40",X"04",X"00",X"44",X"40",X"40",X"40",X"44",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"40",X"40",X"40",X"40",
		X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"44",X"04",X"04",X"40",X"00",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",X"00",X"44",
		X"04",X"04",X"04",X"00",X"00",X"44",X"40",X"40",X"04",X"00",X"00",X"44",X"04",X"04",X"40",X"00",
		X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"04",X"40",X"04",X"44",X"00",X"44",X"04",X"40",
		X"04",X"44",X"00",X"44",X"04",X"04",X"04",X"04",X"00",X"44",X"04",X"04",X"40",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"00",X"44",X"40",X"40",X"40",X"04",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"40",X"44",X"40",X"00",X"04",X"40",X"40",X"40",X"40",X"04",X"44",X"40",X"40",X"40",X"44",
		X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"44",X"40",X"40",X"40",X"44",X"00",X"44",X"00",X"00",
		X"00",X"44",X"00",X"00",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"04",
		X"04",X"40",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"44",X"40",X"40",X"04",X"00",X"00",X"44",
		X"04",X"04",X"04",X"44",X"00",X"44",X"04",X"04",X"04",X"40",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"04",X"44",X"04",X"00",X"40",X"04",X"04",X"04",X"00",X"00",X"44",X"04",X"04",X"04",X"44",
		X"00",X"44",X"04",X"04",X"40",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"40",X"44",X"40",
		X"00",X"44",X"40",X"40",X"40",X"44",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",
		X"00",X"00",X"00",X"44",X"40",X"40",X"40",X"40",X"00",X"44",X"00",X"00",X"04",X"40",X"00",X"44",
		X"04",X"04",X"04",X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"00",X"00",X"40",X"40",X"00",X"44",
		X"40",X"40",X"40",X"44",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"44",X"04",X"04",X"00",X"00",
		X"00",X"44",X"40",X"40",X"04",X"00",X"00",X"44",X"04",X"04",X"04",X"04",X"00",X"04",X"44",X"04",
		X"00",X"44",X"04",X"04",X"04",X"04",X"00",X"44",X"00",X"00",X"00",X"44",X"00",X"04",X"04",X"44",
		X"04",X"04",X"00",X"44",X"04",X"04",X"04",X"04",X"00",X"44",X"04",X"04",X"40",X"00",X"00",X"CE",
		X"D7",X"CE",X"DE",X"CE",X"E5",X"CE",X"EC",X"D0",X"58",X"92",X"2A",X"BF",X"9B",X"0C",X"D0",X"5B",
		X"92",X"5A",X"A0",X"AE",X"08",X"D0",X"61",X"92",X"86",X"BF",X"9A",X"0A",X"D0",X"5E",X"92",X"CD",
		X"BF",X"AA",X"0A",X"CF",X"16",X"43",X"B5",X"44",X"CF",X"1A",X"43",X"D0",X"44",X"CF",X"1F",X"43",
		X"73",X"22",X"CF",X"23",X"43",X"90",X"22",X"CF",X"28",X"43",X"55",X"44",X"CF",X"2C",X"43",X"19",
		X"22",X"CF",X"2F",X"43",X"30",X"22",X"05",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"FF",X"01",
		X"00",X"00",X"FF",X"01",X"00",X"00",X"00",X"FF",X"01",X"00",X"00",X"FF",X"02",X"05",X"FF",X"02",
		X"05",X"00",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"0F",X"0F",X"0F",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"FF",X"F0",
		X"F0",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"FF",
		X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"FF",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"00",
		X"00",X"F0",X"F0",X"FF",X"F0",X"00",X"00",X"0F",X"0F",X"FF",X"00",X"00",X"0F",X"0F",X"0F",X"FF",
		X"FF",X"00",X"FF",X"FF",X"00",X"F0",X"F0",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"00",
		X"FF",X"F0",X"F0",X"F0",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",X"FF",X"0F",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"0F",X"00",X"00",X"FF",
		X"0F",X"0F",X"FF",X"00",X"FF",X"FF",X"F0",X"FF",X"FF",X"00",X"F0",X"FF",X"F0",X"FF",X"F0",X"00",
		X"00",X"FF",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",
		X"FF",X"00",X"FF",X"0F",X"0F",X"0F",X"FF",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"11",X"11",X"22",X"AA",X"00",X"00",X"AA",X"AA",X"11",X"22",X"00",X"A0",X"AA",X"2A",
		X"B6",X"BF",X"AB",X"8E",X"C0",X"08",X"6E",X"96",X"C0",X"10",X"C0",X"39",X"C0",X"50",X"C0",X"70",
		X"BD",X"C0",X"67",X"26",X"23",X"BD",X"C0",X"78",X"CC",X"02",X"E0",X"DD",X"69",X"CC",X"02",X"10",
		X"B7",X"BF",X"AB",X"F7",X"65",X"E2",X"F7",X"67",X"E2",X"8E",X"C0",X"86",X"E6",X"80",X"27",X"08",
		X"10",X"AE",X"81",X"BD",X"D0",X"47",X"20",X"F4",X"39",X"BD",X"C0",X"67",X"26",X"FA",X"BD",X"C0",
		X"78",X"CC",X"03",X"80",X"DD",X"69",X"86",X"04",X"B7",X"BF",X"AB",X"8E",X"C1",X"CB",X"20",X"DC",
		X"BD",X"C0",X"67",X"26",X"E3",X"BD",X"C0",X"78",X"CC",X"01",X"80",X"DD",X"69",X"86",X"06",X"B7",
		X"BF",X"AB",X"8E",X"C3",X"3B",X"20",X"C5",X"9E",X"69",X"30",X"1F",X"27",X"02",X"9F",X"69",X"39",
		X"86",X"10",X"97",X"63",X"7F",X"BF",X"AB",X"39",X"CC",X"00",X"00",X"8E",X"80",X"00",X"ED",X"83",
		X"8C",X"24",X"00",X"26",X"F9",X"39",X"44",X"78",X"60",X"43",X"4F",X"4C",X"4F",X"4E",X"59",X"40",
		X"37",X"00",X"11",X"6E",X"10",X"44",X"45",X"46",X"45",X"4E",X"44",X"40",X"43",X"4F",X"4C",X"4F",
		X"4E",X"59",X"40",X"37",X"40",X"46",X"52",X"4F",X"4D",X"40",X"45",X"4E",X"45",X"4D",X"49",X"45",
		X"53",X"5A",X"00",X"11",X"64",X"20",X"59",X"4F",X"55",X"52",X"40",X"41",X"52",X"53",X"45",X"4E",
		X"41",X"4C",X"40",X"43",X"4F",X"4E",X"53",X"49",X"53",X"54",X"53",X"40",X"4F",X"46",X"00",X"88",
		X"5A",X"10",X"4D",X"41",X"49",X"4E",X"40",X"57",X"45",X"41",X"50",X"4F",X"4E",X"52",X"59",X"40",
		X"00",X"11",X"5A",X"80",X"54",X"52",X"49",X"47",X"47",X"45",X"52",X"45",X"44",X"40",X"42",X"59",
		X"00",X"11",X"54",X"10",X"46",X"49",X"52",X"45",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"40",
		X"54",X"4F",X"40",X"45",X"58",X"50",X"4C",X"4F",X"44",X"45",X"40",X"41",X"54",X"00",X"11",X"4E",
		X"10",X"43",X"52",X"4F",X"53",X"53",X"48",X"41",X"49",X"52",X"5A",X"40",X"41",X"49",X"4D",X"40",
		X"57",X"49",X"54",X"48",X"40",X"4A",X"4F",X"59",X"53",X"54",X"49",X"43",X"4B",X"5A",X"00",X"88",
		X"44",X"10",X"4D",X"45",X"47",X"41",X"42",X"4C",X"41",X"53",X"54",X"45",X"52",X"40",X"00",X"11",
		X"44",X"70",X"57",X"49",X"44",X"45",X"40",X"43",X"4F",X"56",X"45",X"52",X"41",X"47",X"45",X"00",
		X"11",X"3E",X"10",X"57",X"45",X"41",X"50",X"4F",X"4E",X"40",X"50",X"4F",X"57",X"45",X"52",X"45",
		X"44",X"40",X"42",X"59",X"40",X"50",X"55",X"4C",X"53",X"41",X"54",X"49",X"4E",X"47",X"00",X"11",
		X"38",X"10",X"46",X"55",X"45",X"4C",X"40",X"43",X"45",X"4C",X"4C",X"53",X"40",X"49",X"4E",X"40",
		X"54",X"48",X"45",X"40",X"43",X"4F",X"4C",X"4F",X"4E",X"59",X"5A",X"00",X"11",X"32",X"10",X"55",
		X"53",X"45",X"44",X"40",X"46",X"55",X"45",X"4C",X"40",X"43",X"45",X"4C",X"4C",X"53",X"40",X"54",
		X"55",X"52",X"4E",X"40",X"42",X"4C",X"55",X"45",X"5A",X"00",X"22",X"28",X"10",X"45",X"4E",X"45",
		X"4D",X"59",X"40",X"46",X"49",X"52",X"45",X"40",X"4D",X"41",X"59",X"40",X"44",X"45",X"53",X"54",
		X"52",X"4F",X"59",X"40",X"43",X"45",X"4C",X"4C",X"53",X"00",X"00",X"44",X"78",X"60",X"43",X"4F",
		X"4C",X"4F",X"4E",X"59",X"40",X"37",X"00",X"11",X"6E",X"10",X"54",X"48",X"45",X"40",X"00",X"88",
		X"6E",X"30",X"45",X"52",X"41",X"44",X"49",X"43",X"41",X"54",X"4F",X"52",X"40",X"00",X"11",X"6E",
		X"88",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"53",X"00",X"11",X"68",X"10",X"41",X"4C",X"4C",
		X"40",X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",X"40",X"41",X"4E",X"44",X"40",X"42",X"4F",X"4D",
		X"42",X"53",X"40",X"4F",X"4E",X"00",X"11",X"62",X"10",X"54",X"48",X"45",X"40",X"53",X"43",X"52",
		X"45",X"45",X"4E",X"5A",X"40",X"49",X"54",X"40",X"57",X"41",X"49",X"54",X"53",X"40",X"4F",X"4E",
		X"00",X"11",X"5C",X"10",X"54",X"48",X"45",X"40",X"50",X"41",X"44",X"40",X"55",X"4E",X"54",X"49",
		X"4C",X"40",X"4C",X"41",X"55",X"4E",X"43",X"48",X"45",X"44",X"5A",X"00",X"11",X"52",X"10",X"45",
		X"4E",X"45",X"4D",X"59",X"40",X"53",X"50",X"41",X"43",X"45",X"43",X"52",X"41",X"46",X"54",X"40",
		X"41",X"54",X"54",X"41",X"43",X"4B",X"40",X"49",X"4E",X"00",X"11",X"4C",X"10",X"53",X"51",X"55",
		X"41",X"44",X"52",X"4F",X"4E",X"53",X"40",X"4F",X"46",X"40",X"33",X"30",X"40",X"46",X"49",X"47",
		X"48",X"54",X"45",X"52",X"53",X"5A",X"00",X"11",X"46",X"10",X"53",X"43",X"4F",X"55",X"54",X"53",
		X"40",X"43",X"41",X"4C",X"4C",X"40",X"4D",X"4F",X"52",X"45",X"40",X"46",X"49",X"47",X"48",X"54",
		X"45",X"52",X"53",X"00",X"11",X"40",X"10",X"55",X"4E",X"54",X"49",X"4C",X"40",X"54",X"48",X"45",
		X"59",X"40",X"41",X"52",X"45",X"40",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"45",X"44",X"5A",
		X"00",X"33",X"36",X"10",X"42",X"4F",X"4E",X"55",X"53",X"40",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"40",X"41",X"52",X"45",X"40",X"41",X"57",X"41",X"52",X"44",X"45",X"44",X"00",X"33",X"30",X"10",
		X"46",X"4F",X"52",X"40",X"42",X"55",X"49",X"4C",X"44",X"49",X"4E",X"47",X"53",X"40",X"53",X"54",
		X"49",X"4C",X"4C",X"40",X"49",X"4E",X"40",X"54",X"48",X"45",X"00",X"33",X"2A",X"10",X"43",X"4F",
		X"4C",X"4F",X"4E",X"59",X"40",X"57",X"48",X"45",X"4E",X"40",X"54",X"48",X"45",X"40",X"4C",X"41",
		X"53",X"54",X"40",X"53",X"48",X"49",X"50",X"40",X"49",X"4E",X"00",X"33",X"24",X"10",X"45",X"41",
		X"43",X"48",X"40",X"53",X"51",X"55",X"41",X"44",X"52",X"4F",X"4E",X"40",X"49",X"53",X"40",X"44",
		X"45",X"53",X"54",X"52",X"4F",X"59",X"45",X"44",X"5A",X"00",X"00",X"44",X"78",X"60",X"43",X"4F",
		X"4C",X"4F",X"4E",X"59",X"40",X"37",X"00",X"11",X"6E",X"20",X"41",X"40",X"54",X"55",X"52",X"4E",
		X"40",X"45",X"4E",X"44",X"53",X"40",X"57",X"48",X"45",X"4E",X"40",X"42",X"4F",X"54",X"48",X"40",
		X"4F",X"46",X"00",X"11",X"68",X"20",X"54",X"48",X"45",X"40",X"43",X"41",X"4E",X"4E",X"4F",X"4E",
		X"53",X"40",X"41",X"52",X"45",X"40",X"42",X"4C",X"4F",X"57",X"4E",X"40",X"55",X"50",X"00",X"11",
		X"62",X"20",X"4F",X"52",X"40",X"41",X"4C",X"4C",X"40",X"4F",X"46",X"40",X"54",X"48",X"45",X"40",
		X"43",X"4F",X"4C",X"4F",X"4E",X"59",X"40",X"49",X"53",X"00",X"11",X"5C",X"20",X"44",X"45",X"53",
		X"54",X"52",X"4F",X"59",X"45",X"44",X"40",X"42",X"59",X"40",X"54",X"48",X"45",X"40",X"45",X"4E",
		X"45",X"4D",X"49",X"45",X"53",X"5A",X"00",X"88",X"48",X"58",X"47",X"4F",X"4F",X"44",X"40",X"40",
		X"4C",X"55",X"43",X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
