-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_1R is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_1R is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_1R_0 : RAMB16_S2
	generic map (
		INIT_00 => x"53FBA9998808B9A8F55560657504677561FFDEFFF0FDCFDCEDE3644440000000",
		INIT_01 => x"0F4461F465760F4453F465760F4441F465760F4673F465760F4661F465760F47",
		INIT_02 => x"C0445576CF465760F4445DF465760F4453F465760F4441F465760F4473F46576",
		INIT_03 => x"A8A46464646461411431411431411431411431413434646464646F64440EDFCD",
		INIT_04 => x"21F465760F8B936CCC88888880095D94F97D96F95D94F97D96F95D94F8A8A8A8",
		INIT_05 => x"0F0033F465760F0021F465760F0013F465760F0001F465760F0233F465760F02",
		INIT_06 => x"300E0010070080060C900F465760F0001DF465760F0013F465760F0001F46576",
		INIT_07 => x"FBFC0DFEFF3310300676067445604754DF44004000000000000000F044F00C00",
		INIT_08 => x"DFABAA90FFF0FD0DDE4FABAA98FFF8FD0DFECFABAA93FFF3FC0DDE7FABAA9BFF",
		INIT_09 => x"FFF2FF0DDE6FABAA9AFFFAFF0DFEEFABAA91FFF1FE0DDE5FABAA99FFF9FE0DFE",
		INIT_0A => x"FCECFCDEF57676467477CFABAA93FFF3FC0DDE7FABAA9BFFFBFC0DFEFFABAA92",
		INIT_0B => x"4448F88844444A88844644446622226222EEFDECFF0CDCEFDDCFF0CDCCFEDFFE",
		INIT_0C => x"000000031313130F03100132103DF44444444AF444444448F44444444AF88844",
		INIT_0D => x"F01F00F03F02F01FFF3F02F01F00F03F02F01FEEEEEEEAAF5F5F5F0C4C4C4C00",
		INIT_0E => x"9F08F0BF0AF09FCF7F06F05F04F07F06F05FEF7F06F05F04F07F06F05FDF3F02",
		INIT_0F => x"0CF0FF0EF0DFCFFF0EF0DF0CF0FF0EF0DFFFBF0AF09F08F0BF0AF09FDFBF0AF0",
		INIT_10 => x"F93F5553E4F1E4EA000FC09393AA4444444400000000938F8989AB0FFF0EF0DF",
		INIT_11 => x"55000AAA38E55500E00E00FF555FF555E79E79E79E79924E6C555B39005AAFC6",
		INIT_12 => x"3A43A4E4E93902A540AAA01500EA8E02AE5B4F1E4E579395000505A93C6A0005",
		INIT_13 => x"04D3C48CCC442BC48C4404F000006CE4C0031B39AAF0003A44E492CFEA6CE90E",
		INIT_14 => x"E66E66ED555545145944AC534577F3F37737D3F7BFFF772BF7BF7737F3CCC044",
		INIT_15 => x"3A8CFFFFFFFFFFFFFEFF7FF4FF40EDDED9ED5FD195D8BC317C312556ED65566E",
		INIT_16 => x"380808080ABC304C4C4EFC3008080ABC384C4EFC38080ABC304EFC300ABC3AFC",
		INIT_17 => x"4C4C4EFC3808080808080ABC304C4C4C4C4EFC30080808080ABC384C4C4C4EFC",
		INIT_18 => x"00000000000000000000003C4C4C4C4C4C4C4EFC0808080808080ABC384C4C4C",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"C848000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"BA00555445533A9AABA9317710000B98BB889A88032116765446745547656220",
		INIT_1D => x"998AAAAA1761191150988073A9A36800133203023112310133020039A3645552",
		INIT_1E => x"00000000FBBBBBBBBB63477577509160670B9A9BB29176747465441176503138",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"54657564CF6744560765554406067059F546706744560655544059FCFDCB0020",
		INIT_21 => x"F4604C58F312320121214AAA666666666666464424202F64440657454CF56EF4",
		INIT_22 => x"23200233135F3123200032127F4604D58F4604C5CF312320F4604C78F4604D54",
		INIT_23 => x"6F3123200233134F3123200032126F4604D79F4604D59F4604D5BF4604C5FF31",
		INIT_24 => x"766586578575FDFFDC0DED0DFD6F4604D7AF4604D58F4604C5EF312320002100",
		INIT_25 => x"0000000000000000000000000000000000000000000000000DD9615D96111575",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"C3FAFF003F000030F0A11000F5F05030CF0000303F00003000A000203C3F2F00",
		INIT_2B => x"B73FB73033333330F0300000B0FA0A00F0A11000E0000000E00002003FC033C0",
		INIT_2C => x"F33333C0F33330C0F30000C0CCCCC00033131310333333300000000033333330",
		INIT_2D => x"F0000000F0000000F0000000F0300300F0300300F0300300F0300300F0300300",
		INIT_2E => x"DF5F0000D3130000DC4C0000A0048C00A0A00000B1B1B1008C048C00B1B1B1C0",
		INIT_2F => x"B5F533C0B13133C0B4C433C005F5F500A0A0A200C5F5F5300010003012200010",
		INIT_30 => x"FFFFA50000003210000000000000000000000A00000013100000000000000000",
		INIT_31 => x"400080034003800280418040791E4791E4791E4791E4791E4791E4791E4791E4",
		INIT_32 => x"4001400040034003400240014000400340034002400140004003400340024001",
		INIT_33 => x"0103020102010102000140034003400340034003400240014000400340034002",
		INIT_34 => x"0003020002020303020302020201020200010103010102010003010002010301",
		INIT_35 => x"0002000102000002000302000002000302000002000102000002000302000002",
		INIT_36 => x"0200030200020200030200020200020200020200020200010200020200010200",
		INIT_37 => x"4100022A2A8143021515C142013F3F0181400003020000020003020003020003",
		INIT_38 => x"AAAA4302040F0F43010450504300026CE4430304FA5A4302010000C001000000",
		INIT_39 => x"01045555410004000041030840404102043333400104999940000444CC400304",
		INIT_3A => x"AA420304AA5542020455004201040A004200040000420304FFFF410204AAAA41",
		INIT_3B => x"08FF0040010800AA40000855FF4303080000430208DDDD43010800FF430004FF",
		INIT_3C => x"986420010B8E6FB1868A24103CFA385C70200E4341000890E4410308048C4102",
		INIT_3D => x"DAFB5040A281070C2799C74610D0B4D6FB1868A24503CFA795450618107CF279",
		INIT_3E => x"94BC36B214D8284943C3AB254D0288947C32BA9454E3090B8E6791458A249034",
		INIT_3F => x"022055700000000000000000000000000000300AF358E0698147C32B294D4280"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1R_1 : RAMB16_S2
	generic map (
		INIT_00 => x"45F4456474054549F57470457605474549FFDCFCC0CEDCCDFCD8313131313130",
		INIT_01 => x"0F6554F575740F6557F575740F6557F575740F5446F575740F5746F575740F54",
		INIT_02 => x"D05664667F575740F65442F575740F6565F575740F6565F575740F6554F57574",
		INIT_03 => x"213302312013091A90993992891890B93B92A91AB090213203102F75570FCEED",
		INIT_04 => x"06F131300F1005331313131313210A10913913813813B12B12A12A1291320310",
		INIT_05 => x"0F2114F131300F2114F131300F2117F131300F2117F131300F1006F131300F13",
		INIT_06 => x"D00357C00075F00353C00F131300F21002F131300F2125F131300F2125F13130",
		INIT_07 => x"38F003300FA89A8000310331110020100F6480460C64C846846440F457B00275",
		INIT_08 => x"1F030019F239F003001F030019F239F003301F030018F238F003000F030018F2",
		INIT_09 => x"F239F003001F030019F239F003301F030019F239F003001F030019F239F00330",
		INIT_0A => x"F002F001F210102033302F030019F239F103001F030019F239F103301F030019",
		INIT_0B => x"444EF00044444D5476547644546464757533F2021000213F2021000213F32302",
		INIT_0C => x"000000001122330F88A9099B8A80F44444444FF44444444FF44444444EF00044",
		INIT_0D => x"C0EC0EC0DC0DC0DC2FEC0EC0EC0EC0DC0DC0DC256745674055AAFF004488CC00",
		INIT_0E => x"EC0EC0DC0DC0DC0FEC0EC0EC0EC0DC0DC0DC3FEC0EC0EC0EC0DC0DC0DC3FEC0E",
		INIT_0F => x"0EC0DC0DC0DC1FEC0EC0EC0EC0DC0DC0DC0FEC0EC0EC0EC0DC0DC0DC0FEC0EC0",
		INIT_10 => x"554000145505550002A5405454008A8A8A8A8A8A8A8A113F565544FFEC0EC0EC",
		INIT_11 => x"00555555965000565565AA555550000001554054054000001655558000055015",
		INIT_12 => x"940940550540000015555540025025555000505550015400AA0000554155AAA0",
		INIT_13 => x"4813C40C00C89FC4CCC44802222255050000505500002A955500001540025550",
		INIT_14 => x"66AA6AE662A624D24D241E4C2443F377F77B13F73F33FB9FF7FFF77B03CC44C4",
		INIT_15 => x"7CF32226A2A62226A2BCCFCCFCC0C0CC00C08FC4C4C0FC793C792662E66EA6EE",
		INIT_16 => x"74CCCCCCCCFC78CCCCCCFC78CCCCCCFC78CCCCFC78CCCCFC7CCCFC7CCCFC7CFC",
		INIT_17 => x"CCCCCCFC70CCCCCCCCCCCCFC74CCCCCCCCCCFC74CCCCCCCCCCFC74CCCCCCCCFC",
		INIT_18 => x"00000000000000000000003CCCCCCCCCCCCCCCFCCCCCCCCCCCCCCCFC70CCCCCC",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"CCCC000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"50138821201000555540000B81523A130111113770108805555645111005431A",
		INIT_1D => x"8111311000008880312575446102AB03AA8111AA111AA0210A91211088899054",
		INIT_1E => x"00000000F44444444460444544505100255750190211811111112339A356011B",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"557545449F7755540445647404047044F677707755540456474044FECDCF3132",
		INIT_21 => x"F7704D52F013300201116222301112311233030010101F75570302211AF64DF5",
		INIT_22 => x"33001330106F0133000100215F7704D4EF7704D5EF01330AF7704D42F7704D42",
		INIT_23 => x"6F0133001330106F0133000100215F7704D42F7704D42F7704D41F7704D51F01",
		INIT_24 => x"767587448576FEECDF0DCC0DFEAF7704D42F7704D42F7704D51F013300010221",
		INIT_25 => x"0000000000000000000000000000000000000000000000000DDD61DD1611D1B6",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"C3F5FF203FFA5030F0A33000FFAA5030CFFA50303FFA5030055A00203C3FBF00",
		INIT_2B => x"5551111011111110F0332000DFFAA550F0A33000E0000AA0E000FAA0FFC033C0",
		INIT_2C => x"FF7B73C0F33333C0F30200C0CCCCCC8073322110333333300000000033333330",
		INIT_2D => x"FF000000FF000000FF000000F0332300F0332300F0332300F0332300F0332300",
		INIT_2E => x"555005505110055054400550AA8888C0055A00E0BB6611C0448888C0BB6611A0",
		INIT_2F => x"5500114051001140540011400FAA55C0055AA2E0CFAA5530303F0E1011220010",
		INIT_30 => x"555555502222111000000000000000000000A550000021100000000000000000",
		INIT_31 => x"000100010001000100010001C01FFC01AAD55FFD55FFD55FFD55FFD55FFD55FF",
		INIT_32 => x"0001000100010001000100010001000100010001000100010001000100010001",
		INIT_33 => x"0000012000010000010000010001000100010001000100010001000100010001",
		INIT_34 => x"0201200201200101000101000101000102200101200101200101000101000001",
		INIT_35 => x"0200020220020220020120020200020100020220020200020200020100020220",
		INIT_36 => x"2002002002222002200002220002000002022002002002022002000002020002",
		INIT_37 => x"0001034040000000404000000040404000000222000221000222000200000202",
		INIT_38 => x"0000000200505000020000000002030100000100000000010055550101004040",
		INIT_39 => x"0000000001000000000103001515010300000001030000000103000011010200",
		INIT_3A => x"0001010000000101000000010100505001010055550100000000010000000001",
		INIT_3B => x"0000000203005500020300000001020000550102000000010200550001020000",
		INIT_3C => x"0C30C31050920000410001450510820820001004020000010002030011110203",
		INIT_3D => x"30C30820001050D30000000411C50920410410C31C50920410000C31450D3082",
		INIT_3E => x"410D30C70C30C31810920860820821C10510410410001050100000820821450D",
		INIT_3F => x"0802002000000000000000000000000000000920450410411810100040000001"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1R_2 : RAMB16_S2
	generic map (
		INIT_00 => x"30F1101001011000F00000110100100010F30100100011010000213203102132",
		INIT_01 => x"0C0131F001010C0130F001010C0130F001010C0130F001010C0030F001010C11",
		INIT_02 => x"103333331F001010C01331F001010C0131F001010C0131F001010C0131F00101",
		INIT_03 => x"11000322110330210210110110110100000000000002110003332F2010000000",
		INIT_04 => x"30F001010C113023203102132310350350250250250240240240240240333222",
		INIT_05 => x"0C0131F001010C0131F001010C0130F001010C0130F001010C0130F001010C00",
		INIT_06 => x"108D10280C00308D03280F001010C01331F001010C0131F001010C0131F00101",
		INIT_07 => x"00F300010F00000001000001110001110F00440340330032002200FE21280E11",
		INIT_08 => x"0F101104F004F300014F101100F000F300010F101104F004F300014F101100F0",
		INIT_09 => x"F004F300014F101100F000F300010F101104F004F300014F101100F000F30001",
		INIT_0A => x"F131F131F210012100000F101104F004F300014F101100F000F300010F101104",
		INIT_0B => x"3331F3333333313203220330132211003323F2321101001F2321101001F00001",
		INIT_0C => x"131313000000000F110000000004F333333331F333333331F000033331F33333",
		INIT_0D => x"C00C00C00C00C00C0F0C00C00C00C00C00C00C02302301331313130000000003",
		INIT_0E => x"0C00C00C00C00C1F0C00C00C00C00C00C00C0F0C00C00C00C00C00C00C0F0C00",
		INIT_0F => x"00C00C00C00C1F0C00C00C00C00C00C00C1F0C00C00C00C00C00C00C1F0C00C0",
		INIT_10 => x"000671EA556AFFD3B1B6F90000E43102132031021320015F1000101F0C00C00C",
		INIT_11 => x"8E18E6F9000E796FFE55139E1AC9E1ACFD5555FD5FFFFD5FEA1ACA95311B6B00",
		INIT_12 => x"01503FFEAA95C713B9E79E646C0B2AE7956AFD5FC06D50399E1B39395FE43A41",
		INIT_13 => x"0053C040048017C000800041278DFEA01B6C0A95C4338603F540A80E4602A57F",
		INIT_14 => x"4404404484C840500100940400C3CC44800053C040048017C000800043C04480",
		INIT_15 => x"B04C4C4C40840C8400FC97C97C8140940540D7C004057CB13CB10C844480C804",
		INIT_16 => x"B0000000007CB00000007CB00000007CB000007CB000007CB0007CB0007CB07C",
		INIT_17 => x"0000007CB00000000000007CB000000000007CB000000000007CB0000000007C",
		INIT_18 => x"00000000000000000000003C000000000000007C000000000000007CB0000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"8880000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"1440244040443040434441000004000404040400004000004040404040440141",
		INIT_1D => x"4404040444020100144400000412002004004004040044040044040000050000",
		INIT_1E => x"00000000F0440404041424040401111210034401300000404040400011130410",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"010010111F0011100110100103010031F100000011100101001031F011104464",
		INIT_21 => x"F3303C35F110000110101765764756464647666554575F201000000011F101F0",
		INIT_22 => x"00000000011F1100000111001F3303C31F3303C31F110001F3303C35F3303C35",
		INIT_23 => x"1F1100000000011F1100000111001F3303C35F3303C35F3303C35F3303C35F11",
		INIT_24 => x"000000000101F10010001001010F3303C35F3303C35F3303C35F110000001001",
		INIT_25 => x"0000000000000000000000000000000000000000000000000C00000040040071",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"0333330003000000302100003130100033000000030000003020212032030300",
		INIT_2B => x"3333333021032100300000000032020030210000000000000020020023333200",
		INIT_2C => x"3000000033030100333330003020000033131310313131303202020031313130",
		INIT_2D => x"3000000030000000300000003000030030000300300003003000030030000300",
		INIT_2E => x"0313000003130000031300002000000020202100202020000000000020202010",
		INIT_2F => x"1131330011313300113133002131312020202200013131000000002000020100",
		INIT_30 => x"3333210000003210000000000000000000000200000013100000000000000000",
		INIT_31 => x"0000020000000000000000001555515555155001550015500155001550015500",
		INIT_32 => x"0200020002200200020002200220022003200320030003000020002000200220",
		INIT_33 => x"0000023000013000002002200220022002200220022002200220022002000200",
		INIT_34 => x"0033000032000003000002000001000020000023000022000033000032000031",
		INIT_35 => x"3020003110003010000310000010000310002010002110002010002310003000",
		INIT_36 => x"3000033000023000033000023000123000122000122000212000222000212000",
		INIT_37 => x"000002FFFF000002FFFF000001FFFF0000000033000030000033000003000003",
		INIT_38 => x"FFFF000000FFFF000000FFFF000002FFFF000000FFFF000001FFFF000000FFFF",
		INIT_39 => x"0100FFFF000100FFFF000000FFFF000000FFFF000000FFFF000000FFFF000000",
		INIT_3A => x"FF000100FFFF000100FFFF000100FFFF000100FFFF000100FFFF000100FFFF00",
		INIT_3B => x"00FFFF000100FFFF000100FFFF000100FFFF000100FFFF000100FFFF000100FF",
		INIT_3C => x"000000000000000000000000000000000000FFFF000200FFFF000100FFFF0001",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0080AA0000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1R_3 : RAMB16_S2
	generic map (
		INIT_00 => x"00F1111111011110F11110111101111110F01111101111111110DDCCCFFFEEDD",
		INIT_01 => x"0C1100F111110C1100F111110C1100F111110C1100F111110C1100F111110C11",
		INIT_02 => x"100000000F111110C11000F111110C1100F111110C1100F111110C1100F11111",
		INIT_03 => x"CCCAA99999988080080080080080080080080080080FFFFFFEEEEF0111011111",
		INIT_04 => x"00F111110C1100DCCCFFFEEDDCC080080080080080080080080080080DCCCCCC",
		INIT_05 => x"0C1100F111110C1100F111110C1100F111110C1100F111110C1100F111110C11",
		INIT_06 => x"184FEE044EDD140FCF000F111110C11000F111110C1100F111110C1100F11111",
		INIT_07 => x"10F001110F11111001110111111011110FDD88CF88EE88DD88CC88FFCC0CCEFF",
		INIT_08 => x"0F111110F110F001110F111110F110F001110F111110F110F001110F111110F1",
		INIT_09 => x"F110F001110F111110F110F001110F111110F110F001110F111110F110F00111",
		INIT_0A => x"F100F100F011110111110F111110F110F001110F111110F110F001110F111110",
		INIT_0B => x"0000F000000000CCCFFEEDDEDCFEDCCFDCFEF0001101110F0001101110F11110",
		INIT_0C => x"112233000000000F111101111110F000000000F000000000F000000000F00000",
		INIT_0D => x"C00C00C00C00C00C0F0C00C00C00C00C00C00C0FEEDCCFE01122330000000000",
		INIT_0E => x"0C00C00C00C00C0F0C00C00C00C00C00C00C0F0C00C00C00C00C00C00C0F0C00",
		INIT_0F => x"00C00C00C00C0F0C00C00C00C00C00C00C0F0C00C00C00C00C00C00C0F0C00C0",
		INIT_10 => x"800005550000555458054000AA55EEEDDCCCFFFEEDDD080F1111110F0C00C00C",
		INIT_11 => x"25025015A80540000555095001650016015000015555540000016555905055AA",
		INIT_12 => x"000A9500055514595554000056A59554000001556A0000155000959550009400",
		INIT_13 => x"4443C444440443C444044443E95001500056A015169940A9500056A540540015",
		INIT_14 => x"B77777BBFFFFC2802C02C0280283C044044443C444440443C444044443C44404",
		INIT_15 => x"30333FFBBB77733333FC03C03C0002802C0283C444443C303C3033FFBBF3FF3B",
		INIT_16 => x"30000000003C300000003C300000003C3000003C3000003C30003C30003C303C",
		INIT_17 => x"0000003C300000000000003C3000000000003C3000000000003C30000000003C",
		INIT_18 => x"00000000000000000000003C000000000000003C000000000000003C30000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"444C000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"0000000000000000000000000000000000000000000001000000000000000000",
		INIT_1D => x"0000000000000000000000000001000000000000000000000000000000000000",
		INIT_1E => x"00000000F0000000001020000000000200000001000000000000000000000010",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"111111110F1111110111111100011000F111101111110111111000F11110EEDC",
		INIT_21 => x"F0000C00F111110111110CCCFFFEEDDEEDDCCCCCFCFFFF011101111110F110F1",
		INIT_22 => x"11101111110F1111100111110F0000C00F0000C00F111110F0000C00F0000C00",
		INIT_23 => x"0F1111101111110F1111100111110F0000C00F0000C00F0000C00F0000C00F11",
		INIT_24 => x"111101110111F11111011101110F0000C00F0000C00F0000C00F111110011111",
		INIT_25 => x"0000000000000000000000000000000000000000000000000C44404444044471",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"0333332023321000302300003322100033321000033210003112210032033300",
		INIT_2B => x"1111111011100000300000001332211030230000000002200322322023333100",
		INIT_2C => x"3312100033232100333333003322000033322110332211003332211033221100",
		INIT_2D => x"3300000033000000330000003000030030000300300003003000030030000300",
		INIT_2E => x"0110011001100110011001102200000001122120332211000000000033221110",
		INIT_2F => x"1100100011001000110010002322111001122020032211003203100010102100",
		INIT_30 => x"1111111022221110000000000000000000002110000021100000000000000000",
		INIT_31 => x"0120012002300230030003002A8FF2A8FF2A8FF2A8FF2A8FF2A8FF2A8FF2A8FF",
		INIT_32 => x"0010001000000010001000100010000000100010002000200100011001100110",
		INIT_33 => x"1000210000210000210000000000000000000000000000000000000000100010",
		INIT_34 => x"0011100011100021100021100021100012100011100011100011100011100011",
		INIT_35 => x"1210001210001210002110002210002110001210001210001210001110001210",
		INIT_36 => x"1000121000121000121000121000121000121000121000121000121000121000",
		INIT_37 => x"203022AAAA000032AAAA002032AAAA0000020002200003200002200012200012",
		INIT_38 => x"AAAA203020AAAA203020AAAA203023AAAA203022AAAA203023AAAA003023AAAA",
		INIT_39 => x"3022AAAA203020AAAA203020AAAA203020AAAA203020AAAA203020AAAA203020",
		INIT_3A => x"AA203022AAAA203022AAAA203022AAAA203022AAAA203022AAAA203022AAAA20",
		INIT_3B => x"20AAAA203020AAAA203020AAAA203020AAAA203020AAAA203020AAAA203022AA",
		INIT_3C => x"000000000000000000000000000000000000AAAA203020AAAA203020AAAA2030",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"00C8FF3000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
