-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "8A252B57FEA42E57908010A2F9CD590AE9257FC0000000000000000000000015";
    attribute INIT_01 of inst : label is "2A16508120110704E4707E685B0013186B25774576F200209005844015C94B00";
    attribute INIT_02 of inst : label is "7FF9D0037314F13A916916BB436B45B5FAA14DC0A4811B184DA40DEED5683104";
    attribute INIT_03 of inst : label is "954872C0001541A08A986A4ACA0E65371A01AE0620257440DF5A0DA3FEF3FCE7";
    attribute INIT_04 of inst : label is "35256B0595DCBA1C2F213336C7F068B2D15F1D1A2E1562E28A4AF503FC803E00";
    attribute INIT_05 of inst : label is "A801513007F27009F7257F869030D3553DFE6407D2F7FFFFFFFFFFFFFFFDAC75";
    attribute INIT_06 of inst : label is "1D738E7ACAFF5E711FD33D177C99C99C55D69C6208811425254764107E4F0818";
    attribute INIT_07 of inst : label is "CD9FF7BE66674BA6464A36325991928C8C93B329495F26C4FFFA7F6E4E737B8F";
    attribute INIT_08 of inst : label is "0000000000000000018304A42BA64C8D50B2221934C9FFD34FFFEDE840008101";
    attribute INIT_09 of inst : label is "7E000000000000000000000DECDEE1ED240249299402320903476303C63B89AB";
    attribute INIT_0A of inst : label is "AAC6AC508E842610000013095957979784C4C4C4C4C4C3FFFFFFFFF7FFFFFFFF";
    attribute INIT_0B of inst : label is "E86567DC277C43447D888BBCF1928449BD44595D6F53C9FBD1FFF351E7259266";
    attribute INIT_0C of inst : label is "F8289C88517028BC57A3000D8A60103EF2B50A95E5E7EE212EF71088E28A0835";
    attribute INIT_0D of inst : label is "7FEFFFEFF9DF22D2055EC58B13F4258362C58A391BBBFA23033D0DB4DB4E0A4A";
    attribute INIT_0E of inst : label is "058313031314840F88914F5F1520A805C42F250F8FFFEFFBFBF7FEFFFDFF3FBF";
    attribute INIT_0F of inst : label is "BFDCFECC826858A4AFCC015E5930F3F75C3C280E069BFE67728EBAFD61280E08";
    attribute INIT_10 of inst : label is "227FB49C60E2A528BF8F0FFFFB787DE3FE3EA00A519FD6FF977F6DFC0552FD52";
    attribute INIT_11 of inst : label is "6833CCFDDDEDB65BC5B85BC5B8405027FBEB6360D8D83636001B718E7790C5F3";
    attribute INIT_12 of inst : label is "A603952A57022E5166B0B4C3514B108487AD0DB6CE6D05830313133890242A2F";
    attribute INIT_13 of inst : label is "A81027E4FD429D924DFA560D0E9144105EC5B41631C33831D5A350EBF9FC00E6";
    attribute INIT_14 of inst : label is "27FE56336E31CEC51DB230C0600C23E2CCDEC9B4959511140A18683DFDF63CB8";
    attribute INIT_15 of inst : label is "D2000C014106C2282950908020501C610389D788FDDDEDB65BC5B85BC5B84050";
    attribute INIT_16 of inst : label is "7E7F1D39FC7F551600D145A268FF3CAE75002A0220835590580B24B2C9690180";
    attribute INIT_17 of inst : label is "C0FE9C008020920026A9A14FE00E0FBA46AB4D7F06A5E011823EA60C4CA7BBB8";
    attribute INIT_18 of inst : label is "578810D9832F2DEDFFEFFFFFFBF9FEAE4F13E067CC7F98EB3B1D8026988F0695";
    attribute INIT_19 of inst : label is "AFF7FFE7FA4DA8DA2FC236C0D10344311B06063ED0FFB4005250550402621141";
    attribute INIT_1A of inst : label is "AB56AB56AB56AEAA8D47904ED1A6D9EFD339C1BEA396D2ABF9EFFFB061F2916E";
    attribute INIT_1B of inst : label is "CE7FA0CE4D3EB001543FD91FDD1BDC3FBA14694A515514557FF801EBD5D5D5D5";
    attribute INIT_1C of inst : label is "599909DDA96F97BC3E5F2DCE700373EFE7BE7FF5B1DBAC1139FF93899CFF59CC";
    attribute INIT_1D of inst : label is "222224CC332BBE6B188D6039F5DCFAEAE5B193275684762380CA82CB9904426E";
    attribute INIT_1E of inst : label is "C0B1B1B3B3FBF3598138184E0675F53FCFFDFE79DCE026B091094B090DD18D0A";
    attribute INIT_1F of inst : label is "061DCE70B3594AABA134EBFDFA40458C24055E4F258E000BBBBA111132953AF1";
    attribute INIT_20 of inst : label is "F64AFD937984D09FF7F3DEEE7FDFC0497A998DEEF6DCE8D48844109590088054";
    attribute INIT_21 of inst : label is "AEEEFFF5DB155BE6FE7FFDED8ABF37FFFD353CFFF3E7FF738701331544D67E0F";
    attribute INIT_22 of inst : label is "1044451114445111111044411111144445110446EEEBBBBEEEFBBBEEEEEEEBBB";
    attribute INIT_23 of inst : label is "E3F8E51D5AA957FEA0055AA92A8555EF76C782B67F2A9F9BFEEFBBBBEEEBBB11";
    attribute INIT_24 of inst : label is "CD4E320C8C8351A7E9F51FE1C4FFBF8DFBFA67B67FCCFE6D12B1FCF9FFF2BF17";
    attribute INIT_25 of inst : label is "FEB4FFC3F75B719B5DD6DC66D775B719B5DD6DC61B5D771B7181D775B7181FFF";
    attribute INIT_26 of inst : label is "F037539EFD198FFFB7FFB5FFDEA9FFDAFFEF0FFED7FED7FF899FBFDFFB77FDAB";
    attribute INIT_27 of inst : label is "9F1AE987F8A7C33AC6678CEB199633AC6658CEF199633F433EC335BCF7C0CC3D";
    attribute INIT_28 of inst : label is "40001BF643266C91A314259A7717D398E2CF1CF30E2FBFBFC84CE47C69E61DE6";
    attribute INIT_29 of inst : label is "000000166666666D5556AA3FFBFFFC1F18FE03F809E79E79E7FAAAAAAF803EC4";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A2A07E0800727C393E964944940793E94010C000000000000000000000000013";
    attribute INIT_01 of inst : label is "2C6CC9389F69205C96D6DF477F497F74A65C098C8245A00008038400060B0A0A";
    attribute INIT_02 of inst : label is "C1ADF99676387A0549FC9FBB91FB677DF647918F575705D1AF4B6F4B862E763F";
    attribute INIT_03 of inst : label is "42931BC979735A48153ED4997C42A8EBB1989E62EE6CBA31AA0C86C41B5BFDF7";
    attribute INIT_04 of inst : label is "51CCC5E3DE0917A24F29FD5F0BF3EF0459EF38846086163BCC19AF2555378A4C";
    attribute INIT_05 of inst : label is "914C02C398058E5900047FB3E99B1DCE6FFC60E04606AAD5AB5AD6AD5AACFF03";
    attribute INIT_06 of inst : label is "B7D5BFFC1900EE6BA020BECD61274261E80265445996F95A4F9D232BB81AF485";
    attribute INIT_07 of inst : label is "50A2FB8FABA92071119F888CF44467E22335DDD28320ADD10038A22BFFFE12DB";
    attribute INIT_08 of inst : label is "0000000000000000019C0A76E60607D4AB03F49840C00D4F701DE61DEDAD1797";
    attribute INIT_09 of inst : label is "007FFFFFFFFEFFFFFFFFEFEDDADD9C50C3BC326469308DCF5C1D68F54B3EA41C";
    attribute INIT_0A of inst : label is "D77DC2CE584FD336CB2C83C39321216128888888888890000000000000000000";
    attribute INIT_0B of inst : label is "D399BDD1B64AD3695B642B64DE304B04EAF52A3BD6E74FFDBC7FF50FBE6E3C93";
    attribute INIT_0C of inst : label is "13E44095440C79D5202C3948A48569E9A452758ECF3FF59C914F2BE507947241";
    attribute INIT_0D of inst : label is "4D9821B9B695C5298CA52A54A802F320952A56577BD1023011D2475D75D4FC19";
    attribute INIT_0E of inst : label is "22223232224EF3D0454CF8A08A99963D32700CD0C410C9B20864D9821936E086";
    attribute INIT_0F of inst : label is "4000408B50D537C19FC1A3D33E44017AFAD69D9CCF3DFE394E3B0790C79D9043";
    attribute INIT_10 of inst : label is "7081312B1D09B66410A1A7E4910A06B9F8CCD6BCCA690C0A2834C8054CE401DB";
    attribute INIT_11 of inst : label is "A54C0708889B6D2472472432466639426DB24A48929324A48CA48D6914061A01";
    attribute INIT_12 of inst : label is "DA2286CDCD8E6E33744B5210ECEACA5A4E94A165A200EA3222223261DED291CB";
    attribute INIT_13 of inst : label is "1C4918C2373BD6E032CF30E4A10296492A0AB90B2C72E73E74F8923DF8FC7CA1";
    attribute INIT_14 of inst : label is "426CE4A491AD229B212ECB1651754C311840D81983B4C33716F1A51C01EA804C";
    attribute INIT_15 of inst : label is "1B6D6A2CB7609849ADA24A52B5DAE58498C3600308889B6D2472472432466639";
    attribute INIT_16 of inst : label is "0AC16147FCFF266644CB148A06FFB6E297664F64F79831478364C24CB28CB633";
    attribute INIT_17 of inst : label is "22D797906133B46EED3093732DA82D2E8D3B84995F98770712FE432A28C88002";
    attribute INIT_18 of inst : label is "A915E30078FF40104D364D134D8A7FFA208831EB687FB8FF5A1F9177F9D7A258";
    attribute INIT_19 of inst : label is "E168B65A290874855294D2EB0074035A6937AC405D0057E23D9D39D3BD9B4E74";
    attribute INIT_1A of inst : label is "CD67339ACE6736CE7516895285EC7C29174D4AF18ED5762FF37FE09A080AD8CA";
    attribute INIT_1B of inst : label is "9920CC99A613000198B67C5F785F78B6F204284A15155199D55155F3E799E799";
    attribute INIT_1C of inst : label is "A666F736B18C37FC8924D2338C5CC924926926943326D23EE4833AD572418920";
    attribute INIT_1D of inst : label is "50000E0180FD0C1BEA4611D65B4B2D03520C38F1BAB10D08246D2527A88BB195";
    attribute INIT_1E of inst : label is "140607040516AD807A2D96C944A6C60080080580804C7C63CE3CA63CBA38C42E";
    attribute INIT_1F of inst : label is "2FA011844C956FB8AC40345A2922F233CB648532D823C01EEEEFEEEE2FFE7B88";
    attribute INIT_20 of inst : label is "091A024705B15620582C0B058160B8E3AA5660522D823F3B64CB394FFCA7A529";
    attribute INIT_21 of inst : label is "14146107B334E45000F032D99A42800646564A00645000E1DFF48334A6782E60";
    attribute INIT_22 of inst : label is "AEBEBEFAFBEBEFAFFAFBEBEFAF91041415050140141050514145051415414505";
    attribute INIT_23 of inst : label is "2F190C83173A66E66463173A4ECCC4C952F7A640806522A00EEBAFAFEBEAFAAF";
    attribute INIT_24 of inst : label is "7F9E86F1E1B81813E40514056000DEE507E4F1CA0001FEC37FF6001601F9FF3B";
    attribute INIT_25 of inst : label is "09CA017804A58E4581296391604A58E458139639658344A58A48344A48A48308";
    attribute INIT_26 of inst : label is "24A0320817503C065E065E0206E4012C01036009600960185061A0D025E012F0";
    attribute INIT_27 of inst : label is "23AD951401C48A01140028205040A01140028205040A0A2A0AAA07B044929011";
    attribute INIT_28 of inst : label is "12D2AD2494386671C91A3165558A266A8532560AA86AA33FD19E87079415516B";
    attribute INIT_29 of inst : label is "000000122222222CCCCEA8BFD36DB95652D403500CB2CB2CB2FAAFFAAD2A1691";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "22285C2E0A3020A8348410229F42834868007FC0000000000000000000000001";
    attribute INIT_01 of inst : label is "2024C8181E69089A80F0FF1417431A143A0F0047038180418807860007D4880A";
    attribute INIT_02 of inst : label is "8717611553287E10B673670191FA557A774E06061431034001034149D164341F";
    attribute INIT_03 of inst : label is "0D831C98889090C805FC0C180C4043C42798A462921406B53C3C86C4762EA95D";
    attribute INIT_04 of inst : label is "DFB46A65DA01158D18DE4472B4091A1C31B3BC0DA0CE7F3860184A6154334A4D";
    attribute INIT_05 of inst : label is "82CEA8449D50B294211BD52CD562FB419FF9BC22744AAA54A94A52A54AACDE4D";
    attribute INIT_06 of inst : label is "3E81B6B418F0913B8E312F9DAB93057174CA1464591F990A0E56830BB890C42D";
    attribute INIT_07 of inst : label is "0A06920826752BF2923C9091E4AC8725643BB33083002545F03288436318281E";
    attribute INIT_08 of inst : label is "000000000000000001050634A33216008118D0C846420B46DE1567C90A0A0406";
    attribute INIT_09 of inst : label is "7E7FFFFFFFFEFFFFFFFFEFD46D46C410C35C9061FA76BFC27551095C589EA02D";
    attribute INIT_0A of inst : label is "088A1EC63E063750904009C3831CFCBCA8EAE2E0E2E0D3FFFFFFFFF7FFFFFFFF";
    attribute INIT_0B of inst : label is "2CB9A6F492DA40005B6D99A68D3013C5E0E50A2002A54B531D540B3C10D63C34";
    attribute INIT_0C of inst : label is "13A07E268A1B248501939CA0A031DCC71529CF7A4B2D43C56EB808E945965BEE";
    attribute INIT_0D of inst : label is "FBDED7FF7E63C99B84718B162E018120C58B168F570CFDB1DB88FC71C712EC18";
    attribute INIT_0E of inst : label is "02B3A3838344A1CBC6DC61978DB88E19D0360C4BC76BFF7FB5FFBDED7FEFFB5F";
    attribute INIT_0F of inst : label is "E0EC7977C0C551C18FC2619D19443126288B8C0C0739557A7FEB3FFC440C0080";
    attribute INIT_10 of inst : label is "70BD73A7DCA5B66003F73D4348BE5C6F5032118CC2C3FBDCB3D9AF8544647052";
    attribute INIT_11 of inst : label is "A10AC75EFEDDF734E3CF34A3CB332B6FFEDF6F69DBDA76F6CCB795AA35060209";
    attribute INIT_12 of inst : label is "3F22F9E2DB2648634631D01F9C434202067423B7C66FE703B383A378D694AAC2";
    attribute INIT_13 of inst : label is "0C0009234A0AE6E246A52C74218082D92B83290155F57F55F0F1EFDD55A818BF";
    attribute INIT_14 of inst : label is "6FF6BEB7FAB5468265B41BD750751AF15402D019812450730C69A11C01EAE17C";
    attribute INIT_15 of inst : label is "40016A1981408A28296206948456A1240B5BE3835EEECDF776E7EF76A7EB332B";
    attribute INIT_16 of inst : label is "169F4F5BA86A07240E81C0E0AEFF80E1F102436436081575D07EABCE28A10685";
    attribute INIT_17 of inst : label is "232F0F388239960E65A08044692E329EC5A28423573D67A51AB4A00E2AE95DDA";
    attribute INIT_18 of inst : label is "24A5201DBBFB4FAB966F16459BCF80000088B186CDD52BB4337619551947E29C";
    attribute INIT_19 of inst : label is "A0A450281085DC5DC4A4906A1B746F744800AA049A116621169A09A0A4F28268";
    attribute INIT_1A of inst : label is "F17A3E1F0F87C6F23DC2801CF0B44FAEF673729CA71747C3FCFFC01A08E29062";
    attribute INIT_1B of inst : label is "DAAA00FA1737F3F9E017490B490B481692046942155110DE599199C3F99F87E1";
    attribute INIT_1C of inst : label is "135BDB50002037684A8509AF7C36D545028AAA42A152F60B6AA83B51B55089A0";
    attribute INIT_1D of inst : label is "17776AEFBB5F0C91AA07F0C828441408283DEBF6BC21E94803014902AC86D8D2";
    attribute INIT_1E of inst : label is "F415141D1C0A141DF8341A8D66BAE55E61E6F29E6F2C3E22062062207DB8C50A";
    attribute INIT_1F of inst : label is "074EF6B456C149A80846D42910A0E9AF6A34020149ADC00AAAAAAAAAA52E7A82";
    attribute INIT_20 of inst : label is "801EE007702104273B9CE7739CEE783382037C20149ADDBDE05200435001000C";
    attribute INIT_21 of inst : label is "01546951EA143622F2F089F50A2117CE536364789223E00008A22A04622C0E47";
    attribute INIT_22 of inst : label is "5401540550154055055015405511040401004014015005501540550154154055";
    attribute INIT_23 of inst : label is "28130C0EBF05785B4BC6BF0570796B49AEE7A600C269B421F441010040100500";
    attribute INIT_24 of inst : label is "729E06C1C1B49D0AA0003F00F0609FCACFD4E3F6380103A7581DC488F9F0DE1B";
    attribute INIT_25 of inst : label is "F4E3FE8FF37BB3B83CDEEDEE0F37BB7B83CDEACEF83CB33BB3BAEB37BB3BAB08";
    attribute INIT_26 of inst : label is "34955AF69A48ADF981F983F918E7BCC0FC8C3DE607E607F5B3BF5F2FD817EC1B";
    attribute INIT_27 of inst : label is "9BF6DCD208E209585232A541488A91052A2A4654ACA91829582911D7B0FA44EC";
    attribute INIT_28 of inst : label is "9B6349BF62ED44A4A71C90B73FDFF7F343BF7DB9A42E19EA909E36DADB7249FD";
    attribute INIT_29 of inst : label is "000000122222222C4446A8EA9E9251E47C984A612B8E38E38E3AAAAAA9C57599";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "082D75D20A30228D131141741994C11168805400000000000000000000000041";
    attribute INIT_01 of inst : label is "C63061D8FCB62254A5757017242B1120DA4B08DB0184C0200003064017FFD554";
    attribute INIT_02 of inst : label is "671095D3BA9D074A93C93CFDC08D56C974E7E04286B28642A048E000B2D1530B";
    attribute INIT_03 of inst : label is "26415B75012627A404A9AE0B87050310364091125059D0659A3E41D67421FEC2";
    attribute INIT_04 of inst : label is "2741CC66938C10A24B0845AB44058B7C4920B986AD775360260B48C6A85E1568";
    attribute INIT_05 of inst : label is "BACD50149AA00AE94209FF94A8A1141ED9FE15A0340555AB56B52952A554C955";
    attribute INIT_06 of inst : label is "5E7439C68B0811138110C6AA8342FC7D47D2479FCD5A6C0904D8624FE69F90AC";
    attribute INIT_07 of inst : label is "08141041098A738EBE9074F583A7A41D7D64CC3841705C8408062260BDE6982E";
    attribute INIT_08 of inst : label is "00000000000000000207823023B00616A5181544360086C0810A26294A51C5C6";
    attribute INIT_09 of inst : label is "0000000000000000000000303F077060A2FE082DC6863C2001701714298B8C2B";
    attribute INIT_0A of inst : label is "66D79A583327841000490800C17CBCBCA2C0C0C0D0D0C0000000000000000000";
    attribute INIT_0B of inst : label is "4562D96EFBEE9269FDF7D6C96E90C2413EE1780EFE3341FDE97F90B32CB39A06";
    attribute INIT_0C of inst : label is "896D12278C2B155C7093F5618E14A525910D7653C127F2FDC5660AC91453416E";
    attribute INIT_0D of inst : label is "7FCEF7CFF873298254708D1A33018194468D1B4A9DCD0C1587C97B6DB6D2F60B";
    attribute INIT_0E of inst : label is "19D35353530611CB4410639688228F1DE92D05CB477BEFFBBDF7FCEF7DFF3BDF";
    attribute INIT_0F of inst : label is "D0EC44ED60737C60BFFDF1DC18303127BCCA0C0C9599FEF771AB32FC748D2000";
    attribute INIT_10 of inst : label is "3082D1A548C53B2D03160FF388B05852FE3CD7965855B2EC96DB2DC101D00808";
    attribute INIT_11 of inst : label is "EC0AC2E677769295A95B95B95ABAA7679E7DA92B6A4ADA131BF2B48A2082930A";
    attribute INIT_12 of inst : label is "2A9C3952ADCDEE2E7E35F606146FC283263D82DA470D1E535353530AC6118BA0";
    attribute INIT_13 of inst : label is "0E241B7E580A801A4581A56D8080BB6DB482FC840900B41905D3C493FB55030C";
    attribute INIT_14 of inst : label is "67923216D2914412B6971952586C02D0C421586C85A1F6EF8FEDEC1FDFDE0C20";
    attribute INIT_15 of inst : label is "430DA30A810016E1847242B4AD5682958B18F3C4E7666692B4AB4BB4BB4ABAA7";
    attribute INIT_16 of inst : label is "165E2F1B549526B64CCB8DC642FF5D62D225E0DE0C011116D04A28A29A218486";
    attribute INIT_17 of inst : label is "4E2B695679BD32EF4898B51C619EE2DE5893C5E30938270550CA7E7E81415DDA";
    attribute INIT_18 of inst : label is "37850519832104DDB64BB66D92E32AAC0280751E9F3FDE48F7C95D3A54C06049";
    attribute INIT_19 of inst : label is "67A9C4E371A58658673ABA53D30F4CC75D50CEF683DDA0711A4B0CB0A168C36C";
    attribute INIT_1A of inst : label is "FF823FE20FFA06FEFD8FB8CEE3FEAECAB447C37F9A37B44FF6CFF8B020184455";
    attribute INIT_1B of inst : label is "CBAAD2CAA53E9400007FAD3FAD3FAC7F5BF7EF7BDDDDDDC061F21FFDC19FF981";
    attribute INIT_1C of inst : label is "A5AE295677BD9016CAA552B7BE1A5D751AEBAACC5356AF0D2EA20B0597518182";
    attribute INIT_1D of inst : label is "166660CC330A8A3958C5387EEB7F7519EA39C326160032420301030008C3416E";
    attribute INIT_1E of inst : label is "C4747C7C747A75999130994CA66FC65E45E6F2DE6F2E1A36C32C232436B0856A";
    attribute INIT_1F of inst : label is "D86ED6B43A6C23598034CDEA71B192B7B4C98E27518CAAEAAAAAAAAB210F239A";
    attribute INIT_20 of inst : label is "420D10828C00C0172B96C562D8AC5C2684C508E37598CA9681435A468D63EB1F";
    attribute INIT_21 of inst : label is "1554CA4B9729B2231E4C89CB94C118AC9339644C92225015482A6339B34AB900";
    attribute INIT_22 of inst : label is "5555555555555555555155455504515154555555555555555555555555554555";
    attribute INIT_23 of inst : label is "EC43E582BF002AFF4012BF002AFD401C6D4F9CE2232CBF914114545515555555";
    attribute INIT_24 of inst : label is "D2491C555551BB8964448894C01000EF022641A40444FE691FE224889401503E";
    attribute INIT_25 of inst : label is "035AC06B00444441B00111106C0044441B01111101B060044044A60044454E10";
    attribute INIT_26 of inst : label is "1D3194930A98CC84110413044155820A8220AC1054105400398010184118209C";
    attribute INIT_27 of inst : label is "8D965D970CDF331F263E4D7C9AF135F263E4C589AB935193119319449874D726";
    attribute INIT_28 of inst : label is "9BFBF640019B24C6CA4A779773C9B1B0F1894C9BAF27CCFFC4CD8E4A59375CA5";
    attribute INIT_29 of inst : label is "000000144444444BBBBEA8FFE32491FB80E04B812861861861DAAAAAAE000B99";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "D4A077F14B72562C36124916105AC36110A2954000000000000000000000002A";
    attribute INIT_01 of inst : label is "0470E918BAB8201213030C15340924309702A94AA154204110078200057D1477";
    attribute INIT_02 of inst : label is "510119931019661303C83C288440328FF5FA000A021380C1FB68FB685260622D";
    attribute INIT_03 of inst : label is "A1D31881050286EC34798E9917408A19B4201480414089EF8BA6C0D11602AA84";
    attribute INIT_04 of inst : label is "724084E2822040A1490AED0D1875AB2E042230805C1613832C010805FCB24E58";
    attribute INIT_05 of inst : label is "114EA8039D5006452108D5552AAD450A09FA14942AAAAA54A94A52A54AACE122";
    attribute INIT_06 of inst : label is "C00714A4815401B1C2836E03B1268A388972E304F397484240CA89298699A2AC";
    attribute INIT_07 of inst : label is "A950414514457095B5B0A0AD8565642B2B2AA2B2902AFDA055140381B5AC65E1";
    attribute INIT_08 of inst : label is "000000000000000001158B7B4E9B0740A91D15EC33406BD6C6D76ECD7B732DA6";
    attribute INIT_09 of inst : label is "0000000000000000000000071071108AC10C920448948C72401982060DD00412";
    attribute INIT_0A of inst : label is "1110D008544E486400000D149020000000829092808280000000000000000000";
    attribute INIT_0B of inst : label is "31040049009125B20240248001B04A9A90823A839CA103552C5544A114530248";
    attribute INIT_0C of inst : label is "5B642534106E9A4D20047BD3A40F2B600021144A420D5034B3026BD45575D709";
    attribute INIT_0D of inst : label is "208400841000252418A13E5CB8A2D2049D2A55C017405114208745D75D700401";
    attribute INIT_0E of inst : label is "590A024A420A12900B2094201643172E824A40900A0044110022084008821002";
    attribute INIT_0F of inst : label is "6A00A88871AF2B4812D472E820750698B3C0152C91055435A1140448BC952082";
    attribute INIT_10 of inst : label is "3395F4601F39720460C14550060F840055439CE6C801248960805925A0811609";
    attribute INIT_11 of inst : label is "8454088EEECDB7EE2E62EE3E6233216D36DB6B7EDADEB736BFBCC5AAB1201AAF";
    attribute INIT_12 of inst : label is "CDD54E5CBE5D4BFB5873C28864BC4EDA06D089B6C50138CA0A4202135AD7BE8A";
    attribute INIT_13 of inst : label is "96401CCF343B0006C4493A708816B24B7A4B2D8DA81A81AA09C2952150036150";
    attribute INIT_14 of inst : label is "6D7F3FF718B5461BA5B4195B59605402A02004282220D3FF9C61845FC00EE600";
    attribute INIT_15 of inst : label is "8925A33AB682326384F24E529C9A2304C852F8089EFECDFFCE2C62CE3C623321";
    attribute INIT_16 of inst : label is "4341A18101C07FB4DC9B219000FFC2601323C67C670C25610176836830C49713";
    attribute INIT_17 of inst : label is "2E2F6772CBFDF2DD7CB017744D92E2CE5CBA80A21F1D43A670E0D7708A680000";
    attribute INIT_18 of inst : label is "BB554100306A812300B600802D880002A8AA34DAD255548ED491993180D66ACD";
    attribute INIT_19 of inst : label is "636BB7DAE96012013000BF6242C108325E1D8C12014480F328592D92A9284B24";
    attribute INIT_1A of inst : label is "FFFFC2020FFFFF020923C20488E6080A1811C01403040007F04FD2F844484CBA";
    attribute INIT_1B of inst : label is "8964A0893E5327FDFD1E0C8F0C8F0D1E1BF7EF7BDDDDDCDFC1F81FFFFFE18181";
    attribute INIT_1C of inst : label is "2CB021257B5E0000E93C9758C6584B2CDE5964AF0B27CB2C259A9A0512CDC902";
    attribute INIT_1D of inst : label is "54444800804DA6BD9A465977D2BBE9E9D28008609B205B486F6D6F6EC1CB052D";
    attribute INIT_1E of inst : label is "00AE26262636EDC030205108942647860060300603065C564B64A524BB1CE12C";
    attribute INIT_1F of inst : label is "58200000A8342598C81010DAE972B35886E0EDBE9441335FFFFFFFFEAD6F638C";
    attribute INIT_20 of inst : label is "AE1DAB86D62064010080201004020CF2A25411DAE9C4121A448B594A0D656B2B";
    attribute INIT_21 of inst : label is "EAAB6D6710A4B64256CADB88507212CF5B63686AB7436AB07A6F70A4FBAE1942";
    attribute INIT_22 of inst : label is "AAAAAAAAAAAAAAAAAAAEAABAAAEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABAAA";
    attribute INIT_23 of inst : label is "EC03EC82BF002AFF4002BF002AFD40094808446A9B649C357AAAAAAAAAAAAAAA";
    attribute INIT_24 of inst : label is "42010142525498380D06501C6208B1FA923EC3A94B6DAA703D52D5D0D983D07E";
    attribute INIT_25 of inst : label is "40C2080820A64A66A8399299AA0E64E66A829F29A6AA40A64E65040E64E6538C";
    attribute INIT_26 of inst : label is "361524361B0A8C946094629400C40A304A002051825182501005029106048312";
    attribute INIT_27 of inst : label is "9B92D8C28DD08115023805540AE011402BA055408E81140114011201B0D8576C";
    attribute INIT_28 of inst : label is "6404000000009F070C6CA01227DBB3B0559B59B1854C19EA8D8426DA4B6309C4";
    attribute INIT_29 of inst : label is "00000011111111180007FF2A82001E000080020008000000001FFFFFF80000E6";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "03D0280337727E5081134D16548518111806FA4000000000000000000000000B";
    attribute INIT_01 of inst : label is "E46601F95AAB2492D2727A35A4692E2690224D4A052620008800020000800028";
    attribute INIT_02 of inst : label is "C86435D68BB0AE6101981945021032007000100A16121549A54C654C92C7522D";
    attribute INIT_03 of inst : label is "10183A0D4D5282C1B6098CC11C1896187C1D947653549969C2EC18E484C8ABD0";
    attribute INIT_04 of inst : label is "3694C422767829B1620856529B8542A7077D28904A9633136C414A3554166AC8";
    attribute INIT_05 of inst : label is "115EA822BD505245A529D5644B26484DFFFC1488A13EAAD5AB5AD6AD5AAEDC00";
    attribute INIT_06 of inst : label is "1C559EF4C1950F659A403FAFE75FE8F8C94248D54573582620C88D2984DA06B0";
    attribute INIT_07 of inst : label is "E5C841451111B604747022A3811D1C08E8E8003318298A9C94D624E14A521B0E";
    attribute INIT_08 of inst : label is "0000000000000000011D0B7B65D647CEBD3B16593AC85F63CABDF7472933048F";
    attribute INIT_09 of inst : label is "000000000000000000000004EC4EC491450CD3070088642B43B7620DFBB2049A";
    attribute INIT_0A of inst : label is "3308B0C8516E4832496D9B089823030301839193818380000000000000000000";
    attribute INIT_0B of inst : label is "30C00049240000049240001225025A02F58E2054AC60815448D54CE114460609";
    attribute INIT_0C of inst : label is "70448D15042AA2B023044256046842B8E0950CD620055C24B2C22BD49C51C1D9";
    attribute INIT_0D of inst : label is "24052804819C65240CA00C187292F30204083371157195F23DA14555555C2C41";
    attribute INIT_0E of inst : label is "254E460E060F92940320D0680241962C8B6A60B4029404814A024052809014A0";
    attribute INIT_0F of inst : label is "63102110520120CC12D7E2C83040C09831F014924F0755952109E048F4949249";
    attribute INIT_10 of inst : label is "B4657B5865295604AC080D5CF240218354CE14AC090124880082492F9480D449";
    attribute INIT_11 of inst : label is "846D008AAA8925042042042043AAA96D24925A48969324246AA0858E53305A99";
    attribute INIT_12 of inst : label is "0E4F0840AF377AAAD475C2C004FA4ADB6F508D248B98080E4E0646035A569A8E";
    attribute INIT_13 of inst : label is "1C6D2842102B80048810AB708E02D24932DB68351611410617C68B0156A863C0";
    attribute INIT_14 of inst : label is "6D24242410B1CA5B29252F9F71206500A401A5F8332CF3331575847FC0081480";
    attribute INIT_15 of inst : label is "0925E628B7A5B65BE4FA4A7394DA58D4EE20B4008AAA8925042042042043AAA9";
    attribute INIT_16 of inst : label is "206030A0A9AA7BBCD599FCFEEEFFB4F7A226C66C6512358289C1441441049C12";
    attribute INIT_17 of inst : label is "BAD70516DB5560F7583117728D89AD0C183688941D5DEBB736F467E8CDE62220";
    attribute INIT_18 of inst : label is "A1559273060FB21020022008009ED552ED33B94889157A1A42435D689D9AE65D";
    attribute INIT_19 of inst : label is "B1308A4526BB03B01800D2E36481900269328A4129004A6330692F92B22E4BA4";
    attribute INIT_1A of inst : label is "FFFFFFFFF2020602FDFEFBDEFFBCFFEFFF6F7BFFBEF7F7EBFFFFE49C812E4CE2";
    attribute INIT_1B of inst : label is "80011380428847FDFDF7F9FBF9FBF9F7F2042842111111DFC1F81FC1C1818181";
    attribute INIT_1C of inst : label is "C000000A000500429040600004500010282003424A184A28000D562700060F03";
    attribute INIT_1D of inst : label is "5888819866053CDBC04891524D0926194D63060C02A48D696F6D6D6FD98A0804";
    attribute INIT_1E of inst : label is "002DADADAD9126B3046270181C06172182190C2190C4507A4BA4A7E4A019DB2E";
    attribute INIT_1F of inst : label is "C8310840204725ACA999804C26A28000122CB4526B1816C0A0A00A0AB2960369";
    attribute INIT_20 of inst : label is "B8456E10B5A65488C461188C231188B6B65800452231800805CBCB4A0F25392A";
    attribute INIT_21 of inst : label is "155575AE94AC80CC600B124A56466157680A58B324C4A9F3CC2334ACEB52610C";
    attribute INIT_22 of inst : label is "5400015550001555000155500001500554001554000555500015550001555000";
    attribute INIT_23 of inst : label is "8EB7009ABF002AFF4002BF002AFD400B99A06E445405238E9501540055500055";
    attribute INIT_24 of inst : label is "6F012F49C9D6BE1A8496B25760AB2062F03404762A00A8694D4259312B036068";
    attribute INIT_25 of inst : label is "E6F39C8E72106110E4841844392106110E48418410E6925061064921061063CE";
    attribute INIT_26 of inst : label is "A506B32552835F5D1E3D1C3871D71C8C1C38B8E460E460F11F0F67239061C820";
    attribute INIT_27 of inst : label is "13A49020B5C9D062A0C540AE8155063A04540AE81550295029502BD92A94184A";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFC07F070C22415AAA2AC1512D520416A516ABD83FE9692418169";
    attribute INIT_29 of inst : label is "000000100000000800040000020010000080020008000000007FFFFFFC0881BF";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "A8002AAFFF291428144924711BC6914468923FC0000000000000000000000038";
    attribute INIT_01 of inst : label is "93246C9C3C30924DB9E9EC8394E589964E81D1A1D8CC00200802800002028A00";
    attribute INIT_02 of inst : label is "F733B13E607A6A9936DB6D3088578800000000605C584264E198A19868352986";
    attribute INIT_03 of inst : label is "62B191EC2C285D8640DE358C95248918B25447511B1A48E59A1C61A3766755CE";
    attribute INIT_04 of inst : label is "7C8A50A97A28D5E2C4214632D8020498CBB31A62EA4E732E598C63B3545E9BE8";
    attribute INIT_05 of inst : label is "CCBC009958011F3B52CF2AE6473628A7FFFECA101326AA54A94A52A54AAEAA97";
    attribute INIT_06 of inst : label is "7A5D34A58CFF61214F91AC133820C60E18C760044112688085A33AC7A7A91668";
    attribute INIT_07 of inst : label is "B9706186199B33030306111830C8C986464444D6B19FADB4FFCA39608003A93C";
    attribute INIT_08 of inst : label is "000000000000000000C3212913930564C9C90D4C3260F9665FF575FAD6DC9F1E";
    attribute INIT_09 of inst : label is "00000000000000000000001C6DC6C8C61A7D863183063020090909030E909341";
    attribute INIT_0A of inst : label is "B312C8610724C489B6920922B18D8D8D92D0D0D2D2D0C0000000000000000000";
    attribute INIT_0B of inst : label is "B12492000000012492400000121D30C19282898297A04AAF2A2B6411C70A17A4";
    attribute INIT_0C of inst : label is "F0F33CE1860041348D24294E91A529ECB0C61732012AB6361163C68E0C304724";
    attribute INIT_0D of inst : label is "36C6E6C6D8D7786272042C70B7F85818163858594EDBF29CF232020828A6158C";
    attribute INIT_0E of inst : label is "808B030B032248330112192602264284C904C633037366D9B9B36C6E6CDB1B9B";
    attribute INIT_0F of inst : label is "3ECC7E44D8318C58CE4FE84C821230D8B3D842412710AA433090306E2F424104";
    attribute INIT_10 of inst : label is "213F38CCD1CD1A333BA73AB6DB3A1CEEAEC056B4660CB265B2D924FD8A037CA4";
    attribute INIT_11 of inst : label is "30CCC06CCCEDB6319319319318222D65B6DB7370D8D836B698B631BBB86321F9";
    attribute INIT_12 of inst : label is "242591020E844E2277005982922321B1263619B6E50C0C0B0B03031E310C485A";
    attribute INIT_13 of inst : label is "45240160DB860016F6A62466188C5B6DBFF138C31911910914800C82A954C965";
    attribute INIT_14 of inst : label is "65B6B6B6C63777211DB0D7EED414C4C06C001CA8E8C209114061B0D5555A0C20";
    attribute INIT_15 of inst : label is "E492F2804C80410692532129423100064B1913406CCCEDB6319319319318222D";
    attribute INIT_16 of inst : label is "1AD96DD95755C227A6F3FDFEEEFF95767992B22B21C18B38E49871871C7249C8";
    attribute INIT_17 of inst : label is "402E0E21861173845CE6CDD47B0E029A74E3B623341B436C01AB0A2FB8519998";
    attribute INIT_18 of inst : label is "04C26899830A8CDC96CB96E5B2F9AAAFBBEEE82ECDEABBD9737B13E643F6B32B";
    attribute INIT_19 of inst : label is "35C4E0783C21C21C00031A44C3030C198D9097248C996328825C84C84C692172";
    attribute INIT_1A of inst : label is "0102020202020602FDFFFBDEFFFEFFEFFF7FFBFFBFF7F7EFFFFFFF9004F92623";
    attribute INIT_1B of inst : label is "C69E52C7116497FDFDFFFDFFFDFFFDFFFBF7EF7BDDDDDDDFC1F81FFFFFFFFFFF";
    attribute INIT_1C of inst : label is "010908F00005115627838084250334D3C9A69E4238E226811A790B018D3C8580";
    attribute INIT_1D of inst : label is "866660CC330365A909313418700C380470318306061032C498989A9AC4A04A47";
    attribute INIT_1E of inst : label is "C0121213135C3C198432580C164AA918C58CC658CC650713A17A117A0494A091";
    attribute INIT_1F of inst : label is "35CCC630134490CD8630C1713C28008424426783818C0E35DF755DF7452C2418";
    attribute INIT_20 of inst : label is "FD09FF42FC10C2166332CC66598CCA00413198713898C0849331362174D02680";
    attribute INIT_21 of inst : label is "FFFF9EE33382373BFA4FDB99C139DFF9BB61677FB73BFFA14821138263EC2937";
    attribute INIT_22 of inst : label is "FFFFFEAAAAAABFFFFFFEAAAAAABFFAAAABFFFFFEAAAAAAAFFFFFFFAAAAAAAFFF";
    attribute INIT_23 of inst : label is "B861466ABF002AFF4002BF002AFD400E6420651A7E31B695FAABFFFFAAAAAAFF";
    attribute INIT_24 of inst : label is "B289D3E6F6F919C172740FF4427FB025F23C537D3FA056E102B7FDCEFE86D0DA";
    attribute INIT_25 of inst : label is "C94AF92BE4A4CA4799293291E64A4CA479929329279964A4CA4D964A4CA4DCF7";
    attribute INIT_26 of inst : label is "30B981B7185CCDF27BF27BF3E445F93CF9F22FC9E7C9E7DE5D9DBEDF67BFB3DF";
    attribute INIT_27 of inst : label is "CF36DD97FC820BD017A02F445E88BD917B22F605EC0BD60BD68BD82DB8C2E46E";
    attribute INIT_28 of inst : label is "00000000000007F8007F04B6675B3B32F18B19BB2F0D8D957C8A26DADB765DCD";
    attribute INIT_29 of inst : label is "000000100000000800040000020010000080020008000000007000000FFE8780";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "00A80003FE202000048000600BD410483A007FC0000000000000000000000011";
    attribute INIT_01 of inst : label is "A2002810102102C420B0B10604C50D044A01408100A420000800820000888A2A";
    attribute INIT_02 of inst : label is "B292A31C2660081B3713711300150000000000405051068060082008E0160100";
    attribute INIT_03 of inst : label is "021011682830D18001C43080B8059B09E65803600A0C49ED343001A32925550A";
    attribute INIT_04 of inst : label is "449C21B040280D020C630220C8070E985C108422524E6308408063A2007B11EC";
    attribute INIT_05 of inst : label is "0828001070001A28424D2AE64F3669C009F8C809100400000000000000068616";
    attribute INIT_06 of inst : label is "2C54210880FF61010FB185040801440448C31044411030404081080500301420";
    attribute INIT_07 of inst : label is "00006186199B23020206101030888984444CCCC2101F911CFFCE21E0A10A2816";
    attribute INIT_08 of inst : label is "0000000000000000018300202990040489080440B200F0641FE035E210089C1C";
    attribute INIT_09 of inst : label is "00000000000000000000000C24C25C508828820181863020010109010A82010B";
    attribute INIT_0A of inst : label is "B316D8000204CC54920008031004848486C2C6C0C4C0C0000000000000000000";
    attribute INIT_0B of inst : label is "B12000000000000000092492160400C343060023190132AA2C2A6431E78C04AC";
    attribute INIT_0C of inst : label is "E0813D818620E3B0052C6B9C00AD6BC49042361840CAA214136300980C104A2C";
    attribute INIT_0D of inst : label is "36C662C6D8524066040C6CD9E3F00100366CF0886889F2A07633038E30C23880";
    attribute INIT_0E of inst : label is "01830B030B0680310330496206608204C02C4011033166D998B36C662CDB198B";
    attribute INIT_0F of inst : label is "3E443E44C0310C880780604C16001049A78800000004AAE73081306C64000000";
    attribute INIT_10 of inst : label is "203E18C451CD1C011922AAA2C9138A4AAA40D398021DB2ED96C92DFA8C007CC0";
    attribute INIT_11 of inst : label is "004C40E4446493319319319318222D259249313048481292989630A2202001F8";
    attribute INIT_12 of inst : label is "262311020B044422220000829069000006600892470C0403030B0B0800802808";
    attribute INIT_13 of inst : label is "0C000160D900801244222C4009804B6DA4C110071911911915820582AB5408C5";
    attribute INIT_14 of inst : label is "25929292421444011C901EFC10804C40C40088902184011100410058D8D00C60";
    attribute INIT_15 of inst : label is "524BC2000500800AA01200A5214090844B181100E4446493109109109108222D";
    attribute INIT_16 of inst : label is "088844C8541502220441008000FF95B6644AA92A90A51814520A28A28A2920A4";
    attribute INIT_17 of inst : label is "682A18020811660459820005400682B8C181102A00102201020A8C4400888888";
    attribute INIT_18 of inst : label is "0D81249983010DDD92CB92E4B2F1AAAC0300E86524AAA153292A31C2F30088B0";
    attribute INIT_19 of inst : label is "B5A0C0683021821810029A42C3830C014D500AAD88BB222013480580244A0120";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFE0902800480A4080A1001401402040003F04FCF9000FA0061";
    attribute INIT_1B of inst : label is "C61A00C6836DB7FDFC16080B080B081612042842111110C07E13E1FFFFFFFFFF";
    attribute INIT_1C of inst : label is "91090CD210810E5426934884240230C30186180010D06E01986843218C342190";
    attribute INIT_1D of inst : label is "066660CC330628890013701A610D3080613183060E0260000808080808806A46";
    attribute INIT_1E of inst : label is "40101011115A309984B2182C064C01084484424844240632016003600C929002";
    attribute INIT_1F of inst : label is "410442103245006D8030C1683020008420040613098C01E0888A088900041818";
    attribute INIT_20 of inst : label is "F402FD017C00C0522112442248844802021118603418C08CC041400045002800";
    attribute INIT_21 of inst : label is "55559EE421041362FA37C910823B17F9B9232C7F9363FF014001110442C42607";
    attribute INIT_22 of inst : label is "5555555555554000000000000000055555555554000000000000005555555555";
    attribute INIT_23 of inst : label is "0170002ABF002AFF4002BF002AFD400E24A062007E009685F554000000000055";
    attribute INIT_24 of inst : label is "A006108606211BA5497C5BF4407F6F25F1D822563F8054A022A5FCD8FE780F01";
    attribute INIT_25 of inst : label is "C94AF92BE4A68A663929A2998E4A68A663929A29A63964A68A69964A68A69CF7";
    attribute INIT_26 of inst : label is "1031119208188DF663F661F78445BB30FBC22DD987D987CE519CBE5F2637930B";
    attribute INIT_27 of inst : label is "CD124D87F882831106220C40188831006200C401880316031683112C9040C424";
    attribute INIT_28 of inst : label is "00000000000007FFFF80049363491910E0898C9B0E078C957802A64849361CA4";
    attribute INIT_29 of inst : label is "0000001FFFFFFFF800040000020010000080020008000000005000000C09FBC0";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
