library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_arith.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM is
	port (
		ROM_nCS :in  std_logic;
		ROM_nOE :in  std_logic;
		ROM_A   :in  std_logic_vector (16 downto 0); -- Address input
		ROM_D   :out std_logic_vector ( 7 downto 0)  -- Data output
	);
end entity;

architecture behavioral of ROM is
	type mem is array (0 to 131071) of std_logic_vector(7 downto 0);
	constant my_rom : mem := (
		x"3E",x"00",x"32",x"84",x"7D",x"C3",x"66",x"02",x"3A",x"07",x"60",x"0F",x"D0",x"33",x"33",x"C9",
		x"3A",x"00",x"62",x"0F",x"D8",x"33",x"33",x"C9",x"21",x"09",x"60",x"35",x"C8",x"33",x"33",x"C9",
		x"21",x"08",x"60",x"35",x"28",x"F2",x"E1",x"C9",x"87",x"E1",x"5F",x"16",x"00",x"C3",x"32",x"00",
		x"18",x"12",x"19",x"5E",x"23",x"56",x"EB",x"E9",x"11",x"04",x"00",x"06",x"0A",x"79",x"86",x"77",
		x"19",x"10",x"FA",x"C9",x"21",x"27",x"62",x"46",x"0F",x"10",x"FD",x"D8",x"E1",x"C9",x"11",x"08",
		x"69",x"01",x"28",x"00",x"ED",x"B0",x"C9",x"3A",x"18",x"60",x"21",x"1A",x"60",x"86",x"21",x"19",
		x"60",x"86",x"32",x"18",x"60",x"C9",x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"AF",x"32",
		x"84",x"7D",x"3A",x"00",x"7D",x"E6",x"01",x"C2",x"00",x"40",x"21",x"38",x"01",x"CD",x"41",x"01",
		x"3A",x"07",x"60",x"A7",x"C2",x"B5",x"00",x"3A",x"26",x"60",x"A7",x"C2",x"98",x"00",x"3A",x"0E",
		x"60",x"A7",x"3A",x"80",x"7C",x"C2",x"9B",x"00",x"3A",x"00",x"7C",x"47",x"E6",x"0F",x"4F",x"3A",
		x"11",x"60",x"2F",x"A0",x"E6",x"10",x"17",x"17",x"17",x"B1",x"60",x"6F",x"22",x"10",x"60",x"78",
		x"CB",x"77",x"C2",x"00",x"00",x"21",x"1A",x"60",x"35",x"CD",x"57",x"00",x"CD",x"7B",x"01",x"CD",
		x"E0",x"00",x"21",x"D2",x"00",x"E5",x"3A",x"05",x"60",x"EF",x"C3",x"01",x"3C",x"07",x"B2",x"08",
		x"FE",x"06",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"3E",x"01",x"32",x"84",x"7D",x"F1",x"C9",
		x"21",x"80",x"60",x"11",x"00",x"7D",x"3A",x"07",x"60",x"A7",x"C0",x"06",x"08",x"7E",x"A7",x"CA",
		x"F5",x"00",x"35",x"3E",x"01",x"12",x"1C",x"2C",x"10",x"F3",x"21",x"8B",x"60",x"7E",x"A7",x"C2",
		x"08",x"01",x"2D",x"2D",x"7E",x"C3",x"0B",x"01",x"35",x"2D",x"7E",x"32",x"00",x"7C",x"21",x"88",
		x"60",x"AF",x"BE",x"CA",x"18",x"01",x"35",x"3C",x"32",x"80",x"7D",x"C9",x"06",x"08",x"AF",x"21",
		x"00",x"7D",x"11",x"80",x"60",x"77",x"12",x"2C",x"1C",x"10",x"FA",x"06",x"04",x"12",x"1C",x"10",
		x"FC",x"32",x"80",x"7D",x"32",x"00",x"7C",x"C9",x"53",x"00",x"69",x"80",x"41",x"00",x"70",x"80",
		x"81",x"AF",x"32",x"85",x"7D",x"7E",x"32",x"08",x"78",x"23",x"7E",x"32",x"00",x"78",x"23",x"7E",
		x"32",x"00",x"78",x"23",x"7E",x"32",x"01",x"78",x"23",x"7E",x"32",x"01",x"78",x"23",x"7E",x"32",
		x"02",x"78",x"23",x"7E",x"32",x"02",x"78",x"23",x"7E",x"32",x"03",x"78",x"23",x"7E",x"32",x"03",
		x"78",x"3E",x"01",x"32",x"85",x"7D",x"AF",x"32",x"85",x"7D",x"C9",x"3A",x"00",x"7D",x"CB",x"7F",
		x"21",x"03",x"60",x"C2",x"89",x"01",x"36",x"01",x"C9",x"7E",x"A7",x"C8",x"E5",x"3A",x"05",x"60",
		x"FE",x"03",x"CA",x"9D",x"01",x"CD",x"1C",x"01",x"3E",x"03",x"32",x"83",x"60",x"E1",x"36",x"00",
		x"2B",x"34",x"11",x"24",x"60",x"1A",x"96",x"C0",x"77",x"13",x"2B",x"EB",x"1A",x"FE",x"90",x"D0",
		x"86",x"27",x"12",x"11",x"00",x"04",x"CD",x"9F",x"30",x"C9",x"00",x"37",x"00",x"AA",x"AA",x"AA",
		x"50",x"76",x"00",x"CD",x"74",x"08",x"21",x"BA",x"01",x"11",x"B2",x"60",x"01",x"09",x"00",x"ED",
		x"B0",x"3E",x"01",x"32",x"07",x"60",x"32",x"29",x"62",x"32",x"28",x"62",x"CD",x"B8",x"06",x"CD",
		x"07",x"02",x"3E",x"01",x"32",x"82",x"7D",x"32",x"05",x"60",x"32",x"27",x"62",x"AF",x"32",x"0A",
		x"60",x"CD",x"53",x"0A",x"11",x"04",x"03",x"CD",x"9F",x"30",x"11",x"02",x"02",x"CD",x"9F",x"30",
		x"11",x"00",x"02",x"CD",x"9F",x"30",x"C9",x"3A",x"80",x"7D",x"4F",x"21",x"20",x"60",x"E6",x"03",
		x"C6",x"03",x"77",x"23",x"79",x"0F",x"0F",x"E6",x"03",x"47",x"3E",x"07",x"CA",x"26",x"02",x"3E",
		x"05",x"C6",x"05",x"27",x"10",x"FB",x"77",x"23",x"79",x"01",x"01",x"01",x"11",x"02",x"01",x"E6",
		x"70",x"17",x"17",x"17",x"17",x"CA",x"47",x"02",x"DA",x"41",x"02",x"3C",x"4F",x"5A",x"C3",x"47",
		x"02",x"C6",x"02",x"47",x"57",x"87",x"5F",x"72",x"23",x"73",x"23",x"70",x"23",x"71",x"23",x"3A",
		x"80",x"7D",x"07",x"3E",x"01",x"DA",x"59",x"02",x"3D",x"77",x"21",x"65",x"35",x"11",x"00",x"61",
		x"01",x"AA",x"00",x"ED",x"B0",x"C9",x"06",x"10",x"21",x"00",x"60",x"AF",x"4F",x"77",x"23",x"0D",
		x"20",x"FB",x"10",x"F8",x"06",x"04",x"21",x"00",x"70",x"4F",x"77",x"23",x"0D",x"20",x"FB",x"10",
		x"F8",x"06",x"04",x"3E",x"10",x"21",x"00",x"74",x"0E",x"00",x"77",x"23",x"0D",x"20",x"FB",x"10",
		x"F7",x"21",x"C0",x"60",x"06",x"40",x"3E",x"FF",x"77",x"23",x"10",x"FC",x"3E",x"C0",x"32",x"B0",
		x"60",x"32",x"B1",x"60",x"AF",x"32",x"83",x"7D",x"32",x"86",x"7D",x"32",x"87",x"7D",x"3C",x"32",
		x"82",x"7D",x"31",x"00",x"6C",x"CD",x"1C",x"01",x"3E",x"01",x"32",x"84",x"7D",x"26",x"60",x"3A",
		x"B1",x"60",x"6F",x"7E",x"87",x"30",x"1C",x"CD",x"15",x"03",x"CD",x"50",x"03",x"21",x"19",x"60",
		x"34",x"21",x"83",x"63",x"3A",x"1A",x"60",x"BE",x"28",x"E3",x"77",x"CD",x"7F",x"03",x"CD",x"A2",
		x"03",x"18",x"DA",x"E6",x"1F",x"5F",x"16",x"00",x"36",x"FF",x"2C",x"4E",x"36",x"FF",x"2C",x"7D",
		x"FE",x"C0",x"30",x"02",x"3E",x"C0",x"32",x"B1",x"60",x"79",x"21",x"BD",x"02",x"E5",x"21",x"07",
		x"03",x"19",x"5E",x"23",x"56",x"EB",x"E9",x"1C",x"05",x"9B",x"05",x"C6",x"05",x"E9",x"05",x"11",
		x"06",x"2A",x"06",x"B8",x"06",x"3A",x"1A",x"60",x"47",x"E6",x"0F",x"C0",x"CF",x"3A",x"0D",x"60",
		x"CD",x"47",x"03",x"11",x"E0",x"FF",x"CB",x"60",x"28",x"14",x"3E",x"10",x"77",x"19",x"77",x"19",
		x"77",x"3A",x"0F",x"60",x"A7",x"C8",x"3A",x"0D",x"60",x"EE",x"01",x"CD",x"47",x"03",x"3C",x"77",
		x"19",x"36",x"25",x"19",x"36",x"20",x"C9",x"21",x"40",x"77",x"A7",x"C8",x"21",x"E0",x"74",x"C9",
		x"3A",x"2D",x"62",x"A7",x"C0",x"21",x"B3",x"60",x"3A",x"0D",x"60",x"A7",x"28",x"03",x"21",x"B6",
		x"60",x"7E",x"E6",x"F0",x"47",x"23",x"7E",x"E6",x"0F",x"B0",x"0F",x"0F",x"0F",x"0F",x"21",x"21",
		x"60",x"BE",x"D8",x"3E",x"01",x"32",x"2D",x"62",x"21",x"28",x"62",x"34",x"C3",x"B8",x"06",x"21",
		x"84",x"63",x"7E",x"34",x"A7",x"C0",x"21",x"81",x"63",x"7E",x"47",x"34",x"E6",x"07",x"C0",x"78",
		x"0F",x"0F",x"0F",x"47",x"3A",x"29",x"62",x"80",x"FE",x"05",x"38",x"02",x"3E",x"05",x"32",x"80",
		x"63",x"C9",x"3E",x"03",x"F7",x"D7",x"3A",x"50",x"63",x"0F",x"D8",x"21",x"B8",x"62",x"35",x"C0",
		x"36",x"04",x"3A",x"B9",x"62",x"0F",x"D0",x"21",x"29",x"6A",x"06",x"40",x"DD",x"21",x"A0",x"66",
		x"0F",x"D2",x"E4",x"03",x"DD",x"36",x"09",x"02",x"DD",x"36",x"0A",x"02",x"04",x"04",x"CD",x"F2",
		x"03",x"21",x"BA",x"62",x"35",x"C0",x"3E",x"01",x"32",x"B9",x"62",x"32",x"A0",x"63",x"3E",x"10",
		x"32",x"BA",x"62",x"C9",x"DD",x"36",x"09",x"02",x"DD",x"36",x"0A",x"00",x"CD",x"F2",x"03",x"C3",
		x"DE",x"03",x"70",x"3A",x"19",x"60",x"0F",x"D8",x"04",x"70",x"C9",x"3A",x"27",x"62",x"FE",x"02",
		x"C2",x"13",x"04",x"21",x"08",x"69",x"3A",x"A3",x"63",x"4F",x"FF",x"3A",x"10",x"69",x"D6",x"3B",
		x"32",x"B7",x"63",x"3A",x"91",x"63",x"A7",x"C2",x"26",x"04",x"3A",x"1A",x"60",x"A7",x"C2",x"86",
		x"04",x"3E",x"01",x"32",x"91",x"63",x"21",x"90",x"63",x"34",x"7E",x"FE",x"80",x"CA",x"64",x"04",
		x"3A",x"93",x"63",x"A7",x"C2",x"86",x"04",x"7E",x"47",x"E6",x"1F",x"C2",x"86",x"04",x"21",x"CF",
		x"39",x"CB",x"68",x"20",x"03",x"21",x"F7",x"39",x"CD",x"4E",x"00",x"3E",x"03",x"32",x"82",x"60",
		x"3A",x"27",x"62",x"0F",x"D2",x"78",x"04",x"0F",x"DA",x"86",x"04",x"21",x"0B",x"69",x"0E",x"FC",
		x"FF",x"C3",x"86",x"04",x"AF",x"77",x"23",x"77",x"3A",x"93",x"63",x"A7",x"C2",x"86",x"04",x"21",
		x"5C",x"38",x"CD",x"4E",x"00",x"C3",x"50",x"04",x"21",x"08",x"69",x"0E",x"44",x"0F",x"D2",x"85",
		x"04",x"3A",x"B7",x"63",x"4F",x"FF",x"3A",x"90",x"63",x"4F",x"11",x"20",x"00",x"3A",x"27",x"62",
		x"FE",x"04",x"CA",x"BE",x"04",x"79",x"A7",x"CA",x"A1",x"04",x"3E",x"EF",x"CB",x"71",x"C2",x"A3",
		x"04",x"3E",x"10",x"21",x"C4",x"75",x"CD",x"14",x"05",x"3A",x"05",x"69",x"32",x"05",x"69",x"CB",
		x"71",x"C8",x"47",x"79",x"E6",x"07",x"C0",x"78",x"EE",x"03",x"32",x"05",x"69",x"C9",x"3E",x"10",
		x"21",x"23",x"76",x"CD",x"14",x"05",x"21",x"83",x"75",x"CD",x"14",x"05",x"CB",x"71",x"CA",x"09",
		x"05",x"3A",x"03",x"62",x"FE",x"80",x"D2",x"F1",x"04",x"3E",x"DF",x"21",x"23",x"76",x"CD",x"14",
		x"05",x"3A",x"01",x"69",x"F6",x"80",x"32",x"01",x"69",x"3A",x"05",x"69",x"F6",x"80",x"C3",x"AC",
		x"04",x"3E",x"EF",x"21",x"83",x"75",x"CD",x"14",x"05",x"3A",x"01",x"69",x"E6",x"7F",x"32",x"01",
		x"69",x"3A",x"05",x"69",x"E6",x"7F",x"C3",x"AC",x"04",x"3A",x"03",x"62",x"FE",x"80",x"D2",x"F9",
		x"04",x"C3",x"E1",x"04",x"06",x"03",x"77",x"19",x"3D",x"10",x"FB",x"C9",x"4F",x"CF",x"CD",x"5F",
		x"05",x"79",x"81",x"81",x"4F",x"21",x"29",x"35",x"06",x"00",x"09",x"A7",x"06",x"03",x"1A",x"8E",
		x"27",x"12",x"13",x"23",x"10",x"F8",x"D5",x"1B",x"3A",x"0D",x"60",x"CD",x"6B",x"05",x"D1",x"1B",
		x"21",x"BA",x"60",x"06",x"03",x"1A",x"BE",x"D8",x"C2",x"50",x"05",x"1B",x"2B",x"10",x"F6",x"C9",
		x"CD",x"5F",x"05",x"21",x"B8",x"60",x"1A",x"77",x"13",x"23",x"10",x"FA",x"C3",x"DA",x"05",x"11",
		x"B2",x"60",x"3A",x"0D",x"60",x"A7",x"C8",x"11",x"B5",x"60",x"C9",x"DD",x"21",x"81",x"77",x"A7",
		x"28",x"0A",x"DD",x"21",x"21",x"75",x"18",x"04",x"DD",x"21",x"41",x"76",x"EB",x"11",x"E0",x"FF",
		x"01",x"04",x"03",x"7E",x"0F",x"0F",x"0F",x"0F",x"CD",x"93",x"05",x"7E",x"CD",x"93",x"05",x"2B",
		x"10",x"F1",x"C9",x"E6",x"0F",x"DD",x"77",x"00",x"DD",x"19",x"C9",x"FE",x"03",x"D2",x"BD",x"05",
		x"F5",x"21",x"B2",x"60",x"A7",x"CA",x"AB",x"05",x"21",x"B5",x"60",x"FE",x"02",x"C2",x"B3",x"05",
		x"21",x"B8",x"60",x"AF",x"77",x"23",x"77",x"23",x"77",x"F1",x"C3",x"C6",x"05",x"3D",x"F5",x"CD",
		x"9B",x"05",x"F1",x"C8",x"18",x"F7",x"FE",x"03",x"CA",x"E0",x"05",x"11",x"B4",x"60",x"A7",x"CA",
		x"D5",x"05",x"11",x"B7",x"60",x"FE",x"02",x"C2",x"6B",x"05",x"11",x"BA",x"60",x"C3",x"78",x"05",
		x"3D",x"F5",x"CD",x"C6",x"05",x"F1",x"C8",x"18",x"F7",x"21",x"4B",x"36",x"87",x"F5",x"E6",x"7F",
		x"5F",x"16",x"00",x"19",x"5E",x"23",x"56",x"EB",x"5E",x"23",x"56",x"23",x"01",x"E0",x"FF",x"EB",
		x"1A",x"FE",x"3F",x"CA",x"26",x"00",x"77",x"F1",x"30",x"02",x"36",x"10",x"F5",x"13",x"09",x"18",
		x"EF",x"3A",x"07",x"60",x"0F",x"D0",x"3E",x"05",x"CD",x"E9",x"05",x"21",x"01",x"60",x"11",x"E0",
		x"FF",x"DD",x"21",x"BF",x"74",x"06",x"01",x"C3",x"83",x"05",x"A7",x"CA",x"91",x"06",x"3A",x"8C",
		x"63",x"A7",x"C2",x"A8",x"06",x"3A",x"B8",x"63",x"A7",x"C0",x"3A",x"B0",x"62",x"01",x"0A",x"00",
		x"04",x"91",x"C2",x"40",x"06",x"78",x"07",x"07",x"07",x"07",x"32",x"8C",x"63",x"21",x"4A",x"38",
		x"11",x"65",x"74",x"3E",x"06",x"DD",x"21",x"1D",x"00",x"01",x"03",x"00",x"ED",x"B0",x"DD",x"19",
		x"DD",x"E5",x"D1",x"3D",x"C2",x"55",x"06",x"3A",x"8C",x"63",x"4F",x"E6",x"0F",x"47",x"79",x"0F",
		x"0F",x"0F",x"0F",x"E6",x"0F",x"C2",x"89",x"06",x"3E",x"03",x"32",x"89",x"60",x"3E",x"70",x"32",
		x"86",x"74",x"32",x"A6",x"74",x"80",x"47",x"3E",x"10",x"32",x"E6",x"74",x"78",x"32",x"C6",x"74",
		x"C9",x"3A",x"8C",x"63",x"47",x"E6",x"0F",x"C5",x"CD",x"1C",x"05",x"C1",x"78",x"0F",x"0F",x"0F",
		x"0F",x"E6",x"0F",x"C6",x"0A",x"C3",x"1C",x"05",x"D6",x"01",x"20",x"05",x"21",x"B8",x"63",x"36",
		x"01",x"27",x"32",x"8C",x"63",x"C3",x"6A",x"06",x"4F",x"CF",x"06",x"06",x"11",x"E0",x"FF",x"21",
		x"83",x"77",x"36",x"10",x"19",x"10",x"FB",x"3A",x"28",x"62",x"91",x"CA",x"D7",x"06",x"47",x"21",
		x"83",x"77",x"36",x"FF",x"19",x"10",x"FB",x"21",x"03",x"75",x"36",x"1C",x"21",x"E3",x"74",x"36",
		x"34",x"3A",x"29",x"62",x"FE",x"64",x"38",x"05",x"3E",x"63",x"32",x"29",x"62",x"01",x"0A",x"FF",
		x"04",x"91",x"D2",x"F0",x"06",x"81",x"32",x"A3",x"74",x"78",x"32",x"C3",x"74",x"C9",x"3A",x"0A",
		x"60",x"EF",x"86",x"09",x"AB",x"09",x"D6",x"09",x"FE",x"09",x"1B",x"0A",x"37",x"0A",x"63",x"0A",
		x"76",x"0A",x"DA",x"0B",x"00",x"00",x"91",x"0C",x"3C",x"12",x"7A",x"19",x"7C",x"12",x"F2",x"12",
		x"44",x"13",x"8F",x"13",x"A1",x"13",x"AA",x"13",x"BB",x"13",x"1E",x"14",x"86",x"14",x"15",x"16",
		x"6B",x"19",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"0A",x"60",x"3A",
		x"01",x"60",x"A7",x"C2",x"5C",x"07",x"7E",x"EF",x"79",x"07",x"63",x"07",x"3C",x"12",x"77",x"19",
		x"7C",x"12",x"C3",x"07",x"CB",x"07",x"4B",x"08",x"00",x"00",x"00",x"00",x"36",x"00",x"21",x"05",
		x"60",x"34",x"C9",x"E7",x"AF",x"32",x"92",x"63",x"32",x"A0",x"63",x"3E",x"01",x"32",x"27",x"62",
		x"32",x"29",x"62",x"32",x"28",x"62",x"C3",x"92",x"0C",x"21",x"86",x"7D",x"36",x"00",x"23",x"36",
		x"00",x"11",x"1B",x"03",x"CD",x"9F",x"30",x"1C",x"CD",x"9F",x"30",x"CD",x"65",x"09",x"21",x"09",
		x"60",x"36",x"02",x"23",x"34",x"CD",x"74",x"08",x"CD",x"53",x"0A",x"3A",x"0F",x"60",x"FE",x"01",
		x"CC",x"EE",x"09",x"ED",x"5B",x"22",x"60",x"21",x"6C",x"75",x"CD",x"AD",x"07",x"73",x"23",x"23",
		x"72",x"7A",x"D6",x"0A",x"C2",x"BC",x"07",x"77",x"3C",x"32",x"8E",x"75",x"11",x"01",x"02",x"21",
		x"8C",x"76",x"C9",x"CD",x"74",x"08",x"21",x"0A",x"60",x"34",x"C9",x"3A",x"8A",x"63",x"FE",x"00",
		x"C2",x"2D",x"08",x"3E",x"60",x"32",x"8A",x"63",x"0E",x"5F",x"FE",x"00",x"CA",x"3B",x"08",x"21",
		x"86",x"7D",x"36",x"00",x"79",x"CB",x"07",x"30",x"02",x"36",x"01",x"23",x"36",x"00",x"CB",x"07",
		x"30",x"02",x"36",x"01",x"32",x"8B",x"63",x"21",x"08",x"3D",x"3E",x"B0",x"46",x"23",x"5E",x"23",
		x"56",x"12",x"13",x"10",x"FC",x"23",x"7E",x"FE",x"00",x"C2",x"FA",x"07",x"11",x"1E",x"03",x"CD",
		x"9F",x"30",x"13",x"CD",x"9F",x"30",x"21",x"CF",x"39",x"CD",x"4E",x"00",x"CD",x"24",x"3F",x"00",
		x"21",x"08",x"69",x"0E",x"44",x"FF",x"21",x"0B",x"69",x"0E",x"78",x"FF",x"C9",x"3A",x"8B",x"63",
		x"4F",x"3A",x"8A",x"63",x"3D",x"32",x"8A",x"63",x"C3",x"DA",x"07",x"21",x"09",x"60",x"36",x"02",
		x"23",x"34",x"21",x"8A",x"63",x"36",x"00",x"23",x"36",x"00",x"C9",x"E7",x"21",x"0A",x"60",x"36",
		x"00",x"C9",x"21",x"00",x"74",x"0E",x"04",x"06",x"00",x"3E",x"10",x"77",x"23",x"10",x"FC",x"0D",
		x"C2",x"57",x"08",x"21",x"00",x"69",x"0E",x"02",x"06",x"C0",x"AF",x"77",x"23",x"10",x"FC",x"0D",
		x"C2",x"68",x"08",x"C9",x"21",x"04",x"74",x"0E",x"20",x"06",x"1C",x"3E",x"10",x"11",x"04",x"00",
		x"77",x"23",x"10",x"FC",x"19",x"0D",x"C2",x"79",x"08",x"21",x"22",x"75",x"11",x"20",x"00",x"0E",
		x"02",x"3E",x"10",x"06",x"0E",x"77",x"19",x"10",x"FC",x"21",x"23",x"75",x"0D",x"C2",x"93",x"08",
		x"21",x"00",x"69",x"06",x"00",x"3E",x"00",x"77",x"23",x"10",x"FC",x"06",x"80",x"77",x"23",x"10",
		x"FC",x"C9",x"3A",x"0A",x"60",x"EF",x"BA",x"08",x"F8",x"08",x"CD",x"74",x"08",x"AF",x"32",x"07",
		x"60",x"11",x"0C",x"03",x"CD",x"9F",x"30",x"21",x"0A",x"60",x"34",x"CD",x"65",x"09",x"AF",x"21",
		x"86",x"7D",x"77",x"2C",x"77",x"06",x"04",x"1E",x"09",x"3A",x"01",x"60",x"FE",x"01",x"CA",x"E4",
		x"08",x"06",x"0C",x"1C",x"3A",x"1A",x"60",x"E6",x"07",x"C2",x"F3",x"08",x"7B",x"CD",x"E9",x"05",
		x"CD",x"16",x"06",x"3A",x"00",x"7D",x"A0",x"C9",x"CD",x"D5",x"08",x"FE",x"04",x"CA",x"06",x"09",
		x"FE",x"08",x"CA",x"19",x"09",x"C9",x"CD",x"77",x"09",x"21",x"48",x"60",x"06",x"08",x"AF",x"77",
		x"2C",x"10",x"FC",x"21",x"00",x"00",x"C3",x"38",x"09",x"CD",x"77",x"09",x"CD",x"77",x"09",x"11",
		x"48",x"60",x"3A",x"20",x"60",x"12",x"1C",x"21",x"5E",x"09",x"01",x"07",x"00",x"ED",x"B0",x"11",
		x"01",x"01",x"CD",x"9F",x"30",x"21",x"00",x"01",x"22",x"0E",x"60",x"CD",x"74",x"08",x"11",x"40",
		x"60",x"3A",x"20",x"60",x"12",x"1C",x"21",x"5E",x"09",x"01",x"07",x"00",x"ED",x"B0",x"11",x"00",
		x"01",x"CD",x"9F",x"30",x"AF",x"32",x"0A",x"60",x"3E",x"03",x"32",x"05",x"60",x"C9",x"01",x"65",
		x"3A",x"01",x"00",x"00",x"00",x"11",x"00",x"04",x"CD",x"9F",x"30",x"11",x"14",x"03",x"06",x"06",
		x"CD",x"9F",x"30",x"1C",x"10",x"FA",x"C9",x"21",x"01",x"60",x"3E",x"99",x"86",x"27",x"77",x"11",
		x"00",x"04",x"CD",x"9F",x"30",x"C9",x"CD",x"52",x"08",x"CD",x"1C",x"01",x"11",x"82",x"7D",x"3E",
		x"01",x"12",x"21",x"0A",x"60",x"3A",x"0E",x"60",x"A7",x"C2",x"9F",x"09",x"36",x"01",x"C9",x"3A",
		x"26",x"60",x"3D",x"CA",x"A8",x"09",x"AF",x"12",x"36",x"03",x"C9",x"21",x"40",x"60",x"11",x"28",
		x"62",x"01",x"08",x"00",x"ED",x"B0",x"2A",x"2A",x"62",x"7E",x"32",x"27",x"62",x"3A",x"0F",x"60",
		x"A7",x"21",x"09",x"60",x"11",x"0A",x"60",x"CA",x"D0",x"09",x"36",x"78",x"EB",x"36",x"02",x"C9",
		x"36",x"01",x"EB",x"36",x"05",x"C9",x"AF",x"32",x"86",x"7D",x"32",x"87",x"7D",x"11",x"02",x"03",
		x"CD",x"9F",x"30",x"11",x"01",x"02",x"CD",x"9F",x"30",x"3E",x"05",x"32",x"0A",x"60",x"3E",x"02",
		x"32",x"E0",x"74",x"3E",x"25",x"32",x"C0",x"74",x"3E",x"20",x"32",x"A0",x"74",x"C9",x"21",x"48",
		x"60",x"11",x"28",x"62",x"01",x"08",x"00",x"ED",x"B0",x"2A",x"2A",x"62",x"7E",x"32",x"27",x"62",
		x"3E",x"78",x"32",x"09",x"60",x"3E",x"04",x"32",x"0A",x"60",x"C9",x"AF",x"32",x"86",x"7D",x"32",
		x"87",x"7D",x"11",x"03",x"03",x"CD",x"9F",x"30",x"11",x"01",x"02",x"CD",x"9F",x"30",x"CD",x"EE",
		x"09",x"3E",x"05",x"32",x"0A",x"60",x"C9",x"11",x"04",x"03",x"CD",x"9F",x"30",x"11",x"02",x"02",
		x"CD",x"9F",x"30",x"11",x"00",x"02",x"CD",x"9F",x"30",x"11",x"00",x"06",x"CD",x"9F",x"30",x"21",
		x"0A",x"60",x"34",x"3E",x"01",x"32",x"40",x"77",x"3E",x"25",x"32",x"20",x"77",x"3E",x"20",x"32",
		x"00",x"77",x"C9",x"DF",x"CD",x"74",x"08",x"21",x"09",x"60",x"36",x"01",x"2C",x"34",x"11",x"2C",
		x"62",x"1A",x"A7",x"C0",x"34",x"C9",x"3A",x"85",x"63",x"EF",x"8A",x"0A",x"BF",x"0A",x"E8",x"0A",
		x"69",x"30",x"06",x"0B",x"69",x"30",x"68",x"0B",x"B3",x"0B",x"AF",x"32",x"86",x"7D",x"3C",x"32",
		x"87",x"7D",x"11",x"0D",x"38",x"CD",x"A7",x"0D",x"3E",x"10",x"32",x"A3",x"76",x"32",x"63",x"76",
		x"3E",x"D4",x"32",x"AA",x"75",x"AF",x"32",x"AF",x"62",x"21",x"B4",x"38",x"22",x"C2",x"63",x"21",
		x"CB",x"38",x"22",x"C4",x"63",x"3E",x"40",x"32",x"09",x"60",x"21",x"85",x"63",x"34",x"C9",x"DF",
		x"21",x"8C",x"38",x"CD",x"4E",x"00",x"21",x"08",x"69",x"0E",x"30",x"FF",x"21",x"0B",x"69",x"0E",
		x"99",x"FF",x"3E",x"1F",x"32",x"8E",x"63",x"AF",x"32",x"0C",x"69",x"21",x"8A",x"60",x"36",x"01",
		x"23",x"36",x"03",x"21",x"85",x"63",x"34",x"C9",x"CD",x"6F",x"30",x"3A",x"AF",x"62",x"E6",x"0F",
		x"CC",x"4A",x"30",x"3A",x"0B",x"69",x"FE",x"5D",x"D0",x"3E",x"20",x"32",x"09",x"60",x"21",x"85",
		x"63",x"34",x"22",x"C0",x"63",x"C9",x"3A",x"1A",x"60",x"0F",x"D8",x"2A",x"C2",x"63",x"7E",x"FE",
		x"7F",x"CA",x"1E",x"0B",x"23",x"22",x"C2",x"63",x"4F",x"21",x"0B",x"69",x"FF",x"C9",x"21",x"5C",
		x"38",x"CD",x"4E",x"00",x"11",x"00",x"69",x"01",x"08",x"00",x"ED",x"B0",x"21",x"08",x"69",x"0E",
		x"50",x"FF",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"CD",x"4A",x"30",x"3A",x"8E",x"63",x"FE",x"0A",
		x"C2",x"38",x"0B",x"3E",x"03",x"32",x"82",x"60",x"11",x"2C",x"39",x"CD",x"A7",x"0D",x"3E",x"10",
		x"32",x"AA",x"74",x"32",x"8A",x"74",x"3E",x"05",x"32",x"8D",x"63",x"3E",x"20",x"32",x"09",x"60",
		x"21",x"85",x"63",x"34",x"22",x"C0",x"63",x"C9",x"3A",x"1A",x"60",x"0F",x"D8",x"2A",x"C4",x"63",
		x"7E",x"FE",x"7F",x"CA",x"86",x"0B",x"23",x"22",x"C4",x"63",x"21",x"0B",x"69",x"4F",x"FF",x"21",
		x"08",x"69",x"0E",x"FF",x"FF",x"C9",x"21",x"CB",x"38",x"22",x"C4",x"63",x"3E",x"03",x"32",x"82",
		x"60",x"21",x"DC",x"38",x"3A",x"8D",x"63",x"3D",x"07",x"07",x"07",x"07",x"5F",x"16",x"00",x"19",
		x"EB",x"CD",x"A7",x"0D",x"21",x"8D",x"63",x"35",x"C0",x"3E",x"B0",x"32",x"09",x"60",x"21",x"85",
		x"63",x"34",x"C9",x"21",x"8A",x"60",x"3A",x"09",x"60",x"FE",x"90",x"20",x"0B",x"36",x"0F",x"23",
		x"36",x"03",x"21",x"19",x"69",x"34",x"18",x"09",x"FE",x"18",x"20",x"05",x"21",x"19",x"69",x"35",
		x"00",x"DF",x"AF",x"32",x"85",x"63",x"34",x"23",x"34",x"C9",x"CD",x"1C",x"01",x"DF",x"CD",x"74",
		x"08",x"16",x"06",x"3A",x"00",x"62",x"5F",x"CD",x"9F",x"30",x"21",x"86",x"7D",x"36",x"01",x"23",
		x"36",x"00",x"21",x"8A",x"60",x"36",x"02",x"23",x"36",x"03",x"21",x"A7",x"63",x"36",x"00",x"21",
		x"DC",x"76",x"22",x"A8",x"63",x"3A",x"2E",x"62",x"FE",x"06",x"38",x"05",x"3E",x"05",x"32",x"2E",
		x"62",x"3A",x"2F",x"62",x"47",x"3A",x"2A",x"62",x"B8",x"28",x"04",x"21",x"2E",x"62",x"34",x"32",
		x"2F",x"62",x"3A",x"2E",x"62",x"47",x"21",x"BC",x"75",x"0E",x"50",x"71",x"0C",x"2B",x"71",x"0C",
		x"2B",x"71",x"0C",x"2B",x"71",x"79",x"FE",x"67",x"CA",x"43",x"0C",x"0C",x"11",x"23",x"00",x"19",
		x"C3",x"2B",x"0C",x"3A",x"A7",x"63",x"3C",x"32",x"A7",x"63",x"3D",x"CB",x"27",x"CB",x"27",x"E5",
		x"21",x"F0",x"3C",x"C5",x"DD",x"2A",x"A8",x"63",x"4F",x"06",x"00",x"09",x"7E",x"DD",x"77",x"60",
		x"23",x"7E",x"DD",x"77",x"40",x"23",x"7E",x"DD",x"77",x"20",x"DD",x"36",x"E0",x"8B",x"C1",x"DD",
		x"E5",x"E1",x"11",x"FC",x"FF",x"19",x"22",x"A8",x"63",x"E1",x"11",x"5F",x"FF",x"19",x"05",x"C2",
		x"29",x"0C",x"11",x"07",x"03",x"CD",x"9F",x"30",x"21",x"09",x"60",x"36",x"A0",x"23",x"34",x"34",
		x"C9",x"DF",x"CD",x"74",x"08",x"AF",x"32",x"8C",x"63",x"11",x"01",x"05",x"CD",x"9F",x"30",x"21",
		x"86",x"7D",x"36",x"00",x"23",x"36",x"01",x"3A",x"27",x"62",x"3D",x"CA",x"D4",x"0C",x"3D",x"CA",
		x"DF",x"0C",x"3D",x"CA",x"F2",x"0C",x"CD",x"43",x"0D",x"21",x"86",x"7D",x"36",x"01",x"3E",x"0B",
		x"32",x"89",x"60",x"11",x"8B",x"3C",x"CD",x"A7",x"0D",x"3A",x"27",x"62",x"FE",x"04",x"CC",x"00",
		x"0D",x"C3",x"A0",x"3F",x"11",x"E4",x"3A",x"3E",x"08",x"32",x"89",x"60",x"C3",x"C6",x"0C",x"11",
		x"5D",x"3B",x"21",x"86",x"7D",x"36",x"01",x"23",x"36",x"00",x"3E",x"09",x"32",x"89",x"60",x"C3",
		x"C6",x"0C",x"CD",x"27",x"0D",x"3E",x"0A",x"32",x"89",x"60",x"11",x"E5",x"3B",x"C3",x"C6",x"0C",
		x"06",x"08",x"21",x"17",x"0D",x"3E",x"B8",x"0E",x"02",x"5E",x"23",x"56",x"23",x"12",x"3D",x"13",
		x"0D",x"C2",x"0D",x"0D",x"10",x"EF",x"C9",x"CA",x"76",x"CF",x"76",x"D4",x"76",x"D9",x"76",x"2A",
		x"75",x"2F",x"75",x"34",x"75",x"39",x"75",x"21",x"0D",x"77",x"CD",x"30",x"0D",x"21",x"0D",x"76",
		x"06",x"11",x"36",x"FD",x"23",x"10",x"FB",x"11",x"0F",x"00",x"19",x"06",x"11",x"36",x"FC",x"23",
		x"10",x"FB",x"C9",x"21",x"87",x"76",x"CD",x"4C",x"0D",x"21",x"47",x"75",x"06",x"04",x"36",x"FD",
		x"23",x"10",x"FB",x"11",x"1C",x"00",x"19",x"06",x"04",x"36",x"FC",x"23",x"10",x"FB",x"C9",x"CD",
		x"56",x"0F",x"CD",x"41",x"24",x"21",x"09",x"60",x"36",x"40",x"23",x"34",x"21",x"5C",x"38",x"CD",
		x"4E",x"00",x"11",x"00",x"69",x"01",x"08",x"00",x"ED",x"B0",x"3A",x"27",x"62",x"FE",x"04",x"28",
		x"0A",x"0F",x"0F",x"D8",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"C9",x"21",x"08",x"69",x"0E",x"44",
		x"FF",x"11",x"04",x"00",x"01",x"10",x"02",x"21",x"00",x"69",x"CD",x"3D",x"00",x"01",x"F8",x"02",
		x"21",x"03",x"69",x"CD",x"3D",x"00",x"C9",x"1A",x"32",x"B3",x"63",x"FE",x"AA",x"C8",x"13",x"1A",
		x"67",x"44",x"13",x"1A",x"6F",x"4D",x"D5",x"CD",x"F0",x"2F",x"D1",x"22",x"AB",x"63",x"78",x"E6",
		x"07",x"32",x"B4",x"63",x"79",x"E6",x"07",x"32",x"AF",x"63",x"13",x"1A",x"67",x"90",x"D2",x"D3",
		x"0D",x"ED",x"44",x"32",x"B1",x"63",x"13",x"1A",x"6F",x"91",x"32",x"B2",x"63",x"1A",x"E6",x"07",
		x"32",x"B0",x"63",x"D5",x"CD",x"F0",x"2F",x"D1",x"22",x"AD",x"63",x"3A",x"B3",x"63",x"FE",x"02",
		x"F2",x"4F",x"0E",x"3A",x"B2",x"63",x"D6",x"10",x"47",x"3A",x"AF",x"63",x"80",x"32",x"B2",x"63",
		x"3A",x"AF",x"63",x"C6",x"F0",x"2A",x"AB",x"63",x"77",x"2C",x"D6",x"30",x"77",x"3A",x"B3",x"63",
		x"FE",x"01",x"C2",x"19",x"0E",x"AF",x"32",x"B2",x"63",x"3A",x"B2",x"63",x"D6",x"08",x"32",x"B2",
		x"63",x"DA",x"2A",x"0E",x"2C",x"36",x"C0",x"C3",x"19",x"0E",x"3A",x"B0",x"63",x"C6",x"D0",x"2A",
		x"AD",x"63",x"77",x"3A",x"B3",x"63",x"FE",x"01",x"C2",x"3F",x"0E",x"2D",x"36",x"C0",x"2C",x"3A",
		x"B0",x"63",x"FE",x"00",x"CA",x"4B",x"0E",x"C6",x"E0",x"2C",x"77",x"13",x"C3",x"A7",x"0D",x"3A",
		x"B3",x"63",x"FE",x"02",x"C2",x"E8",x"0E",x"3A",x"AF",x"63",x"C6",x"F0",x"32",x"B5",x"63",x"2A",
		x"AB",x"63",x"3A",x"B5",x"63",x"77",x"23",x"7D",x"E6",x"1F",x"CA",x"78",x"0E",x"3A",x"B5",x"63",
		x"FE",x"F0",x"CA",x"78",x"0E",x"D6",x"10",x"77",x"01",x"1F",x"00",x"09",x"3A",x"B1",x"63",x"D6",
		x"08",x"DA",x"CF",x"0E",x"32",x"B1",x"63",x"3A",x"B2",x"63",x"FE",x"00",x"CA",x"62",x"0E",x"3A",
		x"B5",x"63",x"77",x"23",x"7D",x"E6",x"1F",x"CA",x"A0",x"0E",x"3A",x"B5",x"63",x"D6",x"10",x"77",
		x"01",x"1F",x"00",x"09",x"3A",x"B1",x"63",x"D6",x"08",x"DA",x"CF",x"0E",x"32",x"B1",x"63",x"3A",
		x"B2",x"63",x"CB",x"7F",x"C2",x"D3",x"0E",x"3A",x"B5",x"63",x"3C",x"32",x"B5",x"63",x"FE",x"F8",
		x"C2",x"C9",x"0E",x"23",x"3E",x"F0",x"32",x"B5",x"63",x"7D",x"E6",x"1F",x"C2",x"62",x"0E",x"13",
		x"C3",x"A7",x"0D",x"3A",x"B5",x"63",x"3D",x"32",x"B5",x"63",x"FE",x"F0",x"F2",x"E5",x"0E",x"2B",
		x"3E",x"F7",x"32",x"B5",x"63",x"C3",x"62",x"0E",x"3A",x"B3",x"63",x"FE",x"03",x"C2",x"1B",x"0F",
		x"2A",x"AB",x"63",x"3E",x"B3",x"77",x"01",x"20",x"00",x"09",x"3A",x"B1",x"63",x"D6",x"10",x"DA",
		x"14",x"0F",x"32",x"B1",x"63",x"3E",x"B1",x"77",x"01",x"20",x"00",x"09",x"3A",x"B1",x"63",x"D6",
		x"08",x"C3",x"FF",x"0E",x"3E",x"B2",x"77",x"13",x"C3",x"A7",x"0D",x"3A",x"B3",x"63",x"FE",x"07",
		x"F2",x"CF",x"0E",x"FE",x"04",x"CA",x"4C",x"0F",x"FE",x"05",x"CA",x"51",x"0F",x"3E",x"FE",x"32",
		x"B5",x"63",x"2A",x"AB",x"63",x"3A",x"B5",x"63",x"77",x"01",x"20",x"00",x"09",x"3A",x"B1",x"63",
		x"D6",x"08",x"32",x"B1",x"63",x"D2",x"35",x"0F",x"13",x"C3",x"A7",x"0D",x"3E",x"E0",x"C3",x"2F",
		x"0F",x"3E",x"B0",x"C3",x"2F",x"0F",x"06",x"27",x"21",x"00",x"62",x"AF",x"77",x"2C",x"10",x"FC",
		x"0E",x"11",x"16",x"80",x"21",x"80",x"62",x"42",x"77",x"23",x"10",x"FC",x"0D",x"20",x"F8",x"21",
		x"9C",x"3D",x"11",x"80",x"62",x"01",x"40",x"00",x"ED",x"B0",x"3A",x"29",x"62",x"47",x"A7",x"17",
		x"A7",x"17",x"A7",x"17",x"80",x"80",x"C6",x"28",x"FE",x"51",x"38",x"02",x"3E",x"50",x"21",x"B0",
		x"62",x"06",x"03",x"77",x"2C",x"10",x"FC",x"87",x"47",x"3E",x"DC",x"90",x"FE",x"28",x"30",x"02",
		x"3E",x"28",x"77",x"2C",x"77",x"21",x"09",x"62",x"36",x"04",x"2C",x"36",x"08",x"3A",x"27",x"62",
		x"4F",x"CB",x"57",x"20",x"16",x"21",x"00",x"6A",x"3E",x"4F",x"06",x"03",x"77",x"2C",x"36",x"3A",
		x"2C",x"36",x"0F",x"2C",x"36",x"18",x"2C",x"C6",x"10",x"10",x"F1",x"79",x"EF",x"00",x"00",x"D7",
		x"0F",x"1F",x"10",x"87",x"10",x"31",x"11",x"21",x"DC",x"3D",x"11",x"A8",x"69",x"01",x"10",x"00",
		x"ED",x"B0",x"21",x"EC",x"3D",x"11",x"07",x"64",x"0E",x"1C",x"06",x"05",x"CD",x"2A",x"12",x"21",
		x"F4",x"3D",x"CD",x"FA",x"11",x"21",x"00",x"3E",x"11",x"FC",x"69",x"01",x"04",x"00",x"ED",x"B0",
		x"21",x"0C",x"3E",x"CD",x"A6",x"11",x"21",x"1B",x"10",x"11",x"07",x"67",x"01",x"1C",x"08",x"CD",
		x"2A",x"12",x"11",x"07",x"68",x"06",x"02",x"CD",x"2A",x"12",x"C9",x"00",x"00",x"02",x"02",x"21",
		x"EC",x"3D",x"11",x"07",x"64",x"01",x"1C",x"05",x"CD",x"2A",x"12",x"CD",x"86",x"11",x"21",x"18",
		x"3E",x"11",x"A7",x"65",x"01",x"0C",x"06",x"CD",x"2A",x"12",x"DD",x"21",x"A0",x"65",x"21",x"B8",
		x"69",x"11",x"10",x"00",x"06",x"06",x"CD",x"D3",x"11",x"21",x"FA",x"3D",x"CD",x"FA",x"11",x"21",
		x"04",x"3E",x"11",x"FC",x"69",x"01",x"04",x"00",x"ED",x"B0",x"21",x"1C",x"3E",x"11",x"44",x"69",
		x"01",x"08",x"00",x"ED",x"B0",x"21",x"24",x"3E",x"11",x"E4",x"69",x"01",x"18",x"00",x"ED",x"B0",
		x"21",x"10",x"3E",x"CD",x"A6",x"11",x"21",x"3C",x"3E",x"11",x"0C",x"6A",x"01",x"0C",x"00",x"ED",
		x"B0",x"3E",x"01",x"32",x"B9",x"62",x"C9",x"21",x"EC",x"3D",x"11",x"07",x"64",x"01",x"1C",x"05",
		x"CD",x"2A",x"12",x"CD",x"86",x"11",x"21",x"00",x"66",x"11",x"10",x"00",x"3E",x"01",x"06",x"06",
		x"77",x"19",x"10",x"FC",x"0E",x"02",x"3E",x"08",x"06",x"03",x"21",x"0D",x"66",x"77",x"19",x"10",
		x"FC",x"3E",x"08",x"0D",x"C2",x"A8",x"10",x"21",x"64",x"3E",x"11",x"03",x"66",x"01",x"0E",x"06",
		x"CD",x"EC",x"11",x"21",x"60",x"3E",x"11",x"07",x"66",x"01",x"0C",x"06",x"CD",x"2A",x"12",x"DD",
		x"21",x"00",x"66",x"21",x"58",x"69",x"06",x"06",x"11",x"10",x"00",x"CD",x"D3",x"11",x"21",x"48",
		x"3E",x"11",x"0C",x"6A",x"01",x"0C",x"00",x"ED",x"B0",x"DD",x"21",x"00",x"64",x"DD",x"36",x"00",
		x"01",x"DD",x"36",x"03",x"58",x"DD",x"36",x"0E",x"58",x"DD",x"36",x"05",x"80",x"DD",x"36",x"0F",
		x"80",x"DD",x"36",x"20",x"01",x"DD",x"36",x"23",x"EB",x"DD",x"36",x"2E",x"EB",x"DD",x"36",x"25",
		x"60",x"DD",x"36",x"2F",x"60",x"11",x"70",x"69",x"21",x"21",x"11",x"01",x"10",x"00",x"ED",x"B0",
		x"C9",x"37",x"45",x"0F",x"60",x"37",x"45",x"8F",x"F7",x"77",x"45",x"0F",x"60",x"77",x"45",x"8F",
		x"F7",x"21",x"F0",x"3D",x"11",x"07",x"64",x"01",x"1C",x"05",x"CD",x"2A",x"12",x"21",x"14",x"3E",
		x"CD",x"A6",x"11",x"21",x"54",x"3E",x"11",x"0C",x"6A",x"01",x"0C",x"00",x"ED",x"B0",x"21",x"82",
		x"11",x"11",x"A3",x"64",x"01",x"1E",x"02",x"CD",x"EC",x"11",x"21",x"7E",x"11",x"11",x"A7",x"64",
		x"01",x"1C",x"02",x"CD",x"2A",x"12",x"DD",x"21",x"A0",x"64",x"DD",x"36",x"00",x"01",x"DD",x"36",
		x"20",x"01",x"21",x"50",x"69",x"06",x"02",x"11",x"20",x"00",x"CD",x"D3",x"11",x"C9",x"3F",x"0C",
		x"08",x"08",x"73",x"50",x"8D",x"50",x"21",x"A2",x"11",x"11",x"07",x"65",x"01",x"0C",x"0A",x"CD",
		x"2A",x"12",x"DD",x"21",x"00",x"65",x"21",x"80",x"69",x"06",x"0A",x"11",x"10",x"00",x"CD",x"D3",
		x"11",x"C9",x"3B",x"00",x"02",x"02",x"11",x"83",x"66",x"01",x"0E",x"02",x"CD",x"EC",x"11",x"21",
		x"08",x"3E",x"11",x"87",x"66",x"01",x"0C",x"02",x"CD",x"2A",x"12",x"DD",x"21",x"80",x"66",x"DD",
		x"36",x"00",x"01",x"DD",x"36",x"10",x"01",x"21",x"18",x"6A",x"06",x"02",x"11",x"10",x"00",x"CD",
		x"D3",x"11",x"C9",x"DD",x"7E",x"03",x"77",x"2C",x"DD",x"7E",x"07",x"77",x"2C",x"DD",x"7E",x"08",
		x"77",x"2C",x"DD",x"7E",x"05",x"77",x"2C",x"DD",x"19",x"10",x"E8",x"C9",x"7E",x"12",x"23",x"1C",
		x"1C",x"7E",x"12",x"23",x"7B",x"81",x"5F",x"10",x"F3",x"C9",x"DD",x"21",x"A0",x"66",x"11",x"28",
		x"6A",x"DD",x"36",x"00",x"01",x"7E",x"DD",x"77",x"03",x"12",x"1C",x"23",x"7E",x"DD",x"77",x"07",
		x"12",x"1C",x"23",x"7E",x"DD",x"77",x"08",x"12",x"1C",x"23",x"7E",x"DD",x"77",x"05",x"12",x"23",
		x"7E",x"DD",x"77",x"09",x"23",x"7E",x"DD",x"77",x"0A",x"C9",x"E5",x"C5",x"06",x"04",x"7E",x"12",
		x"23",x"1C",x"10",x"FA",x"C1",x"E1",x"7B",x"81",x"5F",x"10",x"EF",x"C9",x"DF",x"3A",x"27",x"62",
		x"FE",x"03",x"01",x"16",x"E0",x"CA",x"4B",x"12",x"01",x"3F",x"F0",x"DD",x"21",x"00",x"62",x"21",
		x"4C",x"69",x"DD",x"36",x"00",x"01",x"DD",x"71",x"03",x"71",x"2C",x"DD",x"36",x"07",x"80",x"36",
		x"80",x"2C",x"DD",x"36",x"08",x"02",x"36",x"02",x"2C",x"DD",x"70",x"05",x"70",x"DD",x"36",x"0F",
		x"01",x"21",x"0A",x"60",x"34",x"11",x"01",x"06",x"CD",x"9F",x"30",x"C9",x"CD",x"BD",x"1D",x"3A",
		x"9D",x"63",x"EF",x"8B",x"12",x"AC",x"12",x"DE",x"12",x"00",x"00",x"DF",x"21",x"4D",x"69",x"3E",
		x"F0",x"CB",x"16",x"1F",x"77",x"21",x"9D",x"63",x"34",x"3E",x"0D",x"32",x"9E",x"63",x"3E",x"08",
		x"32",x"09",x"60",x"CD",x"BD",x"30",x"3E",x"03",x"32",x"88",x"60",x"C9",x"DF",x"3E",x"08",x"32",
		x"09",x"60",x"21",x"9E",x"63",x"35",x"CA",x"CB",x"12",x"21",x"4D",x"69",x"7E",x"1F",x"3E",x"02",
		x"1F",x"47",x"AE",x"77",x"2C",x"78",x"E6",x"80",x"AE",x"77",x"C9",x"21",x"4D",x"69",x"3E",x"F4",
		x"CB",x"16",x"1F",x"77",x"21",x"9D",x"63",x"34",x"3E",x"80",x"32",x"09",x"60",x"C9",x"DF",x"CD",
		x"DB",x"30",x"21",x"0A",x"60",x"3A",x"0E",x"60",x"A7",x"CA",x"ED",x"12",x"34",x"34",x"2B",x"36",
		x"01",x"C9",x"CD",x"1C",x"01",x"AF",x"32",x"2C",x"62",x"21",x"28",x"62",x"35",x"7E",x"11",x"40",
		x"60",x"01",x"08",x"00",x"ED",x"B0",x"A7",x"C2",x"34",x"13",x"3E",x"01",x"21",x"B2",x"60",x"CD",
		x"CA",x"13",x"21",x"D4",x"76",x"3A",x"0F",x"60",x"A7",x"28",x"07",x"11",x"02",x"03",x"CD",x"9F",
		x"30",x"2B",x"CD",x"26",x"18",x"11",x"00",x"03",x"CD",x"9F",x"30",x"21",x"09",x"60",x"36",x"C0",
		x"23",x"36",x"10",x"C9",x"0E",x"08",x"3A",x"0F",x"60",x"A7",x"CA",x"3F",x"13",x"0E",x"17",x"79",
		x"32",x"0A",x"60",x"C9",x"CD",x"1C",x"01",x"AF",x"32",x"2C",x"62",x"21",x"28",x"62",x"35",x"7E",
		x"11",x"48",x"60",x"01",x"08",x"00",x"ED",x"B0",x"A7",x"C2",x"7F",x"13",x"3E",x"03",x"21",x"B5",
		x"60",x"CD",x"CA",x"13",x"11",x"03",x"03",x"CD",x"9F",x"30",x"11",x"00",x"03",x"CD",x"9F",x"30",
		x"21",x"D3",x"76",x"CD",x"26",x"18",x"21",x"09",x"60",x"36",x"C0",x"23",x"36",x"11",x"C9",x"0E",
		x"17",x"3A",x"40",x"60",x"A7",x"C2",x"8A",x"13",x"0E",x"08",x"79",x"32",x"0A",x"60",x"C9",x"DF",
		x"0E",x"17",x"3A",x"48",x"60",x"34",x"A7",x"C2",x"9C",x"13",x"0E",x"14",x"79",x"32",x"0A",x"60",
		x"C9",x"DF",x"0E",x"17",x"3A",x"40",x"60",x"C3",x"95",x"13",x"3A",x"26",x"60",x"32",x"82",x"7D",
		x"AF",x"32",x"0A",x"60",x"21",x"01",x"01",x"22",x"0D",x"60",x"C9",x"AF",x"32",x"0D",x"60",x"32",
		x"0E",x"60",x"32",x"0A",x"60",x"3C",x"32",x"82",x"7D",x"C9",x"11",x"C6",x"61",x"12",x"CF",x"13",
		x"01",x"03",x"00",x"ED",x"B0",x"06",x"03",x"21",x"B1",x"61",x"1B",x"1A",x"0F",x"0F",x"0F",x"0F",
		x"E6",x"0F",x"77",x"23",x"1A",x"E6",x"0F",x"77",x"23",x"10",x"EF",x"06",x"0E",x"36",x"10",x"23",
		x"10",x"FB",x"36",x"3F",x"06",x"05",x"21",x"A5",x"61",x"11",x"C7",x"61",x"1A",x"96",x"23",x"13",
		x"1A",x"9E",x"23",x"13",x"1A",x"9E",x"D8",x"C5",x"06",x"19",x"4E",x"1A",x"77",x"79",x"12",x"2B",
		x"1B",x"10",x"F7",x"01",x"F5",x"FF",x"09",x"EB",x"09",x"EB",x"C1",x"10",x"DF",x"C9",x"CD",x"16",
		x"06",x"DF",x"CD",x"74",x"08",x"3E",x"00",x"32",x"0E",x"60",x"32",x"0D",x"60",x"21",x"1C",x"61",
		x"11",x"22",x"00",x"06",x"05",x"3E",x"01",x"BE",x"CA",x"59",x"14",x"19",x"10",x"F9",x"21",x"1C",
		x"61",x"06",x"05",x"3E",x"03",x"BE",x"CA",x"4F",x"14",x"19",x"10",x"F9",x"C3",x"75",x"14",x"3E",
		x"01",x"32",x"0E",x"60",x"32",x"0D",x"60",x"3E",x"00",x"21",x"26",x"60",x"B6",x"32",x"82",x"7D",
		x"3E",x"00",x"32",x"09",x"60",x"21",x"0A",x"60",x"34",x"11",x"0D",x"03",x"06",x"0C",x"CD",x"9F",
		x"30",x"13",x"10",x"FA",x"C9",x"3E",x"01",x"32",x"82",x"7D",x"32",x"05",x"60",x"32",x"07",x"60",
		x"3E",x"00",x"32",x"0A",x"60",x"C9",x"CD",x"16",x"06",x"21",x"09",x"60",x"7E",x"A7",x"C2",x"DC",
		x"14",x"32",x"86",x"7D",x"32",x"87",x"7D",x"36",x"01",x"21",x"30",x"60",x"36",x"0A",x"23",x"36",
		x"00",x"23",x"36",x"10",x"23",x"36",x"1E",x"23",x"36",x"3E",x"23",x"36",x"00",x"21",x"E8",x"75",
		x"22",x"36",x"60",x"21",x"1C",x"61",x"3A",x"0E",x"60",x"07",x"3C",x"4F",x"11",x"22",x"00",x"06",
		x"04",x"7E",x"B9",x"CA",x"C9",x"14",x"19",x"10",x"F8",x"22",x"38",x"60",x"11",x"F3",x"FF",x"19",
		x"22",x"3A",x"60",x"06",x"00",x"3A",x"35",x"60",x"4F",x"CD",x"FA",x"15",x"21",x"34",x"60",x"35",
		x"C2",x"FC",x"14",x"36",x"3E",x"2B",x"35",x"CA",x"C6",x"15",x"7E",x"06",x"FF",x"04",x"D6",x"0A",
		x"D2",x"ED",x"14",x"C6",x"0A",x"32",x"52",x"75",x"78",x"32",x"72",x"75",x"21",x"30",x"60",x"46",
		x"36",x"0A",x"3A",x"10",x"60",x"CB",x"7F",x"C2",x"46",x"15",x"E6",x"03",x"C2",x"14",x"15",x"3C",
		x"77",x"C3",x"8A",x"15",x"05",x"CA",x"1D",x"15",x"78",x"77",x"C3",x"8A",x"15",x"CB",x"4F",x"C2",
		x"39",x"15",x"3A",x"35",x"60",x"3C",x"FE",x"1E",x"C2",x"2D",x"15",x"3E",x"00",x"32",x"35",x"60",
		x"4F",x"06",x"00",x"CD",x"FA",x"15",x"C3",x"8A",x"15",x"3A",x"35",x"60",x"D6",x"01",x"F2",x"2D",
		x"15",x"3E",x"1D",x"C3",x"2D",x"15",x"3A",x"35",x"60",x"FE",x"1C",x"CA",x"6D",x"15",x"FE",x"1D",
		x"CA",x"C6",x"15",x"2A",x"36",x"60",x"01",x"88",x"75",x"A7",x"ED",x"42",x"CA",x"8A",x"15",x"09",
		x"C6",x"11",x"77",x"01",x"E0",x"FF",x"09",x"22",x"36",x"60",x"C3",x"8A",x"15",x"2A",x"36",x"60",
		x"01",x"20",x"00",x"09",x"A7",x"01",x"08",x"76",x"ED",x"42",x"C2",x"86",x"15",x"21",x"E8",x"75",
		x"3E",x"10",x"77",x"C3",x"67",x"15",x"09",x"C3",x"80",x"15",x"21",x"32",x"60",x"35",x"C2",x"F9",
		x"15",x"3A",x"31",x"60",x"A7",x"C2",x"B8",x"15",x"3E",x"01",x"32",x"31",x"60",x"11",x"BF",x"01",
		x"FD",x"2A",x"38",x"60",x"FD",x"6E",x"04",x"FD",x"66",x"05",x"E5",x"DD",x"E1",x"CD",x"7C",x"05",
		x"3E",x"10",x"32",x"32",x"60",x"C3",x"F9",x"15",x"AF",x"32",x"31",x"60",x"ED",x"5B",x"38",x"60",
		x"13",x"13",x"13",x"C3",x"A0",x"15",x"ED",x"5B",x"38",x"60",x"AF",x"12",x"21",x"09",x"60",x"36",
		x"80",x"23",x"35",x"06",x"0C",x"21",x"E8",x"75",x"FD",x"2A",x"3A",x"60",x"11",x"E0",x"FF",x"7E",
		x"FD",x"77",x"00",x"FD",x"23",x"19",x"10",x"F7",x"06",x"05",x"11",x"14",x"03",x"CD",x"9F",x"30",
		x"13",x"10",x"FA",x"11",x"1A",x"03",x"CD",x"9F",x"30",x"C9",x"D5",x"E5",x"CB",x"21",x"21",x"0F",
		x"36",x"09",x"EB",x"21",x"74",x"69",x"1A",x"13",x"77",x"23",x"36",x"72",x"23",x"36",x"0C",x"23",
		x"1A",x"77",x"E1",x"D1",x"C9",x"CD",x"BD",x"30",x"3A",x"27",x"62",x"0F",x"D2",x"2F",x"16",x"3A",
		x"88",x"63",x"EF",x"54",x"16",x"70",x"16",x"8A",x"16",x"32",x"17",x"57",x"17",x"8E",x"17",x"0F",
		x"D2",x"41",x"16",x"3A",x"88",x"63",x"EF",x"A3",x"16",x"BB",x"16",x"32",x"17",x"57",x"17",x"8E",
		x"17",x"CD",x"BD",x"1D",x"3A",x"88",x"63",x"EF",x"B6",x"17",x"69",x"30",x"39",x"18",x"6F",x"18",
		x"80",x"18",x"C6",x"18",x"CD",x"08",x"17",x"21",x"5C",x"38",x"CD",x"4E",x"00",x"3E",x"20",x"32",
		x"09",x"60",x"21",x"88",x"63",x"34",x"3E",x"01",x"F7",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"C9",
		x"DF",x"21",x"32",x"39",x"CD",x"4E",x"00",x"3E",x"20",x"32",x"09",x"60",x"21",x"88",x"63",x"34",
		x"3E",x"04",x"F7",x"21",x"0B",x"69",x"0E",x"04",x"FF",x"C9",x"DF",x"21",x"8C",x"38",x"CD",x"4E",
		x"00",x"3E",x"66",x"32",x"0C",x"69",x"AF",x"32",x"24",x"69",x"32",x"2C",x"69",x"32",x"AF",x"62",
		x"C3",x"62",x"16",x"CD",x"08",x"17",x"3A",x"10",x"69",x"D6",x"3B",x"21",x"5C",x"38",x"CD",x"4E",
		x"00",x"21",x"08",x"69",x"4F",x"FF",x"21",x"88",x"63",x"34",x"C9",x"AF",x"32",x"A0",x"62",x"3A",
		x"A3",x"63",x"4F",x"3A",x"10",x"69",x"FE",x"5A",x"D2",x"E1",x"16",x"CB",x"79",x"CA",x"D5",x"16",
		x"3E",x"01",x"32",x"A0",x"62",x"CD",x"02",x"26",x"3A",x"A3",x"63",x"4F",x"21",x"08",x"69",x"FF",
		x"C9",x"FE",x"5D",x"DA",x"EE",x"16",x"CB",x"79",x"CA",x"D0",x"16",x"C3",x"D5",x"16",x"21",x"8C",
		x"38",x"CD",x"4E",x"00",x"3E",x"66",x"32",x"0C",x"69",x"AF",x"32",x"24",x"69",x"32",x"2C",x"69",
		x"32",x"AF",x"62",x"21",x"88",x"63",x"34",x"C9",x"CD",x"1C",x"01",x"21",x"20",x"6A",x"36",x"80",
		x"23",x"36",x"76",x"23",x"36",x"09",x"23",x"36",x"20",x"21",x"05",x"69",x"36",x"13",x"21",x"C4",
		x"75",x"11",x"20",x"00",x"3E",x"10",x"CD",x"14",x"05",x"21",x"8A",x"60",x"36",x"07",x"23",x"36",
		x"03",x"C9",x"CD",x"6F",x"30",x"3A",x"13",x"69",x"FE",x"2C",x"D0",x"AF",x"32",x"00",x"69",x"32",
		x"04",x"69",x"32",x"0C",x"69",x"3E",x"6B",x"32",x"24",x"69",x"3D",x"32",x"2C",x"69",x"21",x"21",
		x"6A",x"34",x"21",x"88",x"63",x"34",x"C9",x"CD",x"6F",x"30",x"CD",x"6C",x"17",x"23",x"13",x"CD",
		x"83",x"17",x"3E",x"40",x"32",x"09",x"60",x"21",x"88",x"63",x"34",x"C9",x"11",x"03",x"00",x"21",
		x"2F",x"69",x"06",x"0A",x"A7",x"7E",x"ED",x"52",x"FE",x"19",x"D2",x"7F",x"17",x"36",x"00",x"2B",
		x"10",x"F2",x"C9",x"06",x"0A",x"7E",x"A7",x"C2",x"26",x"00",x"19",x"10",x"F8",x"C9",x"DF",x"2A",
		x"2A",x"62",x"23",x"7E",x"FE",x"7F",x"C2",x"9D",x"17",x"21",x"73",x"3A",x"7E",x"22",x"2A",x"62",
		x"32",x"27",x"62",x"11",x"00",x"05",x"CD",x"9F",x"30",x"AF",x"32",x"88",x"63",x"21",x"09",x"60",
		x"36",x"30",x"23",x"36",x"08",x"C9",x"00",x"CD",x"1C",x"01",x"21",x"8A",x"60",x"36",x"0E",x"23",
		x"36",x"03",x"3E",x"10",x"11",x"20",x"00",x"21",x"23",x"76",x"CD",x"14",x"05",x"21",x"83",x"75",
		x"CD",x"14",x"05",x"21",x"DA",x"76",x"CD",x"26",x"18",x"11",x"47",x"3A",x"CD",x"A7",x"0D",x"21",
		x"D5",x"76",x"CD",x"26",x"18",x"11",x"4D",x"3A",x"CD",x"A7",x"0D",x"21",x"D0",x"76",x"CD",x"26",
		x"18",x"11",x"53",x"3A",x"CD",x"A7",x"0D",x"21",x"CB",x"76",x"CD",x"26",x"18",x"11",x"59",x"3A",
		x"CD",x"A7",x"0D",x"21",x"5C",x"38",x"CD",x"4E",x"00",x"21",x"08",x"69",x"0E",x"44",x"FF",x"21",
		x"05",x"69",x"36",x"13",x"3E",x"20",x"32",x"09",x"60",x"3E",x"80",x"32",x"90",x"63",x"21",x"88",
		x"63",x"34",x"22",x"C0",x"63",x"C9",x"11",x"DB",x"FF",x"0E",x"0E",x"3E",x"10",x"06",x"05",x"77",
		x"23",x"10",x"FC",x"19",x"0D",x"C2",x"2D",x"18",x"C9",x"21",x"90",x"63",x"34",x"CA",x"59",x"18",
		x"7E",x"E6",x"07",x"C0",x"11",x"CF",x"39",x"CB",x"5E",x"20",x"03",x"11",x"F7",x"39",x"EB",x"CD",
		x"4E",x"00",x"21",x"08",x"69",x"0E",x"44",x"FF",x"C9",x"21",x"5C",x"38",x"CD",x"4E",x"00",x"21",
		x"08",x"69",x"0E",x"44",x"FF",x"3E",x"20",x"32",x"09",x"60",x"21",x"88",x"63",x"34",x"C9",x"DF",
		x"21",x"1F",x"3A",x"CD",x"4E",x"00",x"3E",x"03",x"32",x"84",x"60",x"21",x"88",x"63",x"34",x"C9",
		x"21",x"0B",x"69",x"0E",x"01",x"FF",x"3A",x"1B",x"69",x"FE",x"D0",x"C0",x"3E",x"20",x"32",x"19",
		x"69",x"21",x"24",x"6A",x"36",x"7F",x"2C",x"36",x"39",x"2C",x"36",x"01",x"2C",x"36",x"D8",x"21",
		x"C6",x"76",x"CD",x"26",x"18",x"11",x"5F",x"3A",x"CD",x"A7",x"0D",x"11",x"04",x"00",x"01",x"28",
		x"02",x"21",x"03",x"69",x"CD",x"3D",x"00",x"3E",x"00",x"32",x"AF",x"62",x"3E",x"03",x"32",x"82",
		x"60",x"21",x"88",x"63",x"34",x"C9",x"21",x"AF",x"62",x"35",x"CA",x"3D",x"19",x"7E",x"E6",x"07",
		x"C0",x"21",x"25",x"6A",x"7E",x"EE",x"80",x"77",x"21",x"19",x"69",x"46",x"CB",x"A8",x"AF",x"CD",
		x"09",x"30",x"F6",x"20",x"77",x"21",x"AF",x"62",x"7E",x"FE",x"E0",x"C2",x"10",x"19",x"3E",x"50",
		x"32",x"4F",x"69",x"3E",x"00",x"32",x"4D",x"69",x"3E",x"9F",x"32",x"4C",x"69",x"3A",x"03",x"62",
		x"FE",x"80",x"D2",x"0F",x"19",x"3E",x"80",x"32",x"4D",x"69",x"3E",x"5F",x"32",x"4C",x"69",x"7E",
		x"FE",x"C0",x"C0",x"21",x"8A",x"60",x"36",x"0C",x"3A",x"29",x"62",x"0F",x"38",x"02",x"36",x"05",
		x"23",x"36",x"03",x"21",x"23",x"6A",x"36",x"40",x"2B",x"36",x"09",x"2B",x"36",x"76",x"2B",x"36",
		x"8F",x"3A",x"03",x"62",x"FE",x"80",x"D0",x"3E",x"6F",x"32",x"20",x"6A",x"C9",x"2A",x"2A",x"62",
		x"23",x"7E",x"FE",x"7F",x"C2",x"4B",x"19",x"21",x"73",x"3A",x"7E",x"22",x"2A",x"62",x"32",x"27",
		x"62",x"21",x"29",x"62",x"34",x"11",x"00",x"05",x"CD",x"9F",x"30",x"AF",x"32",x"2E",x"62",x"32",
		x"88",x"63",x"21",x"09",x"60",x"36",x"E0",x"23",x"36",x"08",x"C9",x"CD",x"52",x"08",x"3A",x"0E",
		x"60",x"C6",x"12",x"32",x"0A",x"60",x"C9",x"CD",x"EE",x"21",x"CD",x"BD",x"1D",x"CD",x"8C",x"1E",
		x"CD",x"C3",x"1A",x"CD",x"72",x"1F",x"CD",x"8F",x"2C",x"CD",x"03",x"2C",x"CD",x"ED",x"30",x"CD",
		x"04",x"2E",x"CD",x"EA",x"24",x"CD",x"DB",x"2D",x"CD",x"D4",x"2E",x"CD",x"07",x"22",x"CD",x"33",
		x"1A",x"CD",x"85",x"2A",x"CD",x"46",x"1F",x"CD",x"FA",x"26",x"CD",x"F2",x"25",x"CD",x"DA",x"19",
		x"CD",x"FB",x"03",x"CD",x"08",x"28",x"CD",x"1D",x"28",x"CD",x"57",x"1E",x"CD",x"07",x"1A",x"CD",
		x"CB",x"2F",x"00",x"00",x"00",x"3A",x"00",x"62",x"A7",x"C0",x"CD",x"1C",x"01",x"21",x"82",x"60",
		x"36",x"03",x"21",x"0A",x"60",x"34",x"2B",x"36",x"40",x"C9",x"3A",x"03",x"62",x"06",x"03",x"21",
		x"0C",x"6A",x"BE",x"CA",x"ED",x"19",x"2C",x"2C",x"2C",x"2C",x"10",x"F6",x"C9",x"3A",x"05",x"62",
		x"2C",x"2C",x"2C",x"BE",x"C0",x"2D",x"2D",x"CB",x"5E",x"C0",x"2D",x"22",x"43",x"63",x"AF",x"32",
		x"42",x"63",x"3C",x"32",x"40",x"63",x"C9",x"3A",x"86",x"63",x"EF",x"1E",x"1A",x"15",x"1A",x"1F",
		x"1A",x"2A",x"1A",x"00",x"00",x"AF",x"32",x"87",x"63",x"3E",x"02",x"32",x"86",x"63",x"C9",x"21",
		x"87",x"63",x"35",x"C0",x"3E",x"03",x"32",x"86",x"63",x"C9",x"3A",x"16",x"62",x"A7",x"C0",x"E1",
		x"C3",x"D2",x"19",x"3E",x"08",x"F7",x"3A",x"03",x"62",x"FE",x"4B",x"CA",x"4B",x"1A",x"FE",x"B3",
		x"CA",x"4B",x"1A",x"3A",x"91",x"62",x"3D",x"CA",x"51",x"1A",x"C9",x"3E",x"01",x"32",x"91",x"62",
		x"C9",x"32",x"91",x"62",x"47",x"3A",x"05",x"62",x"3D",x"FE",x"D0",x"D0",x"07",x"D2",x"62",x"1A",
		x"CB",x"D0",x"07",x"07",x"D2",x"69",x"1A",x"CB",x"C8",x"E6",x"07",x"FE",x"06",x"C2",x"72",x"1A",
		x"CB",x"C8",x"3A",x"03",x"62",x"07",x"D2",x"7B",x"1A",x"CB",x"C0",x"21",x"92",x"62",x"78",x"85",
		x"6F",x"7E",x"A7",x"C8",x"36",x"00",x"21",x"90",x"62",x"35",x"78",x"01",x"05",x"00",x"1F",x"DA",
		x"BD",x"1A",x"21",x"CB",x"02",x"A7",x"CA",x"9E",x"1A",x"09",x"3D",x"C2",x"99",x"1A",x"01",x"00",
		x"74",x"09",x"3E",x"10",x"77",x"2D",x"77",x"2C",x"2C",x"77",x"3E",x"01",x"32",x"40",x"63",x"32",
		x"42",x"63",x"32",x"25",x"62",x"3A",x"16",x"62",x"A7",x"CC",x"95",x"1D",x"C9",x"21",x"2B",x"01",
		x"C3",x"95",x"1A",x"3A",x"16",x"62",x"3D",x"CA",x"B2",x"1B",x"3A",x"1E",x"62",x"A7",x"C2",x"55",
		x"1B",x"3A",x"17",x"62",x"3D",x"CA",x"E6",x"1A",x"3A",x"15",x"62",x"3D",x"CA",x"38",x"1B",x"3A",
		x"10",x"60",x"17",x"DA",x"6E",x"1B",x"CD",x"1F",x"24",x"3A",x"10",x"60",x"1D",x"CA",x"F5",x"1A",
		x"CB",x"47",x"C2",x"8F",x"1C",x"15",x"CA",x"FE",x"1A",x"CB",x"4F",x"C2",x"AB",x"1C",x"3A",x"17",
		x"62",x"3D",x"C8",x"3A",x"05",x"62",x"C6",x"08",x"57",x"3A",x"03",x"62",x"F6",x"03",x"CB",x"97",
		x"01",x"15",x"00",x"CD",x"6E",x"23",x"F5",x"21",x"07",x"62",x"7E",x"E6",x"80",x"F6",x"06",x"77",
		x"21",x"1A",x"62",x"3E",x"04",x"B9",x"36",x"01",x"D2",x"2C",x"1B",x"35",x"F1",x"A7",x"CA",x"4E",
		x"1B",x"7E",x"A7",x"C0",x"2C",x"72",x"2C",x"70",x"3A",x"10",x"60",x"CB",x"5F",x"C2",x"F2",x"1C",
		x"3A",x"15",x"62",x"A7",x"C8",x"3A",x"10",x"60",x"CB",x"57",x"C2",x"03",x"1D",x"C9",x"2C",x"70",
		x"2C",x"72",x"C3",x"45",x"1B",x"21",x"1E",x"62",x"35",x"C0",x"3A",x"18",x"62",x"32",x"17",x"62",
		x"21",x"07",x"62",x"7E",x"E6",x"80",x"77",x"AF",x"32",x"02",x"62",x"C3",x"A6",x"1D",x"3E",x"01",
		x"32",x"16",x"62",x"21",x"10",x"62",x"3A",x"10",x"60",x"01",x"80",x"00",x"1F",x"DA",x"8A",x"1B",
		x"01",x"80",x"FF",x"1F",x"DA",x"8A",x"1B",x"01",x"00",x"00",x"AF",x"70",x"2C",x"71",x"2C",x"36",
		x"01",x"2C",x"36",x"48",x"2C",x"77",x"32",x"04",x"62",x"32",x"06",x"62",x"3A",x"07",x"62",x"E6",
		x"80",x"F6",x"0E",x"32",x"07",x"62",x"3A",x"05",x"62",x"32",x"0E",x"62",x"21",x"81",x"60",x"36",
		x"03",x"C9",x"DD",x"21",x"00",x"62",x"3A",x"03",x"62",x"DD",x"77",x"0B",x"3A",x"05",x"62",x"DD",
		x"77",x"0C",x"CD",x"9C",x"23",x"CD",x"1F",x"24",x"15",x"C2",x"F2",x"1B",x"DD",x"36",x"10",x"00",
		x"DD",x"36",x"11",x"80",x"DD",x"CB",x"07",x"FE",x"3A",x"20",x"62",x"3D",x"CA",x"EC",x"1B",x"CD",
		x"07",x"24",x"DD",x"74",x"12",x"DD",x"75",x"13",x"DD",x"36",x"14",x"00",x"CD",x"9C",x"23",x"C3",
		x"05",x"1C",x"1D",x"C2",x"05",x"1C",x"DD",x"36",x"10",x"FF",x"DD",x"36",x"11",x"80",x"DD",x"CB",
		x"07",x"BE",x"C3",x"D8",x"1B",x"CD",x"1C",x"2B",x"3D",x"CA",x"3A",x"1C",x"3A",x"1F",x"62",x"3D",
		x"CA",x"76",x"1C",x"3A",x"14",x"62",x"D6",x"14",x"C2",x"33",x"1C",x"3E",x"01",x"32",x"1F",x"62",
		x"CD",x"53",x"28",x"A7",x"CA",x"A6",x"1D",x"32",x"42",x"63",x"3E",x"01",x"32",x"40",x"63",x"32",
		x"25",x"62",x"00",x"3C",x"CC",x"54",x"29",x"C3",x"A6",x"1D",x"05",x"CA",x"4F",x"1C",x"3C",x"32",
		x"1F",x"62",x"AF",x"21",x"10",x"62",x"06",x"05",x"77",x"2C",x"10",x"FC",x"C3",x"A6",x"1D",x"32",
		x"16",x"62",x"3A",x"20",x"62",x"EE",x"01",x"32",x"00",x"62",x"21",x"07",x"62",x"7E",x"E6",x"80",
		x"F6",x"0F",x"77",x"3E",x"04",x"32",x"1E",x"62",x"AF",x"32",x"1F",x"62",x"3A",x"25",x"62",x"3D",
		x"CC",x"95",x"1D",x"C3",x"A6",x"1D",x"3A",x"05",x"62",x"21",x"0E",x"62",x"D6",x"0F",x"BE",x"DA",
		x"A6",x"1D",x"3E",x"01",x"32",x"20",x"62",x"21",x"84",x"60",x"36",x"03",x"C3",x"A6",x"1D",x"06",
		x"01",x"3A",x"0F",x"62",x"A7",x"C2",x"D2",x"1C",x"3A",x"02",x"62",x"47",x"3E",x"05",x"CD",x"09",
		x"30",x"32",x"02",x"62",x"E6",x"03",x"F6",x"80",x"C3",x"C2",x"1C",x"06",x"FF",x"3A",x"0F",x"62",
		x"A7",x"C2",x"D2",x"1C",x"3A",x"02",x"62",x"47",x"3E",x"01",x"CD",x"09",x"30",x"32",x"02",x"62",
		x"E6",x"03",x"21",x"07",x"62",x"77",x"1F",x"DC",x"8F",x"1D",x"3E",x"02",x"32",x"0F",x"62",x"C3",
		x"A6",x"1D",x"21",x"03",x"62",x"7E",x"80",x"77",x"3A",x"27",x"62",x"3D",x"C2",x"EB",x"1C",x"66",
		x"3A",x"05",x"62",x"6F",x"CD",x"33",x"23",x"7D",x"32",x"05",x"62",x"21",x"0F",x"62",x"35",x"C3",
		x"A6",x"1D",x"3A",x"0F",x"62",x"A7",x"C2",x"8A",x"1D",x"3E",x"03",x"32",x"0F",x"62",x"3E",x"02",
		x"C3",x"11",x"1D",x"3A",x"0F",x"62",x"A7",x"C2",x"76",x"1D",x"3E",x"04",x"32",x"0F",x"62",x"3E",
		x"FE",x"21",x"05",x"62",x"86",x"77",x"47",x"3A",x"22",x"62",x"EE",x"01",x"32",x"22",x"62",x"C2",
		x"51",x"1D",x"78",x"C6",x"08",x"21",x"1C",x"62",x"BE",x"CA",x"67",x"1D",x"2D",x"96",x"CA",x"67",
		x"1D",x"06",x"05",x"D6",x"08",x"CA",x"3F",x"1D",x"05",x"D6",x"04",x"CA",x"3F",x"1D",x"05",x"3E",
		x"80",x"21",x"07",x"62",x"A6",x"EE",x"80",x"B0",x"77",x"3E",x"01",x"32",x"15",x"62",x"C3",x"A6",
		x"1D",x"2D",x"2D",x"7E",x"F6",x"03",x"CB",x"97",x"77",x"3A",x"24",x"62",x"EE",x"01",x"32",x"24",
		x"62",x"CC",x"8F",x"1D",x"C3",x"49",x"1D",x"3E",x"06",x"32",x"07",x"62",x"AF",x"32",x"19",x"62",
		x"32",x"15",x"62",x"C3",x"A6",x"1D",x"3A",x"1A",x"62",x"A7",x"CA",x"8A",x"1D",x"32",x"19",x"62",
		x"3A",x"1C",x"62",x"D6",x"13",x"21",x"05",x"62",x"BE",x"D0",x"21",x"0F",x"62",x"35",x"C9",x"3E",
		x"03",x"32",x"80",x"60",x"C9",x"32",x"25",x"62",x"3A",x"27",x"62",x"3D",x"C8",x"21",x"8A",x"60",
		x"36",x"0D",x"2C",x"36",x"03",x"C9",x"21",x"4C",x"69",x"3A",x"03",x"62",x"77",x"3A",x"07",x"62",
		x"2C",x"77",x"3A",x"08",x"62",x"2C",x"77",x"3A",x"05",x"62",x"2C",x"77",x"C9",x"3A",x"40",x"63",
		x"EF",x"49",x"1E",x"C9",x"1D",x"4A",x"1E",x"00",x"00",x"3E",x"40",x"32",x"41",x"63",x"3E",x"02",
		x"32",x"40",x"63",x"3A",x"42",x"63",x"1F",x"DA",x"70",x"3E",x"1F",x"DA",x"00",x"1E",x"1F",x"DA",
		x"F5",x"1D",x"21",x"85",x"60",x"36",x"03",x"3A",x"29",x"62",x"3D",x"CA",x"00",x"1E",x"3D",x"CA",
		x"08",x"1E",x"C3",x"10",x"1E",x"3A",x"18",x"60",x"1F",x"DA",x"08",x"1E",x"1F",x"DA",x"10",x"1E",
		x"06",x"7D",x"11",x"03",x"00",x"C3",x"15",x"1E",x"06",x"7E",x"11",x"05",x"00",x"C3",x"15",x"1E",
		x"06",x"7F",x"11",x"08",x"00",x"CD",x"9F",x"30",x"2A",x"43",x"63",x"7E",x"36",x"00",x"2C",x"2C",
		x"2C",x"4E",x"C3",x"36",x"1E",x"11",x"01",x"00",x"CD",x"9F",x"30",x"3A",x"05",x"62",x"C6",x"14",
		x"4F",x"3A",x"03",x"62",x"00",x"00",x"21",x"30",x"6A",x"77",x"2C",x"70",x"2C",x"36",x"07",x"2C",
		x"71",x"3E",x"05",x"F7",x"21",x"85",x"60",x"36",x"03",x"C9",x"21",x"41",x"63",x"35",x"C0",x"AF",
		x"32",x"30",x"6A",x"32",x"40",x"63",x"C9",x"3A",x"27",x"62",x"CB",x"57",x"C2",x"80",x"1E",x"1F",
		x"3A",x"05",x"62",x"DA",x"7A",x"1E",x"FE",x"51",x"D0",x"3A",x"03",x"62",x"17",x"3E",x"00",x"DA",
		x"74",x"1E",x"3E",x"80",x"32",x"4D",x"69",x"C3",x"85",x"1E",x"FE",x"31",x"D0",x"C3",x"6D",x"1E",
		x"3A",x"90",x"62",x"A7",x"C0",x"3E",x"16",x"32",x"0A",x"60",x"E1",x"C9",x"3A",x"50",x"63",x"A7",
		x"C8",x"CD",x"96",x"1E",x"E1",x"C9",x"3A",x"45",x"63",x"EF",x"A0",x"1E",x"09",x"1F",x"23",x"1F",
		x"3A",x"52",x"63",x"FE",x"65",x"21",x"B8",x"69",x"CA",x"B4",x"1E",x"21",x"D0",x"69",x"DA",x"B4",
		x"1E",x"21",x"80",x"69",x"DD",x"2A",x"51",x"63",x"16",x"00",x"3A",x"53",x"63",x"5F",x"01",x"04",
		x"00",x"3A",x"54",x"63",x"A7",x"CA",x"CF",x"1E",x"09",x"DD",x"19",x"3D",x"C2",x"C8",x"1E",x"DD",
		x"36",x"00",x"00",x"DD",x"7E",x"15",x"A7",x"3E",x"02",x"CA",x"DE",x"1E",x"3E",x"04",x"32",x"42",
		x"63",x"01",x"2C",x"6A",x"7E",x"36",x"00",x"02",x"0C",x"2C",x"3E",x"60",x"02",x"0C",x"2C",x"3E",
		x"0C",x"02",x"0C",x"2C",x"7E",x"02",x"21",x"45",x"63",x"34",x"2C",x"36",x"06",x"2C",x"36",x"05",
		x"21",x"8A",x"60",x"36",x"06",x"2C",x"36",x"03",x"C9",x"21",x"46",x"63",x"35",x"C0",x"36",x"06",
		x"2C",x"35",x"CA",x"1D",x"1F",x"21",x"2D",x"6A",x"7E",x"EE",x"01",x"77",x"C9",x"36",x"04",x"2D",
		x"2D",x"34",x"C9",x"21",x"46",x"63",x"35",x"C0",x"36",x"0C",x"2C",x"35",x"CA",x"34",x"1F",x"21",
		x"2D",x"6A",x"34",x"C9",x"2D",x"2D",x"AF",x"77",x"32",x"50",x"63",x"3C",x"32",x"40",x"63",x"21",
		x"2C",x"6A",x"22",x"43",x"63",x"C9",x"3A",x"21",x"62",x"A7",x"C8",x"AF",x"32",x"04",x"62",x"32",
		x"06",x"62",x"32",x"21",x"62",x"32",x"10",x"62",x"32",x"11",x"62",x"32",x"12",x"62",x"32",x"13",
		x"62",x"32",x"14",x"62",x"3C",x"32",x"16",x"62",x"32",x"1F",x"62",x"3A",x"05",x"62",x"32",x"0E",
		x"62",x"C9",x"3A",x"27",x"62",x"3D",x"C0",x"DD",x"21",x"00",x"67",x"21",x"80",x"69",x"11",x"20",
		x"00",x"06",x"0A",x"DD",x"7E",x"00",x"3D",x"CA",x"93",x"1F",x"2C",x"2C",x"2C",x"2C",x"DD",x"19",
		x"10",x"F1",x"C9",x"DD",x"7E",x"01",x"3D",x"CA",x"EC",x"20",x"DD",x"7E",x"02",x"1F",x"DA",x"AC",
		x"1F",x"1F",x"DA",x"E5",x"1F",x"1F",x"DA",x"EF",x"1F",x"C3",x"53",x"20",x"D9",x"DD",x"34",x"05",
		x"DD",x"7E",x"17",x"DD",x"BE",x"05",x"C2",x"CE",x"1F",x"DD",x"7E",x"15",x"07",x"07",x"C6",x"15",
		x"DD",x"77",x"07",x"DD",x"7E",x"02",x"EE",x"07",x"DD",x"77",x"02",x"C3",x"BA",x"21",x"DD",x"7E",
		x"0F",x"3D",x"C2",x"DF",x"1F",x"DD",x"7E",x"07",x"EE",x"01",x"DD",x"77",x"07",x"3E",x"04",x"DD",
		x"77",x"0F",x"C3",x"BA",x"21",x"D9",x"01",x"00",x"01",x"DD",x"34",x"03",x"C3",x"F6",x"1F",x"D9",
		x"01",x"04",x"FF",x"DD",x"35",x"03",x"DD",x"66",x"03",x"DD",x"6E",x"05",x"7C",x"E6",x"07",x"FE",
		x"03",x"CA",x"5F",x"21",x"2D",x"2D",x"2D",x"CD",x"33",x"23",x"2C",x"2C",x"2C",x"7D",x"DD",x"77",
		x"05",x"CD",x"DE",x"23",x"CD",x"B4",x"24",x"DD",x"7E",x"03",x"FE",x"1C",x"DA",x"2F",x"20",x"FE",
		x"E4",x"DA",x"BA",x"21",x"AF",x"DD",x"77",x"10",x"DD",x"36",x"11",x"60",x"C3",x"38",x"20",x"AF",
		x"DD",x"36",x"10",x"FF",x"DD",x"36",x"11",x"A0",x"DD",x"36",x"12",x"FF",x"DD",x"36",x"13",x"F0",
		x"DD",x"77",x"14",x"DD",x"77",x"0E",x"DD",x"77",x"04",x"DD",x"77",x"06",x"DD",x"36",x"02",x"08",
		x"C3",x"BA",x"21",x"D9",x"CD",x"9C",x"23",x"CD",x"2F",x"2A",x"A7",x"C2",x"83",x"20",x"DD",x"7E",
		x"03",x"C6",x"08",x"FE",x"10",x"DA",x"79",x"20",x"CD",x"B4",x"24",x"DD",x"7E",x"10",x"E6",x"01",
		x"07",x"07",x"4F",x"CD",x"DE",x"23",x"C3",x"BA",x"21",x"AF",x"DD",x"77",x"00",x"DD",x"77",x"03",
		x"C3",x"BA",x"21",x"DD",x"34",x"0E",x"DD",x"7E",x"0E",x"3D",x"CA",x"A2",x"20",x"3D",x"CA",x"C3",
		x"20",x"DD",x"7E",x"10",x"3D",x"3E",x"04",x"C2",x"9C",x"20",x"3E",x"02",x"DD",x"77",x"02",x"C3",
		x"BA",x"21",x"DD",x"7E",x"15",x"A7",x"C2",x"B5",x"20",x"21",x"05",x"62",x"DD",x"7E",x"05",x"D6",
		x"16",x"BE",x"D2",x"C3",x"20",x"DD",x"7E",x"10",x"A7",x"C2",x"E1",x"20",x"DD",x"77",x"11",x"DD",
		x"36",x"10",x"FF",x"CD",x"07",x"24",x"CB",x"3C",x"CB",x"1D",x"CB",x"3C",x"CB",x"1D",x"DD",x"74",
		x"12",x"DD",x"75",x"13",x"AF",x"DD",x"77",x"14",x"DD",x"77",x"04",x"DD",x"77",x"06",x"C3",x"BA",
		x"21",x"DD",x"36",x"10",x"01",x"DD",x"36",x"11",x"00",x"C3",x"C3",x"20",x"D9",x"CD",x"9C",x"23",
		x"7C",x"D6",x"1A",x"DD",x"46",x"19",x"B8",x"DA",x"04",x"21",x"CD",x"2F",x"2A",x"A7",x"C2",x"18",
		x"21",x"CD",x"B4",x"24",x"DD",x"7E",x"03",x"C6",x"08",x"FE",x"10",x"D2",x"CE",x"1F",x"AF",x"DD",
		x"77",x"00",x"DD",x"77",x"03",x"C3",x"BA",x"21",x"DD",x"7E",x"05",x"FE",x"E0",x"DA",x"46",x"21",
		x"DD",x"7E",x"07",x"E6",x"FC",x"F6",x"01",x"DD",x"77",x"07",x"AF",x"DD",x"77",x"01",x"DD",x"77",
		x"02",x"DD",x"36",x"10",x"FF",x"DD",x"77",x"11",x"DD",x"77",x"12",x"DD",x"36",x"13",x"B0",x"DD",
		x"36",x"0E",x"01",x"C3",x"53",x"21",x"CD",x"07",x"24",x"CD",x"CB",x"22",x"DD",x"7E",x"05",x"DD",
		x"77",x"19",x"AF",x"DD",x"77",x"14",x"DD",x"77",x"04",x"DD",x"77",x"06",x"C3",x"BA",x"21",x"7D",
		x"C6",x"05",x"57",x"7C",x"01",x"15",x"00",x"CD",x"6D",x"21",x"C3",x"BA",x"21",x"CD",x"6E",x"23",
		x"3D",x"C0",x"78",x"D6",x"05",x"DD",x"77",x"17",x"3A",x"48",x"63",x"A7",x"CA",x"B2",x"21",x"3A",
		x"05",x"62",x"D6",x"04",x"BA",x"D8",x"3A",x"80",x"63",x"1F",x"3C",x"47",x"3A",x"18",x"60",x"4F",
		x"E6",x"03",x"B8",x"D0",x"21",x"10",x"60",x"3A",x"03",x"62",x"BB",x"CA",x"B2",x"21",x"D2",x"A9",
		x"21",x"CB",x"46",x"CA",x"AE",x"21",x"C3",x"B2",x"21",x"CB",x"4E",x"C2",x"B2",x"21",x"79",x"E6",
		x"18",x"C0",x"DD",x"34",x"07",x"DD",x"CB",x"02",x"C6",x"C9",x"D9",x"DD",x"7E",x"03",x"77",x"2C",
		x"DD",x"7E",x"07",x"77",x"2C",x"DD",x"7E",x"08",x"77",x"2C",x"DD",x"7E",x"05",x"77",x"C3",x"8D",
		x"1F",x"80",x"FE",x"01",x"C0",x"04",x"50",x"02",x"10",x"82",x"60",x"02",x"10",x"82",x"CA",x"01",
		x"10",x"81",x"FF",x"02",x"38",x"01",x"80",x"02",x"FF",x"04",x"80",x"04",x"60",x"80",x"11",x"D1",
		x"21",x"21",x"CC",x"63",x"7E",x"07",x"83",x"5F",x"1A",x"32",x"10",x"60",x"2C",x"7E",x"35",x"A7",
		x"C0",x"1C",x"1A",x"77",x"2D",x"34",x"C9",x"3E",x"02",x"F7",x"3A",x"1A",x"60",x"1F",x"21",x"80",
		x"62",x"7E",x"DA",x"19",x"22",x"21",x"88",x"62",x"7E",x"E5",x"EF",x"27",x"22",x"59",x"22",x"99",
		x"22",x"A2",x"22",x"00",x"00",x"00",x"00",x"E1",x"2C",x"35",x"C2",x"3A",x"22",x"2D",x"34",x"2C",
		x"2C",x"CD",x"43",x"22",x"3E",x"01",x"32",x"1A",x"62",x"C9",x"2C",x"CD",x"43",x"22",x"AF",x"32",
		x"1A",x"62",x"C9",x"3A",x"05",x"62",x"FE",x"7A",x"D2",x"57",x"22",x"3A",x"16",x"62",x"A7",x"C2",
		x"57",x"22",x"3A",x"03",x"62",x"BE",x"C8",x"E1",x"C9",x"E1",x"2C",x"2C",x"2C",x"2C",x"35",x"C0",
		x"3E",x"04",x"77",x"2D",x"34",x"CD",x"BD",x"22",x"3E",x"78",x"BE",x"C2",x"75",x"22",x"2D",x"2D",
		x"2D",x"34",x"2C",x"2C",x"2C",x"2D",x"CD",x"43",x"22",x"3A",x"05",x"62",x"FE",x"68",x"D2",x"8A",
		x"22",x"21",x"05",x"62",x"34",x"CD",x"C0",x"3F",x"34",x"C9",x"1F",x"DA",x"81",x"22",x"1F",x"3E",
		x"01",x"DA",x"95",x"22",x"AF",x"32",x"22",x"62",x"C9",x"E1",x"3A",x"18",x"60",x"E6",x"3C",x"C0",
		x"34",x"C9",x"E1",x"2C",x"2C",x"2C",x"2C",x"35",x"C0",x"36",x"02",x"2D",x"35",x"CD",x"BD",x"22",
		x"3E",x"68",x"BE",x"C0",x"AF",x"06",x"80",x"2D",x"2D",x"70",x"2D",x"77",x"C9",x"7E",x"CB",x"5D",
		x"11",x"4B",x"69",x"C2",x"C9",x"22",x"11",x"47",x"69",x"12",x"C9",x"3A",x"48",x"63",x"A7",x"CA",
		x"E1",x"22",x"3A",x"80",x"63",x"3D",x"EF",x"F6",x"22",x"F6",x"22",x"03",x"23",x"03",x"23",x"1A",
		x"23",x"3A",x"29",x"62",x"47",x"05",x"3E",x"01",x"CA",x"F9",x"22",x"05",x"3E",x"B1",x"CA",x"F9",
		x"22",x"3E",x"E9",x"C3",x"F9",x"22",x"3A",x"18",x"60",x"DD",x"77",x"11",x"E6",x"01",x"3D",x"DD",
		x"77",x"10",x"C9",x"3A",x"18",x"60",x"DD",x"77",x"11",x"3A",x"03",x"62",x"DD",x"BE",x"03",x"3E",
		x"01",x"D2",x"16",x"23",x"3D",x"3D",x"DD",x"77",x"10",x"C9",x"3A",x"03",x"62",x"DD",x"96",x"03",
		x"0E",x"FF",x"DA",x"26",x"23",x"0C",x"07",x"CB",x"11",x"07",x"CB",x"11",x"DD",x"71",x"10",x"DD",
		x"77",x"11",x"C9",x"3E",x"0F",x"A4",x"05",x"CA",x"42",x"23",x"FE",x"0F",x"D8",x"06",x"FF",x"C3",
		x"47",x"23",x"FE",x"01",x"D0",x"06",x"01",x"3E",x"F0",x"BD",x"CA",x"60",x"23",x"3E",x"4C",x"BD",
		x"CA",x"66",x"23",x"7D",x"CB",x"6F",x"CA",x"5C",x"23",x"90",x"6F",x"C9",x"80",x"C3",x"5A",x"23",
		x"CB",x"7C",x"C2",x"59",x"23",x"C9",x"7C",x"FE",x"98",x"D8",x"7D",x"C3",x"5C",x"23",x"21",x"00",
		x"63",x"ED",x"B1",x"C2",x"9A",x"23",x"E5",x"C5",x"01",x"14",x"00",x"09",x"0C",x"5F",x"7A",x"BE",
		x"CA",x"8F",x"23",x"09",x"BE",x"CA",x"95",x"23",x"57",x"7B",x"C1",x"E1",x"C3",x"71",x"23",x"09",
		x"3E",x"01",x"C3",x"98",x"23",x"AF",x"ED",x"42",x"C1",x"46",x"E1",x"C9",x"DD",x"7E",x"04",x"DD",
		x"86",x"11",x"DD",x"77",x"04",x"DD",x"7E",x"03",x"DD",x"8E",x"10",x"DD",x"77",x"03",x"DD",x"7E",
		x"06",x"DD",x"96",x"13",x"6F",x"DD",x"7E",x"05",x"DD",x"9E",x"12",x"67",x"DD",x"7E",x"14",x"A7",
		x"17",x"3C",x"06",x"00",x"CB",x"10",x"CB",x"27",x"CB",x"10",x"CB",x"27",x"CB",x"10",x"CB",x"27",
		x"CB",x"10",x"4F",x"09",x"DD",x"74",x"05",x"DD",x"75",x"06",x"DD",x"34",x"14",x"C9",x"DD",x"7E",
		x"0F",x"3D",x"C2",x"03",x"24",x"AF",x"DD",x"CB",x"07",x"26",x"17",x"DD",x"CB",x"08",x"26",x"17",
		x"47",x"3E",x"03",x"B1",x"CD",x"09",x"30",x"1F",x"DD",x"CB",x"08",x"1E",x"1F",x"DD",x"CB",x"07",
		x"1E",x"3E",x"04",x"DD",x"77",x"0F",x"C9",x"DD",x"7E",x"14",x"07",x"07",x"07",x"07",x"4F",x"E6",
		x"0F",x"67",x"79",x"E6",x"F0",x"6F",x"DD",x"4E",x"13",x"DD",x"46",x"12",x"ED",x"42",x"C9",x"11",
		x"00",x"01",x"3A",x"03",x"62",x"FE",x"16",x"D8",x"15",x"1C",x"FE",x"EA",x"D0",x"1D",x"3A",x"27",
		x"62",x"0F",x"D0",x"3A",x"05",x"62",x"FE",x"58",x"D0",x"3A",x"03",x"62",x"FE",x"6C",x"D0",x"14",
		x"C9",x"21",x"0C",x"3F",x"3E",x"5E",x"06",x"06",x"86",x"23",x"10",x"FC",x"FD",x"21",x"10",x"63",
		x"A7",x"CA",x"56",x"24",x"FD",x"23",x"3A",x"27",x"62",x"3D",x"21",x"E4",x"3A",x"CA",x"71",x"24",
		x"3D",x"21",x"5D",x"3B",x"CA",x"71",x"24",x"3D",x"21",x"E5",x"3B",x"CA",x"71",x"24",x"21",x"8B",
		x"3C",x"DD",x"21",x"00",x"63",x"11",x"05",x"00",x"7E",x"A7",x"CA",x"88",x"24",x"3D",x"CA",x"9E",
		x"24",x"FE",x"A9",x"C8",x"19",x"C3",x"78",x"24",x"23",x"7E",x"DD",x"77",x"00",x"23",x"7E",x"DD",
		x"77",x"15",x"23",x"23",x"7E",x"DD",x"77",x"2A",x"DD",x"23",x"23",x"C3",x"78",x"24",x"23",x"7E",
		x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77",x"15",x"23",x"23",x"7E",x"FD",x"77",x"2A",x"FD",x"23",
		x"23",x"C3",x"78",x"24",x"DD",x"7E",x"05",x"FE",x"E8",x"D8",x"DD",x"7E",x"03",x"FE",x"2A",x"D0",
		x"FE",x"20",x"D8",x"DD",x"7E",x"15",x"A7",x"CA",x"D0",x"24",x"3E",x"03",x"32",x"B9",x"62",x"AF",
		x"DD",x"77",x"00",x"DD",x"77",x"03",x"21",x"82",x"60",x"36",x"03",x"E1",x"3A",x"48",x"63",x"A7",
		x"C2",x"BA",x"21",x"3C",x"32",x"48",x"63",x"C3",x"BA",x"21",x"3E",x"02",x"F7",x"CD",x"23",x"25",
		x"CD",x"91",x"25",x"DD",x"21",x"A0",x"65",x"06",x"06",x"21",x"B8",x"69",x"DD",x"7E",x"00",x"A7",
		x"CA",x"1C",x"25",x"DD",x"7E",x"03",x"77",x"2C",x"DD",x"7E",x"07",x"77",x"2C",x"DD",x"7E",x"08",
		x"77",x"2C",x"DD",x"7E",x"05",x"77",x"2C",x"DD",x"19",x"10",x"E1",x"C9",x"7D",x"C6",x"04",x"6F",
		x"C3",x"17",x"25",x"21",x"9B",x"63",x"7E",x"A7",x"C2",x"8F",x"25",x"3A",x"9A",x"63",x"A7",x"C8",
		x"06",x"06",x"11",x"10",x"00",x"DD",x"21",x"A0",x"65",x"DD",x"CB",x"00",x"46",x"CA",x"45",x"25",
		x"DD",x"19",x"10",x"F5",x"C9",x"CD",x"57",x"00",x"FE",x"60",x"DD",x"36",x"05",x"7C",x"DA",x"58",
		x"25",x"3A",x"A3",x"62",x"3D",x"C2",x"6E",x"25",x"DD",x"36",x"05",x"CC",x"3A",x"A6",x"62",x"07",
		x"DD",x"36",x"03",x"07",x"D2",x"76",x"25",x"DD",x"36",x"03",x"F8",x"C3",x"76",x"25",x"CD",x"57",
		x"00",x"FE",x"68",x"C3",x"60",x"25",x"DD",x"36",x"00",x"01",x"DD",x"36",x"07",x"4B",x"DD",x"36",
		x"09",x"08",x"DD",x"36",x"0A",x"03",x"3E",x"7C",x"32",x"9B",x"63",x"AF",x"32",x"9A",x"63",x"35",
		x"C9",x"DD",x"21",x"A0",x"65",x"11",x"10",x"00",x"06",x"06",x"DD",x"CB",x"00",x"46",x"CA",x"BB",
		x"25",x"DD",x"7E",x"03",x"67",x"C6",x"07",x"FE",x"0E",x"DA",x"D6",x"25",x"DD",x"7E",x"05",x"FE",
		x"7C",x"CA",x"C0",x"25",x"3A",x"A6",x"63",x"84",x"DD",x"77",x"03",x"DD",x"19",x"10",x"DB",x"C9",
		x"7C",x"FE",x"80",x"CA",x"D6",x"25",x"3A",x"A5",x"63",x"D2",x"CF",x"25",x"3A",x"A4",x"63",x"84",
		x"DD",x"77",x"03",x"C3",x"BB",x"25",x"21",x"B8",x"69",x"3E",x"06",x"90",x"CA",x"E7",x"25",x"2C",
		x"2C",x"2C",x"2C",x"3D",x"C3",x"DC",x"25",x"AF",x"DD",x"77",x"00",x"DD",x"77",x"03",x"77",x"C3",
		x"BB",x"25",x"3E",x"02",x"F7",x"CD",x"02",x"26",x"CD",x"2F",x"26",x"CD",x"79",x"26",x"CD",x"D3",
		x"2A",x"C9",x"3A",x"1A",x"60",x"0F",x"DA",x"16",x"26",x"21",x"A0",x"62",x"35",x"C2",x"16",x"26",
		x"36",x"80",x"2C",x"CD",x"DE",x"26",x"21",x"A1",x"62",x"CD",x"E9",x"26",x"32",x"A3",x"63",x"3A",
		x"1A",x"60",x"E6",x"1F",x"FE",x"01",x"C0",x"11",x"E4",x"69",x"EB",x"CD",x"A6",x"26",x"C9",x"21",
		x"A3",x"62",x"3A",x"05",x"62",x"FE",x"C0",x"DA",x"6F",x"26",x"3A",x"1A",x"60",x"0F",x"DA",x"4C",
		x"26",x"2D",x"35",x"C2",x"4C",x"26",x"36",x"C0",x"2C",x"CD",x"DE",x"26",x"21",x"A3",x"62",x"CD",
		x"E9",x"26",x"32",x"A5",x"63",x"ED",x"44",x"32",x"A4",x"63",x"3A",x"1A",x"60",x"E6",x"1F",x"C0",
		x"2D",x"11",x"EC",x"69",x"EB",x"CD",x"A6",x"26",x"E6",x"7F",x"21",x"ED",x"69",x"77",x"C9",x"CB",
		x"7E",x"C2",x"4C",x"26",x"36",x"FF",x"C3",x"4C",x"26",x"3A",x"1A",x"60",x"0F",x"DA",x"8D",x"26",
		x"21",x"A5",x"62",x"35",x"C2",x"8D",x"26",x"36",x"FF",x"2C",x"CD",x"DE",x"26",x"21",x"A6",x"62",
		x"CD",x"E9",x"26",x"32",x"A6",x"63",x"3A",x"1A",x"60",x"E6",x"1F",x"FE",x"02",x"C0",x"11",x"F4",
		x"69",x"EB",x"CD",x"A6",x"26",x"C9",x"2C",x"1A",x"17",x"DA",x"C5",x"26",x"7E",x"3C",x"FE",x"53",
		x"C2",x"B5",x"26",x"3E",x"50",x"77",x"7D",x"C6",x"04",x"6F",x"7E",x"3D",x"FE",x"CF",x"C2",x"C3",
		x"26",x"3E",x"D2",x"77",x"C9",x"7E",x"3D",x"FE",x"4F",x"C2",x"CE",x"26",x"3E",x"52",x"77",x"7D",
		x"C6",x"04",x"6F",x"7E",x"3C",x"FE",x"D3",x"C2",x"DC",x"26",x"3E",x"D0",x"77",x"C9",x"CB",x"7E",
		x"CA",x"E6",x"26",x"36",x"02",x"C9",x"36",x"FE",x"C9",x"3A",x"1A",x"60",x"E6",x"01",x"C8",x"CB",
		x"7E",x"3E",x"FF",x"C2",x"F8",x"26",x"3E",x"01",x"77",x"C9",x"3E",x"04",x"F7",x"3A",x"05",x"62",
		x"FE",x"F0",x"D2",x"7F",x"27",x"3A",x"29",x"62",x"3D",x"3A",x"1A",x"60",x"C2",x"1A",x"27",x"E6",
		x"03",x"FE",x"01",x"CA",x"1E",x"27",x"DA",x"22",x"27",x"C9",x"0F",x"DA",x"22",x"27",x"CD",x"45",
		x"27",x"C9",x"CD",x"97",x"27",x"CD",x"DA",x"27",x"06",x"06",x"11",x"10",x"00",x"21",x"58",x"69",
		x"DD",x"21",x"00",x"66",x"DD",x"7E",x"03",x"77",x"2C",x"2C",x"2C",x"DD",x"7E",x"05",x"77",x"2C",
		x"DD",x"19",x"10",x"F0",x"C9",x"3A",x"98",x"63",x"A7",x"C8",x"3A",x"16",x"62",x"A7",x"C0",x"3A",
		x"03",x"62",x"FE",x"2C",x"DA",x"66",x"27",x"FE",x"43",x"DA",x"6F",x"27",x"FE",x"6C",x"DA",x"66",
		x"27",x"FE",x"83",x"DA",x"87",x"27",x"AF",x"32",x"98",x"63",x"3C",x"32",x"21",x"62",x"C9",x"3A",
		x"05",x"62",x"FE",x"71",x"DA",x"7F",x"27",x"3D",x"32",x"05",x"62",x"32",x"4F",x"69",x"C9",x"AF",
		x"32",x"00",x"62",x"32",x"98",x"63",x"C9",x"3A",x"05",x"62",x"FE",x"E8",x"D2",x"7F",x"27",x"3C",
		x"32",x"05",x"62",x"32",x"4F",x"69",x"C9",x"06",x"06",x"11",x"10",x"00",x"DD",x"21",x"00",x"66",
		x"DD",x"CB",x"00",x"46",x"CA",x"C2",x"27",x"DD",x"CB",x"0D",x"5E",x"CA",x"C7",x"27",x"DD",x"7E",
		x"05",x"3D",x"DD",x"77",x"05",x"FE",x"60",x"C2",x"C2",x"27",x"DD",x"36",x"03",x"77",x"DD",x"36",
		x"0D",x"04",x"DD",x"19",x"10",x"DA",x"C9",x"DD",x"7E",x"05",x"3C",x"DD",x"77",x"05",x"FE",x"F8",
		x"C2",x"C2",x"27",x"DD",x"36",x"00",x"00",x"C3",x"C2",x"27",x"21",x"A7",x"62",x"7E",x"A7",x"C2",
		x"06",x"28",x"06",x"06",x"DD",x"21",x"00",x"66",x"DD",x"CB",x"00",x"46",x"CA",x"F4",x"27",x"DD",
		x"19",x"10",x"F5",x"C9",x"DD",x"36",x"00",x"01",x"DD",x"36",x"03",x"37",x"DD",x"36",x"05",x"F8",
		x"DD",x"36",x"0D",x"08",x"36",x"34",x"35",x"C9",x"FD",x"21",x"00",x"62",x"3A",x"05",x"62",x"4F",
		x"21",x"07",x"04",x"CD",x"6F",x"28",x"A7",x"C8",x"3D",x"32",x"00",x"62",x"C9",x"06",x"02",x"11",
		x"10",x"00",x"FD",x"21",x"80",x"66",x"FD",x"CB",x"01",x"46",x"C2",x"32",x"28",x"FD",x"19",x"10",
		x"F5",x"C9",x"FD",x"4E",x"05",x"FD",x"66",x"09",x"FD",x"6E",x"0A",x"CD",x"6F",x"28",x"A7",x"C8",
		x"32",x"50",x"63",x"3A",x"B9",x"63",x"90",x"32",x"54",x"63",x"7B",x"32",x"53",x"63",x"DD",x"22",
		x"51",x"63",x"C9",x"FD",x"21",x"00",x"62",x"3A",x"05",x"62",x"C6",x"0C",x"4F",x"3A",x"10",x"60",
		x"E6",x"03",x"21",x"08",x"05",x"CA",x"6B",x"28",x"21",x"08",x"13",x"CD",x"88",x"3E",x"C9",x"3A",
		x"27",x"62",x"E5",x"EF",x"00",x"00",x"80",x"28",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",
		x"E1",x"06",x"0A",x"78",x"32",x"B9",x"63",x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"13",
		x"29",x"06",x"05",x"78",x"32",x"B9",x"63",x"1E",x"20",x"DD",x"21",x"00",x"64",x"CD",x"13",x"29",
		x"06",x"01",x"78",x"32",x"B9",x"63",x"1E",x"00",x"DD",x"21",x"A0",x"66",x"CD",x"13",x"29",x"C9",
		x"E1",x"06",x"05",x"78",x"32",x"B9",x"63",x"11",x"20",x"00",x"DD",x"21",x"00",x"64",x"CD",x"13",
		x"29",x"06",x"06",x"78",x"32",x"B9",x"63",x"1E",x"10",x"DD",x"21",x"A0",x"65",x"CD",x"13",x"29",
		x"06",x"01",x"78",x"32",x"B9",x"63",x"1E",x"00",x"DD",x"21",x"A0",x"66",x"CD",x"13",x"29",x"C9",
		x"E1",x"06",x"05",x"78",x"32",x"B9",x"63",x"11",x"20",x"00",x"DD",x"21",x"00",x"64",x"CD",x"13",
		x"29",x"06",x"0A",x"78",x"32",x"B9",x"63",x"1E",x"10",x"DD",x"21",x"00",x"65",x"CD",x"13",x"29",
		x"C9",x"E1",x"06",x"07",x"78",x"32",x"B9",x"63",x"11",x"20",x"00",x"DD",x"21",x"00",x"64",x"CD",
		x"13",x"29",x"C9",x"DD",x"E5",x"DD",x"CB",x"00",x"46",x"CA",x"4C",x"29",x"79",x"DD",x"96",x"05",
		x"D2",x"25",x"29",x"ED",x"44",x"3C",x"95",x"DA",x"30",x"29",x"DD",x"96",x"0A",x"D2",x"4C",x"29",
		x"FD",x"7E",x"03",x"DD",x"96",x"03",x"D2",x"3B",x"29",x"ED",x"44",x"94",x"DA",x"45",x"29",x"DD",
		x"96",x"09",x"D2",x"4C",x"29",x"3E",x"01",x"DD",x"E1",x"33",x"33",x"C9",x"DD",x"19",x"10",x"C5",
		x"AF",x"DD",x"E1",x"C9",x"3E",x"0B",x"F7",x"CD",x"74",x"29",x"32",x"18",x"62",x"0F",x"0F",x"32",
		x"85",x"60",x"78",x"A7",x"C8",x"FE",x"01",x"CA",x"6F",x"29",x"DD",x"36",x"01",x"01",x"C9",x"DD",
		x"36",x"11",x"01",x"C9",x"FD",x"21",x"00",x"62",x"3A",x"05",x"62",x"4F",x"21",x"08",x"04",x"06",
		x"02",x"11",x"10",x"00",x"DD",x"21",x"80",x"66",x"CD",x"13",x"29",x"C9",x"2A",x"C8",x"63",x"7D",
		x"C6",x"0E",x"6F",x"56",x"2C",x"7E",x"C6",x"0C",x"5F",x"EB",x"CD",x"F0",x"2F",x"7E",x"FE",x"B0",
		x"DA",x"AC",x"29",x"E6",x"0F",x"FE",x"08",x"D2",x"AC",x"29",x"AF",x"C9",x"3E",x"01",x"C9",x"3E",
		x"04",x"F7",x"FD",x"21",x"00",x"62",x"3A",x"05",x"62",x"4F",x"21",x"08",x"04",x"CD",x"22",x"2A",
		x"A7",x"CA",x"20",x"2A",x"3E",x"06",x"90",x"CA",x"D0",x"29",x"DD",x"19",x"3D",x"C3",x"C7",x"29",
		x"DD",x"7E",x"05",x"D6",x"04",x"57",x"3A",x"0C",x"62",x"C6",x"05",x"BA",x"D2",x"EE",x"29",x"7A",
		x"D6",x"08",x"32",x"05",x"62",x"3E",x"01",x"47",x"32",x"98",x"63",x"33",x"33",x"C9",x"3A",x"0C",
		x"62",x"D6",x"0E",x"BA",x"D2",x"1B",x"2A",x"3A",x"10",x"62",x"A7",x"3A",x"03",x"62",x"CA",x"08",
		x"2A",x"F6",x"07",x"D6",x"04",x"C3",x"0E",x"2A",x"D6",x"08",x"F6",x"07",x"C6",x"04",x"32",x"03",
		x"62",x"32",x"4C",x"69",x"3E",x"01",x"06",x"00",x"33",x"33",x"C9",x"AF",x"32",x"00",x"62",x"C9",
		x"47",x"C9",x"06",x"06",x"11",x"10",x"00",x"DD",x"21",x"00",x"66",x"CD",x"13",x"29",x"C9",x"DD",
		x"7E",x"03",x"67",x"DD",x"7E",x"05",x"C6",x"04",x"6F",x"E5",x"CD",x"F0",x"2F",x"D1",x"7E",x"FE",
		x"B0",x"DA",x"7B",x"2A",x"E6",x"0F",x"FE",x"08",x"D2",x"7B",x"2A",x"7E",x"FE",x"C0",x"CA",x"7B",
		x"2A",x"DA",x"69",x"2A",x"FE",x"D0",x"DA",x"6E",x"2A",x"FE",x"E0",x"DA",x"63",x"2A",x"FE",x"F0",
		x"DA",x"6E",x"2A",x"E6",x"0F",x"3D",x"C3",x"72",x"2A",x"3E",x"FF",x"C3",x"72",x"2A",x"E6",x"0F",
		x"D6",x"09",x"4F",x"7B",x"E6",x"F8",x"81",x"BB",x"DA",x"7D",x"2A",x"AF",x"C9",x"D6",x"04",x"DD",
		x"77",x"05",x"3E",x"01",x"C9",x"3A",x"15",x"62",x"A7",x"C0",x"3A",x"16",x"62",x"A7",x"C0",x"3A",
		x"98",x"63",x"FE",x"01",x"C8",x"3A",x"03",x"62",x"D6",x"03",x"67",x"3A",x"05",x"62",x"C6",x"0C",
		x"6F",x"E5",x"CD",x"F0",x"2F",x"D1",x"7E",x"FE",x"B0",x"DA",x"B4",x"2A",x"E6",x"0F",x"FE",x"08",
		x"D2",x"B4",x"2A",x"C9",x"7A",x"E6",x"07",x"CA",x"CD",x"2A",x"01",x"20",x"00",x"ED",x"42",x"7E",
		x"FE",x"B0",x"DA",x"CD",x"2A",x"E6",x"0F",x"FE",x"08",x"D2",x"CD",x"2A",x"C9",x"3E",x"01",x"32",
		x"21",x"62",x"C9",x"3A",x"03",x"62",x"47",x"3A",x"05",x"62",x"FE",x"50",x"CA",x"EA",x"2A",x"FE",
		x"78",x"CA",x"F6",x"2A",x"FE",x"C8",x"CA",x"F0",x"2A",x"C9",x"3A",x"A3",x"63",x"C3",x"02",x"2B",
		x"3A",x"A6",x"63",x"C3",x"02",x"2B",x"78",x"FE",x"80",x"3A",x"A5",x"63",x"D2",x"02",x"2B",x"3A",
		x"A4",x"63",x"80",x"32",x"03",x"62",x"32",x"4C",x"69",x"CD",x"1F",x"24",x"21",x"03",x"62",x"1D",
		x"CA",x"18",x"2B",x"15",x"CA",x"1A",x"2B",x"C9",x"35",x"C9",x"34",x"C9",x"DD",x"21",x"00",x"62",
		x"CD",x"29",x"2B",x"CD",x"AF",x"29",x"AF",x"47",x"C9",x"3A",x"27",x"62",x"3D",x"C2",x"53",x"2B",
		x"3A",x"03",x"62",x"67",x"3A",x"05",x"62",x"C6",x"07",x"6F",x"CD",x"9B",x"2B",x"A7",x"CA",x"51",
		x"2B",x"7B",x"91",x"FE",x"04",x"D2",x"74",x"2B",x"79",x"D6",x"07",x"32",x"05",x"62",x"3E",x"01",
		x"47",x"E1",x"C9",x"3A",x"03",x"62",x"D6",x"03",x"67",x"3A",x"05",x"62",x"C6",x"07",x"6F",x"CD",
		x"9B",x"2B",x"FE",x"02",x"CA",x"7A",x"2B",x"7A",x"C6",x"07",x"67",x"6B",x"CD",x"9B",x"2B",x"A7",
		x"C8",x"C3",x"7A",x"2B",x"3E",x"00",x"06",x"00",x"E1",x"C9",x"3A",x"10",x"62",x"A7",x"3A",x"03",
		x"62",x"CA",x"8B",x"2B",x"F6",x"07",x"D6",x"04",x"C3",x"91",x"2B",x"D6",x"08",x"F6",x"07",x"C6",
		x"04",x"32",x"03",x"62",x"32",x"4C",x"69",x"3E",x"01",x"E1",x"C9",x"E5",x"CD",x"F0",x"2F",x"D1",
		x"7E",x"FE",x"B0",x"DA",x"D9",x"2B",x"E6",x"0F",x"FE",x"08",x"D2",x"D9",x"2B",x"7E",x"FE",x"C0",
		x"CA",x"D9",x"2B",x"DA",x"DC",x"2B",x"FE",x"D0",x"DA",x"CB",x"2B",x"FE",x"E0",x"DA",x"C5",x"2B",
		x"FE",x"F0",x"DA",x"CB",x"2B",x"E6",x"0F",x"3D",x"C3",x"CF",x"2B",x"E6",x"0F",x"D6",x"09",x"4F",
		x"7B",x"E6",x"F8",x"81",x"4F",x"BB",x"DA",x"E1",x"2B",x"AF",x"47",x"C9",x"7B",x"E6",x"F8",x"3D",
		x"4F",x"3A",x"0C",x"62",x"DD",x"96",x"05",x"83",x"B9",x"CA",x"EF",x"2B",x"D2",x"F8",x"2B",x"79",
		x"D6",x"07",x"32",x"05",x"62",x"C3",x"FD",x"2B",x"3E",x"02",x"06",x"00",x"C9",x"3E",x"01",x"47",
		x"E1",x"E1",x"C9",x"3E",x"01",x"F7",x"D7",x"3A",x"93",x"63",x"0F",x"D8",x"3A",x"B1",x"62",x"A7",
		x"C8",x"4F",x"3A",x"B0",x"62",x"D6",x"02",x"B9",x"DA",x"7B",x"2C",x"3A",x"82",x"63",x"CB",x"4F",
		x"C2",x"86",x"2C",x"3A",x"80",x"63",x"47",x"3A",x"1A",x"60",x"E6",x"1F",x"B8",x"CA",x"33",x"2C",
		x"10",x"FA",x"C9",x"3A",x"B0",x"62",x"CB",x"3F",x"B9",x"DA",x"41",x"2C",x"3A",x"19",x"60",x"0F",
		x"D0",x"CD",x"57",x"00",x"E6",x"0F",x"C2",x"86",x"2C",x"3E",x"01",x"32",x"82",x"63",x"3C",x"32",
		x"8F",x"63",x"3E",x"01",x"32",x"92",x"63",x"3A",x"B2",x"62",x"B9",x"C0",x"D6",x"08",x"32",x"B2",
		x"62",x"11",x"20",x"00",x"21",x"00",x"64",x"06",x"05",x"7E",x"A7",x"CA",x"72",x"2C",x"19",x"10",
		x"F8",x"C9",x"3A",x"82",x"63",x"F6",x"80",x"32",x"82",x"63",x"C9",x"C6",x"02",x"B9",x"CA",x"49",
		x"2C",x"3E",x"02",x"C3",x"4B",x"2C",x"AF",x"32",x"82",x"63",x"3E",x"03",x"C3",x"4F",x"2C",x"3E",
		x"01",x"F7",x"D7",x"3A",x"93",x"63",x"0F",x"DA",x"15",x"2D",x"3A",x"92",x"63",x"0F",x"D0",x"DD",
		x"21",x"00",x"67",x"11",x"20",x"00",x"06",x"0A",x"DD",x"7E",x"00",x"0F",x"DA",x"B3",x"2C",x"0F",
		x"D2",x"B8",x"2C",x"DD",x"19",x"10",x"F1",x"C9",x"DD",x"22",x"AA",x"62",x"DD",x"36",x"00",x"02",
		x"16",x"00",x"3E",x"0A",x"90",x"87",x"87",x"5F",x"21",x"80",x"69",x"19",x"22",x"AC",x"62",x"3E",
		x"01",x"32",x"93",x"63",x"11",x"01",x"05",x"CD",x"9F",x"30",x"21",x"B1",x"62",x"35",x"C2",x"E6",
		x"2C",x"3E",x"01",x"32",x"86",x"63",x"7E",x"FE",x"04",x"D2",x"F6",x"2C",x"21",x"A8",x"69",x"87",
		x"87",x"5F",x"16",x"00",x"19",x"72",x"DD",x"36",x"07",x"15",x"DD",x"36",x"08",x"0B",x"DD",x"36",
		x"15",x"00",x"3A",x"82",x"63",x"07",x"D2",x"15",x"2D",x"DD",x"36",x"07",x"19",x"DD",x"36",x"08",
		x"0C",x"DD",x"36",x"15",x"01",x"21",x"AF",x"62",x"35",x"C0",x"36",x"18",x"3A",x"8F",x"63",x"A7",
		x"CA",x"51",x"2D",x"4F",x"21",x"32",x"39",x"3A",x"82",x"63",x"0F",x"DA",x"2F",x"2D",x"0D",x"79",
		x"87",x"87",x"87",x"4F",x"87",x"87",x"81",x"5F",x"16",x"00",x"19",x"CD",x"4E",x"00",x"21",x"8F",
		x"63",x"35",x"C2",x"51",x"2D",x"3E",x"01",x"32",x"AF",x"62",x"3A",x"82",x"63",x"0F",x"DA",x"83",
		x"2D",x"2A",x"A8",x"62",x"7E",x"DD",x"2A",x"AA",x"62",x"ED",x"5B",x"AC",x"62",x"FE",x"7F",x"CA",
		x"8C",x"2D",x"4F",x"E6",x"7F",x"12",x"DD",x"7E",x"07",x"CB",x"79",x"CA",x"70",x"2D",x"EE",x"03",
		x"13",x"12",x"DD",x"77",x"07",x"DD",x"7E",x"08",x"13",x"12",x"23",x"7E",x"13",x"12",x"23",x"22",
		x"A8",x"62",x"C9",x"21",x"CC",x"39",x"22",x"A8",x"62",x"C3",x"54",x"2D",x"21",x"C3",x"39",x"22",
		x"A8",x"62",x"DD",x"36",x"01",x"01",x"3A",x"82",x"63",x"0F",x"DA",x"A5",x"2D",x"DD",x"36",x"01",
		x"00",x"DD",x"36",x"02",x"02",x"DD",x"36",x"00",x"01",x"DD",x"36",x"0F",x"01",x"AF",x"DD",x"77",
		x"10",x"DD",x"77",x"11",x"DD",x"77",x"12",x"DD",x"77",x"13",x"DD",x"77",x"14",x"32",x"93",x"63",
		x"32",x"92",x"63",x"1A",x"DD",x"77",x"03",x"13",x"13",x"13",x"1A",x"DD",x"77",x"05",x"21",x"5C",
		x"38",x"CD",x"4E",x"00",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"C9",x"3E",x"0A",x"F7",x"D7",x"3A",
		x"80",x"63",x"3C",x"A7",x"1F",x"47",x"3A",x"27",x"62",x"FE",x"02",x"20",x"01",x"04",x"3E",x"FE",
		x"37",x"1F",x"A7",x"10",x"FC",x"47",x"3A",x"1A",x"60",x"A0",x"C0",x"3E",x"01",x"32",x"A0",x"63",
		x"32",x"9A",x"63",x"C9",x"3E",x"04",x"F7",x"D7",x"DD",x"21",x"00",x"65",x"FD",x"21",x"80",x"69",
		x"06",x"0A",x"DD",x"7E",x"00",x"0F",x"D2",x"A7",x"2E",x"3A",x"1A",x"60",x"E6",x"0F",x"C2",x"29",
		x"2E",x"FD",x"7E",x"01",x"EE",x"07",x"FD",x"77",x"01",x"DD",x"7E",x"0D",x"FE",x"04",x"CA",x"84",
		x"2E",x"DD",x"34",x"03",x"DD",x"34",x"03",x"DD",x"6E",x"0E",x"DD",x"66",x"0F",x"7E",x"4F",x"FE",
		x"7F",x"CA",x"9C",x"2E",x"23",x"DD",x"86",x"05",x"DD",x"77",x"05",x"DD",x"75",x"0E",x"DD",x"74",
		x"0F",x"DD",x"7E",x"03",x"FE",x"B7",x"DA",x"6C",x"2E",x"79",x"FE",x"7F",x"C2",x"6C",x"2E",x"DD",
		x"36",x"0D",x"04",x"AF",x"32",x"83",x"60",x"3E",x"03",x"32",x"84",x"60",x"DD",x"7E",x"03",x"FD",
		x"77",x"00",x"DD",x"7E",x"05",x"FD",x"77",x"03",x"11",x"10",x"00",x"DD",x"19",x"1E",x"04",x"FD",
		x"19",x"10",x"8F",x"C9",x"3E",x"03",x"DD",x"86",x"05",x"DD",x"77",x"05",x"FE",x"F8",x"DA",x"6C",
		x"2E",x"DD",x"36",x"03",x"00",x"DD",x"36",x"00",x"00",x"C3",x"6C",x"2E",x"21",x"AA",x"39",x"3E",
		x"03",x"32",x"83",x"60",x"C3",x"4B",x"2E",x"3A",x"96",x"63",x"0F",x"D2",x"78",x"2E",x"AF",x"32",
		x"96",x"63",x"DD",x"36",x"05",x"50",x"DD",x"36",x"0D",x"01",x"CD",x"57",x"00",x"E6",x"0F",x"C6",
		x"F8",x"DD",x"77",x"03",x"DD",x"36",x"00",x"01",x"21",x"AA",x"39",x"DD",x"75",x"0E",x"DD",x"74",
		x"0F",x"C3",x"78",x"2E",x"3E",x"0B",x"F7",x"D7",x"11",x"18",x"6A",x"DD",x"21",x"80",x"66",x"DD",
		x"7E",x"01",x"0F",x"DA",x"ED",x"2E",x"11",x"1C",x"6A",x"DD",x"21",x"90",x"66",x"DD",x"36",x"0E",
		x"00",x"DD",x"36",x"0F",x"F0",x"3A",x"17",x"62",x"0F",x"D2",x"97",x"2F",x"AF",x"32",x"18",x"62",
		x"21",x"89",x"60",x"36",x"04",x"DD",x"36",x"09",x"06",x"DD",x"36",x"0A",x"03",x"06",x"1E",x"3A",
		x"07",x"62",x"CB",x"27",x"D2",x"1B",x"2F",x"F6",x"80",x"CB",x"F8",x"F6",x"08",x"4F",x"3A",x"94",
		x"63",x"CB",x"5F",x"CA",x"43",x"2F",x"CB",x"C0",x"CB",x"C1",x"DD",x"36",x"09",x"05",x"DD",x"36",
		x"0A",x"06",x"DD",x"36",x"0F",x"00",x"DD",x"36",x"0E",x"F0",x"CB",x"79",x"CA",x"43",x"2F",x"DD",
		x"36",x"0E",x"10",x"79",x"32",x"4D",x"69",x"0E",x"07",x"21",x"94",x"63",x"34",x"C2",x"B7",x"2F",
		x"21",x"95",x"63",x"34",x"7E",x"FE",x"02",x"C2",x"BE",x"2F",x"AF",x"32",x"95",x"63",x"32",x"17",
		x"62",x"DD",x"77",x"01",x"3A",x"03",x"62",x"ED",x"44",x"DD",x"77",x"0E",x"3A",x"07",x"62",x"32",
		x"4D",x"69",x"DD",x"36",x"00",x"00",x"3A",x"89",x"63",x"32",x"89",x"60",x"EB",x"3A",x"03",x"62",
		x"DD",x"86",x"0E",x"77",x"DD",x"77",x"03",x"23",x"70",x"23",x"71",x"23",x"3A",x"05",x"62",x"DD",
		x"86",x"0F",x"77",x"DD",x"77",x"05",x"C9",x"3A",x"18",x"62",x"0F",x"D0",x"DD",x"36",x"09",x"06",
		x"DD",x"36",x"0A",x"03",x"3A",x"07",x"62",x"07",x"3E",x"3C",x"1F",x"47",x"0E",x"07",x"3A",x"89",
		x"60",x"32",x"89",x"63",x"C3",x"7C",x"2F",x"3A",x"95",x"63",x"A7",x"CA",x"7C",x"2F",x"3A",x"1A",
		x"60",x"CB",x"5F",x"CA",x"7C",x"2F",x"0E",x"01",x"C3",x"7C",x"2F",x"3E",x"0E",x"F7",x"21",x"B4",
		x"62",x"35",x"C0",x"3E",x"03",x"32",x"B9",x"62",x"32",x"96",x"63",x"11",x"01",x"05",x"CD",x"9F",
		x"30",x"3A",x"B3",x"62",x"77",x"21",x"B1",x"62",x"35",x"C0",x"3E",x"01",x"32",x"86",x"63",x"C9",
		x"7D",x"0F",x"0F",x"0F",x"E6",x"1F",x"6F",x"7C",x"2F",x"E6",x"F8",x"5F",x"AF",x"67",x"CB",x"13",
		x"17",x"CB",x"13",x"17",x"C6",x"74",x"57",x"19",x"C9",x"57",x"0F",x"DA",x"22",x"30",x"0E",x"93",
		x"0F",x"0F",x"D2",x"17",x"30",x"0E",x"6C",x"07",x"DA",x"31",x"30",x"79",x"E6",x"F0",x"4F",x"C3",
		x"31",x"30",x"0E",x"B4",x"0F",x"0F",x"D2",x"2B",x"30",x"0E",x"1E",x"CB",x"50",x"CA",x"31",x"30",
		x"05",x"79",x"0F",x"0F",x"4F",x"E6",x"03",x"B8",x"C2",x"31",x"30",x"79",x"0F",x"0F",x"E6",x"03",
		x"FE",x"03",x"C0",x"CB",x"92",x"15",x"C0",x"3E",x"04",x"C9",x"11",x"E0",x"FF",x"3A",x"8E",x"63",
		x"4F",x"06",x"00",x"21",x"00",x"76",x"CD",x"64",x"30",x"21",x"C0",x"75",x"CD",x"64",x"30",x"21",
		x"8E",x"63",x"35",x"C9",x"09",x"7E",x"19",x"77",x"C9",x"DF",x"2A",x"C0",x"63",x"34",x"C9",x"21",
		x"AF",x"62",x"34",x"7E",x"E6",x"07",x"C0",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"0E",x"81",x"21",
		x"09",x"69",x"CD",x"96",x"30",x"21",x"1D",x"69",x"CD",x"96",x"30",x"CD",x"57",x"00",x"E6",x"80",
		x"21",x"2D",x"69",x"AE",x"77",x"C9",x"06",x"02",x"79",x"AE",x"77",x"19",x"10",x"FA",x"C9",x"E5",
		x"21",x"C0",x"60",x"3A",x"B0",x"60",x"6F",x"CB",x"7E",x"CA",x"BB",x"30",x"72",x"2C",x"73",x"2C",
		x"7D",x"FE",x"C0",x"D2",x"B8",x"30",x"3E",x"C0",x"32",x"B0",x"60",x"E1",x"C9",x"21",x"50",x"69",
		x"06",x"02",x"CD",x"E4",x"30",x"2E",x"80",x"06",x"0A",x"CD",x"E4",x"30",x"2E",x"B8",x"06",x"0B",
		x"CD",x"E4",x"30",x"21",x"0C",x"6A",x"06",x"05",x"C3",x"E4",x"30",x"21",x"4C",x"69",x"36",x"00",
		x"2E",x"58",x"06",x"06",x"7D",x"36",x"00",x"C6",x"04",x"6F",x"10",x"F9",x"C9",x"CD",x"FA",x"30",
		x"CD",x"3C",x"31",x"CD",x"B1",x"31",x"CD",x"F3",x"34",x"C9",x"3A",x"80",x"63",x"FE",x"06",x"38",
		x"02",x"3E",x"05",x"EF",x"10",x"31",x"10",x"31",x"1B",x"31",x"26",x"31",x"26",x"31",x"31",x"31",
		x"3A",x"1A",x"60",x"E6",x"01",x"FE",x"01",x"C8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"07",
		x"FE",x"05",x"F8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"03",x"FE",x"03",x"F8",x"33",x"33",
		x"C9",x"3A",x"1A",x"60",x"E6",x"07",x"FE",x"07",x"F8",x"33",x"33",x"C9",x"DD",x"21",x"00",x"64",
		x"AF",x"32",x"A1",x"63",x"06",x"05",x"11",x"20",x"00",x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"7C",
		x"31",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"3E",x"01",x"DD",x"77",x"08",x"3A",x"17",x"62",
		x"FE",x"01",x"C2",x"6A",x"31",x"3E",x"00",x"DD",x"77",x"08",x"DD",x"19",x"10",x"DB",x"21",x"A0",
		x"63",x"36",x"00",x"3A",x"A1",x"63",x"FE",x"00",x"C0",x"33",x"33",x"C9",x"3A",x"A1",x"63",x"FE",
		x"05",x"CA",x"6A",x"31",x"3A",x"27",x"62",x"FE",x"02",x"C2",x"95",x"31",x"3A",x"A1",x"63",x"4F",
		x"3A",x"80",x"63",x"B9",x"C8",x"3A",x"A0",x"63",x"FE",x"01",x"C2",x"6A",x"31",x"DD",x"77",x"00",
		x"DD",x"77",x"18",x"AF",x"32",x"A0",x"63",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"C3",x"6A",
		x"31",x"CD",x"DD",x"31",x"AF",x"32",x"A2",x"63",x"21",x"E0",x"63",x"22",x"C8",x"63",x"2A",x"C8",
		x"63",x"01",x"20",x"00",x"09",x"22",x"C8",x"63",x"7E",x"A7",x"CA",x"D0",x"31",x"CD",x"02",x"32",
		x"3A",x"A2",x"63",x"3C",x"32",x"A2",x"63",x"FE",x"05",x"C2",x"BE",x"31",x"C9",x"3A",x"80",x"63",
		x"FE",x"03",x"F8",x"CD",x"F6",x"31",x"FE",x"01",x"C0",x"21",x"39",x"64",x"3E",x"02",x"77",x"21",
		x"79",x"64",x"3E",x"02",x"77",x"C9",x"3A",x"18",x"60",x"E6",x"03",x"FE",x"01",x"C0",x"3A",x"1A",
		x"60",x"C9",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"18",x"FE",x"01",x"CA",x"7A",x"32",x"DD",x"7E",
		x"0D",x"FE",x"04",x"F2",x"30",x"32",x"DD",x"7E",x"19",x"FE",x"02",x"CA",x"7E",x"32",x"CD",x"0F",
		x"33",x"3A",x"18",x"60",x"E6",x"03",x"C2",x"33",x"32",x"DD",x"7E",x"0D",x"A7",x"CA",x"57",x"32",
		x"CD",x"3D",x"33",x"DD",x"7E",x"0D",x"FE",x"04",x"F2",x"91",x"32",x"CD",x"AD",x"33",x"CD",x"8C",
		x"29",x"FE",x"01",x"CA",x"97",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0E",x"FE",x"10",x"DA",
		x"8C",x"32",x"FE",x"F0",x"D2",x"84",x"32",x"DD",x"7E",x"13",x"FE",x"00",x"C2",x"B9",x"32",x"3E",
		x"11",x"DD",x"77",x"13",x"16",x"00",x"5F",x"21",x"7A",x"3A",x"19",x"7E",x"DD",x"46",x"0E",x"DD",
		x"70",x"03",x"DD",x"4E",x"0F",x"81",x"DD",x"77",x"05",x"C9",x"CD",x"BD",x"32",x"C9",x"CD",x"D6",
		x"32",x"C3",x"29",x"32",x"3E",x"02",x"DD",x"77",x"0D",x"C3",x"57",x"32",x"3E",x"01",x"C3",x"86",
		x"32",x"CD",x"E7",x"33",x"C3",x"57",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0D",x"FE",x"01",
		x"C2",x"B1",x"32",x"3E",x"02",x"DD",x"35",x"0E",x"DD",x"77",x"0D",x"CD",x"C3",x"33",x"C3",x"57",
		x"32",x"3E",x"01",x"DD",x"34",x"0E",x"C3",x"A8",x"32",x"3D",x"C3",x"61",x"32",x"3A",x"27",x"62",
		x"FE",x"01",x"CA",x"CE",x"32",x"FE",x"02",x"CA",x"D2",x"32",x"CD",x"B9",x"34",x"C9",x"CD",x"2C",
		x"34",x"C9",x"CD",x"78",x"34",x"C9",x"DD",x"7E",x"1C",x"FE",x"00",x"C2",x"FD",x"32",x"DD",x"7E",
		x"1D",x"FE",x"01",x"C2",x"0B",x"33",x"DD",x"36",x"1D",x"00",x"3A",x"05",x"62",x"DD",x"46",x"0F",
		x"90",x"DA",x"03",x"33",x"DD",x"36",x"1C",x"FF",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"35",x"1C",
		x"C2",x"F8",x"32",x"DD",x"36",x"19",x"00",x"DD",x"36",x"1C",x"00",x"CD",x"0F",x"33",x"C9",x"DD",
		x"7E",x"16",x"FE",x"00",x"C2",x"32",x"33",x"DD",x"36",x"16",x"2B",x"DD",x"36",x"0D",x"00",x"3A",
		x"18",x"60",x"0F",x"D2",x"32",x"33",x"DD",x"7E",x"0D",x"FE",x"01",x"CA",x"36",x"33",x"DD",x"36",
		x"0D",x"01",x"DD",x"35",x"16",x"C9",x"DD",x"36",x"0D",x"02",x"C3",x"32",x"33",x"DD",x"7E",x"0D",
		x"FE",x"08",x"CA",x"71",x"33",x"FE",x"04",x"CA",x"8A",x"33",x"CD",x"A1",x"33",x"DD",x"7E",x"0F",
		x"C6",x"08",x"57",x"DD",x"7E",x"0E",x"01",x"15",x"00",x"CD",x"6E",x"23",x"A7",x"CA",x"99",x"33",
		x"DD",x"70",x"1F",x"3A",x"05",x"62",x"47",x"DD",x"7E",x"0F",x"90",x"D0",x"DD",x"36",x"0D",x"04",
		x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"DD",
		x"7E",x"19",x"FE",x"02",x"C0",x"DD",x"36",x"1D",x"01",x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",
		x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"70",x"1F",x"DD",x"36",x"0D",x"08",
		x"C9",x"3E",x"07",x"F7",x"DD",x"7E",x"0F",x"FE",x"59",x"D0",x"33",x"33",x"C9",x"DD",x"7E",x"0D",
		x"FE",x"01",x"CA",x"D9",x"33",x"DD",x"7E",x"07",x"E6",x"7F",x"DD",x"77",x"07",x"DD",x"35",x"0E",
		x"CD",x"09",x"34",x"3A",x"27",x"62",x"FE",x"01",x"C0",x"DD",x"66",x"0E",x"DD",x"6E",x"0F",x"DD",
		x"46",x"0D",x"CD",x"33",x"23",x"DD",x"75",x"0F",x"C9",x"DD",x"7E",x"07",x"F6",x"80",x"DD",x"77",
		x"07",x"DD",x"34",x"0E",x"C3",x"C0",x"33",x"CD",x"09",x"34",x"DD",x"7E",x"0D",x"FE",x"08",x"C2",
		x"05",x"34",x"DD",x"7E",x"14",x"A7",x"C2",x"01",x"34",x"DD",x"36",x"14",x"02",x"DD",x"35",x"0F",
		x"C9",x"DD",x"35",x"14",x"C9",x"DD",x"34",x"0F",x"C9",x"DD",x"7E",x"15",x"A7",x"C2",x"28",x"34",
		x"DD",x"36",x"15",x"02",x"DD",x"34",x"07",x"DD",x"7E",x"07",x"E6",x"0F",x"FE",x"0F",x"C0",x"DD",
		x"7E",x"07",x"EE",x"02",x"DD",x"77",x"07",x"C9",x"DD",x"35",x"15",x"C9",x"DD",x"6E",x"1A",x"DD",
		x"66",x"1B",x"AF",x"01",x"00",x"00",x"ED",x"4A",x"C2",x"42",x"34",x"21",x"8C",x"3A",x"DD",x"36",
		x"03",x"26",x"DD",x"34",x"03",x"7E",x"FE",x"AA",x"CA",x"56",x"34",x"DD",x"77",x"05",x"23",x"DD",
		x"75",x"1A",x"DD",x"74",x"1B",x"C9",x"AF",x"DD",x"77",x"13",x"DD",x"77",x"18",x"DD",x"77",x"0D",
		x"DD",x"77",x"1C",x"DD",x"7E",x"03",x"DD",x"77",x"0E",x"DD",x"7E",x"05",x"DD",x"77",x"0F",x"DD",
		x"36",x"1A",x"00",x"DD",x"36",x"1B",x"00",x"C9",x"DD",x"6E",x"1A",x"DD",x"66",x"1B",x"AF",x"01",
		x"00",x"00",x"ED",x"4A",x"C2",x"9A",x"34",x"21",x"AC",x"3A",x"3A",x"03",x"62",x"CB",x"7F",x"CA",
		x"A8",x"34",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"03",x"7E",x"DD",x"7E",x"0D",x"FE",x"01",x"C2",
		x"B3",x"34",x"DD",x"34",x"03",x"C3",x"45",x"34",x"DD",x"36",x"0D",x"02",x"DD",x"36",x"03",x"80",
		x"C3",x"9A",x"34",x"DD",x"35",x"03",x"C3",x"45",x"34",x"3A",x"27",x"62",x"FE",x"03",x"C8",x"3A",
		x"03",x"62",x"CB",x"7F",x"C2",x"ED",x"34",x"21",x"C4",x"3A",x"06",x"00",x"3A",x"19",x"60",x"E6",
		x"06",x"4F",x"09",x"7E",x"DD",x"77",x"03",x"DD",x"77",x"0E",x"23",x"7E",x"DD",x"77",x"05",x"DD",
		x"77",x"0F",x"AF",x"DD",x"77",x"0D",x"DD",x"77",x"18",x"DD",x"77",x"1C",x"C9",x"21",x"D4",x"3A",
		x"C3",x"CA",x"34",x"21",x"00",x"64",x"11",x"D0",x"69",x"06",x"05",x"7E",x"A7",x"CA",x"1E",x"35",
		x"2C",x"2C",x"2C",x"7E",x"12",x"3E",x"04",x"85",x"6F",x"1C",x"7E",x"12",x"2C",x"1C",x"7E",x"12",
		x"2D",x"2D",x"2D",x"1C",x"7E",x"12",x"13",x"3E",x"1B",x"85",x"6F",x"10",x"DE",x"C9",x"3E",x"05",
		x"85",x"6F",x"3E",x"04",x"83",x"5F",x"C3",x"17",x"35",x"00",x"00",x"00",x"00",x"01",x"00",x"00",
		x"02",x"00",x"00",x"03",x"00",x"00",x"04",x"00",x"00",x"05",x"00",x"00",x"06",x"00",x"00",x"07",
		x"00",x"00",x"08",x"00",x"00",x"09",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",
		x"00",x"30",x"00",x"00",x"40",x"00",x"00",x"50",x"00",x"00",x"60",x"00",x"00",x"70",x"00",x"00",
		x"80",x"00",x"00",x"90",x"00",x"94",x"77",x"01",x"23",x"24",x"10",x"10",x"00",x"00",x"07",x"06",
		x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3F",x"00",x"50",x"76",x"00",x"F4",x"76",x"96",x"77",x"02",x"1E",x"14",x"10",x"10",x"00",x"00",
		x"06",x"01",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"3F",x"00",x"00",x"61",x"00",x"F6",x"76",x"98",x"77",x"03",x"22",x"14",x"10",x"10",
		x"00",x"00",x"05",x"09",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"59",x"00",x"F8",x"76",x"9A",x"77",x"04",x"24",x"18",
		x"10",x"10",x"00",x"00",x"05",x"00",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"50",x"00",x"FA",x"76",x"9C",x"77",x"05",
		x"24",x"18",x"10",x"10",x"00",x"00",x"04",x"03",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"00",x"43",x"00",x"FC",x"76",x"3B",
		x"5C",x"4B",x"5C",x"5B",x"5C",x"6B",x"5C",x"7B",x"5C",x"8B",x"5C",x"9B",x"5C",x"AB",x"5C",x"BB",
		x"5C",x"CB",x"5C",x"3B",x"6C",x"4B",x"6C",x"5B",x"6C",x"6B",x"6C",x"7B",x"6C",x"8B",x"6C",x"9B",
		x"6C",x"AB",x"6C",x"BB",x"6C",x"CB",x"6C",x"3B",x"7C",x"4B",x"7C",x"5B",x"7C",x"6B",x"7C",x"7B",
		x"7C",x"8B",x"7C",x"9B",x"7C",x"AB",x"7C",x"BB",x"7C",x"CB",x"7C",x"8B",x"36",x"01",x"00",x"98",
		x"36",x"A5",x"36",x"B2",x"36",x"BF",x"36",x"06",x"00",x"CC",x"36",x"08",x"00",x"E6",x"36",x"FD",
		x"36",x"0B",x"00",x"15",x"37",x"1C",x"37",x"30",x"37",x"38",x"37",x"47",x"37",x"5D",x"37",x"73",
		x"37",x"8B",x"37",x"00",x"61",x"22",x"61",x"44",x"61",x"66",x"61",x"88",x"61",x"9E",x"37",x"B6",
		x"37",x"D2",x"37",x"E1",x"37",x"1D",x"00",x"00",x"3F",x"09",x"3F",x"96",x"76",x"17",x"11",x"1D",
		x"15",x"10",x"10",x"1F",x"26",x"15",x"22",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",
		x"10",x"30",x"32",x"31",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"30",x"33",
		x"31",x"3F",x"80",x"76",x"18",x"19",x"17",x"18",x"10",x"23",x"13",x"1F",x"22",x"15",x"3F",x"9F",
		x"75",x"13",x"22",x"15",x"14",x"19",x"24",x"10",x"10",x"10",x"10",x"3F",x"5E",x"77",x"18",x"1F",
		x"27",x"10",x"18",x"19",x"17",x"18",x"10",x"13",x"11",x"1E",x"10",x"29",x"1F",x"25",x"10",x"17",
		x"15",x"24",x"10",x"FB",x"10",x"3F",x"29",x"77",x"1F",x"1E",x"1C",x"29",x"10",x"01",x"10",x"20",
		x"1C",x"11",x"29",x"15",x"22",x"10",x"12",x"25",x"24",x"24",x"1F",x"1E",x"3F",x"29",x"77",x"01",
		x"10",x"1F",x"22",x"10",x"02",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"23",x"10",x"12",x"25",
		x"24",x"24",x"1F",x"1E",x"3F",x"27",x"76",x"20",x"25",x"23",x"18",x"3F",x"06",x"77",x"1E",x"11",
		x"1D",x"15",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"22",x"11",x"24",x"19",x"1F",x"1E",x"3F",
		x"88",x"76",x"1E",x"11",x"1D",x"15",x"2E",x"3F",x"E9",x"75",x"2D",x"2D",x"2D",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"0B",x"77",x"11",x"10",x"12",x"10",x"13",x"10",x"14",
		x"10",x"15",x"10",x"16",x"10",x"17",x"10",x"18",x"10",x"19",x"10",x"1A",x"3F",x"0D",x"77",x"1B",
		x"10",x"1C",x"10",x"1D",x"10",x"1E",x"10",x"1F",x"10",x"20",x"10",x"21",x"10",x"22",x"10",x"23",
		x"10",x"24",x"3F",x"0F",x"77",x"25",x"10",x"26",x"10",x"27",x"10",x"28",x"10",x"29",x"10",x"2A",
		x"10",x"2B",x"10",x"2C",x"44",x"45",x"46",x"47",x"48",x"10",x"3F",x"F2",x"76",x"22",x"15",x"17",
		x"19",x"10",x"24",x"19",x"1D",x"15",x"10",x"10",x"30",x"03",x"00",x"31",x"10",x"3F",x"92",x"77",
		x"22",x"11",x"1E",x"1B",x"10",x"10",x"23",x"13",x"1F",x"22",x"15",x"10",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"10",x"10",x"10",x"3F",x"72",x"77",x"29",x"1F",x"25",x"22",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"27",x"11",x"23",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"15",x"22",x"15",x"14",
		x"42",x"3F",x"A7",x"76",x"19",x"1E",x"23",x"15",x"22",x"24",x"10",x"13",x"1F",x"19",x"1E",x"10",
		x"3F",x"0A",x"77",x"10",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"10",x"10",x"10",x"13",
		x"1F",x"19",x"1E",x"3F",x"FC",x"76",x"49",x"4A",x"10",x"1E",x"19",x"1E",x"24",x"15",x"1E",x"14",
		x"1F",x"10",x"10",x"10",x"10",x"3F",x"7C",x"75",x"01",x"09",x"08",x"01",x"3F",x"02",x"97",x"38",
		x"68",x"38",x"02",x"DF",x"54",x"10",x"54",x"02",x"EF",x"6D",x"20",x"6D",x"02",x"DF",x"8E",x"10",
		x"8E",x"02",x"EF",x"AF",x"20",x"AF",x"02",x"DF",x"D0",x"10",x"D0",x"02",x"EF",x"F1",x"10",x"F1",
		x"00",x"53",x"18",x"53",x"54",x"00",x"63",x"18",x"63",x"54",x"00",x"93",x"38",x"93",x"54",x"00",
		x"83",x"54",x"83",x"F1",x"00",x"93",x"54",x"93",x"F1",x"AA",x"8D",x"7D",x"8C",x"6F",x"00",x"7C",
		x"6E",x"00",x"7C",x"6D",x"00",x"7C",x"6C",x"00",x"7C",x"8F",x"7F",x"8E",x"47",x"27",x"08",x"50",
		x"2F",x"A7",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"23",x"07",x"40",
		x"46",x"A9",x"08",x"44",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",x"70",x"08",x"48",
		x"00",x"70",x"0A",x"48",x"6F",x"10",x"09",x"23",x"6F",x"11",x"0A",x"33",x"50",x"34",x"08",x"3C",
		x"00",x"35",x"08",x"3C",x"53",x"32",x"08",x"40",x"63",x"33",x"08",x"40",x"00",x"70",x"08",x"48",
		x"53",x"36",x"08",x"50",x"63",x"37",x"08",x"50",x"6B",x"31",x"08",x"41",x"00",x"70",x"08",x"48",
		x"6A",x"14",x"0A",x"48",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"7F",x"04",x"7F",x"F0",x"10",
		x"F0",x"02",x"DF",x"F2",x"70",x"F8",x"02",x"6F",x"F8",x"10",x"F8",x"AA",x"04",x"DF",x"D0",x"90",
		x"D0",x"02",x"DF",x"DC",x"20",x"D1",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"04",x"DF",x"A8",x"20",
		x"A8",x"04",x"5F",x"B0",x"20",x"B0",x"02",x"DF",x"B0",x"20",x"BB",x"AA",x"04",x"DF",x"88",x"30",
		x"88",x"04",x"DF",x"90",x"B0",x"90",x"02",x"DF",x"9A",x"20",x"8F",x"AA",x"04",x"BF",x"68",x"20",
		x"68",x"04",x"3F",x"70",x"20",x"70",x"02",x"DF",x"6E",x"20",x"79",x"AA",x"02",x"DF",x"58",x"A0",
		x"55",x"AA",x"00",x"70",x"08",x"44",x"2B",x"AC",x"08",x"4C",x"3B",x"AE",x"08",x"4C",x"3B",x"AF",
		x"08",x"3C",x"4B",x"B0",x"07",x"3C",x"4B",x"AD",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"47",x"27",x"08",x"4C",x"2F",x"A7",
		x"08",x"4C",x"3B",x"25",x"08",x"4C",x"00",x"70",x"08",x"44",x"3B",x"23",x"07",x"3C",x"4B",x"2A",
		x"08",x"3C",x"4B",x"2B",x"08",x"4C",x"2B",x"AA",x"08",x"3C",x"2B",x"AB",x"08",x"4C",x"00",x"70",
		x"0A",x"44",x"00",x"70",x"08",x"44",x"4B",x"2C",x"08",x"4C",x"3B",x"2E",x"08",x"4C",x"3B",x"2F",
		x"08",x"3C",x"2B",x"30",x"07",x"3C",x"2B",x"2D",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"02",x"02",x"02",x"02",x"03",
		x"03",x"03",x"7F",x"1E",x"4E",x"BB",x"4C",x"D8",x"4E",x"59",x"4E",x"7F",x"BB",x"4D",x"7F",x"47",
		x"27",x"08",x"50",x"2D",x"26",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",
		x"24",x"07",x"40",x"4B",x"28",x"08",x"40",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",
		x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"49",x"A6",x"08",x"50",x"2F",x"A7",x"08",x"50",x"3B",
		x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"24",x"07",x"40",x"46",x"A9",x"08",x"44",x"00",
		x"70",x"08",x"48",x"2B",x"A8",x"08",x"40",x"00",x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"73",
		x"A7",x"88",x"60",x"8B",x"27",x"88",x"60",x"7F",x"25",x"88",x"60",x"00",x"70",x"88",x"68",x"7F",
		x"24",x"87",x"70",x"74",x"29",x"88",x"6C",x"00",x"70",x"88",x"68",x"8A",x"A9",x"88",x"6C",x"00",
		x"70",x"88",x"68",x"00",x"70",x"8A",x"68",x"05",x"AF",x"F0",x"50",x"F0",x"AA",x"05",x"AF",x"E8",
		x"50",x"E8",x"AA",x"05",x"AF",x"E0",x"50",x"E0",x"AA",x"05",x"AF",x"D8",x"50",x"D8",x"AA",x"05",
		x"B7",x"58",x"48",x"58",x"AA",x"01",x"04",x"01",x"03",x"04",x"01",x"02",x"03",x"04",x"01",x"02",
		x"01",x"03",x"04",x"01",x"02",x"01",x"03",x"01",x"04",x"7F",x"FF",x"00",x"FF",x"FF",x"FE",x"FE",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"00",x"E8",x"E5",x"E3",x"E2",
		x"E1",x"E0",x"DF",x"DE",x"DD",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DE",x"DF",
		x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E7",x"E9",x"EB",x"ED",x"F0",x"AA",x"80",x"7B",x"78",x"76",
		x"74",x"73",x"72",x"71",x"70",x"70",x"6F",x"6F",x"6F",x"70",x"70",x"71",x"72",x"73",x"74",x"75",
		x"76",x"77",x"78",x"AA",x"EE",x"F0",x"DB",x"A0",x"E6",x"C8",x"D6",x"78",x"EB",x"F0",x"DB",x"A0",
		x"E6",x"C8",x"E6",x"C8",x"1B",x"C8",x"23",x"A0",x"2B",x"78",x"12",x"F0",x"1B",x"C8",x"23",x"A0",
		x"12",x"F0",x"1B",x"C8",x"02",x"97",x"38",x"68",x"38",x"02",x"9F",x"54",x"10",x"54",x"02",x"DF",
		x"58",x"A0",x"55",x"02",x"EF",x"6D",x"20",x"79",x"02",x"DF",x"9A",x"10",x"8E",x"02",x"EF",x"AF",
		x"20",x"BB",x"02",x"DF",x"DC",x"10",x"D0",x"02",x"FF",x"F0",x"80",x"F7",x"02",x"7F",x"F8",x"00",
		x"F8",x"00",x"CB",x"57",x"CB",x"6F",x"00",x"CB",x"99",x"CB",x"B1",x"00",x"CB",x"DB",x"CB",x"F3",
		x"00",x"63",x"18",x"63",x"54",x"01",x"63",x"D5",x"63",x"F8",x"00",x"33",x"78",x"33",x"90",x"00",
		x"33",x"BA",x"33",x"D2",x"00",x"53",x"18",x"53",x"54",x"01",x"53",x"92",x"53",x"B8",x"00",x"5B",
		x"76",x"5B",x"92",x"00",x"73",x"B6",x"73",x"D6",x"00",x"83",x"95",x"83",x"B5",x"00",x"93",x"38",
		x"93",x"54",x"01",x"BB",x"70",x"BB",x"98",x"01",x"6B",x"54",x"6B",x"75",x"AA",x"06",x"8F",x"90",
		x"70",x"90",x"06",x"8F",x"98",x"70",x"98",x"06",x"8F",x"A0",x"70",x"A0",x"00",x"63",x"18",x"63",
		x"58",x"00",x"63",x"80",x"63",x"A8",x"00",x"63",x"D0",x"63",x"F8",x"00",x"53",x"18",x"53",x"58",
		x"00",x"53",x"A8",x"53",x"D0",x"00",x"9B",x"80",x"9B",x"A8",x"00",x"9B",x"D0",x"9B",x"F8",x"01",
		x"23",x"58",x"23",x"80",x"01",x"DB",x"58",x"DB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"A3",x"A8",x"A3",x"D0",x"00",x"2B",x"D0",x"2B",x"F8",x"00",x"D3",x"D0",
		x"D3",x"F8",x"00",x"93",x"38",x"93",x"58",x"02",x"97",x"38",x"68",x"38",x"03",x"EF",x"58",x"10",
		x"58",x"03",x"F7",x"80",x"88",x"80",x"03",x"77",x"80",x"08",x"80",x"02",x"A7",x"A8",x"50",x"A8",
		x"02",x"E7",x"A8",x"B8",x"A8",x"02",x"3F",x"A8",x"18",x"A8",x"03",x"EF",x"D0",x"10",x"D0",x"02",
		x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"63",x"18",x"63",x"58",x"00",x"63",x"88",x"63",x"D0",x"00",
		x"53",x"18",x"53",x"58",x"00",x"53",x"88",x"53",x"D0",x"00",x"E3",x"68",x"E3",x"90",x"00",x"E3",
		x"B8",x"E3",x"D0",x"00",x"CB",x"90",x"CB",x"B0",x"00",x"B3",x"58",x"B3",x"78",x"00",x"9B",x"80",
		x"9B",x"A0",x"00",x"93",x"38",x"93",x"58",x"00",x"23",x"88",x"23",x"C0",x"00",x"1B",x"C0",x"1B",
		x"E8",x"02",x"97",x"38",x"68",x"38",x"02",x"B7",x"58",x"10",x"58",x"02",x"EF",x"68",x"E0",x"68",
		x"02",x"D7",x"70",x"C8",x"70",x"02",x"BF",x"78",x"B0",x"78",x"02",x"A7",x"80",x"90",x"80",x"02",
		x"67",x"88",x"48",x"88",x"02",x"27",x"88",x"10",x"88",x"02",x"EF",x"90",x"C8",x"90",x"02",x"A7",
		x"A0",x"98",x"A0",x"02",x"BF",x"A8",x"B0",x"A8",x"02",x"D7",x"B0",x"C8",x"B0",x"02",x"EF",x"B8",
		x"E0",x"B8",x"02",x"27",x"C0",x"10",x"C0",x"02",x"EF",x"D0",x"D8",x"D0",x"02",x"67",x"D0",x"50",
		x"D0",x"02",x"CF",x"D8",x"C0",x"D8",x"02",x"B7",x"E0",x"A8",x"E0",x"02",x"9F",x"E8",x"88",x"E8",
		x"02",x"27",x"E8",x"10",x"E8",x"02",x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"7B",x"80",x"7B",x"A8",
		x"00",x"7B",x"D0",x"7B",x"F8",x"00",x"33",x"58",x"33",x"80",x"00",x"53",x"58",x"53",x"80",x"00",
		x"AB",x"58",x"AB",x"80",x"00",x"CB",x"58",x"CB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"23",x"A8",x"23",x"D0",x"00",x"5B",x"A8",x"5B",x"D0",x"00",x"A3",x"A8",
		x"A3",x"D0",x"00",x"DB",x"A8",x"DB",x"D0",x"00",x"1B",x"D0",x"1B",x"F8",x"00",x"E3",x"D0",x"E3",
		x"F8",x"05",x"B7",x"30",x"48",x"30",x"05",x"CF",x"58",x"30",x"58",x"05",x"D7",x"80",x"28",x"80",
		x"05",x"DF",x"A8",x"20",x"A8",x"05",x"E7",x"D0",x"18",x"D0",x"05",x"EF",x"F8",x"10",x"F8",x"AA",
		x"10",x"82",x"85",x"8B",x"10",x"85",x"80",x"8B",x"10",x"87",x"85",x"8B",x"81",x"80",x"80",x"8B",
		x"81",x"82",x"85",x"8B",x"81",x"85",x"80",x"8B",x"05",x"88",x"77",x"01",x"68",x"77",x"01",x"6C",
		x"77",x"03",x"49",x"77",x"05",x"08",x"77",x"01",x"E8",x"76",x"01",x"EC",x"76",x"05",x"C8",x"76",
		x"05",x"88",x"76",x"02",x"69",x"76",x"02",x"4A",x"76",x"05",x"28",x"76",x"05",x"E8",x"75",x"01",
		x"CA",x"75",x"03",x"A9",x"75",x"01",x"88",x"75",x"01",x"8C",x"75",x"05",x"48",x"75",x"01",x"28",
		x"75",x"01",x"2A",x"75",x"01",x"2C",x"75",x"01",x"08",x"75",x"01",x"0A",x"75",x"01",x"0C",x"75",
		x"03",x"C8",x"74",x"03",x"AA",x"74",x"03",x"88",x"74",x"05",x"2F",x"77",x"05",x"0F",x"77",x"02",
		x"F0",x"76",x"02",x"CF",x"76",x"02",x"D2",x"76",x"05",x"8F",x"76",x"05",x"6F",x"76",x"01",x"4F",
		x"76",x"01",x"53",x"76",x"05",x"2F",x"76",x"05",x"EF",x"75",x"02",x"D0",x"75",x"02",x"B1",x"75",
		x"05",x"8F",x"75",x"03",x"50",x"75",x"05",x"2F",x"75",x"01",x"0F",x"75",x"01",x"13",x"75",x"01",
		x"EF",x"74",x"01",x"F1",x"74",x"01",x"F3",x"74",x"02",x"D1",x"74",x"00",x"00",x"00",x"23",x"68",
		x"01",x"11",x"00",x"00",x"00",x"10",x"DB",x"68",x"01",x"40",x"00",x"00",x"08",x"01",x"01",x"01",
		x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"01",x"C0",x"FF",
		x"01",x"FF",x"FF",x"34",x"C3",x"39",x"00",x"67",x"80",x"69",x"1A",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"0B",x"4B",
		x"14",x"18",x"0B",x"4B",x"1E",x"18",x"0B",x"3B",x"14",x"18",x"0B",x"3B",x"3D",x"01",x"03",x"02",
		x"4D",x"01",x"04",x"01",x"27",x"70",x"01",x"E0",x"00",x"00",x"7F",x"40",x"01",x"78",x"02",x"00",
		x"27",x"49",x"0C",x"F0",x"7F",x"49",x"0C",x"88",x"1E",x"07",x"03",x"09",x"24",x"64",x"BB",x"C0",
		x"23",x"8D",x"7B",x"B4",x"1B",x"8C",x"7C",x"64",x"4B",x"0E",x"04",x"02",x"23",x"46",x"03",x"68",
		x"DB",x"46",x"03",x"68",x"17",x"50",x"00",x"5C",x"E7",x"D0",x"00",x"5C",x"8C",x"50",x"00",x"84",
		x"73",x"D0",x"00",x"84",x"17",x"50",x"00",x"D4",x"E7",x"D0",x"00",x"D4",x"53",x"73",x"0A",x"A0",
		x"8B",x"74",x"0A",x"F0",x"DB",x"75",x"0A",x"A0",x"5B",x"73",x"0A",x"C8",x"E3",x"74",x"0A",x"60",
		x"1B",x"75",x"0A",x"80",x"DB",x"73",x"0A",x"C8",x"93",x"74",x"0A",x"F0",x"33",x"75",x"0A",x"50",
		x"44",x"03",x"08",x"04",x"37",x"F4",x"37",x"C0",x"37",x"8C",x"77",x"70",x"77",x"A4",x"77",x"D8",
		x"11",x"01",x"00",x"06",x"7B",x"1F",x"D2",x"28",x"1E",x"1E",x"03",x"06",x"7D",x"1F",x"D2",x"28",
		x"1E",x"1E",x"05",x"06",x"7F",x"C3",x"28",x"1E",x"3A",x"27",x"62",x"E5",x"EF",x"00",x"00",x"99",
		x"3E",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",x"E1",x"AF",x"32",x"60",x"60",x"06",x"0A",
		x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"C3",x"3E",x"06",x"05",x"DD",x"21",x"00",x"64",
		x"CD",x"C3",x"3E",x"3A",x"60",x"60",x"A7",x"C8",x"FE",x"01",x"C8",x"FE",x"03",x"3E",x"03",x"D8",
		x"3E",x"07",x"C9",x"DD",x"CB",x"00",x"46",x"CA",x"FA",x"3E",x"79",x"DD",x"96",x"05",x"D2",x"D3",
		x"3E",x"ED",x"44",x"3C",x"95",x"DA",x"DE",x"3E",x"DD",x"96",x"0A",x"D2",x"FA",x"3E",x"FD",x"7E",
		x"03",x"DD",x"96",x"03",x"D2",x"E9",x"3E",x"ED",x"44",x"94",x"DA",x"F3",x"3E",x"DD",x"96",x"09",
		x"D2",x"FA",x"3E",x"3A",x"60",x"60",x"3C",x"32",x"60",x"60",x"DD",x"19",x"10",x"C5",x"C9",x"00",
		x"5C",x"76",x"49",x"4A",x"01",x"09",x"08",x"01",x"3F",x"7D",x"77",x"1E",x"19",x"1E",x"24",x"15",
		x"1E",x"14",x"1F",x"10",x"1F",x"16",x"10",x"11",x"1D",x"15",x"22",x"19",x"13",x"11",x"10",x"19",
		x"1E",x"13",x"2B",x"3F",x"21",x"AF",x"74",x"11",x"E0",x"FF",x"36",x"9F",x"19",x"36",x"9E",x"C9",
		x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"2C",x"57",x"45",x"20",x"57",x"4F",x"55",x"4C",x"44",
		x"20",x"54",x"45",x"41",x"43",x"48",x"20",x"59",x"4F",x"55",x"2E",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"54",x"45",x"4C",x"2E",x"54",x"4F",x"4B",x"59",x"4F",x"2D",x"4A",x"41",x"50",x"41",x"4E",x"20",
		x"30",x"34",x"34",x"28",x"32",x"34",x"34",x"29",x"32",x"31",x"35",x"31",x"20",x"20",x"20",x"20",
		x"45",x"58",x"54",x"45",x"4E",x"54",x"49",x"4F",x"4E",x"20",x"33",x"30",x"34",x"20",x"20",x"20",
		x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"44",x"45",x"53",x"49",x"47",x"4E",x"20",x"20",x"20",
		x"49",x"4B",x"45",x"47",x"41",x"4D",x"49",x"20",x"43",x"4F",x"2E",x"20",x"4C",x"49",x"4D",x"2E",
		x"CD",x"A6",x"3F",x"C3",x"5F",x"0D",x"3E",x"02",x"F7",x"06",x"02",x"21",x"6C",x"77",x"36",x"10",
		x"23",x"23",x"36",x"C0",x"21",x"8C",x"74",x"10",x"F5",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"4D",x"69",x"36",x"03",x"2C",x"2C",x"C9",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"7F",x"7F",x"18",x"3C",x"76",x"63",x"41",x"00",x"00",x"7F",x"7F",x"49",x"49",x"49",x"41",
		x"00",x"1C",x"3E",x"63",x"41",x"49",x"79",x"79",x"00",x"7C",x"7E",x"13",x"11",x"13",x"7E",x"7C",
		x"00",x"7F",x"7F",x"0E",x"1C",x"0E",x"7F",x"7F",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"17",x"CB",x"13",x"17",x"C6",x"74",x"57",x"19",x"C9",x"57",x"0F",x"DA",x"22",x"30",x"0E",x"93",
		x"0F",x"0F",x"D2",x"17",x"30",x"0E",x"6C",x"07",x"DA",x"31",x"30",x"79",x"E6",x"F0",x"4F",x"C3",
		x"31",x"30",x"0E",x"B4",x"0F",x"0F",x"D2",x"2B",x"30",x"0E",x"1E",x"CB",x"50",x"CA",x"31",x"30",
		x"05",x"79",x"0F",x"0F",x"4F",x"E6",x"03",x"B8",x"C2",x"31",x"30",x"79",x"0F",x"0F",x"E6",x"03",
		x"FE",x"03",x"C0",x"CB",x"92",x"15",x"C0",x"3E",x"04",x"C9",x"11",x"E0",x"FF",x"3A",x"8E",x"63",
		x"4F",x"06",x"00",x"21",x"00",x"76",x"CD",x"64",x"30",x"21",x"C0",x"75",x"CD",x"64",x"30",x"21",
		x"8E",x"63",x"35",x"C9",x"09",x"7E",x"19",x"77",x"C9",x"DF",x"2A",x"C0",x"63",x"34",x"C9",x"21",
		x"AF",x"62",x"34",x"7E",x"E6",x"07",x"C0",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"0E",x"81",x"21",
		x"09",x"69",x"CD",x"96",x"30",x"21",x"1D",x"69",x"CD",x"96",x"30",x"CD",x"57",x"00",x"E6",x"80",
		x"21",x"2D",x"69",x"AE",x"77",x"C9",x"06",x"02",x"79",x"AE",x"77",x"19",x"10",x"FA",x"C9",x"E5",
		x"21",x"C0",x"60",x"3A",x"B0",x"60",x"6F",x"CB",x"7E",x"CA",x"BB",x"30",x"72",x"2C",x"73",x"2C",
		x"7D",x"FE",x"C0",x"D2",x"B8",x"30",x"3E",x"C0",x"32",x"B0",x"60",x"E1",x"C9",x"21",x"50",x"69",
		x"06",x"02",x"CD",x"E4",x"30",x"2E",x"80",x"06",x"0A",x"CD",x"E4",x"30",x"2E",x"B8",x"06",x"0B",
		x"CD",x"E4",x"30",x"21",x"0C",x"6A",x"06",x"05",x"C3",x"E4",x"30",x"21",x"4C",x"69",x"36",x"00",
		x"2E",x"58",x"06",x"06",x"7D",x"36",x"00",x"C6",x"04",x"6F",x"10",x"F9",x"C9",x"CD",x"FA",x"30",
		x"CD",x"3C",x"31",x"CD",x"B1",x"31",x"CD",x"F3",x"34",x"C9",x"3A",x"80",x"63",x"FE",x"06",x"38",
		x"02",x"3E",x"05",x"EF",x"10",x"31",x"10",x"31",x"1B",x"31",x"26",x"31",x"26",x"31",x"31",x"31",
		x"3A",x"1A",x"60",x"E6",x"01",x"FE",x"01",x"C8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"07",
		x"FE",x"05",x"F8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"03",x"FE",x"03",x"F8",x"33",x"33",
		x"C9",x"3A",x"1A",x"60",x"E6",x"07",x"FE",x"07",x"F8",x"33",x"33",x"C9",x"DD",x"21",x"00",x"64",
		x"AF",x"32",x"A1",x"63",x"06",x"05",x"11",x"20",x"00",x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"7C",
		x"31",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"3E",x"01",x"DD",x"77",x"08",x"3A",x"17",x"62",
		x"FE",x"01",x"C2",x"6A",x"31",x"3E",x"00",x"DD",x"77",x"08",x"DD",x"19",x"10",x"DB",x"21",x"A0",
		x"63",x"36",x"00",x"3A",x"A1",x"63",x"FE",x"00",x"C0",x"33",x"33",x"C9",x"3A",x"A1",x"63",x"FE",
		x"05",x"CA",x"6A",x"31",x"3A",x"27",x"62",x"FE",x"02",x"C2",x"95",x"31",x"3A",x"A1",x"63",x"4F",
		x"3A",x"80",x"63",x"B9",x"C8",x"3A",x"A0",x"63",x"FE",x"01",x"C2",x"6A",x"31",x"DD",x"77",x"00",
		x"DD",x"77",x"18",x"AF",x"32",x"A0",x"63",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"C3",x"6A",
		x"31",x"CD",x"DD",x"31",x"AF",x"32",x"A2",x"63",x"21",x"E0",x"63",x"22",x"C8",x"63",x"2A",x"C8",
		x"63",x"01",x"20",x"00",x"09",x"22",x"C8",x"63",x"7E",x"A7",x"CA",x"D0",x"31",x"CD",x"02",x"32",
		x"3A",x"A2",x"63",x"3C",x"32",x"A2",x"63",x"FE",x"05",x"C2",x"BE",x"31",x"C9",x"3A",x"80",x"63",
		x"FE",x"03",x"F8",x"CD",x"F6",x"31",x"FE",x"01",x"C0",x"21",x"39",x"64",x"3E",x"02",x"77",x"21",
		x"79",x"64",x"3E",x"02",x"77",x"C9",x"3A",x"18",x"60",x"E6",x"03",x"FE",x"01",x"C0",x"3A",x"1A",
		x"60",x"C9",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"18",x"FE",x"01",x"CA",x"7A",x"32",x"DD",x"7E",
		x"0D",x"FE",x"04",x"F2",x"30",x"32",x"DD",x"7E",x"19",x"FE",x"02",x"CA",x"7E",x"32",x"CD",x"0F",
		x"33",x"3A",x"18",x"60",x"E6",x"03",x"C2",x"33",x"32",x"DD",x"7E",x"0D",x"A7",x"CA",x"57",x"32",
		x"CD",x"3D",x"33",x"DD",x"7E",x"0D",x"FE",x"04",x"F2",x"91",x"32",x"CD",x"AD",x"33",x"CD",x"8C",
		x"29",x"FE",x"01",x"CA",x"97",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0E",x"FE",x"10",x"DA",
		x"8C",x"32",x"FE",x"F0",x"D2",x"84",x"32",x"DD",x"7E",x"13",x"FE",x"00",x"C2",x"B9",x"32",x"3E",
		x"11",x"DD",x"77",x"13",x"16",x"00",x"5F",x"21",x"7A",x"3A",x"19",x"7E",x"DD",x"46",x"0E",x"DD",
		x"70",x"03",x"DD",x"4E",x"0F",x"81",x"DD",x"77",x"05",x"C9",x"CD",x"BD",x"32",x"C9",x"CD",x"D6",
		x"32",x"C3",x"29",x"32",x"3E",x"02",x"DD",x"77",x"0D",x"C3",x"57",x"32",x"3E",x"01",x"C3",x"86",
		x"32",x"CD",x"E7",x"33",x"C3",x"57",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0D",x"FE",x"01",
		x"C2",x"B1",x"32",x"3E",x"02",x"DD",x"35",x"0E",x"DD",x"77",x"0D",x"CD",x"C3",x"33",x"C3",x"57",
		x"32",x"3E",x"01",x"DD",x"34",x"0E",x"C3",x"A8",x"32",x"3D",x"C3",x"61",x"32",x"3A",x"27",x"62",
		x"FE",x"01",x"CA",x"CE",x"32",x"FE",x"02",x"CA",x"D2",x"32",x"CD",x"B9",x"34",x"C9",x"CD",x"2C",
		x"34",x"C9",x"CD",x"78",x"34",x"C9",x"DD",x"7E",x"1C",x"FE",x"00",x"C2",x"FD",x"32",x"DD",x"7E",
		x"1D",x"FE",x"01",x"C2",x"0B",x"33",x"DD",x"36",x"1D",x"00",x"3A",x"05",x"62",x"DD",x"46",x"0F",
		x"90",x"DA",x"03",x"33",x"DD",x"36",x"1C",x"FF",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"35",x"1C",
		x"C2",x"F8",x"32",x"DD",x"36",x"19",x"00",x"DD",x"36",x"1C",x"00",x"CD",x"0F",x"33",x"C9",x"DD",
		x"7E",x"16",x"FE",x"00",x"C2",x"32",x"33",x"DD",x"36",x"16",x"2B",x"DD",x"36",x"0D",x"00",x"3A",
		x"18",x"60",x"0F",x"D2",x"32",x"33",x"DD",x"7E",x"0D",x"FE",x"01",x"CA",x"36",x"33",x"DD",x"36",
		x"0D",x"01",x"DD",x"35",x"16",x"C9",x"DD",x"36",x"0D",x"02",x"C3",x"32",x"33",x"DD",x"7E",x"0D",
		x"FE",x"08",x"CA",x"71",x"33",x"FE",x"04",x"CA",x"8A",x"33",x"CD",x"A1",x"33",x"DD",x"7E",x"0F",
		x"C6",x"08",x"57",x"DD",x"7E",x"0E",x"01",x"15",x"00",x"CD",x"6E",x"23",x"A7",x"CA",x"99",x"33",
		x"DD",x"70",x"1F",x"3A",x"05",x"62",x"47",x"DD",x"7E",x"0F",x"90",x"D0",x"DD",x"36",x"0D",x"04",
		x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"DD",
		x"7E",x"19",x"FE",x"02",x"C0",x"DD",x"36",x"1D",x"01",x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",
		x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"70",x"1F",x"DD",x"36",x"0D",x"08",
		x"C9",x"3E",x"07",x"F7",x"DD",x"7E",x"0F",x"FE",x"59",x"D0",x"33",x"33",x"C9",x"DD",x"7E",x"0D",
		x"FE",x"01",x"CA",x"D9",x"33",x"DD",x"7E",x"07",x"E6",x"7F",x"DD",x"77",x"07",x"DD",x"35",x"0E",
		x"CD",x"09",x"34",x"3A",x"27",x"62",x"FE",x"01",x"C0",x"DD",x"66",x"0E",x"DD",x"6E",x"0F",x"DD",
		x"46",x"0D",x"CD",x"33",x"23",x"DD",x"75",x"0F",x"C9",x"DD",x"7E",x"07",x"F6",x"80",x"DD",x"77",
		x"07",x"DD",x"34",x"0E",x"C3",x"C0",x"33",x"CD",x"09",x"34",x"DD",x"7E",x"0D",x"FE",x"08",x"C2",
		x"05",x"34",x"DD",x"7E",x"14",x"A7",x"C2",x"01",x"34",x"DD",x"36",x"14",x"02",x"DD",x"35",x"0F",
		x"C9",x"DD",x"35",x"14",x"C9",x"DD",x"34",x"0F",x"C9",x"DD",x"7E",x"15",x"A7",x"C2",x"28",x"34",
		x"DD",x"36",x"15",x"02",x"DD",x"34",x"07",x"DD",x"7E",x"07",x"E6",x"0F",x"FE",x"0F",x"C0",x"DD",
		x"7E",x"07",x"EE",x"02",x"DD",x"77",x"07",x"C9",x"DD",x"35",x"15",x"C9",x"DD",x"6E",x"1A",x"DD",
		x"66",x"1B",x"AF",x"01",x"00",x"00",x"ED",x"4A",x"C2",x"42",x"34",x"21",x"8C",x"3A",x"DD",x"36",
		x"03",x"26",x"DD",x"34",x"03",x"7E",x"FE",x"AA",x"CA",x"56",x"34",x"DD",x"77",x"05",x"23",x"DD",
		x"75",x"1A",x"DD",x"74",x"1B",x"C9",x"AF",x"DD",x"77",x"13",x"DD",x"77",x"18",x"DD",x"77",x"0D",
		x"DD",x"77",x"1C",x"DD",x"7E",x"03",x"DD",x"77",x"0E",x"DD",x"7E",x"05",x"DD",x"77",x"0F",x"DD",
		x"36",x"1A",x"00",x"DD",x"36",x"1B",x"00",x"C9",x"DD",x"6E",x"1A",x"DD",x"66",x"1B",x"AF",x"01",
		x"00",x"00",x"ED",x"4A",x"C2",x"9A",x"34",x"21",x"AC",x"3A",x"3A",x"03",x"62",x"CB",x"7F",x"CA",
		x"A8",x"34",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"03",x"7E",x"DD",x"7E",x"0D",x"FE",x"01",x"C2",
		x"B3",x"34",x"DD",x"34",x"03",x"C3",x"45",x"34",x"DD",x"36",x"0D",x"02",x"DD",x"36",x"03",x"80",
		x"C3",x"9A",x"34",x"DD",x"35",x"03",x"C3",x"45",x"34",x"3A",x"27",x"62",x"FE",x"03",x"C8",x"3A",
		x"03",x"62",x"CB",x"7F",x"C2",x"ED",x"34",x"21",x"C4",x"3A",x"06",x"00",x"3A",x"19",x"60",x"E6",
		x"06",x"4F",x"09",x"7E",x"DD",x"77",x"03",x"DD",x"77",x"0E",x"23",x"7E",x"DD",x"77",x"05",x"DD",
		x"77",x"0F",x"AF",x"DD",x"77",x"0D",x"DD",x"77",x"18",x"DD",x"77",x"1C",x"C9",x"21",x"D4",x"3A",
		x"C3",x"CA",x"34",x"21",x"00",x"64",x"11",x"D0",x"69",x"06",x"05",x"7E",x"A7",x"CA",x"1E",x"35",
		x"2C",x"2C",x"2C",x"7E",x"12",x"3E",x"04",x"85",x"6F",x"1C",x"7E",x"12",x"2C",x"1C",x"7E",x"12",
		x"2D",x"2D",x"2D",x"1C",x"7E",x"12",x"13",x"3E",x"1B",x"85",x"6F",x"10",x"DE",x"C9",x"3E",x"05",
		x"85",x"6F",x"3E",x"04",x"83",x"5F",x"C3",x"17",x"35",x"00",x"00",x"00",x"00",x"01",x"00",x"00",
		x"02",x"00",x"00",x"03",x"00",x"00",x"04",x"00",x"00",x"05",x"00",x"00",x"06",x"00",x"00",x"07",
		x"00",x"00",x"08",x"00",x"00",x"09",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",
		x"00",x"30",x"00",x"00",x"40",x"00",x"00",x"50",x"00",x"00",x"60",x"00",x"00",x"70",x"00",x"00",
		x"80",x"00",x"00",x"90",x"00",x"94",x"77",x"01",x"23",x"24",x"10",x"10",x"00",x"00",x"07",x"06",
		x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3F",x"00",x"50",x"76",x"00",x"F4",x"76",x"96",x"77",x"02",x"1E",x"14",x"10",x"10",x"00",x"00",
		x"06",x"01",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"3F",x"00",x"00",x"61",x"00",x"F6",x"76",x"98",x"77",x"03",x"22",x"14",x"10",x"10",
		x"00",x"00",x"05",x"09",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"59",x"00",x"F8",x"76",x"9A",x"77",x"04",x"24",x"18",
		x"10",x"10",x"00",x"00",x"05",x"00",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"50",x"00",x"FA",x"76",x"9C",x"77",x"05",
		x"24",x"18",x"10",x"10",x"00",x"00",x"04",x"03",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"00",x"43",x"00",x"FC",x"76",x"3B",
		x"5C",x"4B",x"5C",x"5B",x"5C",x"6B",x"5C",x"7B",x"5C",x"8B",x"5C",x"9B",x"5C",x"AB",x"5C",x"BB",
		x"5C",x"CB",x"5C",x"3B",x"6C",x"4B",x"6C",x"5B",x"6C",x"6B",x"6C",x"7B",x"6C",x"8B",x"6C",x"9B",
		x"6C",x"AB",x"6C",x"BB",x"6C",x"CB",x"6C",x"3B",x"7C",x"4B",x"7C",x"5B",x"7C",x"6B",x"7C",x"7B",
		x"7C",x"8B",x"7C",x"9B",x"7C",x"AB",x"7C",x"BB",x"7C",x"CB",x"7C",x"8B",x"36",x"01",x"00",x"98",
		x"36",x"A5",x"36",x"B2",x"36",x"BF",x"36",x"06",x"00",x"CC",x"36",x"08",x"00",x"E6",x"36",x"FD",
		x"36",x"0B",x"00",x"15",x"37",x"1C",x"37",x"30",x"37",x"38",x"37",x"47",x"37",x"5D",x"37",x"73",
		x"37",x"8B",x"37",x"00",x"61",x"22",x"61",x"44",x"61",x"66",x"61",x"88",x"61",x"9E",x"37",x"B6",
		x"37",x"D2",x"37",x"E1",x"37",x"1D",x"00",x"00",x"3F",x"09",x"3F",x"96",x"76",x"17",x"11",x"1D",
		x"15",x"10",x"10",x"1F",x"26",x"15",x"22",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",
		x"10",x"30",x"32",x"31",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"30",x"33",
		x"31",x"3F",x"80",x"76",x"18",x"19",x"17",x"18",x"10",x"23",x"13",x"1F",x"22",x"15",x"3F",x"9F",
		x"75",x"13",x"22",x"15",x"14",x"19",x"24",x"10",x"10",x"10",x"10",x"3F",x"5E",x"77",x"18",x"1F",
		x"27",x"10",x"18",x"19",x"17",x"18",x"10",x"13",x"11",x"1E",x"10",x"29",x"1F",x"25",x"10",x"17",
		x"15",x"24",x"10",x"FB",x"10",x"3F",x"29",x"77",x"1F",x"1E",x"1C",x"29",x"10",x"01",x"10",x"20",
		x"1C",x"11",x"29",x"15",x"22",x"10",x"12",x"25",x"24",x"24",x"1F",x"1E",x"3F",x"29",x"77",x"01",
		x"10",x"1F",x"22",x"10",x"02",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"23",x"10",x"12",x"25",
		x"24",x"24",x"1F",x"1E",x"3F",x"27",x"76",x"20",x"25",x"23",x"18",x"3F",x"06",x"77",x"1E",x"11",
		x"1D",x"15",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"22",x"11",x"24",x"19",x"1F",x"1E",x"3F",
		x"88",x"76",x"1E",x"11",x"1D",x"15",x"2E",x"3F",x"E9",x"75",x"2D",x"2D",x"2D",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"0B",x"77",x"11",x"10",x"12",x"10",x"13",x"10",x"14",
		x"10",x"15",x"10",x"16",x"10",x"17",x"10",x"18",x"10",x"19",x"10",x"1A",x"3F",x"0D",x"77",x"1B",
		x"10",x"1C",x"10",x"1D",x"10",x"1E",x"10",x"1F",x"10",x"20",x"10",x"21",x"10",x"22",x"10",x"23",
		x"10",x"24",x"3F",x"0F",x"77",x"25",x"10",x"26",x"10",x"27",x"10",x"28",x"10",x"29",x"10",x"2A",
		x"10",x"2B",x"10",x"2C",x"44",x"45",x"46",x"47",x"48",x"10",x"3F",x"F2",x"76",x"22",x"15",x"17",
		x"19",x"10",x"24",x"19",x"1D",x"15",x"10",x"10",x"30",x"03",x"00",x"31",x"10",x"3F",x"92",x"77",
		x"22",x"11",x"1E",x"1B",x"10",x"10",x"23",x"13",x"1F",x"22",x"15",x"10",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"10",x"10",x"10",x"3F",x"72",x"77",x"29",x"1F",x"25",x"22",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"27",x"11",x"23",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"15",x"22",x"15",x"14",
		x"42",x"3F",x"A7",x"76",x"19",x"1E",x"23",x"15",x"22",x"24",x"10",x"13",x"1F",x"19",x"1E",x"10",
		x"3F",x"0A",x"77",x"10",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"10",x"10",x"10",x"13",
		x"1F",x"19",x"1E",x"3F",x"FC",x"76",x"49",x"4A",x"10",x"1E",x"19",x"1E",x"24",x"15",x"1E",x"14",
		x"1F",x"10",x"10",x"10",x"10",x"3F",x"7C",x"75",x"01",x"09",x"08",x"01",x"3F",x"02",x"97",x"38",
		x"68",x"38",x"02",x"DF",x"54",x"10",x"54",x"02",x"EF",x"6D",x"20",x"6D",x"02",x"DF",x"8E",x"10",
		x"8E",x"02",x"EF",x"AF",x"20",x"AF",x"02",x"DF",x"D0",x"10",x"D0",x"02",x"EF",x"F1",x"10",x"F1",
		x"00",x"53",x"18",x"53",x"54",x"00",x"63",x"18",x"63",x"54",x"00",x"93",x"38",x"93",x"54",x"00",
		x"83",x"54",x"83",x"F1",x"00",x"93",x"54",x"93",x"F1",x"AA",x"8D",x"7D",x"8C",x"6F",x"00",x"7C",
		x"6E",x"00",x"7C",x"6D",x"00",x"7C",x"6C",x"00",x"7C",x"8F",x"7F",x"8E",x"47",x"27",x"08",x"50",
		x"2F",x"A7",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"23",x"07",x"40",
		x"46",x"A9",x"08",x"44",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",x"70",x"08",x"48",
		x"00",x"70",x"0A",x"48",x"6F",x"10",x"09",x"23",x"6F",x"11",x"0A",x"33",x"50",x"34",x"08",x"3C",
		x"00",x"35",x"08",x"3C",x"53",x"32",x"08",x"40",x"63",x"33",x"08",x"40",x"00",x"70",x"08",x"48",
		x"53",x"36",x"08",x"50",x"63",x"37",x"08",x"50",x"6B",x"31",x"08",x"41",x"00",x"70",x"08",x"48",
		x"6A",x"14",x"0A",x"48",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"7F",x"04",x"7F",x"F0",x"10",
		x"F0",x"02",x"DF",x"F2",x"70",x"F8",x"02",x"6F",x"F8",x"10",x"F8",x"AA",x"04",x"DF",x"D0",x"90",
		x"D0",x"02",x"DF",x"DC",x"20",x"D1",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"04",x"DF",x"A8",x"20",
		x"A8",x"04",x"5F",x"B0",x"20",x"B0",x"02",x"DF",x"B0",x"20",x"BB",x"AA",x"04",x"DF",x"88",x"30",
		x"88",x"04",x"DF",x"90",x"B0",x"90",x"02",x"DF",x"9A",x"20",x"8F",x"AA",x"04",x"BF",x"68",x"20",
		x"68",x"04",x"3F",x"70",x"20",x"70",x"02",x"DF",x"6E",x"20",x"79",x"AA",x"02",x"DF",x"58",x"A0",
		x"55",x"AA",x"00",x"70",x"08",x"44",x"2B",x"AC",x"08",x"4C",x"3B",x"AE",x"08",x"4C",x"3B",x"AF",
		x"08",x"3C",x"4B",x"B0",x"07",x"3C",x"4B",x"AD",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"47",x"27",x"08",x"4C",x"2F",x"A7",
		x"08",x"4C",x"3B",x"25",x"08",x"4C",x"00",x"70",x"08",x"44",x"3B",x"23",x"07",x"3C",x"4B",x"2A",
		x"08",x"3C",x"4B",x"2B",x"08",x"4C",x"2B",x"AA",x"08",x"3C",x"2B",x"AB",x"08",x"4C",x"00",x"70",
		x"0A",x"44",x"00",x"70",x"08",x"44",x"4B",x"2C",x"08",x"4C",x"3B",x"2E",x"08",x"4C",x"3B",x"2F",
		x"08",x"3C",x"2B",x"30",x"07",x"3C",x"2B",x"2D",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"02",x"02",x"02",x"02",x"03",
		x"03",x"03",x"7F",x"1E",x"4E",x"BB",x"4C",x"D8",x"4E",x"59",x"4E",x"7F",x"BB",x"4D",x"7F",x"47",
		x"27",x"08",x"50",x"2D",x"26",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",
		x"24",x"07",x"40",x"4B",x"28",x"08",x"40",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",
		x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"49",x"A6",x"08",x"50",x"2F",x"A7",x"08",x"50",x"3B",
		x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"24",x"07",x"40",x"46",x"A9",x"08",x"44",x"00",
		x"70",x"08",x"48",x"2B",x"A8",x"08",x"40",x"00",x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"73",
		x"A7",x"88",x"60",x"8B",x"27",x"88",x"60",x"7F",x"25",x"88",x"60",x"00",x"70",x"88",x"68",x"7F",
		x"24",x"87",x"70",x"74",x"29",x"88",x"6C",x"00",x"70",x"88",x"68",x"8A",x"A9",x"88",x"6C",x"00",
		x"70",x"88",x"68",x"00",x"70",x"8A",x"68",x"05",x"AF",x"F0",x"50",x"F0",x"AA",x"05",x"AF",x"E8",
		x"50",x"E8",x"AA",x"05",x"AF",x"E0",x"50",x"E0",x"AA",x"05",x"AF",x"D8",x"50",x"D8",x"AA",x"05",
		x"B7",x"58",x"48",x"58",x"AA",x"01",x"04",x"01",x"03",x"04",x"01",x"02",x"03",x"04",x"01",x"02",
		x"01",x"03",x"04",x"01",x"02",x"01",x"03",x"01",x"04",x"7F",x"FF",x"00",x"FF",x"FF",x"FE",x"FE",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"00",x"E8",x"E5",x"E3",x"E2",
		x"E1",x"E0",x"DF",x"DE",x"DD",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DE",x"DF",
		x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E7",x"E9",x"EB",x"ED",x"F0",x"AA",x"80",x"7B",x"78",x"76",
		x"74",x"73",x"72",x"71",x"70",x"70",x"6F",x"6F",x"6F",x"70",x"70",x"71",x"72",x"73",x"74",x"75",
		x"76",x"77",x"78",x"AA",x"EE",x"F0",x"DB",x"A0",x"E6",x"C8",x"D6",x"78",x"EB",x"F0",x"DB",x"A0",
		x"E6",x"C8",x"E6",x"C8",x"1B",x"C8",x"23",x"A0",x"2B",x"78",x"12",x"F0",x"1B",x"C8",x"23",x"A0",
		x"12",x"F0",x"1B",x"C8",x"02",x"97",x"38",x"68",x"38",x"02",x"9F",x"54",x"10",x"54",x"02",x"DF",
		x"58",x"A0",x"55",x"02",x"EF",x"6D",x"20",x"79",x"02",x"DF",x"9A",x"10",x"8E",x"02",x"EF",x"AF",
		x"20",x"BB",x"02",x"DF",x"DC",x"10",x"D0",x"02",x"FF",x"F0",x"80",x"F7",x"02",x"7F",x"F8",x"00",
		x"F8",x"00",x"CB",x"57",x"CB",x"6F",x"00",x"CB",x"99",x"CB",x"B1",x"00",x"CB",x"DB",x"CB",x"F3",
		x"00",x"63",x"18",x"63",x"54",x"01",x"63",x"D5",x"63",x"F8",x"00",x"33",x"78",x"33",x"90",x"00",
		x"33",x"BA",x"33",x"D2",x"00",x"53",x"18",x"53",x"54",x"01",x"53",x"92",x"53",x"B8",x"00",x"5B",
		x"76",x"5B",x"92",x"00",x"73",x"B6",x"73",x"D6",x"00",x"83",x"95",x"83",x"B5",x"00",x"93",x"38",
		x"93",x"54",x"01",x"BB",x"70",x"BB",x"98",x"01",x"6B",x"54",x"6B",x"75",x"AA",x"06",x"8F",x"90",
		x"70",x"90",x"06",x"8F",x"98",x"70",x"98",x"06",x"8F",x"A0",x"70",x"A0",x"00",x"63",x"18",x"63",
		x"58",x"00",x"63",x"80",x"63",x"A8",x"00",x"63",x"D0",x"63",x"F8",x"00",x"53",x"18",x"53",x"58",
		x"00",x"53",x"A8",x"53",x"D0",x"00",x"9B",x"80",x"9B",x"A8",x"00",x"9B",x"D0",x"9B",x"F8",x"01",
		x"23",x"58",x"23",x"80",x"01",x"DB",x"58",x"DB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"A3",x"A8",x"A3",x"D0",x"00",x"2B",x"D0",x"2B",x"F8",x"00",x"D3",x"D0",
		x"D3",x"F8",x"00",x"93",x"38",x"93",x"58",x"02",x"97",x"38",x"68",x"38",x"03",x"EF",x"58",x"10",
		x"58",x"03",x"F7",x"80",x"88",x"80",x"03",x"77",x"80",x"08",x"80",x"02",x"A7",x"A8",x"50",x"A8",
		x"02",x"E7",x"A8",x"B8",x"A8",x"02",x"3F",x"A8",x"18",x"A8",x"03",x"EF",x"D0",x"10",x"D0",x"02",
		x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"63",x"18",x"63",x"58",x"00",x"63",x"88",x"63",x"D0",x"00",
		x"53",x"18",x"53",x"58",x"00",x"53",x"88",x"53",x"D0",x"00",x"E3",x"68",x"E3",x"90",x"00",x"E3",
		x"B8",x"E3",x"D0",x"00",x"CB",x"90",x"CB",x"B0",x"00",x"B3",x"58",x"B3",x"78",x"00",x"9B",x"80",
		x"9B",x"A0",x"00",x"93",x"38",x"93",x"58",x"00",x"23",x"88",x"23",x"C0",x"00",x"1B",x"C0",x"1B",
		x"E8",x"02",x"97",x"38",x"68",x"38",x"02",x"B7",x"58",x"10",x"58",x"02",x"EF",x"68",x"E0",x"68",
		x"02",x"D7",x"70",x"C8",x"70",x"02",x"BF",x"78",x"B0",x"78",x"02",x"A7",x"80",x"90",x"80",x"02",
		x"67",x"88",x"48",x"88",x"02",x"27",x"88",x"10",x"88",x"02",x"EF",x"90",x"C8",x"90",x"02",x"A7",
		x"A0",x"98",x"A0",x"02",x"BF",x"A8",x"B0",x"A8",x"02",x"D7",x"B0",x"C8",x"B0",x"02",x"EF",x"B8",
		x"E0",x"B8",x"02",x"27",x"C0",x"10",x"C0",x"02",x"EF",x"D0",x"D8",x"D0",x"02",x"67",x"D0",x"50",
		x"D0",x"02",x"CF",x"D8",x"C0",x"D8",x"02",x"B7",x"E0",x"A8",x"E0",x"02",x"9F",x"E8",x"88",x"E8",
		x"02",x"27",x"E8",x"10",x"E8",x"02",x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"7B",x"80",x"7B",x"A8",
		x"00",x"7B",x"D0",x"7B",x"F8",x"00",x"33",x"58",x"33",x"80",x"00",x"53",x"58",x"53",x"80",x"00",
		x"AB",x"58",x"AB",x"80",x"00",x"CB",x"58",x"CB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"23",x"A8",x"23",x"D0",x"00",x"5B",x"A8",x"5B",x"D0",x"00",x"A3",x"A8",
		x"A3",x"D0",x"00",x"DB",x"A8",x"DB",x"D0",x"00",x"1B",x"D0",x"1B",x"F8",x"00",x"E3",x"D0",x"E3",
		x"F8",x"05",x"B7",x"30",x"48",x"30",x"05",x"CF",x"58",x"30",x"58",x"05",x"D7",x"80",x"28",x"80",
		x"05",x"DF",x"A8",x"20",x"A8",x"05",x"E7",x"D0",x"18",x"D0",x"05",x"EF",x"F8",x"10",x"F8",x"AA",
		x"10",x"82",x"85",x"8B",x"10",x"85",x"80",x"8B",x"10",x"87",x"85",x"8B",x"81",x"80",x"80",x"8B",
		x"81",x"82",x"85",x"8B",x"81",x"85",x"80",x"8B",x"05",x"88",x"77",x"01",x"68",x"77",x"01",x"6C",
		x"77",x"03",x"49",x"77",x"05",x"08",x"77",x"01",x"E8",x"76",x"01",x"EC",x"76",x"05",x"C8",x"76",
		x"05",x"88",x"76",x"02",x"69",x"76",x"02",x"4A",x"76",x"05",x"28",x"76",x"05",x"E8",x"75",x"01",
		x"CA",x"75",x"03",x"A9",x"75",x"01",x"88",x"75",x"01",x"8C",x"75",x"05",x"48",x"75",x"01",x"28",
		x"75",x"01",x"2A",x"75",x"01",x"2C",x"75",x"01",x"08",x"75",x"01",x"0A",x"75",x"01",x"0C",x"75",
		x"03",x"C8",x"74",x"03",x"AA",x"74",x"03",x"88",x"74",x"05",x"2F",x"77",x"05",x"0F",x"77",x"02",
		x"F0",x"76",x"02",x"CF",x"76",x"02",x"D2",x"76",x"05",x"8F",x"76",x"05",x"6F",x"76",x"01",x"4F",
		x"76",x"01",x"53",x"76",x"05",x"2F",x"76",x"05",x"EF",x"75",x"02",x"D0",x"75",x"02",x"B1",x"75",
		x"05",x"8F",x"75",x"03",x"50",x"75",x"05",x"2F",x"75",x"01",x"0F",x"75",x"01",x"13",x"75",x"01",
		x"EF",x"74",x"01",x"F1",x"74",x"01",x"F3",x"74",x"02",x"D1",x"74",x"00",x"00",x"00",x"23",x"68",
		x"01",x"11",x"00",x"00",x"00",x"10",x"DB",x"68",x"01",x"40",x"00",x"00",x"08",x"01",x"01",x"01",
		x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"01",x"C0",x"FF",
		x"01",x"FF",x"FF",x"34",x"C3",x"39",x"00",x"67",x"80",x"69",x"1A",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"0B",x"4B",
		x"14",x"18",x"0B",x"4B",x"1E",x"18",x"0B",x"3B",x"14",x"18",x"0B",x"3B",x"3D",x"01",x"03",x"02",
		x"4D",x"01",x"04",x"01",x"27",x"70",x"01",x"E0",x"00",x"00",x"7F",x"40",x"01",x"78",x"02",x"00",
		x"27",x"49",x"0C",x"F0",x"7F",x"49",x"0C",x"88",x"1E",x"07",x"03",x"09",x"24",x"64",x"BB",x"C0",
		x"23",x"8D",x"7B",x"B4",x"1B",x"8C",x"7C",x"64",x"4B",x"0E",x"04",x"02",x"23",x"46",x"03",x"68",
		x"DB",x"46",x"03",x"68",x"17",x"50",x"00",x"5C",x"E7",x"D0",x"00",x"5C",x"8C",x"50",x"00",x"84",
		x"73",x"D0",x"00",x"84",x"17",x"50",x"00",x"D4",x"E7",x"D0",x"00",x"D4",x"53",x"73",x"0A",x"A0",
		x"8B",x"74",x"0A",x"F0",x"DB",x"75",x"0A",x"A0",x"5B",x"73",x"0A",x"C8",x"E3",x"74",x"0A",x"60",
		x"1B",x"75",x"0A",x"80",x"DB",x"73",x"0A",x"C8",x"93",x"74",x"0A",x"F0",x"33",x"75",x"0A",x"50",
		x"44",x"03",x"08",x"04",x"37",x"F4",x"37",x"C0",x"37",x"8C",x"77",x"70",x"77",x"A4",x"77",x"D8",
		x"11",x"01",x"00",x"06",x"7B",x"1F",x"D2",x"28",x"1E",x"1E",x"03",x"06",x"7D",x"1F",x"D2",x"28",
		x"1E",x"1E",x"05",x"06",x"7F",x"C3",x"28",x"1E",x"3A",x"27",x"62",x"E5",x"EF",x"00",x"00",x"99",
		x"3E",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",x"E1",x"AF",x"32",x"60",x"60",x"06",x"0A",
		x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"C3",x"3E",x"06",x"05",x"DD",x"21",x"00",x"64",
		x"CD",x"C3",x"3E",x"3A",x"60",x"60",x"A7",x"C8",x"FE",x"01",x"C8",x"FE",x"03",x"3E",x"03",x"D8",
		x"3E",x"07",x"C9",x"DD",x"CB",x"00",x"46",x"CA",x"FA",x"3E",x"79",x"DD",x"96",x"05",x"D2",x"D3",
		x"3E",x"ED",x"44",x"3C",x"95",x"DA",x"DE",x"3E",x"DD",x"96",x"0A",x"D2",x"FA",x"3E",x"FD",x"7E",
		x"03",x"DD",x"96",x"03",x"D2",x"E9",x"3E",x"ED",x"44",x"94",x"DA",x"F3",x"3E",x"DD",x"96",x"09",
		x"D2",x"FA",x"3E",x"3A",x"60",x"60",x"3C",x"32",x"60",x"60",x"DD",x"19",x"10",x"C5",x"C9",x"00",
		x"5C",x"76",x"49",x"4A",x"01",x"09",x"08",x"01",x"3F",x"7D",x"77",x"1E",x"19",x"1E",x"24",x"15",
		x"1E",x"14",x"1F",x"10",x"1F",x"16",x"10",x"11",x"1D",x"15",x"22",x"19",x"13",x"11",x"10",x"19",
		x"1E",x"13",x"2B",x"3F",x"21",x"AF",x"74",x"11",x"E0",x"FF",x"36",x"9F",x"19",x"36",x"9E",x"C9",
		x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"2C",x"57",x"45",x"20",x"57",x"4F",x"55",x"4C",x"44",
		x"20",x"54",x"45",x"41",x"43",x"48",x"20",x"59",x"4F",x"55",x"2E",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"54",x"45",x"4C",x"2E",x"54",x"4F",x"4B",x"59",x"4F",x"2D",x"4A",x"41",x"50",x"41",x"4E",x"20",
		x"30",x"34",x"34",x"28",x"32",x"34",x"34",x"29",x"32",x"31",x"35",x"31",x"20",x"20",x"20",x"20",
		x"45",x"58",x"54",x"45",x"4E",x"54",x"49",x"4F",x"4E",x"20",x"33",x"30",x"34",x"20",x"20",x"20",
		x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"44",x"45",x"53",x"49",x"47",x"4E",x"20",x"20",x"20",
		x"49",x"4B",x"45",x"47",x"41",x"4D",x"49",x"20",x"43",x"4F",x"2E",x"20",x"4C",x"49",x"4D",x"2E",
		x"CD",x"A6",x"3F",x"C3",x"5F",x"0D",x"3E",x"02",x"F7",x"06",x"02",x"21",x"6C",x"77",x"36",x"10",
		x"23",x"23",x"36",x"C0",x"21",x"8C",x"74",x"10",x"F5",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"4D",x"69",x"36",x"03",x"2C",x"2C",x"C9",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"7F",x"7F",x"18",x"3C",x"76",x"63",x"41",x"00",x"00",x"7F",x"7F",x"49",x"49",x"49",x"41",
		x"00",x"1C",x"3E",x"63",x"41",x"49",x"79",x"79",x"00",x"7C",x"7E",x"13",x"11",x"13",x"7E",x"7C",
		x"00",x"7F",x"7F",x"0E",x"1C",x"0E",x"7F",x"7F",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"17",x"CB",x"13",x"17",x"C6",x"74",x"57",x"19",x"C9",x"57",x"0F",x"DA",x"22",x"30",x"0E",x"93",
		x"0F",x"0F",x"D2",x"17",x"30",x"0E",x"6C",x"07",x"DA",x"31",x"30",x"79",x"E6",x"F0",x"4F",x"C3",
		x"31",x"30",x"0E",x"B4",x"0F",x"0F",x"D2",x"2B",x"30",x"0E",x"1E",x"CB",x"50",x"CA",x"31",x"30",
		x"05",x"79",x"0F",x"0F",x"4F",x"E6",x"03",x"B8",x"C2",x"31",x"30",x"79",x"0F",x"0F",x"E6",x"03",
		x"FE",x"03",x"C0",x"CB",x"92",x"15",x"C0",x"3E",x"04",x"C9",x"11",x"E0",x"FF",x"3A",x"8E",x"63",
		x"4F",x"06",x"00",x"21",x"00",x"76",x"CD",x"64",x"30",x"21",x"C0",x"75",x"CD",x"64",x"30",x"21",
		x"8E",x"63",x"35",x"C9",x"09",x"7E",x"19",x"77",x"C9",x"DF",x"2A",x"C0",x"63",x"34",x"C9",x"21",
		x"AF",x"62",x"34",x"7E",x"E6",x"07",x"C0",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"0E",x"81",x"21",
		x"09",x"69",x"CD",x"96",x"30",x"21",x"1D",x"69",x"CD",x"96",x"30",x"CD",x"57",x"00",x"E6",x"80",
		x"21",x"2D",x"69",x"AE",x"77",x"C9",x"06",x"02",x"79",x"AE",x"77",x"19",x"10",x"FA",x"C9",x"E5",
		x"21",x"C0",x"60",x"3A",x"B0",x"60",x"6F",x"CB",x"7E",x"CA",x"BB",x"30",x"72",x"2C",x"73",x"2C",
		x"7D",x"FE",x"C0",x"D2",x"B8",x"30",x"3E",x"C0",x"32",x"B0",x"60",x"E1",x"C9",x"21",x"50",x"69",
		x"06",x"02",x"CD",x"E4",x"30",x"2E",x"80",x"06",x"0A",x"CD",x"E4",x"30",x"2E",x"B8",x"06",x"0B",
		x"CD",x"E4",x"30",x"21",x"0C",x"6A",x"06",x"05",x"C3",x"E4",x"30",x"21",x"4C",x"69",x"36",x"00",
		x"2E",x"58",x"06",x"06",x"7D",x"36",x"00",x"C6",x"04",x"6F",x"10",x"F9",x"C9",x"CD",x"FA",x"30",
		x"CD",x"3C",x"31",x"CD",x"B1",x"31",x"CD",x"F3",x"34",x"C9",x"3A",x"80",x"63",x"FE",x"06",x"38",
		x"02",x"3E",x"05",x"EF",x"10",x"31",x"10",x"31",x"1B",x"31",x"26",x"31",x"26",x"31",x"31",x"31",
		x"3A",x"1A",x"60",x"E6",x"01",x"FE",x"01",x"C8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"07",
		x"FE",x"05",x"F8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"03",x"FE",x"03",x"F8",x"33",x"33",
		x"C9",x"3A",x"1A",x"60",x"E6",x"07",x"FE",x"07",x"F8",x"33",x"33",x"C9",x"DD",x"21",x"00",x"64",
		x"AF",x"32",x"A1",x"63",x"06",x"05",x"11",x"20",x"00",x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"7C",
		x"31",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"3E",x"01",x"DD",x"77",x"08",x"3A",x"17",x"62",
		x"FE",x"01",x"C2",x"6A",x"31",x"3E",x"00",x"DD",x"77",x"08",x"DD",x"19",x"10",x"DB",x"21",x"A0",
		x"63",x"36",x"00",x"3A",x"A1",x"63",x"FE",x"00",x"C0",x"33",x"33",x"C9",x"3A",x"A1",x"63",x"FE",
		x"05",x"CA",x"6A",x"31",x"3A",x"27",x"62",x"FE",x"02",x"C2",x"95",x"31",x"3A",x"A1",x"63",x"4F",
		x"3A",x"80",x"63",x"B9",x"C8",x"3A",x"A0",x"63",x"FE",x"01",x"C2",x"6A",x"31",x"DD",x"77",x"00",
		x"DD",x"77",x"18",x"AF",x"32",x"A0",x"63",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"C3",x"6A",
		x"31",x"CD",x"DD",x"31",x"AF",x"32",x"A2",x"63",x"21",x"E0",x"63",x"22",x"C8",x"63",x"2A",x"C8",
		x"63",x"01",x"20",x"00",x"09",x"22",x"C8",x"63",x"7E",x"A7",x"CA",x"D0",x"31",x"CD",x"02",x"32",
		x"3A",x"A2",x"63",x"3C",x"32",x"A2",x"63",x"FE",x"05",x"C2",x"BE",x"31",x"C9",x"3A",x"80",x"63",
		x"FE",x"03",x"F8",x"CD",x"F6",x"31",x"FE",x"01",x"C0",x"21",x"39",x"64",x"3E",x"02",x"77",x"21",
		x"79",x"64",x"3E",x"02",x"77",x"C9",x"3A",x"18",x"60",x"E6",x"03",x"FE",x"01",x"C0",x"3A",x"1A",
		x"60",x"C9",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"18",x"FE",x"01",x"CA",x"7A",x"32",x"DD",x"7E",
		x"0D",x"FE",x"04",x"F2",x"30",x"32",x"DD",x"7E",x"19",x"FE",x"02",x"CA",x"7E",x"32",x"CD",x"0F",
		x"33",x"3A",x"18",x"60",x"E6",x"03",x"C2",x"33",x"32",x"DD",x"7E",x"0D",x"A7",x"CA",x"57",x"32",
		x"CD",x"3D",x"33",x"DD",x"7E",x"0D",x"FE",x"04",x"F2",x"91",x"32",x"CD",x"AD",x"33",x"CD",x"8C",
		x"29",x"FE",x"01",x"CA",x"97",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0E",x"FE",x"10",x"DA",
		x"8C",x"32",x"FE",x"F0",x"D2",x"84",x"32",x"DD",x"7E",x"13",x"FE",x"00",x"C2",x"B9",x"32",x"3E",
		x"11",x"DD",x"77",x"13",x"16",x"00",x"5F",x"21",x"7A",x"3A",x"19",x"7E",x"DD",x"46",x"0E",x"DD",
		x"70",x"03",x"DD",x"4E",x"0F",x"81",x"DD",x"77",x"05",x"C9",x"CD",x"BD",x"32",x"C9",x"CD",x"D6",
		x"32",x"C3",x"29",x"32",x"3E",x"02",x"DD",x"77",x"0D",x"C3",x"57",x"32",x"3E",x"01",x"C3",x"86",
		x"32",x"CD",x"E7",x"33",x"C3",x"57",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0D",x"FE",x"01",
		x"C2",x"B1",x"32",x"3E",x"02",x"DD",x"35",x"0E",x"DD",x"77",x"0D",x"CD",x"C3",x"33",x"C3",x"57",
		x"32",x"3E",x"01",x"DD",x"34",x"0E",x"C3",x"A8",x"32",x"3D",x"C3",x"61",x"32",x"3A",x"27",x"62",
		x"FE",x"01",x"CA",x"CE",x"32",x"FE",x"02",x"CA",x"D2",x"32",x"CD",x"B9",x"34",x"C9",x"CD",x"2C",
		x"34",x"C9",x"CD",x"78",x"34",x"C9",x"DD",x"7E",x"1C",x"FE",x"00",x"C2",x"FD",x"32",x"DD",x"7E",
		x"1D",x"FE",x"01",x"C2",x"0B",x"33",x"DD",x"36",x"1D",x"00",x"3A",x"05",x"62",x"DD",x"46",x"0F",
		x"90",x"DA",x"03",x"33",x"DD",x"36",x"1C",x"FF",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"35",x"1C",
		x"C2",x"F8",x"32",x"DD",x"36",x"19",x"00",x"DD",x"36",x"1C",x"00",x"CD",x"0F",x"33",x"C9",x"DD",
		x"7E",x"16",x"FE",x"00",x"C2",x"32",x"33",x"DD",x"36",x"16",x"2B",x"DD",x"36",x"0D",x"00",x"3A",
		x"18",x"60",x"0F",x"D2",x"32",x"33",x"DD",x"7E",x"0D",x"FE",x"01",x"CA",x"36",x"33",x"DD",x"36",
		x"0D",x"01",x"DD",x"35",x"16",x"C9",x"DD",x"36",x"0D",x"02",x"C3",x"32",x"33",x"DD",x"7E",x"0D",
		x"FE",x"08",x"CA",x"71",x"33",x"FE",x"04",x"CA",x"8A",x"33",x"CD",x"A1",x"33",x"DD",x"7E",x"0F",
		x"C6",x"08",x"57",x"DD",x"7E",x"0E",x"01",x"15",x"00",x"CD",x"6E",x"23",x"A7",x"CA",x"99",x"33",
		x"DD",x"70",x"1F",x"3A",x"05",x"62",x"47",x"DD",x"7E",x"0F",x"90",x"D0",x"DD",x"36",x"0D",x"04",
		x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"DD",
		x"7E",x"19",x"FE",x"02",x"C0",x"DD",x"36",x"1D",x"01",x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",
		x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"70",x"1F",x"DD",x"36",x"0D",x"08",
		x"C9",x"3E",x"07",x"F7",x"DD",x"7E",x"0F",x"FE",x"59",x"D0",x"33",x"33",x"C9",x"DD",x"7E",x"0D",
		x"FE",x"01",x"CA",x"D9",x"33",x"DD",x"7E",x"07",x"E6",x"7F",x"DD",x"77",x"07",x"DD",x"35",x"0E",
		x"CD",x"09",x"34",x"3A",x"27",x"62",x"FE",x"01",x"C0",x"DD",x"66",x"0E",x"DD",x"6E",x"0F",x"DD",
		x"46",x"0D",x"CD",x"33",x"23",x"DD",x"75",x"0F",x"C9",x"DD",x"7E",x"07",x"F6",x"80",x"DD",x"77",
		x"07",x"DD",x"34",x"0E",x"C3",x"C0",x"33",x"CD",x"09",x"34",x"DD",x"7E",x"0D",x"FE",x"08",x"C2",
		x"05",x"34",x"DD",x"7E",x"14",x"A7",x"C2",x"01",x"34",x"DD",x"36",x"14",x"02",x"DD",x"35",x"0F",
		x"C9",x"DD",x"35",x"14",x"C9",x"DD",x"34",x"0F",x"C9",x"DD",x"7E",x"15",x"A7",x"C2",x"28",x"34",
		x"DD",x"36",x"15",x"02",x"DD",x"34",x"07",x"DD",x"7E",x"07",x"E6",x"0F",x"FE",x"0F",x"C0",x"DD",
		x"7E",x"07",x"EE",x"02",x"DD",x"77",x"07",x"C9",x"DD",x"35",x"15",x"C9",x"DD",x"6E",x"1A",x"DD",
		x"66",x"1B",x"AF",x"01",x"00",x"00",x"ED",x"4A",x"C2",x"42",x"34",x"21",x"8C",x"3A",x"DD",x"36",
		x"03",x"26",x"DD",x"34",x"03",x"7E",x"FE",x"AA",x"CA",x"56",x"34",x"DD",x"77",x"05",x"23",x"DD",
		x"75",x"1A",x"DD",x"74",x"1B",x"C9",x"AF",x"DD",x"77",x"13",x"DD",x"77",x"18",x"DD",x"77",x"0D",
		x"DD",x"77",x"1C",x"DD",x"7E",x"03",x"DD",x"77",x"0E",x"DD",x"7E",x"05",x"DD",x"77",x"0F",x"DD",
		x"36",x"1A",x"00",x"DD",x"36",x"1B",x"00",x"C9",x"DD",x"6E",x"1A",x"DD",x"66",x"1B",x"AF",x"01",
		x"00",x"00",x"ED",x"4A",x"C2",x"9A",x"34",x"21",x"AC",x"3A",x"3A",x"03",x"62",x"CB",x"7F",x"CA",
		x"A8",x"34",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"03",x"7E",x"DD",x"7E",x"0D",x"FE",x"01",x"C2",
		x"B3",x"34",x"DD",x"34",x"03",x"C3",x"45",x"34",x"DD",x"36",x"0D",x"02",x"DD",x"36",x"03",x"80",
		x"C3",x"9A",x"34",x"DD",x"35",x"03",x"C3",x"45",x"34",x"3A",x"27",x"62",x"FE",x"03",x"C8",x"3A",
		x"03",x"62",x"CB",x"7F",x"C2",x"ED",x"34",x"21",x"C4",x"3A",x"06",x"00",x"3A",x"19",x"60",x"E6",
		x"06",x"4F",x"09",x"7E",x"DD",x"77",x"03",x"DD",x"77",x"0E",x"23",x"7E",x"DD",x"77",x"05",x"DD",
		x"77",x"0F",x"AF",x"DD",x"77",x"0D",x"DD",x"77",x"18",x"DD",x"77",x"1C",x"C9",x"21",x"D4",x"3A",
		x"C3",x"CA",x"34",x"21",x"00",x"64",x"11",x"D0",x"69",x"06",x"05",x"7E",x"A7",x"CA",x"1E",x"35",
		x"2C",x"2C",x"2C",x"7E",x"12",x"3E",x"04",x"85",x"6F",x"1C",x"7E",x"12",x"2C",x"1C",x"7E",x"12",
		x"2D",x"2D",x"2D",x"1C",x"7E",x"12",x"13",x"3E",x"1B",x"85",x"6F",x"10",x"DE",x"C9",x"3E",x"05",
		x"85",x"6F",x"3E",x"04",x"83",x"5F",x"C3",x"17",x"35",x"00",x"00",x"00",x"00",x"01",x"00",x"00",
		x"02",x"00",x"00",x"03",x"00",x"00",x"04",x"00",x"00",x"05",x"00",x"00",x"06",x"00",x"00",x"07",
		x"00",x"00",x"08",x"00",x"00",x"09",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",
		x"00",x"30",x"00",x"00",x"40",x"00",x"00",x"50",x"00",x"00",x"60",x"00",x"00",x"70",x"00",x"00",
		x"80",x"00",x"00",x"90",x"00",x"94",x"77",x"01",x"23",x"24",x"10",x"10",x"00",x"00",x"07",x"06",
		x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3F",x"00",x"50",x"76",x"00",x"F4",x"76",x"96",x"77",x"02",x"1E",x"14",x"10",x"10",x"00",x"00",
		x"06",x"01",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"3F",x"00",x"00",x"61",x"00",x"F6",x"76",x"98",x"77",x"03",x"22",x"14",x"10",x"10",
		x"00",x"00",x"05",x"09",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"59",x"00",x"F8",x"76",x"9A",x"77",x"04",x"24",x"18",
		x"10",x"10",x"00",x"00",x"05",x"00",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"50",x"00",x"FA",x"76",x"9C",x"77",x"05",
		x"24",x"18",x"10",x"10",x"00",x"00",x"04",x"03",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"00",x"43",x"00",x"FC",x"76",x"3B",
		x"5C",x"4B",x"5C",x"5B",x"5C",x"6B",x"5C",x"7B",x"5C",x"8B",x"5C",x"9B",x"5C",x"AB",x"5C",x"BB",
		x"5C",x"CB",x"5C",x"3B",x"6C",x"4B",x"6C",x"5B",x"6C",x"6B",x"6C",x"7B",x"6C",x"8B",x"6C",x"9B",
		x"6C",x"AB",x"6C",x"BB",x"6C",x"CB",x"6C",x"3B",x"7C",x"4B",x"7C",x"5B",x"7C",x"6B",x"7C",x"7B",
		x"7C",x"8B",x"7C",x"9B",x"7C",x"AB",x"7C",x"BB",x"7C",x"CB",x"7C",x"8B",x"36",x"01",x"00",x"98",
		x"36",x"A5",x"36",x"B2",x"36",x"BF",x"36",x"06",x"00",x"CC",x"36",x"08",x"00",x"E6",x"36",x"FD",
		x"36",x"0B",x"00",x"15",x"37",x"1C",x"37",x"30",x"37",x"38",x"37",x"47",x"37",x"5D",x"37",x"73",
		x"37",x"8B",x"37",x"00",x"61",x"22",x"61",x"44",x"61",x"66",x"61",x"88",x"61",x"9E",x"37",x"B6",
		x"37",x"D2",x"37",x"E1",x"37",x"1D",x"00",x"00",x"3F",x"09",x"3F",x"96",x"76",x"17",x"11",x"1D",
		x"15",x"10",x"10",x"1F",x"26",x"15",x"22",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",
		x"10",x"30",x"32",x"31",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"30",x"33",
		x"31",x"3F",x"80",x"76",x"18",x"19",x"17",x"18",x"10",x"23",x"13",x"1F",x"22",x"15",x"3F",x"9F",
		x"75",x"13",x"22",x"15",x"14",x"19",x"24",x"10",x"10",x"10",x"10",x"3F",x"5E",x"77",x"18",x"1F",
		x"27",x"10",x"18",x"19",x"17",x"18",x"10",x"13",x"11",x"1E",x"10",x"29",x"1F",x"25",x"10",x"17",
		x"15",x"24",x"10",x"FB",x"10",x"3F",x"29",x"77",x"1F",x"1E",x"1C",x"29",x"10",x"01",x"10",x"20",
		x"1C",x"11",x"29",x"15",x"22",x"10",x"12",x"25",x"24",x"24",x"1F",x"1E",x"3F",x"29",x"77",x"01",
		x"10",x"1F",x"22",x"10",x"02",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"23",x"10",x"12",x"25",
		x"24",x"24",x"1F",x"1E",x"3F",x"27",x"76",x"20",x"25",x"23",x"18",x"3F",x"06",x"77",x"1E",x"11",
		x"1D",x"15",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"22",x"11",x"24",x"19",x"1F",x"1E",x"3F",
		x"88",x"76",x"1E",x"11",x"1D",x"15",x"2E",x"3F",x"E9",x"75",x"2D",x"2D",x"2D",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"0B",x"77",x"11",x"10",x"12",x"10",x"13",x"10",x"14",
		x"10",x"15",x"10",x"16",x"10",x"17",x"10",x"18",x"10",x"19",x"10",x"1A",x"3F",x"0D",x"77",x"1B",
		x"10",x"1C",x"10",x"1D",x"10",x"1E",x"10",x"1F",x"10",x"20",x"10",x"21",x"10",x"22",x"10",x"23",
		x"10",x"24",x"3F",x"0F",x"77",x"25",x"10",x"26",x"10",x"27",x"10",x"28",x"10",x"29",x"10",x"2A",
		x"10",x"2B",x"10",x"2C",x"44",x"45",x"46",x"47",x"48",x"10",x"3F",x"F2",x"76",x"22",x"15",x"17",
		x"19",x"10",x"24",x"19",x"1D",x"15",x"10",x"10",x"30",x"03",x"00",x"31",x"10",x"3F",x"92",x"77",
		x"22",x"11",x"1E",x"1B",x"10",x"10",x"23",x"13",x"1F",x"22",x"15",x"10",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"10",x"10",x"10",x"3F",x"72",x"77",x"29",x"1F",x"25",x"22",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"27",x"11",x"23",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"15",x"22",x"15",x"14",
		x"42",x"3F",x"A7",x"76",x"19",x"1E",x"23",x"15",x"22",x"24",x"10",x"13",x"1F",x"19",x"1E",x"10",
		x"3F",x"0A",x"77",x"10",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"10",x"10",x"10",x"13",
		x"1F",x"19",x"1E",x"3F",x"FC",x"76",x"49",x"4A",x"10",x"1E",x"19",x"1E",x"24",x"15",x"1E",x"14",
		x"1F",x"10",x"10",x"10",x"10",x"3F",x"7C",x"75",x"01",x"09",x"08",x"01",x"3F",x"02",x"97",x"38",
		x"68",x"38",x"02",x"DF",x"54",x"10",x"54",x"02",x"EF",x"6D",x"20",x"6D",x"02",x"DF",x"8E",x"10",
		x"8E",x"02",x"EF",x"AF",x"20",x"AF",x"02",x"DF",x"D0",x"10",x"D0",x"02",x"EF",x"F1",x"10",x"F1",
		x"00",x"53",x"18",x"53",x"54",x"00",x"63",x"18",x"63",x"54",x"00",x"93",x"38",x"93",x"54",x"00",
		x"83",x"54",x"83",x"F1",x"00",x"93",x"54",x"93",x"F1",x"AA",x"8D",x"7D",x"8C",x"6F",x"00",x"7C",
		x"6E",x"00",x"7C",x"6D",x"00",x"7C",x"6C",x"00",x"7C",x"8F",x"7F",x"8E",x"47",x"27",x"08",x"50",
		x"2F",x"A7",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"23",x"07",x"40",
		x"46",x"A9",x"08",x"44",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",x"70",x"08",x"48",
		x"00",x"70",x"0A",x"48",x"6F",x"10",x"09",x"23",x"6F",x"11",x"0A",x"33",x"50",x"34",x"08",x"3C",
		x"00",x"35",x"08",x"3C",x"53",x"32",x"08",x"40",x"63",x"33",x"08",x"40",x"00",x"70",x"08",x"48",
		x"53",x"36",x"08",x"50",x"63",x"37",x"08",x"50",x"6B",x"31",x"08",x"41",x"00",x"70",x"08",x"48",
		x"6A",x"14",x"0A",x"48",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"7F",x"04",x"7F",x"F0",x"10",
		x"F0",x"02",x"DF",x"F2",x"70",x"F8",x"02",x"6F",x"F8",x"10",x"F8",x"AA",x"04",x"DF",x"D0",x"90",
		x"D0",x"02",x"DF",x"DC",x"20",x"D1",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"04",x"DF",x"A8",x"20",
		x"A8",x"04",x"5F",x"B0",x"20",x"B0",x"02",x"DF",x"B0",x"20",x"BB",x"AA",x"04",x"DF",x"88",x"30",
		x"88",x"04",x"DF",x"90",x"B0",x"90",x"02",x"DF",x"9A",x"20",x"8F",x"AA",x"04",x"BF",x"68",x"20",
		x"68",x"04",x"3F",x"70",x"20",x"70",x"02",x"DF",x"6E",x"20",x"79",x"AA",x"02",x"DF",x"58",x"A0",
		x"55",x"AA",x"00",x"70",x"08",x"44",x"2B",x"AC",x"08",x"4C",x"3B",x"AE",x"08",x"4C",x"3B",x"AF",
		x"08",x"3C",x"4B",x"B0",x"07",x"3C",x"4B",x"AD",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"47",x"27",x"08",x"4C",x"2F",x"A7",
		x"08",x"4C",x"3B",x"25",x"08",x"4C",x"00",x"70",x"08",x"44",x"3B",x"23",x"07",x"3C",x"4B",x"2A",
		x"08",x"3C",x"4B",x"2B",x"08",x"4C",x"2B",x"AA",x"08",x"3C",x"2B",x"AB",x"08",x"4C",x"00",x"70",
		x"0A",x"44",x"00",x"70",x"08",x"44",x"4B",x"2C",x"08",x"4C",x"3B",x"2E",x"08",x"4C",x"3B",x"2F",
		x"08",x"3C",x"2B",x"30",x"07",x"3C",x"2B",x"2D",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"02",x"02",x"02",x"02",x"03",
		x"03",x"03",x"7F",x"1E",x"4E",x"BB",x"4C",x"D8",x"4E",x"59",x"4E",x"7F",x"BB",x"4D",x"7F",x"47",
		x"27",x"08",x"50",x"2D",x"26",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",
		x"24",x"07",x"40",x"4B",x"28",x"08",x"40",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",
		x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"49",x"A6",x"08",x"50",x"2F",x"A7",x"08",x"50",x"3B",
		x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"24",x"07",x"40",x"46",x"A9",x"08",x"44",x"00",
		x"70",x"08",x"48",x"2B",x"A8",x"08",x"40",x"00",x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"73",
		x"A7",x"88",x"60",x"8B",x"27",x"88",x"60",x"7F",x"25",x"88",x"60",x"00",x"70",x"88",x"68",x"7F",
		x"24",x"87",x"70",x"74",x"29",x"88",x"6C",x"00",x"70",x"88",x"68",x"8A",x"A9",x"88",x"6C",x"00",
		x"70",x"88",x"68",x"00",x"70",x"8A",x"68",x"05",x"AF",x"F0",x"50",x"F0",x"AA",x"05",x"AF",x"E8",
		x"50",x"E8",x"AA",x"05",x"AF",x"E0",x"50",x"E0",x"AA",x"05",x"AF",x"D8",x"50",x"D8",x"AA",x"05",
		x"B7",x"58",x"48",x"58",x"AA",x"01",x"04",x"01",x"03",x"04",x"01",x"02",x"03",x"04",x"01",x"02",
		x"01",x"03",x"04",x"01",x"02",x"01",x"03",x"01",x"04",x"7F",x"FF",x"00",x"FF",x"FF",x"FE",x"FE",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"00",x"E8",x"E5",x"E3",x"E2",
		x"E1",x"E0",x"DF",x"DE",x"DD",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DE",x"DF",
		x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E7",x"E9",x"EB",x"ED",x"F0",x"AA",x"80",x"7B",x"78",x"76",
		x"74",x"73",x"72",x"71",x"70",x"70",x"6F",x"6F",x"6F",x"70",x"70",x"71",x"72",x"73",x"74",x"75",
		x"76",x"77",x"78",x"AA",x"EE",x"F0",x"DB",x"A0",x"E6",x"C8",x"D6",x"78",x"EB",x"F0",x"DB",x"A0",
		x"E6",x"C8",x"E6",x"C8",x"1B",x"C8",x"23",x"A0",x"2B",x"78",x"12",x"F0",x"1B",x"C8",x"23",x"A0",
		x"12",x"F0",x"1B",x"C8",x"02",x"97",x"38",x"68",x"38",x"02",x"9F",x"54",x"10",x"54",x"02",x"DF",
		x"58",x"A0",x"55",x"02",x"EF",x"6D",x"20",x"79",x"02",x"DF",x"9A",x"10",x"8E",x"02",x"EF",x"AF",
		x"20",x"BB",x"02",x"DF",x"DC",x"10",x"D0",x"02",x"FF",x"F0",x"80",x"F7",x"02",x"7F",x"F8",x"00",
		x"F8",x"00",x"CB",x"57",x"CB",x"6F",x"00",x"CB",x"99",x"CB",x"B1",x"00",x"CB",x"DB",x"CB",x"F3",
		x"00",x"63",x"18",x"63",x"54",x"01",x"63",x"D5",x"63",x"F8",x"00",x"33",x"78",x"33",x"90",x"00",
		x"33",x"BA",x"33",x"D2",x"00",x"53",x"18",x"53",x"54",x"01",x"53",x"92",x"53",x"B8",x"00",x"5B",
		x"76",x"5B",x"92",x"00",x"73",x"B6",x"73",x"D6",x"00",x"83",x"95",x"83",x"B5",x"00",x"93",x"38",
		x"93",x"54",x"01",x"BB",x"70",x"BB",x"98",x"01",x"6B",x"54",x"6B",x"75",x"AA",x"06",x"8F",x"90",
		x"70",x"90",x"06",x"8F",x"98",x"70",x"98",x"06",x"8F",x"A0",x"70",x"A0",x"00",x"63",x"18",x"63",
		x"58",x"00",x"63",x"80",x"63",x"A8",x"00",x"63",x"D0",x"63",x"F8",x"00",x"53",x"18",x"53",x"58",
		x"00",x"53",x"A8",x"53",x"D0",x"00",x"9B",x"80",x"9B",x"A8",x"00",x"9B",x"D0",x"9B",x"F8",x"01",
		x"23",x"58",x"23",x"80",x"01",x"DB",x"58",x"DB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"A3",x"A8",x"A3",x"D0",x"00",x"2B",x"D0",x"2B",x"F8",x"00",x"D3",x"D0",
		x"D3",x"F8",x"00",x"93",x"38",x"93",x"58",x"02",x"97",x"38",x"68",x"38",x"03",x"EF",x"58",x"10",
		x"58",x"03",x"F7",x"80",x"88",x"80",x"03",x"77",x"80",x"08",x"80",x"02",x"A7",x"A8",x"50",x"A8",
		x"02",x"E7",x"A8",x"B8",x"A8",x"02",x"3F",x"A8",x"18",x"A8",x"03",x"EF",x"D0",x"10",x"D0",x"02",
		x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"63",x"18",x"63",x"58",x"00",x"63",x"88",x"63",x"D0",x"00",
		x"53",x"18",x"53",x"58",x"00",x"53",x"88",x"53",x"D0",x"00",x"E3",x"68",x"E3",x"90",x"00",x"E3",
		x"B8",x"E3",x"D0",x"00",x"CB",x"90",x"CB",x"B0",x"00",x"B3",x"58",x"B3",x"78",x"00",x"9B",x"80",
		x"9B",x"A0",x"00",x"93",x"38",x"93",x"58",x"00",x"23",x"88",x"23",x"C0",x"00",x"1B",x"C0",x"1B",
		x"E8",x"02",x"97",x"38",x"68",x"38",x"02",x"B7",x"58",x"10",x"58",x"02",x"EF",x"68",x"E0",x"68",
		x"02",x"D7",x"70",x"C8",x"70",x"02",x"BF",x"78",x"B0",x"78",x"02",x"A7",x"80",x"90",x"80",x"02",
		x"67",x"88",x"48",x"88",x"02",x"27",x"88",x"10",x"88",x"02",x"EF",x"90",x"C8",x"90",x"02",x"A7",
		x"A0",x"98",x"A0",x"02",x"BF",x"A8",x"B0",x"A8",x"02",x"D7",x"B0",x"C8",x"B0",x"02",x"EF",x"B8",
		x"E0",x"B8",x"02",x"27",x"C0",x"10",x"C0",x"02",x"EF",x"D0",x"D8",x"D0",x"02",x"67",x"D0",x"50",
		x"D0",x"02",x"CF",x"D8",x"C0",x"D8",x"02",x"B7",x"E0",x"A8",x"E0",x"02",x"9F",x"E8",x"88",x"E8",
		x"02",x"27",x"E8",x"10",x"E8",x"02",x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"7B",x"80",x"7B",x"A8",
		x"00",x"7B",x"D0",x"7B",x"F8",x"00",x"33",x"58",x"33",x"80",x"00",x"53",x"58",x"53",x"80",x"00",
		x"AB",x"58",x"AB",x"80",x"00",x"CB",x"58",x"CB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"23",x"A8",x"23",x"D0",x"00",x"5B",x"A8",x"5B",x"D0",x"00",x"A3",x"A8",
		x"A3",x"D0",x"00",x"DB",x"A8",x"DB",x"D0",x"00",x"1B",x"D0",x"1B",x"F8",x"00",x"E3",x"D0",x"E3",
		x"F8",x"05",x"B7",x"30",x"48",x"30",x"05",x"CF",x"58",x"30",x"58",x"05",x"D7",x"80",x"28",x"80",
		x"05",x"DF",x"A8",x"20",x"A8",x"05",x"E7",x"D0",x"18",x"D0",x"05",x"EF",x"F8",x"10",x"F8",x"AA",
		x"10",x"82",x"85",x"8B",x"10",x"85",x"80",x"8B",x"10",x"87",x"85",x"8B",x"81",x"80",x"80",x"8B",
		x"81",x"82",x"85",x"8B",x"81",x"85",x"80",x"8B",x"05",x"88",x"77",x"01",x"68",x"77",x"01",x"6C",
		x"77",x"03",x"49",x"77",x"05",x"08",x"77",x"01",x"E8",x"76",x"01",x"EC",x"76",x"05",x"C8",x"76",
		x"05",x"88",x"76",x"02",x"69",x"76",x"02",x"4A",x"76",x"05",x"28",x"76",x"05",x"E8",x"75",x"01",
		x"CA",x"75",x"03",x"A9",x"75",x"01",x"88",x"75",x"01",x"8C",x"75",x"05",x"48",x"75",x"01",x"28",
		x"75",x"01",x"2A",x"75",x"01",x"2C",x"75",x"01",x"08",x"75",x"01",x"0A",x"75",x"01",x"0C",x"75",
		x"03",x"C8",x"74",x"03",x"AA",x"74",x"03",x"88",x"74",x"05",x"2F",x"77",x"05",x"0F",x"77",x"02",
		x"F0",x"76",x"02",x"CF",x"76",x"02",x"D2",x"76",x"05",x"8F",x"76",x"05",x"6F",x"76",x"01",x"4F",
		x"76",x"01",x"53",x"76",x"05",x"2F",x"76",x"05",x"EF",x"75",x"02",x"D0",x"75",x"02",x"B1",x"75",
		x"05",x"8F",x"75",x"03",x"50",x"75",x"05",x"2F",x"75",x"01",x"0F",x"75",x"01",x"13",x"75",x"01",
		x"EF",x"74",x"01",x"F1",x"74",x"01",x"F3",x"74",x"02",x"D1",x"74",x"00",x"00",x"00",x"23",x"68",
		x"01",x"11",x"00",x"00",x"00",x"10",x"DB",x"68",x"01",x"40",x"00",x"00",x"08",x"01",x"01",x"01",
		x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"01",x"C0",x"FF",
		x"01",x"FF",x"FF",x"34",x"C3",x"39",x"00",x"67",x"80",x"69",x"1A",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"0B",x"4B",
		x"14",x"18",x"0B",x"4B",x"1E",x"18",x"0B",x"3B",x"14",x"18",x"0B",x"3B",x"3D",x"01",x"03",x"02",
		x"4D",x"01",x"04",x"01",x"27",x"70",x"01",x"E0",x"00",x"00",x"7F",x"40",x"01",x"78",x"02",x"00",
		x"27",x"49",x"0C",x"F0",x"7F",x"49",x"0C",x"88",x"1E",x"07",x"03",x"09",x"24",x"64",x"BB",x"C0",
		x"23",x"8D",x"7B",x"B4",x"1B",x"8C",x"7C",x"64",x"4B",x"0E",x"04",x"02",x"23",x"46",x"03",x"68",
		x"DB",x"46",x"03",x"68",x"17",x"50",x"00",x"5C",x"E7",x"D0",x"00",x"5C",x"8C",x"50",x"00",x"84",
		x"73",x"D0",x"00",x"84",x"17",x"50",x"00",x"D4",x"E7",x"D0",x"00",x"D4",x"53",x"73",x"0A",x"A0",
		x"8B",x"74",x"0A",x"F0",x"DB",x"75",x"0A",x"A0",x"5B",x"73",x"0A",x"C8",x"E3",x"74",x"0A",x"60",
		x"1B",x"75",x"0A",x"80",x"DB",x"73",x"0A",x"C8",x"93",x"74",x"0A",x"F0",x"33",x"75",x"0A",x"50",
		x"44",x"03",x"08",x"04",x"37",x"F4",x"37",x"C0",x"37",x"8C",x"77",x"70",x"77",x"A4",x"77",x"D8",
		x"11",x"01",x"00",x"06",x"7B",x"1F",x"D2",x"28",x"1E",x"1E",x"03",x"06",x"7D",x"1F",x"D2",x"28",
		x"1E",x"1E",x"05",x"06",x"7F",x"C3",x"28",x"1E",x"3A",x"27",x"62",x"E5",x"EF",x"00",x"00",x"99",
		x"3E",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",x"E1",x"AF",x"32",x"60",x"60",x"06",x"0A",
		x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"C3",x"3E",x"06",x"05",x"DD",x"21",x"00",x"64",
		x"CD",x"C3",x"3E",x"3A",x"60",x"60",x"A7",x"C8",x"FE",x"01",x"C8",x"FE",x"03",x"3E",x"03",x"D8",
		x"3E",x"07",x"C9",x"DD",x"CB",x"00",x"46",x"CA",x"FA",x"3E",x"79",x"DD",x"96",x"05",x"D2",x"D3",
		x"3E",x"ED",x"44",x"3C",x"95",x"DA",x"DE",x"3E",x"DD",x"96",x"0A",x"D2",x"FA",x"3E",x"FD",x"7E",
		x"03",x"DD",x"96",x"03",x"D2",x"E9",x"3E",x"ED",x"44",x"94",x"DA",x"F3",x"3E",x"DD",x"96",x"09",
		x"D2",x"FA",x"3E",x"3A",x"60",x"60",x"3C",x"32",x"60",x"60",x"DD",x"19",x"10",x"C5",x"C9",x"00",
		x"5C",x"76",x"49",x"4A",x"01",x"09",x"08",x"01",x"3F",x"7D",x"77",x"1E",x"19",x"1E",x"24",x"15",
		x"1E",x"14",x"1F",x"10",x"1F",x"16",x"10",x"11",x"1D",x"15",x"22",x"19",x"13",x"11",x"10",x"19",
		x"1E",x"13",x"2B",x"3F",x"21",x"AF",x"74",x"11",x"E0",x"FF",x"36",x"9F",x"19",x"36",x"9E",x"C9",
		x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"2C",x"57",x"45",x"20",x"57",x"4F",x"55",x"4C",x"44",
		x"20",x"54",x"45",x"41",x"43",x"48",x"20",x"59",x"4F",x"55",x"2E",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"54",x"45",x"4C",x"2E",x"54",x"4F",x"4B",x"59",x"4F",x"2D",x"4A",x"41",x"50",x"41",x"4E",x"20",
		x"30",x"34",x"34",x"28",x"32",x"34",x"34",x"29",x"32",x"31",x"35",x"31",x"20",x"20",x"20",x"20",
		x"45",x"58",x"54",x"45",x"4E",x"54",x"49",x"4F",x"4E",x"20",x"33",x"30",x"34",x"20",x"20",x"20",
		x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"44",x"45",x"53",x"49",x"47",x"4E",x"20",x"20",x"20",
		x"49",x"4B",x"45",x"47",x"41",x"4D",x"49",x"20",x"43",x"4F",x"2E",x"20",x"4C",x"49",x"4D",x"2E",
		x"CD",x"A6",x"3F",x"C3",x"5F",x"0D",x"3E",x"02",x"F7",x"06",x"02",x"21",x"6C",x"77",x"36",x"10",
		x"23",x"23",x"36",x"C0",x"21",x"8C",x"74",x"10",x"F5",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"4D",x"69",x"36",x"03",x"2C",x"2C",x"C9",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"7F",x"7F",x"18",x"3C",x"76",x"63",x"41",x"00",x"00",x"7F",x"7F",x"49",x"49",x"49",x"41",
		x"00",x"1C",x"3E",x"63",x"41",x"49",x"79",x"79",x"00",x"7C",x"7E",x"13",x"11",x"13",x"7E",x"7C",
		x"00",x"7F",x"7F",x"0E",x"1C",x"0E",x"7F",x"7F",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00",
		x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",
		x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"00",x"00",x"00",x"00",x"28",x"00",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
		x"00",x"00",x"82",x"C6",x"6C",x"38",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"82",x"00",x"00",
		x"00",x"00",x"82",x"FE",x"FE",x"82",x"00",x"00",x"82",x"FE",x"FE",x"82",x"82",x"FE",x"FE",x"82",
		x"00",x"28",x"28",x"28",x"28",x"28",x"28",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"F6",x"F6",x"00",x"00",x"F6",x"F6",x"00",x"00",x"FA",x"FA",x"00",x"00",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"FA",x"FA",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",x"00",x"E0",x"C0",x"00",x"E0",x"C0",x"00",x"00",
		x"00",x"60",x"E0",x"00",x"60",x"E0",x"00",x"00",x"00",x"00",x"C0",x"00",x"C0",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",
		x"38",x"28",x"3E",x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3C",x"02",x"02",x"3C",x"00",x"0E",
		x"22",x"2A",x"3E",x"00",x"00",x"0E",x"3A",x"2A",x"22",x"3E",x"00",x"3E",x"08",x"10",x"3E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"A5",x"BD",x"81",x"42",x"3C",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"A5",x"FE",x"C2",x"82",x"BA",x"44",x"44",x"28",x"10",
		x"10",x"28",x"44",x"44",x"AA",x"BA",x"82",x"C2",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"A3",x"59",x"FD",x"FD",x"9D",x"8C",x"88",x"00",x"00",x"00",x"01",x"03",x"31",x"59",x"28",x"5C",
		x"00",x"00",x"00",x"00",x"80",x"78",x"FC",x"7F",x"00",x"00",x"07",x"0F",x"0E",x"09",x"07",x"00",
		x"40",x"A0",x"50",x"B0",x"D0",x"68",x"B8",x"50",x"3E",x"9E",x"AE",x"DA",x"CA",x"DE",x"CD",x"D1",
		x"3F",x"7B",x"F1",x"FB",x"7F",x"FF",x"FD",x"78",x"00",x"0C",x"1E",x"3F",x"3F",x"3E",x"3E",x"1C",
		x"B8",x"50",x"A8",x"50",x"B0",x"50",x"A0",x"40",x"D1",x"D1",x"CD",x"DE",x"DA",x"AA",x"BE",x"9E",
		x"7D",x"7F",x"FF",x"FE",x"7C",x"FE",x"7F",x"3F",x"1E",x"3C",x"3E",x"3E",x"3F",x"1E",x"0C",x"00",
		x"00",x"88",x"8C",x"9D",x"FD",x"FD",x"59",x"A3",x"AE",x"1C",x"6D",x"19",x"33",x"01",x"00",x"00",
		x"7F",x"FF",x"7E",x"BE",x"1C",x"00",x"00",x"00",x"00",x"07",x"09",x"0E",x"0F",x"07",x"00",x"00",
		x"45",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"3C",x"7E",x"52",x"4A",x"7E",x"3C",x"00",x"00",x"02",x"02",x"7E",x"7E",x"22",x"02",x"00",
		x"00",x"22",x"72",x"5A",x"4E",x"66",x"22",x"00",x"00",x"44",x"6E",x"7A",x"52",x"46",x"44",x"00",
		x"00",x"04",x"7E",x"7E",x"34",x"1C",x"0C",x"00",x"00",x"4C",x"5E",x"52",x"52",x"76",x"74",x"00",
		x"00",x"0C",x"5E",x"52",x"52",x"7E",x"3C",x"00",x"00",x"60",x"70",x"58",x"4E",x"46",x"40",x"00",
		x"00",x"2C",x"7E",x"52",x"52",x"7E",x"2C",x"00",x"00",x"38",x"7C",x"56",x"52",x"72",x"20",x"00",
		x"7E",x"7E",x"30",x"18",x"30",x"7E",x"7E",x"00",x"1E",x"20",x"20",x"1E",x"20",x"20",x"3E",x"00",
		x"00",x"00",x"C0",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"7F",x"80",x"80",x"80",x"00",x"00",
		x"20",x"20",x"20",x"20",x"C0",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"7F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3C",x"42",x"81",x"BD",x"B1",x"9D",x"B1",x"BD",x"81",x"A1",x"BD",x"BD",x"A1",x"81",x"42",x"3C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"7E",x"42",x"42",x"42",x"42",x"42",x"42",x"7E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"41",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"41",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"FF",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"FF",
		x"7F",x"44",x"44",x"44",x"44",x"44",x"44",x"7F",x"3F",x"24",x"24",x"24",x"24",x"24",x"24",x"3F",
		x"1F",x"14",x"14",x"14",x"14",x"14",x"14",x"1F",x"0F",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0F",
		x"07",x"04",x"04",x"04",x"04",x"04",x"04",x"07",x"83",x"82",x"82",x"82",x"82",x"82",x"82",x"83",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"A0",x"20",x"20",x"20",x"20",x"20",x"20",x"A0",
		x"D0",x"50",x"50",x"50",x"50",x"50",x"50",x"D0",x"E8",x"48",x"48",x"48",x"48",x"48",x"48",x"E8",
		x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"FA",x"42",x"42",x"42",x"42",x"42",x"42",x"FA",
		x"FD",x"45",x"45",x"45",x"45",x"45",x"45",x"FD",x"FE",x"44",x"44",x"44",x"44",x"44",x"44",x"FE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"00",x"FE",x"10",x"10",x"FF",x"FF",
		x"00",x"08",x"0C",x"FC",x"FC",x"00",x"A4",x"A6",x"00",x"C0",x"E8",x"00",x"40",x"A0",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"00",x"F0",x"40",x"40",x"E0",x"E0",
		x"00",x"04",x"04",x"FC",x"F8",x"00",x"A8",x"A8",x"E0",x"F8",x"7D",x"01",x"70",x"88",x"FE",x"FE",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"90",x"90",x"8A",x"80",x"40",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"81",x"00",x"00",x"18",x"18",x"00",x"00",x"81",x"24",x"6D",x"CF",x"EE",x"8E",x"DF",x"51",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00",
		x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",
		x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"00",x"00",x"00",x"00",x"28",x"00",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
		x"00",x"00",x"82",x"C6",x"6C",x"38",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"82",x"00",x"00",
		x"00",x"00",x"82",x"FE",x"FE",x"82",x"00",x"00",x"82",x"FE",x"FE",x"82",x"82",x"FE",x"FE",x"82",
		x"00",x"28",x"28",x"28",x"28",x"28",x"28",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"F6",x"F6",x"00",x"00",x"F6",x"F6",x"00",x"00",x"FA",x"FA",x"00",x"00",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"FA",x"FA",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",x"00",x"E0",x"C0",x"00",x"E0",x"C0",x"00",x"00",
		x"00",x"60",x"E0",x"00",x"60",x"E0",x"00",x"00",x"00",x"00",x"C0",x"00",x"C0",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",
		x"38",x"28",x"3E",x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3C",x"02",x"02",x"3C",x"00",x"0E",
		x"22",x"2A",x"3E",x"00",x"00",x"0E",x"3A",x"2A",x"22",x"3E",x"00",x"3E",x"08",x"10",x"3E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"A5",x"BD",x"81",x"42",x"3C",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"A5",x"FE",x"C2",x"82",x"BA",x"44",x"44",x"28",x"10",
		x"10",x"28",x"44",x"44",x"AA",x"BA",x"82",x"C2",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"A3",x"59",x"FD",x"FD",x"9D",x"8C",x"88",x"00",x"00",x"00",x"01",x"03",x"31",x"59",x"28",x"5C",
		x"00",x"00",x"00",x"00",x"80",x"78",x"FC",x"7F",x"00",x"00",x"07",x"0F",x"0E",x"09",x"07",x"00",
		x"40",x"A0",x"50",x"B0",x"D0",x"68",x"B8",x"50",x"3E",x"9E",x"AE",x"DA",x"CA",x"DE",x"CD",x"D1",
		x"3F",x"7B",x"F1",x"FB",x"7F",x"FF",x"FD",x"78",x"00",x"0C",x"1E",x"3F",x"3F",x"3E",x"3E",x"1C",
		x"B8",x"50",x"A8",x"50",x"B0",x"50",x"A0",x"40",x"D1",x"D1",x"CD",x"DE",x"DA",x"AA",x"BE",x"9E",
		x"7D",x"7F",x"FF",x"FE",x"7C",x"FE",x"7F",x"3F",x"1E",x"3C",x"3E",x"3E",x"3F",x"1E",x"0C",x"00",
		x"00",x"88",x"8C",x"9D",x"FD",x"FD",x"59",x"A3",x"AE",x"1C",x"6D",x"19",x"33",x"01",x"00",x"00",
		x"7F",x"FF",x"7E",x"BE",x"1C",x"00",x"00",x"00",x"00",x"07",x"09",x"0E",x"0F",x"07",x"00",x"00",
		x"45",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"3C",x"7E",x"52",x"4A",x"7E",x"3C",x"00",x"00",x"02",x"02",x"7E",x"7E",x"22",x"02",x"00",
		x"00",x"22",x"72",x"5A",x"4E",x"66",x"22",x"00",x"00",x"44",x"6E",x"7A",x"52",x"46",x"44",x"00",
		x"00",x"04",x"7E",x"7E",x"34",x"1C",x"0C",x"00",x"00",x"4C",x"5E",x"52",x"52",x"76",x"74",x"00",
		x"00",x"0C",x"5E",x"52",x"52",x"7E",x"3C",x"00",x"00",x"60",x"70",x"58",x"4E",x"46",x"40",x"00",
		x"00",x"2C",x"7E",x"52",x"52",x"7E",x"2C",x"00",x"00",x"38",x"7C",x"56",x"52",x"72",x"20",x"00",
		x"7E",x"7E",x"30",x"18",x"30",x"7E",x"7E",x"00",x"1E",x"20",x"20",x"1E",x"20",x"20",x"3E",x"00",
		x"00",x"00",x"C0",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"7F",x"80",x"80",x"80",x"00",x"00",
		x"20",x"20",x"20",x"20",x"C0",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"7F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3C",x"42",x"81",x"BD",x"B1",x"9D",x"B1",x"BD",x"81",x"A1",x"BD",x"BD",x"A1",x"81",x"42",x"3C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"7E",x"42",x"42",x"42",x"42",x"42",x"42",x"7E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"41",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"41",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"FF",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"FF",
		x"7F",x"44",x"44",x"44",x"44",x"44",x"44",x"7F",x"3F",x"24",x"24",x"24",x"24",x"24",x"24",x"3F",
		x"1F",x"14",x"14",x"14",x"14",x"14",x"14",x"1F",x"0F",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0F",
		x"07",x"04",x"04",x"04",x"04",x"04",x"04",x"07",x"83",x"82",x"82",x"82",x"82",x"82",x"82",x"83",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"A0",x"20",x"20",x"20",x"20",x"20",x"20",x"A0",
		x"D0",x"50",x"50",x"50",x"50",x"50",x"50",x"D0",x"E8",x"48",x"48",x"48",x"48",x"48",x"48",x"E8",
		x"F4",x"44",x"44",x"44",x"44",x"44",x"44",x"F4",x"FA",x"42",x"42",x"42",x"42",x"42",x"42",x"FA",
		x"FD",x"45",x"45",x"45",x"45",x"45",x"45",x"FD",x"FE",x"44",x"44",x"44",x"44",x"44",x"44",x"FE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"00",x"FE",x"10",x"10",x"FF",x"FF",
		x"00",x"08",x"0C",x"FC",x"FC",x"00",x"A4",x"A6",x"00",x"C0",x"E8",x"00",x"40",x"A0",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"00",x"F0",x"40",x"40",x"E0",x"E0",
		x"00",x"04",x"04",x"FC",x"F8",x"00",x"A8",x"A8",x"E0",x"F8",x"7D",x"01",x"70",x"88",x"FE",x"FE",
		x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"90",x"90",x"8A",x"80",x"40",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"81",x"00",x"00",x"18",x"18",x"00",x"00",x"81",x"24",x"6D",x"CF",x"EE",x"8E",x"DF",x"51",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00",
		x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",
		x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"00",x"00",x"00",x"00",x"28",x"00",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
		x"00",x"00",x"82",x"C6",x"6C",x"38",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"82",x"00",x"00",
		x"00",x"00",x"82",x"FE",x"FE",x"82",x"00",x"00",x"82",x"FE",x"FE",x"82",x"82",x"FE",x"FE",x"82",
		x"00",x"28",x"28",x"28",x"28",x"28",x"28",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"F6",x"F6",x"00",x"00",x"F6",x"F6",x"00",x"00",x"FA",x"FA",x"00",x"00",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"FA",x"FA",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",x"00",x"E0",x"C0",x"00",x"E0",x"C0",x"00",x"00",
		x"00",x"60",x"E0",x"00",x"60",x"E0",x"00",x"00",x"00",x"00",x"C0",x"00",x"C0",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",
		x"38",x"28",x"3E",x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3C",x"02",x"02",x"3C",x"00",x"0E",
		x"22",x"2A",x"3E",x"00",x"00",x"0E",x"3A",x"2A",x"22",x"3E",x"00",x"3E",x"08",x"10",x"3E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"A5",x"BD",x"81",x"42",x"3C",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"A5",x"7C",x"40",x"00",x"38",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"28",x"38",x"00",x"40",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"A2",x"00",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",
		x"00",x"01",x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",
		x"54",x"A6",x"02",x"02",x"62",x"73",x"77",x"FF",x"FF",x"8F",x"76",x"7C",x"4E",x"A6",x"D7",x"A3",
		x"FF",x"FF",x"FE",x"FD",x"7F",x"87",x"03",x"80",x"1F",x"3F",x"78",x"F0",x"F1",x"F6",x"F8",x"6F",
		x"BF",x"5F",x"AF",x"4F",x"2A",x"90",x"40",x"A8",x"C1",x"61",x"51",x"25",x"35",x"A1",x"B2",x"AE",
		x"CE",x"9A",x"31",x"3B",x"BF",x"3F",x"1D",x"08",x"1F",x"33",x"61",x"C0",x"C0",x"C7",x"C7",x"65",
		x"40",x"A8",x"50",x"AA",x"4F",x"AF",x"5F",x"BF",x"AE",x"AE",x"B2",x"A1",x"25",x"55",x"41",x"61",
		x"05",x"07",x"03",x"02",x"80",x"00",x"81",x"C1",x"61",x"C5",x"C7",x"C7",x"C0",x"61",x"33",x"1F",
		x"FF",x"77",x"73",x"62",x"02",x"02",x"A6",x"54",x"51",x"E3",x"92",x"66",x"CC",x"76",x"0F",x"FF",
		x"81",x"00",x"81",x"41",x"E0",x"FE",x"FF",x"FF",x"6F",x"F8",x"F6",x"F1",x"F0",x"78",x"3F",x"1F",
		x"A2",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F0",x"00",
		x"FF",x"FF",x"FF",x"7F",x"1F",x"07",x"01",x"00",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"72",x"02",x"52",x"AA",x"AA",x"FA",x"FA",x"FA",x"FA",x"FA",x"02",x"72",x"8A",x"8A",x"FA",x"FA",
		x"FA",x"FA",x"F2",x"02",x"FA",x"12",x"22",x"7A",x"BA",x"AA",x"EA",x"6A",x"02",x"F2",x"0A",x"0A",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"4E",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"B2",x"B2",x"B2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"3C",x"7E",x"52",x"4A",x"7E",x"3C",x"00",x"00",x"02",x"02",x"7E",x"7E",x"22",x"02",x"00",
		x"00",x"22",x"72",x"5A",x"4E",x"66",x"22",x"00",x"00",x"44",x"6E",x"7A",x"52",x"46",x"44",x"00",
		x"00",x"04",x"7E",x"7E",x"34",x"1C",x"0C",x"00",x"00",x"4C",x"5E",x"52",x"52",x"76",x"74",x"00",
		x"00",x"0C",x"5E",x"52",x"52",x"7E",x"3C",x"00",x"00",x"60",x"70",x"58",x"4E",x"46",x"40",x"00",
		x"00",x"2C",x"7E",x"52",x"52",x"7E",x"2C",x"00",x"00",x"38",x"7C",x"56",x"52",x"72",x"20",x"00",
		x"7E",x"7E",x"30",x"18",x"30",x"7E",x"7E",x"00",x"1E",x"20",x"20",x"1E",x"20",x"20",x"3E",x"00",
		x"00",x"00",x"C0",x"20",x"A0",x"A0",x"A0",x"A0",x"00",x"00",x"7F",x"80",x"83",x"82",x"02",x"B2",
		x"A0",x"A0",x"A0",x"20",x"C0",x"00",x"00",x"00",x"02",x"82",x"83",x"80",x"7F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"BE",x"A6",x"82",x"82",x"82",x"82",x"A6",x"BE",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"86",x"FF",x"FF",x"3F",x"3F",x"FF",x"FF",x"8E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"7F",x"44",x"44",x"44",x"44",x"44",x"44",x"7F",
		x"BF",x"84",x"84",x"84",x"84",x"84",x"84",x"BF",x"DF",x"C4",x"44",x"44",x"44",x"44",x"44",x"DF",
		x"6F",x"E4",x"A4",x"24",x"24",x"24",x"A4",x"EF",x"37",x"74",x"D4",x"94",x"14",x"94",x"D4",x"77",
		x"1B",x"38",x"68",x"C8",x"88",x"C8",x"68",x"3B",x"0D",x"1C",x"34",x"64",x"44",x"64",x"34",x"1D",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"86",x"8E",x"9A",x"B2",x"A2",x"B2",x"9A",x"8E",x"C3",x"47",x"4D",x"59",x"51",x"59",x"4D",x"C7",
		x"E1",x"63",x"66",x"6C",x"68",x"6C",x"66",x"E3",x"F0",x"51",x"53",x"56",x"54",x"56",x"53",x"F1",
		x"F8",x"48",x"49",x"4B",x"4A",x"4B",x"49",x"F8",x"FC",x"44",x"44",x"45",x"45",x"45",x"44",x"FC",
		x"FE",x"46",x"46",x"46",x"46",x"46",x"46",x"FE",x"FF",x"45",x"45",x"45",x"45",x"45",x"45",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"00",x"FE",x"10",x"10",x"FF",x"FF",
		x"00",x"08",x"0C",x"FC",x"FC",x"00",x"A4",x"A6",x"00",x"C0",x"E8",x"00",x"40",x"A0",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"C0",x"C0",x"40",x"40",x"40",x"40",x"40",x"C0",
		x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",x"30",x"70",x"D0",x"90",x"10",x"90",x"D0",x"70",
		x"18",x"38",x"68",x"C8",x"88",x"C8",x"68",x"38",x"0C",x"1C",x"34",x"64",x"44",x"64",x"34",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"00",x"F0",x"40",x"40",x"E0",x"E0",
		x"00",x"04",x"04",x"FC",x"F8",x"00",x"A8",x"A8",x"E0",x"F8",x"7D",x"01",x"70",x"88",x"FE",x"FE",
		x"86",x"8E",x"9A",x"B2",x"A2",x"B2",x"9A",x"8E",x"43",x"47",x"4D",x"59",x"51",x"59",x"4D",x"47",
		x"21",x"23",x"26",x"2C",x"28",x"2C",x"26",x"23",x"10",x"11",x"13",x"16",x"14",x"16",x"13",x"11",
		x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",x"04",x"04",x"04",x"05",x"05",x"05",x"04",x"04",
		x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"90",x"90",x"8A",x"80",x"40",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"42",x"24",x"00",x"00",x"24",x"42",x"00",x"26",x"6F",x"71",x"78",x"78",x"71",x"35",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"F8",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"0C",x"5E",x"D2",x"92",x"92",x"F6",x"64",x"00",
		x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"F8",x"FE",x"1C",x"38",x"1C",x"FE",x"F8",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",
		x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"00",x"00",x"00",x"00",x"28",x"00",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",
		x"00",x"00",x"82",x"C6",x"6C",x"38",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"82",x"00",x"00",
		x"00",x"00",x"82",x"FE",x"FE",x"82",x"00",x"00",x"82",x"FE",x"FE",x"82",x"82",x"FE",x"FE",x"82",
		x"00",x"28",x"28",x"28",x"28",x"28",x"28",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"F6",x"F6",x"00",x"00",x"F6",x"F6",x"00",x"00",x"FA",x"FA",x"00",x"00",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"FA",x"FA",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",x"00",x"E0",x"C0",x"00",x"E0",x"C0",x"00",x"00",
		x"00",x"60",x"E0",x"00",x"60",x"E0",x"00",x"00",x"00",x"00",x"C0",x"00",x"C0",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",
		x"38",x"28",x"3E",x"00",x"00",x"00",x"00",x"00",x"3E",x"00",x"3C",x"02",x"02",x"3C",x"00",x"0E",
		x"22",x"2A",x"3E",x"00",x"00",x"0E",x"3A",x"2A",x"22",x"3E",x"00",x"3E",x"08",x"10",x"3E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"A5",x"BD",x"81",x"42",x"3C",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"A5",x"7C",x"40",x"00",x"38",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"28",x"38",x"00",x"40",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"A2",x"00",x"F0",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",
		x"00",x"01",x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",
		x"54",x"A6",x"02",x"02",x"62",x"73",x"77",x"FF",x"FF",x"8F",x"76",x"7C",x"4E",x"A6",x"D7",x"A3",
		x"FF",x"FF",x"FE",x"FD",x"7F",x"87",x"03",x"80",x"1F",x"3F",x"78",x"F0",x"F1",x"F6",x"F8",x"6F",
		x"BF",x"5F",x"AF",x"4F",x"2A",x"90",x"40",x"A8",x"C1",x"61",x"51",x"25",x"35",x"A1",x"B2",x"AE",
		x"CE",x"9A",x"31",x"3B",x"BF",x"3F",x"1D",x"08",x"1F",x"33",x"61",x"C0",x"C0",x"C7",x"C7",x"65",
		x"40",x"A8",x"50",x"AA",x"4F",x"AF",x"5F",x"BF",x"AE",x"AE",x"B2",x"A1",x"25",x"55",x"41",x"61",
		x"05",x"07",x"03",x"02",x"80",x"00",x"81",x"C1",x"61",x"C5",x"C7",x"C7",x"C0",x"61",x"33",x"1F",
		x"FF",x"77",x"73",x"62",x"02",x"02",x"A6",x"54",x"51",x"E3",x"92",x"66",x"CC",x"76",x"0F",x"FF",
		x"81",x"00",x"81",x"41",x"E0",x"FE",x"FF",x"FF",x"6F",x"F8",x"F6",x"F1",x"F0",x"78",x"3F",x"1F",
		x"A2",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F0",x"00",
		x"FF",x"FF",x"FF",x"7F",x"1F",x"07",x"01",x"00",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"72",x"02",x"52",x"AA",x"AA",x"FA",x"FA",x"FA",x"FA",x"FA",x"02",x"72",x"8A",x"8A",x"FA",x"FA",
		x"FA",x"FA",x"F2",x"02",x"FA",x"12",x"22",x"7A",x"BA",x"AA",x"EA",x"6A",x"02",x"F2",x"0A",x"0A",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"4E",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"1C",x"BE",x"B2",x"B2",x"B2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"0C",x"6E",x"9A",x"9A",x"B2",x"F2",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"3C",x"7E",x"52",x"4A",x"7E",x"3C",x"00",x"00",x"02",x"02",x"7E",x"7E",x"22",x"02",x"00",
		x"00",x"22",x"72",x"5A",x"4E",x"66",x"22",x"00",x"00",x"44",x"6E",x"7A",x"52",x"46",x"44",x"00",
		x"00",x"04",x"7E",x"7E",x"34",x"1C",x"0C",x"00",x"00",x"4C",x"5E",x"52",x"52",x"76",x"74",x"00",
		x"00",x"0C",x"5E",x"52",x"52",x"7E",x"3C",x"00",x"00",x"60",x"70",x"58",x"4E",x"46",x"40",x"00",
		x"00",x"2C",x"7E",x"52",x"52",x"7E",x"2C",x"00",x"00",x"38",x"7C",x"56",x"52",x"72",x"20",x"00",
		x"7E",x"7E",x"30",x"18",x"30",x"7E",x"7E",x"00",x"1E",x"20",x"20",x"1E",x"20",x"20",x"3E",x"00",
		x"00",x"00",x"C0",x"20",x"A0",x"A0",x"A0",x"A0",x"00",x"00",x"7F",x"80",x"83",x"82",x"02",x"B2",
		x"A0",x"A0",x"A0",x"20",x"C0",x"00",x"00",x"00",x"02",x"82",x"83",x"80",x"7F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"BE",x"A6",x"82",x"82",x"82",x"82",x"A6",x"BE",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"86",x"FF",x"FF",x"3F",x"3F",x"FF",x"FF",x"8E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"7F",x"44",x"44",x"44",x"44",x"44",x"44",x"7F",
		x"BF",x"84",x"84",x"84",x"84",x"84",x"84",x"BF",x"DF",x"C4",x"44",x"44",x"44",x"44",x"44",x"DF",
		x"6F",x"E4",x"A4",x"24",x"24",x"24",x"A4",x"EF",x"37",x"74",x"D4",x"94",x"14",x"94",x"D4",x"77",
		x"1B",x"38",x"68",x"C8",x"88",x"C8",x"68",x"3B",x"0D",x"1C",x"34",x"64",x"44",x"64",x"34",x"1D",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"86",x"8E",x"9A",x"B2",x"A2",x"B2",x"9A",x"8E",x"C3",x"47",x"4D",x"59",x"51",x"59",x"4D",x"C7",
		x"E1",x"63",x"66",x"6C",x"68",x"6C",x"66",x"E3",x"F0",x"51",x"53",x"56",x"54",x"56",x"53",x"F1",
		x"F8",x"48",x"49",x"4B",x"4A",x"4B",x"49",x"F8",x"FC",x"44",x"44",x"45",x"45",x"45",x"44",x"FC",
		x"FE",x"46",x"46",x"46",x"46",x"46",x"46",x"FE",x"FF",x"45",x"45",x"45",x"45",x"45",x"45",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"00",x"FE",x"10",x"10",x"FF",x"FF",
		x"00",x"08",x"0C",x"FC",x"FC",x"00",x"A4",x"A6",x"00",x"C0",x"E8",x"00",x"40",x"A0",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"C0",x"C0",x"40",x"40",x"40",x"40",x"40",x"C0",
		x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",x"30",x"70",x"D0",x"90",x"10",x"90",x"D0",x"70",
		x"18",x"38",x"68",x"C8",x"88",x"C8",x"68",x"38",x"0C",x"1C",x"34",x"64",x"44",x"64",x"34",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"00",x"F0",x"40",x"40",x"E0",x"E0",
		x"00",x"04",x"04",x"FC",x"F8",x"00",x"A8",x"A8",x"E0",x"F8",x"7D",x"01",x"70",x"88",x"FE",x"FE",
		x"86",x"8E",x"9A",x"B2",x"A2",x"B2",x"9A",x"8E",x"43",x"47",x"4D",x"59",x"51",x"59",x"4D",x"47",
		x"21",x"23",x"26",x"2C",x"28",x"2C",x"26",x"23",x"10",x"11",x"13",x"16",x"14",x"16",x"13",x"11",
		x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",x"04",x"04",x"04",x"05",x"05",x"05",x"04",x"04",
		x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"90",x"90",x"8A",x"80",x"40",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"42",x"24",x"00",x"00",x"24",x"42",x"00",x"26",x"6F",x"71",x"78",x"78",x"71",x"35",x"00",
		x"17",x"CB",x"13",x"17",x"C6",x"74",x"57",x"19",x"C9",x"57",x"0F",x"DA",x"22",x"30",x"0E",x"93",
		x"0F",x"0F",x"D2",x"17",x"30",x"0E",x"6C",x"07",x"DA",x"31",x"30",x"79",x"E6",x"F0",x"4F",x"C3",
		x"31",x"30",x"0E",x"B4",x"0F",x"0F",x"D2",x"2B",x"30",x"0E",x"1E",x"CB",x"50",x"CA",x"31",x"30",
		x"05",x"79",x"0F",x"0F",x"4F",x"E6",x"03",x"B8",x"C2",x"31",x"30",x"79",x"0F",x"0F",x"E6",x"03",
		x"FE",x"03",x"C0",x"CB",x"92",x"15",x"C0",x"3E",x"04",x"C9",x"11",x"E0",x"FF",x"3A",x"8E",x"63",
		x"4F",x"06",x"00",x"21",x"00",x"76",x"CD",x"64",x"30",x"21",x"C0",x"75",x"CD",x"64",x"30",x"21",
		x"8E",x"63",x"35",x"C9",x"09",x"7E",x"19",x"77",x"C9",x"DF",x"2A",x"C0",x"63",x"34",x"C9",x"21",
		x"AF",x"62",x"34",x"7E",x"E6",x"07",x"C0",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"0E",x"81",x"21",
		x"09",x"69",x"CD",x"96",x"30",x"21",x"1D",x"69",x"CD",x"96",x"30",x"CD",x"57",x"00",x"E6",x"80",
		x"21",x"2D",x"69",x"AE",x"77",x"C9",x"06",x"02",x"79",x"AE",x"77",x"19",x"10",x"FA",x"C9",x"E5",
		x"21",x"C0",x"60",x"3A",x"B0",x"60",x"6F",x"CB",x"7E",x"CA",x"BB",x"30",x"72",x"2C",x"73",x"2C",
		x"7D",x"FE",x"C0",x"D2",x"B8",x"30",x"3E",x"C0",x"32",x"B0",x"60",x"E1",x"C9",x"21",x"50",x"69",
		x"06",x"02",x"CD",x"E4",x"30",x"2E",x"80",x"06",x"0A",x"CD",x"E4",x"30",x"2E",x"B8",x"06",x"0B",
		x"CD",x"E4",x"30",x"21",x"0C",x"6A",x"06",x"05",x"C3",x"E4",x"30",x"21",x"4C",x"69",x"36",x"00",
		x"2E",x"58",x"06",x"06",x"7D",x"36",x"00",x"C6",x"04",x"6F",x"10",x"F9",x"C9",x"CD",x"FA",x"30",
		x"CD",x"3C",x"31",x"CD",x"B1",x"31",x"CD",x"F3",x"34",x"C9",x"3A",x"80",x"63",x"FE",x"06",x"38",
		x"02",x"3E",x"05",x"EF",x"10",x"31",x"10",x"31",x"1B",x"31",x"26",x"31",x"26",x"31",x"31",x"31",
		x"3A",x"1A",x"60",x"E6",x"01",x"FE",x"01",x"C8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"07",
		x"FE",x"05",x"F8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"03",x"FE",x"03",x"F8",x"33",x"33",
		x"C9",x"3A",x"1A",x"60",x"E6",x"07",x"FE",x"07",x"F8",x"33",x"33",x"C9",x"DD",x"21",x"00",x"64",
		x"AF",x"32",x"A1",x"63",x"06",x"05",x"11",x"20",x"00",x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"7C",
		x"31",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"3E",x"01",x"DD",x"77",x"08",x"3A",x"17",x"62",
		x"FE",x"01",x"C2",x"6A",x"31",x"3E",x"00",x"DD",x"77",x"08",x"DD",x"19",x"10",x"DB",x"21",x"A0",
		x"63",x"36",x"00",x"3A",x"A1",x"63",x"FE",x"00",x"C0",x"33",x"33",x"C9",x"3A",x"A1",x"63",x"FE",
		x"05",x"CA",x"6A",x"31",x"3A",x"27",x"62",x"FE",x"02",x"C2",x"95",x"31",x"3A",x"A1",x"63",x"4F",
		x"3A",x"80",x"63",x"B9",x"C8",x"3A",x"A0",x"63",x"FE",x"01",x"C2",x"6A",x"31",x"DD",x"77",x"00",
		x"DD",x"77",x"18",x"AF",x"32",x"A0",x"63",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"C3",x"6A",
		x"31",x"CD",x"DD",x"31",x"AF",x"32",x"A2",x"63",x"21",x"E0",x"63",x"22",x"C8",x"63",x"2A",x"C8",
		x"63",x"01",x"20",x"00",x"09",x"22",x"C8",x"63",x"7E",x"A7",x"CA",x"D0",x"31",x"CD",x"02",x"32",
		x"3A",x"A2",x"63",x"3C",x"32",x"A2",x"63",x"FE",x"05",x"C2",x"BE",x"31",x"C9",x"3A",x"80",x"63",
		x"FE",x"03",x"F8",x"CD",x"F6",x"31",x"FE",x"01",x"C0",x"21",x"39",x"64",x"3E",x"02",x"77",x"21",
		x"79",x"64",x"3E",x"02",x"77",x"C9",x"3A",x"18",x"60",x"E6",x"03",x"FE",x"01",x"C0",x"3A",x"1A",
		x"60",x"C9",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"18",x"FE",x"01",x"CA",x"7A",x"32",x"DD",x"7E",
		x"0D",x"FE",x"04",x"F2",x"30",x"32",x"DD",x"7E",x"19",x"FE",x"02",x"CA",x"7E",x"32",x"CD",x"0F",
		x"33",x"3A",x"18",x"60",x"E6",x"03",x"C2",x"33",x"32",x"DD",x"7E",x"0D",x"A7",x"CA",x"57",x"32",
		x"CD",x"3D",x"33",x"DD",x"7E",x"0D",x"FE",x"04",x"F2",x"91",x"32",x"CD",x"AD",x"33",x"CD",x"8C",
		x"29",x"FE",x"01",x"CA",x"97",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0E",x"FE",x"10",x"DA",
		x"8C",x"32",x"FE",x"F0",x"D2",x"84",x"32",x"DD",x"7E",x"13",x"FE",x"00",x"C2",x"B9",x"32",x"3E",
		x"11",x"DD",x"77",x"13",x"16",x"00",x"5F",x"21",x"7A",x"3A",x"19",x"7E",x"DD",x"46",x"0E",x"DD",
		x"70",x"03",x"DD",x"4E",x"0F",x"81",x"DD",x"77",x"05",x"C9",x"CD",x"BD",x"32",x"C9",x"CD",x"D6",
		x"32",x"C3",x"29",x"32",x"3E",x"02",x"DD",x"77",x"0D",x"C3",x"57",x"32",x"3E",x"01",x"C3",x"86",
		x"32",x"CD",x"E7",x"33",x"C3",x"57",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0D",x"FE",x"01",
		x"C2",x"B1",x"32",x"3E",x"02",x"DD",x"35",x"0E",x"DD",x"77",x"0D",x"CD",x"C3",x"33",x"C3",x"57",
		x"32",x"3E",x"01",x"DD",x"34",x"0E",x"C3",x"A8",x"32",x"3D",x"C3",x"61",x"32",x"3A",x"27",x"62",
		x"FE",x"01",x"CA",x"CE",x"32",x"FE",x"02",x"CA",x"D2",x"32",x"CD",x"B9",x"34",x"C9",x"CD",x"2C",
		x"34",x"C9",x"CD",x"78",x"34",x"C9",x"DD",x"7E",x"1C",x"FE",x"00",x"C2",x"FD",x"32",x"DD",x"7E",
		x"1D",x"FE",x"01",x"C2",x"0B",x"33",x"DD",x"36",x"1D",x"00",x"3A",x"05",x"62",x"DD",x"46",x"0F",
		x"90",x"DA",x"03",x"33",x"DD",x"36",x"1C",x"FF",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"35",x"1C",
		x"C2",x"F8",x"32",x"DD",x"36",x"19",x"00",x"DD",x"36",x"1C",x"00",x"CD",x"0F",x"33",x"C9",x"DD",
		x"7E",x"16",x"FE",x"00",x"C2",x"32",x"33",x"DD",x"36",x"16",x"2B",x"DD",x"36",x"0D",x"00",x"3A",
		x"18",x"60",x"0F",x"D2",x"32",x"33",x"DD",x"7E",x"0D",x"FE",x"01",x"CA",x"36",x"33",x"DD",x"36",
		x"0D",x"01",x"DD",x"35",x"16",x"C9",x"DD",x"36",x"0D",x"02",x"C3",x"32",x"33",x"DD",x"7E",x"0D",
		x"FE",x"08",x"CA",x"71",x"33",x"FE",x"04",x"CA",x"8A",x"33",x"CD",x"A1",x"33",x"DD",x"7E",x"0F",
		x"C6",x"08",x"57",x"DD",x"7E",x"0E",x"01",x"15",x"00",x"CD",x"6E",x"23",x"A7",x"CA",x"99",x"33",
		x"DD",x"70",x"1F",x"3A",x"05",x"62",x"47",x"DD",x"7E",x"0F",x"90",x"D0",x"DD",x"36",x"0D",x"04",
		x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"DD",
		x"7E",x"19",x"FE",x"02",x"C0",x"DD",x"36",x"1D",x"01",x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",
		x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"70",x"1F",x"DD",x"36",x"0D",x"08",
		x"C9",x"3E",x"07",x"F7",x"DD",x"7E",x"0F",x"FE",x"59",x"D0",x"33",x"33",x"C9",x"DD",x"7E",x"0D",
		x"FE",x"01",x"CA",x"D9",x"33",x"DD",x"7E",x"07",x"E6",x"7F",x"DD",x"77",x"07",x"DD",x"35",x"0E",
		x"CD",x"09",x"34",x"3A",x"27",x"62",x"FE",x"01",x"C0",x"DD",x"66",x"0E",x"DD",x"6E",x"0F",x"DD",
		x"46",x"0D",x"CD",x"33",x"23",x"DD",x"75",x"0F",x"C9",x"DD",x"7E",x"07",x"F6",x"80",x"DD",x"77",
		x"07",x"DD",x"34",x"0E",x"C3",x"C0",x"33",x"CD",x"09",x"34",x"DD",x"7E",x"0D",x"FE",x"08",x"C2",
		x"05",x"34",x"DD",x"7E",x"14",x"A7",x"C2",x"01",x"34",x"DD",x"36",x"14",x"02",x"DD",x"35",x"0F",
		x"C9",x"DD",x"35",x"14",x"C9",x"DD",x"34",x"0F",x"C9",x"DD",x"7E",x"15",x"A7",x"C2",x"28",x"34",
		x"DD",x"36",x"15",x"02",x"DD",x"34",x"07",x"DD",x"7E",x"07",x"E6",x"0F",x"FE",x"0F",x"C0",x"DD",
		x"7E",x"07",x"EE",x"02",x"DD",x"77",x"07",x"C9",x"DD",x"35",x"15",x"C9",x"DD",x"6E",x"1A",x"DD",
		x"66",x"1B",x"AF",x"01",x"00",x"00",x"ED",x"4A",x"C2",x"42",x"34",x"21",x"8C",x"3A",x"DD",x"36",
		x"03",x"26",x"DD",x"34",x"03",x"7E",x"FE",x"AA",x"CA",x"56",x"34",x"DD",x"77",x"05",x"23",x"DD",
		x"75",x"1A",x"DD",x"74",x"1B",x"C9",x"AF",x"DD",x"77",x"13",x"DD",x"77",x"18",x"DD",x"77",x"0D",
		x"DD",x"77",x"1C",x"DD",x"7E",x"03",x"DD",x"77",x"0E",x"DD",x"7E",x"05",x"DD",x"77",x"0F",x"DD",
		x"36",x"1A",x"00",x"DD",x"36",x"1B",x"00",x"C9",x"DD",x"6E",x"1A",x"DD",x"66",x"1B",x"AF",x"01",
		x"00",x"00",x"ED",x"4A",x"C2",x"9A",x"34",x"21",x"AC",x"3A",x"3A",x"03",x"62",x"CB",x"7F",x"CA",
		x"A8",x"34",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"03",x"7E",x"DD",x"7E",x"0D",x"FE",x"01",x"C2",
		x"B3",x"34",x"DD",x"34",x"03",x"C3",x"45",x"34",x"DD",x"36",x"0D",x"02",x"DD",x"36",x"03",x"80",
		x"C3",x"9A",x"34",x"DD",x"35",x"03",x"C3",x"45",x"34",x"3A",x"27",x"62",x"FE",x"03",x"C8",x"3A",
		x"03",x"62",x"CB",x"7F",x"C2",x"ED",x"34",x"21",x"C4",x"3A",x"06",x"00",x"3A",x"19",x"60",x"E6",
		x"06",x"4F",x"09",x"7E",x"DD",x"77",x"03",x"DD",x"77",x"0E",x"23",x"7E",x"DD",x"77",x"05",x"DD",
		x"77",x"0F",x"AF",x"DD",x"77",x"0D",x"DD",x"77",x"18",x"DD",x"77",x"1C",x"C9",x"21",x"D4",x"3A",
		x"C3",x"CA",x"34",x"21",x"00",x"64",x"11",x"D0",x"69",x"06",x"05",x"7E",x"A7",x"CA",x"1E",x"35",
		x"2C",x"2C",x"2C",x"7E",x"12",x"3E",x"04",x"85",x"6F",x"1C",x"7E",x"12",x"2C",x"1C",x"7E",x"12",
		x"2D",x"2D",x"2D",x"1C",x"7E",x"12",x"13",x"3E",x"1B",x"85",x"6F",x"10",x"DE",x"C9",x"3E",x"05",
		x"85",x"6F",x"3E",x"04",x"83",x"5F",x"C3",x"17",x"35",x"00",x"00",x"00",x"00",x"01",x"00",x"00",
		x"02",x"00",x"00",x"03",x"00",x"00",x"04",x"00",x"00",x"05",x"00",x"00",x"06",x"00",x"00",x"07",
		x"00",x"00",x"08",x"00",x"00",x"09",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",
		x"00",x"30",x"00",x"00",x"40",x"00",x"00",x"50",x"00",x"00",x"60",x"00",x"00",x"70",x"00",x"00",
		x"80",x"00",x"00",x"90",x"00",x"94",x"77",x"01",x"23",x"24",x"10",x"10",x"00",x"00",x"07",x"06",
		x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3F",x"00",x"50",x"76",x"00",x"F4",x"76",x"96",x"77",x"02",x"1E",x"14",x"10",x"10",x"00",x"00",
		x"06",x"01",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"3F",x"00",x"00",x"61",x"00",x"F6",x"76",x"98",x"77",x"03",x"22",x"14",x"10",x"10",
		x"00",x"00",x"05",x"09",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"59",x"00",x"F8",x"76",x"9A",x"77",x"04",x"24",x"18",
		x"10",x"10",x"00",x"00",x"05",x"00",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"50",x"00",x"FA",x"76",x"9C",x"77",x"05",
		x"24",x"18",x"10",x"10",x"00",x"00",x"04",x"03",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"00",x"43",x"00",x"FC",x"76",x"3B",
		x"5C",x"4B",x"5C",x"5B",x"5C",x"6B",x"5C",x"7B",x"5C",x"8B",x"5C",x"9B",x"5C",x"AB",x"5C",x"BB",
		x"5C",x"CB",x"5C",x"3B",x"6C",x"4B",x"6C",x"5B",x"6C",x"6B",x"6C",x"7B",x"6C",x"8B",x"6C",x"9B",
		x"6C",x"AB",x"6C",x"BB",x"6C",x"CB",x"6C",x"3B",x"7C",x"4B",x"7C",x"5B",x"7C",x"6B",x"7C",x"7B",
		x"7C",x"8B",x"7C",x"9B",x"7C",x"AB",x"7C",x"BB",x"7C",x"CB",x"7C",x"8B",x"36",x"01",x"00",x"98",
		x"36",x"A5",x"36",x"B2",x"36",x"BF",x"36",x"06",x"00",x"CC",x"36",x"08",x"00",x"E6",x"36",x"FD",
		x"36",x"0B",x"00",x"15",x"37",x"1C",x"37",x"30",x"37",x"38",x"37",x"47",x"37",x"5D",x"37",x"73",
		x"37",x"8B",x"37",x"00",x"61",x"22",x"61",x"44",x"61",x"66",x"61",x"88",x"61",x"9E",x"37",x"B6",
		x"37",x"D2",x"37",x"E1",x"37",x"1D",x"00",x"00",x"3F",x"09",x"3F",x"96",x"76",x"17",x"11",x"1D",
		x"15",x"10",x"10",x"1F",x"26",x"15",x"22",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",
		x"10",x"30",x"32",x"31",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"30",x"33",
		x"31",x"3F",x"80",x"76",x"18",x"19",x"17",x"18",x"10",x"23",x"13",x"1F",x"22",x"15",x"3F",x"9F",
		x"75",x"13",x"22",x"15",x"14",x"19",x"24",x"10",x"10",x"10",x"10",x"3F",x"5E",x"77",x"18",x"1F",
		x"27",x"10",x"18",x"19",x"17",x"18",x"10",x"13",x"11",x"1E",x"10",x"29",x"1F",x"25",x"10",x"17",
		x"15",x"24",x"10",x"FB",x"10",x"3F",x"29",x"77",x"1F",x"1E",x"1C",x"29",x"10",x"01",x"10",x"20",
		x"1C",x"11",x"29",x"15",x"22",x"10",x"12",x"25",x"24",x"24",x"1F",x"1E",x"3F",x"29",x"77",x"01",
		x"10",x"1F",x"22",x"10",x"02",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"23",x"10",x"12",x"25",
		x"24",x"24",x"1F",x"1E",x"3F",x"27",x"76",x"20",x"25",x"23",x"18",x"3F",x"06",x"77",x"1E",x"11",
		x"1D",x"15",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"22",x"11",x"24",x"19",x"1F",x"1E",x"3F",
		x"88",x"76",x"1E",x"11",x"1D",x"15",x"2E",x"3F",x"E9",x"75",x"2D",x"2D",x"2D",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"0B",x"77",x"11",x"10",x"12",x"10",x"13",x"10",x"14",
		x"10",x"15",x"10",x"16",x"10",x"17",x"10",x"18",x"10",x"19",x"10",x"1A",x"3F",x"0D",x"77",x"1B",
		x"10",x"1C",x"10",x"1D",x"10",x"1E",x"10",x"1F",x"10",x"20",x"10",x"21",x"10",x"22",x"10",x"23",
		x"10",x"24",x"3F",x"0F",x"77",x"25",x"10",x"26",x"10",x"27",x"10",x"28",x"10",x"29",x"10",x"2A",
		x"10",x"2B",x"10",x"2C",x"44",x"45",x"46",x"47",x"48",x"10",x"3F",x"F2",x"76",x"22",x"15",x"17",
		x"19",x"10",x"24",x"19",x"1D",x"15",x"10",x"10",x"30",x"03",x"00",x"31",x"10",x"3F",x"92",x"77",
		x"22",x"11",x"1E",x"1B",x"10",x"10",x"23",x"13",x"1F",x"22",x"15",x"10",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"10",x"10",x"10",x"3F",x"72",x"77",x"29",x"1F",x"25",x"22",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"27",x"11",x"23",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"15",x"22",x"15",x"14",
		x"42",x"3F",x"A7",x"76",x"19",x"1E",x"23",x"15",x"22",x"24",x"10",x"13",x"1F",x"19",x"1E",x"10",
		x"3F",x"0A",x"77",x"10",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"10",x"10",x"10",x"13",
		x"1F",x"19",x"1E",x"3F",x"FC",x"76",x"49",x"4A",x"10",x"1E",x"19",x"1E",x"24",x"15",x"1E",x"14",
		x"1F",x"10",x"10",x"10",x"10",x"3F",x"7C",x"75",x"01",x"09",x"08",x"01",x"3F",x"02",x"97",x"38",
		x"68",x"38",x"02",x"DF",x"54",x"10",x"54",x"02",x"EF",x"6D",x"20",x"6D",x"02",x"DF",x"8E",x"10",
		x"8E",x"02",x"EF",x"AF",x"20",x"AF",x"02",x"DF",x"D0",x"10",x"D0",x"02",x"EF",x"F1",x"10",x"F1",
		x"00",x"53",x"18",x"53",x"54",x"00",x"63",x"18",x"63",x"54",x"00",x"93",x"38",x"93",x"54",x"00",
		x"83",x"54",x"83",x"F1",x"00",x"93",x"54",x"93",x"F1",x"AA",x"8D",x"7D",x"8C",x"6F",x"00",x"7C",
		x"6E",x"00",x"7C",x"6D",x"00",x"7C",x"6C",x"00",x"7C",x"8F",x"7F",x"8E",x"47",x"27",x"08",x"50",
		x"2F",x"A7",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"23",x"07",x"40",
		x"46",x"A9",x"08",x"44",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",x"70",x"08",x"48",
		x"00",x"70",x"0A",x"48",x"6F",x"10",x"09",x"23",x"6F",x"11",x"0A",x"33",x"50",x"34",x"08",x"3C",
		x"00",x"35",x"08",x"3C",x"53",x"32",x"08",x"40",x"63",x"33",x"08",x"40",x"00",x"70",x"08",x"48",
		x"53",x"36",x"08",x"50",x"63",x"37",x"08",x"50",x"6B",x"31",x"08",x"41",x"00",x"70",x"08",x"48",
		x"6A",x"14",x"0A",x"48",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"7F",x"04",x"7F",x"F0",x"10",
		x"F0",x"02",x"DF",x"F2",x"70",x"F8",x"02",x"6F",x"F8",x"10",x"F8",x"AA",x"04",x"DF",x"D0",x"90",
		x"D0",x"02",x"DF",x"DC",x"20",x"D1",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"04",x"DF",x"A8",x"20",
		x"A8",x"04",x"5F",x"B0",x"20",x"B0",x"02",x"DF",x"B0",x"20",x"BB",x"AA",x"04",x"DF",x"88",x"30",
		x"88",x"04",x"DF",x"90",x"B0",x"90",x"02",x"DF",x"9A",x"20",x"8F",x"AA",x"04",x"BF",x"68",x"20",
		x"68",x"04",x"3F",x"70",x"20",x"70",x"02",x"DF",x"6E",x"20",x"79",x"AA",x"02",x"DF",x"58",x"A0",
		x"55",x"AA",x"00",x"70",x"08",x"44",x"2B",x"AC",x"08",x"4C",x"3B",x"AE",x"08",x"4C",x"3B",x"AF",
		x"08",x"3C",x"4B",x"B0",x"07",x"3C",x"4B",x"AD",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"47",x"27",x"08",x"4C",x"2F",x"A7",
		x"08",x"4C",x"3B",x"25",x"08",x"4C",x"00",x"70",x"08",x"44",x"3B",x"23",x"07",x"3C",x"4B",x"2A",
		x"08",x"3C",x"4B",x"2B",x"08",x"4C",x"2B",x"AA",x"08",x"3C",x"2B",x"AB",x"08",x"4C",x"00",x"70",
		x"0A",x"44",x"00",x"70",x"08",x"44",x"4B",x"2C",x"08",x"4C",x"3B",x"2E",x"08",x"4C",x"3B",x"2F",
		x"08",x"3C",x"2B",x"30",x"07",x"3C",x"2B",x"2D",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"02",x"02",x"02",x"02",x"03",
		x"03",x"03",x"7F",x"1E",x"4E",x"BB",x"4C",x"D8",x"4E",x"59",x"4E",x"7F",x"BB",x"4D",x"7F",x"47",
		x"27",x"08",x"50",x"2D",x"26",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",
		x"24",x"07",x"40",x"4B",x"28",x"08",x"40",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",
		x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"49",x"A6",x"08",x"50",x"2F",x"A7",x"08",x"50",x"3B",
		x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"24",x"07",x"40",x"46",x"A9",x"08",x"44",x"00",
		x"70",x"08",x"48",x"2B",x"A8",x"08",x"40",x"00",x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"73",
		x"A7",x"88",x"60",x"8B",x"27",x"88",x"60",x"7F",x"25",x"88",x"60",x"00",x"70",x"88",x"68",x"7F",
		x"24",x"87",x"70",x"74",x"29",x"88",x"6C",x"00",x"70",x"88",x"68",x"8A",x"A9",x"88",x"6C",x"00",
		x"70",x"88",x"68",x"00",x"70",x"8A",x"68",x"05",x"AF",x"F0",x"50",x"F0",x"AA",x"05",x"AF",x"E8",
		x"50",x"E8",x"AA",x"05",x"AF",x"E0",x"50",x"E0",x"AA",x"05",x"AF",x"D8",x"50",x"D8",x"AA",x"05",
		x"B7",x"58",x"48",x"58",x"AA",x"01",x"04",x"01",x"03",x"04",x"01",x"02",x"03",x"04",x"01",x"02",
		x"01",x"03",x"04",x"01",x"02",x"01",x"03",x"01",x"04",x"7F",x"FF",x"00",x"FF",x"FF",x"FE",x"FE",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"00",x"E8",x"E5",x"E3",x"E2",
		x"E1",x"E0",x"DF",x"DE",x"DD",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DE",x"DF",
		x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E7",x"E9",x"EB",x"ED",x"F0",x"AA",x"80",x"7B",x"78",x"76",
		x"74",x"73",x"72",x"71",x"70",x"70",x"6F",x"6F",x"6F",x"70",x"70",x"71",x"72",x"73",x"74",x"75",
		x"76",x"77",x"78",x"AA",x"EE",x"F0",x"DB",x"A0",x"E6",x"C8",x"D6",x"78",x"EB",x"F0",x"DB",x"A0",
		x"E6",x"C8",x"E6",x"C8",x"1B",x"C8",x"23",x"A0",x"2B",x"78",x"12",x"F0",x"1B",x"C8",x"23",x"A0",
		x"12",x"F0",x"1B",x"C8",x"02",x"97",x"38",x"68",x"38",x"02",x"9F",x"54",x"10",x"54",x"02",x"DF",
		x"58",x"A0",x"55",x"02",x"EF",x"6D",x"20",x"79",x"02",x"DF",x"9A",x"10",x"8E",x"02",x"EF",x"AF",
		x"20",x"BB",x"02",x"DF",x"DC",x"10",x"D0",x"02",x"FF",x"F0",x"80",x"F7",x"02",x"7F",x"F8",x"00",
		x"F8",x"00",x"CB",x"57",x"CB",x"6F",x"00",x"CB",x"99",x"CB",x"B1",x"00",x"CB",x"DB",x"CB",x"F3",
		x"00",x"63",x"18",x"63",x"54",x"01",x"63",x"D5",x"63",x"F8",x"00",x"33",x"78",x"33",x"90",x"00",
		x"33",x"BA",x"33",x"D2",x"00",x"53",x"18",x"53",x"54",x"01",x"53",x"92",x"53",x"B8",x"00",x"5B",
		x"76",x"5B",x"92",x"00",x"73",x"B6",x"73",x"D6",x"00",x"83",x"95",x"83",x"B5",x"00",x"93",x"38",
		x"93",x"54",x"01",x"BB",x"70",x"BB",x"98",x"01",x"6B",x"54",x"6B",x"75",x"AA",x"06",x"8F",x"90",
		x"70",x"90",x"06",x"8F",x"98",x"70",x"98",x"06",x"8F",x"A0",x"70",x"A0",x"00",x"63",x"18",x"63",
		x"58",x"00",x"63",x"80",x"63",x"A8",x"00",x"63",x"D0",x"63",x"F8",x"00",x"53",x"18",x"53",x"58",
		x"00",x"53",x"A8",x"53",x"D0",x"00",x"9B",x"80",x"9B",x"A8",x"00",x"9B",x"D0",x"9B",x"F8",x"01",
		x"23",x"58",x"23",x"80",x"01",x"DB",x"58",x"DB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"A3",x"A8",x"A3",x"D0",x"00",x"2B",x"D0",x"2B",x"F8",x"00",x"D3",x"D0",
		x"D3",x"F8",x"00",x"93",x"38",x"93",x"58",x"02",x"97",x"38",x"68",x"38",x"03",x"EF",x"58",x"10",
		x"58",x"03",x"F7",x"80",x"88",x"80",x"03",x"77",x"80",x"08",x"80",x"02",x"A7",x"A8",x"50",x"A8",
		x"02",x"E7",x"A8",x"B8",x"A8",x"02",x"3F",x"A8",x"18",x"A8",x"03",x"EF",x"D0",x"10",x"D0",x"02",
		x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"63",x"18",x"63",x"58",x"00",x"63",x"88",x"63",x"D0",x"00",
		x"53",x"18",x"53",x"58",x"00",x"53",x"88",x"53",x"D0",x"00",x"E3",x"68",x"E3",x"90",x"00",x"E3",
		x"B8",x"E3",x"D0",x"00",x"CB",x"90",x"CB",x"B0",x"00",x"B3",x"58",x"B3",x"78",x"00",x"9B",x"80",
		x"9B",x"A0",x"00",x"93",x"38",x"93",x"58",x"00",x"23",x"88",x"23",x"C0",x"00",x"1B",x"C0",x"1B",
		x"E8",x"02",x"97",x"38",x"68",x"38",x"02",x"B7",x"58",x"10",x"58",x"02",x"EF",x"68",x"E0",x"68",
		x"02",x"D7",x"70",x"C8",x"70",x"02",x"BF",x"78",x"B0",x"78",x"02",x"A7",x"80",x"90",x"80",x"02",
		x"67",x"88",x"48",x"88",x"02",x"27",x"88",x"10",x"88",x"02",x"EF",x"90",x"C8",x"90",x"02",x"A7",
		x"A0",x"98",x"A0",x"02",x"BF",x"A8",x"B0",x"A8",x"02",x"D7",x"B0",x"C8",x"B0",x"02",x"EF",x"B8",
		x"E0",x"B8",x"02",x"27",x"C0",x"10",x"C0",x"02",x"EF",x"D0",x"D8",x"D0",x"02",x"67",x"D0",x"50",
		x"D0",x"02",x"CF",x"D8",x"C0",x"D8",x"02",x"B7",x"E0",x"A8",x"E0",x"02",x"9F",x"E8",x"88",x"E8",
		x"02",x"27",x"E8",x"10",x"E8",x"02",x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"7B",x"80",x"7B",x"A8",
		x"00",x"7B",x"D0",x"7B",x"F8",x"00",x"33",x"58",x"33",x"80",x"00",x"53",x"58",x"53",x"80",x"00",
		x"AB",x"58",x"AB",x"80",x"00",x"CB",x"58",x"CB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"23",x"A8",x"23",x"D0",x"00",x"5B",x"A8",x"5B",x"D0",x"00",x"A3",x"A8",
		x"A3",x"D0",x"00",x"DB",x"A8",x"DB",x"D0",x"00",x"1B",x"D0",x"1B",x"F8",x"00",x"E3",x"D0",x"E3",
		x"F8",x"05",x"B7",x"30",x"48",x"30",x"05",x"CF",x"58",x"30",x"58",x"05",x"D7",x"80",x"28",x"80",
		x"05",x"DF",x"A8",x"20",x"A8",x"05",x"E7",x"D0",x"18",x"D0",x"05",x"EF",x"F8",x"10",x"F8",x"AA",
		x"10",x"82",x"85",x"8B",x"10",x"85",x"80",x"8B",x"10",x"87",x"85",x"8B",x"81",x"80",x"80",x"8B",
		x"81",x"82",x"85",x"8B",x"81",x"85",x"80",x"8B",x"05",x"88",x"77",x"01",x"68",x"77",x"01",x"6C",
		x"77",x"03",x"49",x"77",x"05",x"08",x"77",x"01",x"E8",x"76",x"01",x"EC",x"76",x"05",x"C8",x"76",
		x"05",x"88",x"76",x"02",x"69",x"76",x"02",x"4A",x"76",x"05",x"28",x"76",x"05",x"E8",x"75",x"01",
		x"CA",x"75",x"03",x"A9",x"75",x"01",x"88",x"75",x"01",x"8C",x"75",x"05",x"48",x"75",x"01",x"28",
		x"75",x"01",x"2A",x"75",x"01",x"2C",x"75",x"01",x"08",x"75",x"01",x"0A",x"75",x"01",x"0C",x"75",
		x"03",x"C8",x"74",x"03",x"AA",x"74",x"03",x"88",x"74",x"05",x"2F",x"77",x"05",x"0F",x"77",x"02",
		x"F0",x"76",x"02",x"CF",x"76",x"02",x"D2",x"76",x"05",x"8F",x"76",x"05",x"6F",x"76",x"01",x"4F",
		x"76",x"01",x"53",x"76",x"05",x"2F",x"76",x"05",x"EF",x"75",x"02",x"D0",x"75",x"02",x"B1",x"75",
		x"05",x"8F",x"75",x"03",x"50",x"75",x"05",x"2F",x"75",x"01",x"0F",x"75",x"01",x"13",x"75",x"01",
		x"EF",x"74",x"01",x"F1",x"74",x"01",x"F3",x"74",x"02",x"D1",x"74",x"00",x"00",x"00",x"23",x"68",
		x"01",x"11",x"00",x"00",x"00",x"10",x"DB",x"68",x"01",x"40",x"00",x"00",x"08",x"01",x"01",x"01",
		x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"01",x"C0",x"FF",
		x"01",x"FF",x"FF",x"34",x"C3",x"39",x"00",x"67",x"80",x"69",x"1A",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"0B",x"4B",
		x"14",x"18",x"0B",x"4B",x"1E",x"18",x"0B",x"3B",x"14",x"18",x"0B",x"3B",x"3D",x"01",x"03",x"02",
		x"4D",x"01",x"04",x"01",x"27",x"70",x"01",x"E0",x"00",x"00",x"7F",x"40",x"01",x"78",x"02",x"00",
		x"27",x"49",x"0C",x"F0",x"7F",x"49",x"0C",x"88",x"1E",x"07",x"03",x"09",x"24",x"64",x"BB",x"C0",
		x"23",x"8D",x"7B",x"B4",x"1B",x"8C",x"7C",x"64",x"4B",x"0E",x"04",x"02",x"23",x"46",x"03",x"68",
		x"DB",x"46",x"03",x"68",x"17",x"50",x"00",x"5C",x"E7",x"D0",x"00",x"5C",x"8C",x"50",x"00",x"84",
		x"73",x"D0",x"00",x"84",x"17",x"50",x"00",x"D4",x"E7",x"D0",x"00",x"D4",x"53",x"73",x"0A",x"A0",
		x"8B",x"74",x"0A",x"F0",x"DB",x"75",x"0A",x"A0",x"5B",x"73",x"0A",x"C8",x"E3",x"74",x"0A",x"60",
		x"1B",x"75",x"0A",x"80",x"DB",x"73",x"0A",x"C8",x"93",x"74",x"0A",x"F0",x"33",x"75",x"0A",x"50",
		x"44",x"03",x"08",x"04",x"37",x"F4",x"37",x"C0",x"37",x"8C",x"77",x"70",x"77",x"A4",x"77",x"D8",
		x"11",x"01",x"00",x"06",x"7B",x"1F",x"D2",x"28",x"1E",x"1E",x"03",x"06",x"7D",x"1F",x"D2",x"28",
		x"1E",x"1E",x"05",x"06",x"7F",x"C3",x"28",x"1E",x"3A",x"27",x"62",x"E5",x"EF",x"00",x"00",x"99",
		x"3E",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",x"E1",x"AF",x"32",x"60",x"60",x"06",x"0A",
		x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"C3",x"3E",x"06",x"05",x"DD",x"21",x"00",x"64",
		x"CD",x"C3",x"3E",x"3A",x"60",x"60",x"A7",x"C8",x"FE",x"01",x"C8",x"FE",x"03",x"3E",x"03",x"D8",
		x"3E",x"07",x"C9",x"DD",x"CB",x"00",x"46",x"CA",x"FA",x"3E",x"79",x"DD",x"96",x"05",x"D2",x"D3",
		x"3E",x"ED",x"44",x"3C",x"95",x"DA",x"DE",x"3E",x"DD",x"96",x"0A",x"D2",x"FA",x"3E",x"FD",x"7E",
		x"03",x"DD",x"96",x"03",x"D2",x"E9",x"3E",x"ED",x"44",x"94",x"DA",x"F3",x"3E",x"DD",x"96",x"09",
		x"D2",x"FA",x"3E",x"3A",x"60",x"60",x"3C",x"32",x"60",x"60",x"DD",x"19",x"10",x"C5",x"C9",x"00",
		x"5C",x"76",x"49",x"4A",x"01",x"09",x"08",x"01",x"3F",x"7D",x"77",x"1E",x"19",x"1E",x"24",x"15",
		x"1E",x"14",x"1F",x"10",x"1F",x"16",x"10",x"11",x"1D",x"15",x"22",x"19",x"13",x"11",x"10",x"19",
		x"1E",x"13",x"2B",x"3F",x"21",x"AF",x"74",x"11",x"E0",x"FF",x"36",x"9F",x"19",x"36",x"9E",x"C9",
		x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"2C",x"57",x"45",x"20",x"57",x"4F",x"55",x"4C",x"44",
		x"20",x"54",x"45",x"41",x"43",x"48",x"20",x"59",x"4F",x"55",x"2E",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"54",x"45",x"4C",x"2E",x"54",x"4F",x"4B",x"59",x"4F",x"2D",x"4A",x"41",x"50",x"41",x"4E",x"20",
		x"30",x"34",x"34",x"28",x"32",x"34",x"34",x"29",x"32",x"31",x"35",x"31",x"20",x"20",x"20",x"20",
		x"45",x"58",x"54",x"45",x"4E",x"54",x"49",x"4F",x"4E",x"20",x"33",x"30",x"34",x"20",x"20",x"20",
		x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"44",x"45",x"53",x"49",x"47",x"4E",x"20",x"20",x"20",
		x"49",x"4B",x"45",x"47",x"41",x"4D",x"49",x"20",x"43",x"4F",x"2E",x"20",x"4C",x"49",x"4D",x"2E",
		x"CD",x"A6",x"3F",x"C3",x"5F",x"0D",x"3E",x"02",x"F7",x"06",x"02",x"21",x"6C",x"77",x"36",x"10",
		x"23",x"23",x"36",x"C0",x"21",x"8C",x"74",x"10",x"F5",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"4D",x"69",x"36",x"03",x"2C",x"2C",x"C9",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"7F",x"7F",x"18",x"3C",x"76",x"63",x"41",x"00",x"00",x"7F",x"7F",x"49",x"49",x"49",x"41",
		x"00",x"1C",x"3E",x"63",x"41",x"49",x"79",x"79",x"00",x"7C",x"7E",x"13",x"11",x"13",x"7E",x"7C",
		x"00",x"7F",x"7F",x"0E",x"1C",x"0E",x"7F",x"7F",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"17",x"CB",x"13",x"17",x"C6",x"74",x"57",x"19",x"C9",x"57",x"0F",x"DA",x"22",x"30",x"0E",x"93",
		x"0F",x"0F",x"D2",x"17",x"30",x"0E",x"6C",x"07",x"DA",x"31",x"30",x"79",x"E6",x"F0",x"4F",x"C3",
		x"31",x"30",x"0E",x"B4",x"0F",x"0F",x"D2",x"2B",x"30",x"0E",x"1E",x"CB",x"50",x"CA",x"31",x"30",
		x"05",x"79",x"0F",x"0F",x"4F",x"E6",x"03",x"B8",x"C2",x"31",x"30",x"79",x"0F",x"0F",x"E6",x"03",
		x"FE",x"03",x"C0",x"CB",x"92",x"15",x"C0",x"3E",x"04",x"C9",x"11",x"E0",x"FF",x"3A",x"8E",x"63",
		x"4F",x"06",x"00",x"21",x"00",x"76",x"CD",x"64",x"30",x"21",x"C0",x"75",x"CD",x"64",x"30",x"21",
		x"8E",x"63",x"35",x"C9",x"09",x"7E",x"19",x"77",x"C9",x"DF",x"2A",x"C0",x"63",x"34",x"C9",x"21",
		x"AF",x"62",x"34",x"7E",x"E6",x"07",x"C0",x"21",x"0B",x"69",x"0E",x"FC",x"FF",x"0E",x"81",x"21",
		x"09",x"69",x"CD",x"96",x"30",x"21",x"1D",x"69",x"CD",x"96",x"30",x"CD",x"57",x"00",x"E6",x"80",
		x"21",x"2D",x"69",x"AE",x"77",x"C9",x"06",x"02",x"79",x"AE",x"77",x"19",x"10",x"FA",x"C9",x"E5",
		x"21",x"C0",x"60",x"3A",x"B0",x"60",x"6F",x"CB",x"7E",x"CA",x"BB",x"30",x"72",x"2C",x"73",x"2C",
		x"7D",x"FE",x"C0",x"D2",x"B8",x"30",x"3E",x"C0",x"32",x"B0",x"60",x"E1",x"C9",x"21",x"50",x"69",
		x"06",x"02",x"CD",x"E4",x"30",x"2E",x"80",x"06",x"0A",x"CD",x"E4",x"30",x"2E",x"B8",x"06",x"0B",
		x"CD",x"E4",x"30",x"21",x"0C",x"6A",x"06",x"05",x"C3",x"E4",x"30",x"21",x"4C",x"69",x"36",x"00",
		x"2E",x"58",x"06",x"06",x"7D",x"36",x"00",x"C6",x"04",x"6F",x"10",x"F9",x"C9",x"CD",x"FA",x"30",
		x"CD",x"3C",x"31",x"CD",x"B1",x"31",x"CD",x"F3",x"34",x"C9",x"3A",x"80",x"63",x"FE",x"06",x"38",
		x"02",x"3E",x"05",x"EF",x"10",x"31",x"10",x"31",x"1B",x"31",x"26",x"31",x"26",x"31",x"31",x"31",
		x"3A",x"1A",x"60",x"E6",x"01",x"FE",x"01",x"C8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"07",
		x"FE",x"05",x"F8",x"33",x"33",x"C9",x"3A",x"1A",x"60",x"E6",x"03",x"FE",x"03",x"F8",x"33",x"33",
		x"C9",x"3A",x"1A",x"60",x"E6",x"07",x"FE",x"07",x"F8",x"33",x"33",x"C9",x"DD",x"21",x"00",x"64",
		x"AF",x"32",x"A1",x"63",x"06",x"05",x"11",x"20",x"00",x"DD",x"7E",x"00",x"FE",x"00",x"CA",x"7C",
		x"31",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"3E",x"01",x"DD",x"77",x"08",x"3A",x"17",x"62",
		x"FE",x"01",x"C2",x"6A",x"31",x"3E",x"00",x"DD",x"77",x"08",x"DD",x"19",x"10",x"DB",x"21",x"A0",
		x"63",x"36",x"00",x"3A",x"A1",x"63",x"FE",x"00",x"C0",x"33",x"33",x"C9",x"3A",x"A1",x"63",x"FE",
		x"05",x"CA",x"6A",x"31",x"3A",x"27",x"62",x"FE",x"02",x"C2",x"95",x"31",x"3A",x"A1",x"63",x"4F",
		x"3A",x"80",x"63",x"B9",x"C8",x"3A",x"A0",x"63",x"FE",x"01",x"C2",x"6A",x"31",x"DD",x"77",x"00",
		x"DD",x"77",x"18",x"AF",x"32",x"A0",x"63",x"3A",x"A1",x"63",x"3C",x"32",x"A1",x"63",x"C3",x"6A",
		x"31",x"CD",x"DD",x"31",x"AF",x"32",x"A2",x"63",x"21",x"E0",x"63",x"22",x"C8",x"63",x"2A",x"C8",
		x"63",x"01",x"20",x"00",x"09",x"22",x"C8",x"63",x"7E",x"A7",x"CA",x"D0",x"31",x"CD",x"02",x"32",
		x"3A",x"A2",x"63",x"3C",x"32",x"A2",x"63",x"FE",x"05",x"C2",x"BE",x"31",x"C9",x"3A",x"80",x"63",
		x"FE",x"03",x"F8",x"CD",x"F6",x"31",x"FE",x"01",x"C0",x"21",x"39",x"64",x"3E",x"02",x"77",x"21",
		x"79",x"64",x"3E",x"02",x"77",x"C9",x"3A",x"18",x"60",x"E6",x"03",x"FE",x"01",x"C0",x"3A",x"1A",
		x"60",x"C9",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"18",x"FE",x"01",x"CA",x"7A",x"32",x"DD",x"7E",
		x"0D",x"FE",x"04",x"F2",x"30",x"32",x"DD",x"7E",x"19",x"FE",x"02",x"CA",x"7E",x"32",x"CD",x"0F",
		x"33",x"3A",x"18",x"60",x"E6",x"03",x"C2",x"33",x"32",x"DD",x"7E",x"0D",x"A7",x"CA",x"57",x"32",
		x"CD",x"3D",x"33",x"DD",x"7E",x"0D",x"FE",x"04",x"F2",x"91",x"32",x"CD",x"AD",x"33",x"CD",x"8C",
		x"29",x"FE",x"01",x"CA",x"97",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0E",x"FE",x"10",x"DA",
		x"8C",x"32",x"FE",x"F0",x"D2",x"84",x"32",x"DD",x"7E",x"13",x"FE",x"00",x"C2",x"B9",x"32",x"3E",
		x"11",x"DD",x"77",x"13",x"16",x"00",x"5F",x"21",x"7A",x"3A",x"19",x"7E",x"DD",x"46",x"0E",x"DD",
		x"70",x"03",x"DD",x"4E",x"0F",x"81",x"DD",x"77",x"05",x"C9",x"CD",x"BD",x"32",x"C9",x"CD",x"D6",
		x"32",x"C3",x"29",x"32",x"3E",x"02",x"DD",x"77",x"0D",x"C3",x"57",x"32",x"3E",x"01",x"C3",x"86",
		x"32",x"CD",x"E7",x"33",x"C3",x"57",x"32",x"DD",x"2A",x"C8",x"63",x"DD",x"7E",x"0D",x"FE",x"01",
		x"C2",x"B1",x"32",x"3E",x"02",x"DD",x"35",x"0E",x"DD",x"77",x"0D",x"CD",x"C3",x"33",x"C3",x"57",
		x"32",x"3E",x"01",x"DD",x"34",x"0E",x"C3",x"A8",x"32",x"3D",x"C3",x"61",x"32",x"3A",x"27",x"62",
		x"FE",x"01",x"CA",x"CE",x"32",x"FE",x"02",x"CA",x"D2",x"32",x"CD",x"B9",x"34",x"C9",x"CD",x"2C",
		x"34",x"C9",x"CD",x"78",x"34",x"C9",x"DD",x"7E",x"1C",x"FE",x"00",x"C2",x"FD",x"32",x"DD",x"7E",
		x"1D",x"FE",x"01",x"C2",x"0B",x"33",x"DD",x"36",x"1D",x"00",x"3A",x"05",x"62",x"DD",x"46",x"0F",
		x"90",x"DA",x"03",x"33",x"DD",x"36",x"1C",x"FF",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"35",x"1C",
		x"C2",x"F8",x"32",x"DD",x"36",x"19",x"00",x"DD",x"36",x"1C",x"00",x"CD",x"0F",x"33",x"C9",x"DD",
		x"7E",x"16",x"FE",x"00",x"C2",x"32",x"33",x"DD",x"36",x"16",x"2B",x"DD",x"36",x"0D",x"00",x"3A",
		x"18",x"60",x"0F",x"D2",x"32",x"33",x"DD",x"7E",x"0D",x"FE",x"01",x"CA",x"36",x"33",x"DD",x"36",
		x"0D",x"01",x"DD",x"35",x"16",x"C9",x"DD",x"36",x"0D",x"02",x"C3",x"32",x"33",x"DD",x"7E",x"0D",
		x"FE",x"08",x"CA",x"71",x"33",x"FE",x"04",x"CA",x"8A",x"33",x"CD",x"A1",x"33",x"DD",x"7E",x"0F",
		x"C6",x"08",x"57",x"DD",x"7E",x"0E",x"01",x"15",x"00",x"CD",x"6E",x"23",x"A7",x"CA",x"99",x"33",
		x"DD",x"70",x"1F",x"3A",x"05",x"62",x"47",x"DD",x"7E",x"0F",x"90",x"D0",x"DD",x"36",x"0D",x"04",
		x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"DD",
		x"7E",x"19",x"FE",x"02",x"C0",x"DD",x"36",x"1D",x"01",x"C9",x"DD",x"7E",x"0F",x"C6",x"08",x"DD",
		x"46",x"1F",x"B8",x"C0",x"DD",x"36",x"0D",x"00",x"C9",x"DD",x"70",x"1F",x"DD",x"36",x"0D",x"08",
		x"C9",x"3E",x"07",x"F7",x"DD",x"7E",x"0F",x"FE",x"59",x"D0",x"33",x"33",x"C9",x"DD",x"7E",x"0D",
		x"FE",x"01",x"CA",x"D9",x"33",x"DD",x"7E",x"07",x"E6",x"7F",x"DD",x"77",x"07",x"DD",x"35",x"0E",
		x"CD",x"09",x"34",x"3A",x"27",x"62",x"FE",x"01",x"C0",x"DD",x"66",x"0E",x"DD",x"6E",x"0F",x"DD",
		x"46",x"0D",x"CD",x"33",x"23",x"DD",x"75",x"0F",x"C9",x"DD",x"7E",x"07",x"F6",x"80",x"DD",x"77",
		x"07",x"DD",x"34",x"0E",x"C3",x"C0",x"33",x"CD",x"09",x"34",x"DD",x"7E",x"0D",x"FE",x"08",x"C2",
		x"05",x"34",x"DD",x"7E",x"14",x"A7",x"C2",x"01",x"34",x"DD",x"36",x"14",x"02",x"DD",x"35",x"0F",
		x"C9",x"DD",x"35",x"14",x"C9",x"DD",x"34",x"0F",x"C9",x"DD",x"7E",x"15",x"A7",x"C2",x"28",x"34",
		x"DD",x"36",x"15",x"02",x"DD",x"34",x"07",x"DD",x"7E",x"07",x"E6",x"0F",x"FE",x"0F",x"C0",x"DD",
		x"7E",x"07",x"EE",x"02",x"DD",x"77",x"07",x"C9",x"DD",x"35",x"15",x"C9",x"DD",x"6E",x"1A",x"DD",
		x"66",x"1B",x"AF",x"01",x"00",x"00",x"ED",x"4A",x"C2",x"42",x"34",x"21",x"8C",x"3A",x"DD",x"36",
		x"03",x"26",x"DD",x"34",x"03",x"7E",x"FE",x"AA",x"CA",x"56",x"34",x"DD",x"77",x"05",x"23",x"DD",
		x"75",x"1A",x"DD",x"74",x"1B",x"C9",x"AF",x"DD",x"77",x"13",x"DD",x"77",x"18",x"DD",x"77",x"0D",
		x"DD",x"77",x"1C",x"DD",x"7E",x"03",x"DD",x"77",x"0E",x"DD",x"7E",x"05",x"DD",x"77",x"0F",x"DD",
		x"36",x"1A",x"00",x"DD",x"36",x"1B",x"00",x"C9",x"DD",x"6E",x"1A",x"DD",x"66",x"1B",x"AF",x"01",
		x"00",x"00",x"ED",x"4A",x"C2",x"9A",x"34",x"21",x"AC",x"3A",x"3A",x"03",x"62",x"CB",x"7F",x"CA",
		x"A8",x"34",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"03",x"7E",x"DD",x"7E",x"0D",x"FE",x"01",x"C2",
		x"B3",x"34",x"DD",x"34",x"03",x"C3",x"45",x"34",x"DD",x"36",x"0D",x"02",x"DD",x"36",x"03",x"80",
		x"C3",x"9A",x"34",x"DD",x"35",x"03",x"C3",x"45",x"34",x"3A",x"27",x"62",x"FE",x"03",x"C8",x"3A",
		x"03",x"62",x"CB",x"7F",x"C2",x"ED",x"34",x"21",x"C4",x"3A",x"06",x"00",x"3A",x"19",x"60",x"E6",
		x"06",x"4F",x"09",x"7E",x"DD",x"77",x"03",x"DD",x"77",x"0E",x"23",x"7E",x"DD",x"77",x"05",x"DD",
		x"77",x"0F",x"AF",x"DD",x"77",x"0D",x"DD",x"77",x"18",x"DD",x"77",x"1C",x"C9",x"21",x"D4",x"3A",
		x"C3",x"CA",x"34",x"21",x"00",x"64",x"11",x"D0",x"69",x"06",x"05",x"7E",x"A7",x"CA",x"1E",x"35",
		x"2C",x"2C",x"2C",x"7E",x"12",x"3E",x"04",x"85",x"6F",x"1C",x"7E",x"12",x"2C",x"1C",x"7E",x"12",
		x"2D",x"2D",x"2D",x"1C",x"7E",x"12",x"13",x"3E",x"1B",x"85",x"6F",x"10",x"DE",x"C9",x"3E",x"05",
		x"85",x"6F",x"3E",x"04",x"83",x"5F",x"C3",x"17",x"35",x"00",x"00",x"00",x"00",x"01",x"00",x"00",
		x"02",x"00",x"00",x"03",x"00",x"00",x"04",x"00",x"00",x"05",x"00",x"00",x"06",x"00",x"00",x"07",
		x"00",x"00",x"08",x"00",x"00",x"09",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",
		x"00",x"30",x"00",x"00",x"40",x"00",x"00",x"50",x"00",x"00",x"60",x"00",x"00",x"70",x"00",x"00",
		x"80",x"00",x"00",x"90",x"00",x"94",x"77",x"01",x"23",x"24",x"10",x"10",x"00",x"00",x"07",x"06",
		x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3F",x"00",x"50",x"76",x"00",x"F4",x"76",x"96",x"77",x"02",x"1E",x"14",x"10",x"10",x"00",x"00",
		x"06",x"01",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"3F",x"00",x"00",x"61",x"00",x"F6",x"76",x"98",x"77",x"03",x"22",x"14",x"10",x"10",
		x"00",x"00",x"05",x"09",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"59",x"00",x"F8",x"76",x"9A",x"77",x"04",x"24",x"18",
		x"10",x"10",x"00",x"00",x"05",x"00",x"05",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"50",x"50",x"00",x"FA",x"76",x"9C",x"77",x"05",
		x"24",x"18",x"10",x"10",x"00",x"00",x"04",x"03",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"00",x"00",x"43",x"00",x"FC",x"76",x"3B",
		x"5C",x"4B",x"5C",x"5B",x"5C",x"6B",x"5C",x"7B",x"5C",x"8B",x"5C",x"9B",x"5C",x"AB",x"5C",x"BB",
		x"5C",x"CB",x"5C",x"3B",x"6C",x"4B",x"6C",x"5B",x"6C",x"6B",x"6C",x"7B",x"6C",x"8B",x"6C",x"9B",
		x"6C",x"AB",x"6C",x"BB",x"6C",x"CB",x"6C",x"3B",x"7C",x"4B",x"7C",x"5B",x"7C",x"6B",x"7C",x"7B",
		x"7C",x"8B",x"7C",x"9B",x"7C",x"AB",x"7C",x"BB",x"7C",x"CB",x"7C",x"8B",x"36",x"01",x"00",x"98",
		x"36",x"A5",x"36",x"B2",x"36",x"BF",x"36",x"06",x"00",x"CC",x"36",x"08",x"00",x"E6",x"36",x"FD",
		x"36",x"0B",x"00",x"15",x"37",x"1C",x"37",x"30",x"37",x"38",x"37",x"47",x"37",x"5D",x"37",x"73",
		x"37",x"8B",x"37",x"00",x"61",x"22",x"61",x"44",x"61",x"66",x"61",x"88",x"61",x"9E",x"37",x"B6",
		x"37",x"D2",x"37",x"E1",x"37",x"1D",x"00",x"00",x"3F",x"09",x"3F",x"96",x"76",x"17",x"11",x"1D",
		x"15",x"10",x"10",x"1F",x"26",x"15",x"22",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",
		x"10",x"30",x"32",x"31",x"3F",x"94",x"76",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"30",x"33",
		x"31",x"3F",x"80",x"76",x"18",x"19",x"17",x"18",x"10",x"23",x"13",x"1F",x"22",x"15",x"3F",x"9F",
		x"75",x"13",x"22",x"15",x"14",x"19",x"24",x"10",x"10",x"10",x"10",x"3F",x"5E",x"77",x"18",x"1F",
		x"27",x"10",x"18",x"19",x"17",x"18",x"10",x"13",x"11",x"1E",x"10",x"29",x"1F",x"25",x"10",x"17",
		x"15",x"24",x"10",x"FB",x"10",x"3F",x"29",x"77",x"1F",x"1E",x"1C",x"29",x"10",x"01",x"10",x"20",
		x"1C",x"11",x"29",x"15",x"22",x"10",x"12",x"25",x"24",x"24",x"1F",x"1E",x"3F",x"29",x"77",x"01",
		x"10",x"1F",x"22",x"10",x"02",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"23",x"10",x"12",x"25",
		x"24",x"24",x"1F",x"1E",x"3F",x"27",x"76",x"20",x"25",x"23",x"18",x"3F",x"06",x"77",x"1E",x"11",
		x"1D",x"15",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"22",x"11",x"24",x"19",x"1F",x"1E",x"3F",
		x"88",x"76",x"1E",x"11",x"1D",x"15",x"2E",x"3F",x"E9",x"75",x"2D",x"2D",x"2D",x"10",x"10",x"10",
		x"10",x"10",x"10",x"10",x"10",x"10",x"3F",x"0B",x"77",x"11",x"10",x"12",x"10",x"13",x"10",x"14",
		x"10",x"15",x"10",x"16",x"10",x"17",x"10",x"18",x"10",x"19",x"10",x"1A",x"3F",x"0D",x"77",x"1B",
		x"10",x"1C",x"10",x"1D",x"10",x"1E",x"10",x"1F",x"10",x"20",x"10",x"21",x"10",x"22",x"10",x"23",
		x"10",x"24",x"3F",x"0F",x"77",x"25",x"10",x"26",x"10",x"27",x"10",x"28",x"10",x"29",x"10",x"2A",
		x"10",x"2B",x"10",x"2C",x"44",x"45",x"46",x"47",x"48",x"10",x"3F",x"F2",x"76",x"22",x"15",x"17",
		x"19",x"10",x"24",x"19",x"1D",x"15",x"10",x"10",x"30",x"03",x"00",x"31",x"10",x"3F",x"92",x"77",
		x"22",x"11",x"1E",x"1B",x"10",x"10",x"23",x"13",x"1F",x"22",x"15",x"10",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"10",x"10",x"10",x"3F",x"72",x"77",x"29",x"1F",x"25",x"22",x"10",x"1E",x"11",x"1D",
		x"15",x"10",x"27",x"11",x"23",x"10",x"22",x"15",x"17",x"19",x"23",x"24",x"15",x"22",x"15",x"14",
		x"42",x"3F",x"A7",x"76",x"19",x"1E",x"23",x"15",x"22",x"24",x"10",x"13",x"1F",x"19",x"1E",x"10",
		x"3F",x"0A",x"77",x"10",x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10",x"10",x"10",x"10",x"13",
		x"1F",x"19",x"1E",x"3F",x"FC",x"76",x"49",x"4A",x"10",x"1E",x"19",x"1E",x"24",x"15",x"1E",x"14",
		x"1F",x"10",x"10",x"10",x"10",x"3F",x"7C",x"75",x"01",x"09",x"08",x"01",x"3F",x"02",x"97",x"38",
		x"68",x"38",x"02",x"DF",x"54",x"10",x"54",x"02",x"EF",x"6D",x"20",x"6D",x"02",x"DF",x"8E",x"10",
		x"8E",x"02",x"EF",x"AF",x"20",x"AF",x"02",x"DF",x"D0",x"10",x"D0",x"02",x"EF",x"F1",x"10",x"F1",
		x"00",x"53",x"18",x"53",x"54",x"00",x"63",x"18",x"63",x"54",x"00",x"93",x"38",x"93",x"54",x"00",
		x"83",x"54",x"83",x"F1",x"00",x"93",x"54",x"93",x"F1",x"AA",x"8D",x"7D",x"8C",x"6F",x"00",x"7C",
		x"6E",x"00",x"7C",x"6D",x"00",x"7C",x"6C",x"00",x"7C",x"8F",x"7F",x"8E",x"47",x"27",x"08",x"50",
		x"2F",x"A7",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"23",x"07",x"40",
		x"46",x"A9",x"08",x"44",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",x"70",x"08",x"48",
		x"00",x"70",x"0A",x"48",x"6F",x"10",x"09",x"23",x"6F",x"11",x"0A",x"33",x"50",x"34",x"08",x"3C",
		x"00",x"35",x"08",x"3C",x"53",x"32",x"08",x"40",x"63",x"33",x"08",x"40",x"00",x"70",x"08",x"48",
		x"53",x"36",x"08",x"50",x"63",x"37",x"08",x"50",x"6B",x"31",x"08",x"41",x"00",x"70",x"08",x"48",
		x"6A",x"14",x"0A",x"48",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"7F",x"04",x"7F",x"F0",x"10",
		x"F0",x"02",x"DF",x"F2",x"70",x"F8",x"02",x"6F",x"F8",x"10",x"F8",x"AA",x"04",x"DF",x"D0",x"90",
		x"D0",x"02",x"DF",x"DC",x"20",x"D1",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"04",x"DF",x"A8",x"20",
		x"A8",x"04",x"5F",x"B0",x"20",x"B0",x"02",x"DF",x"B0",x"20",x"BB",x"AA",x"04",x"DF",x"88",x"30",
		x"88",x"04",x"DF",x"90",x"B0",x"90",x"02",x"DF",x"9A",x"20",x"8F",x"AA",x"04",x"BF",x"68",x"20",
		x"68",x"04",x"3F",x"70",x"20",x"70",x"02",x"DF",x"6E",x"20",x"79",x"AA",x"02",x"DF",x"58",x"A0",
		x"55",x"AA",x"00",x"70",x"08",x"44",x"2B",x"AC",x"08",x"4C",x"3B",x"AE",x"08",x"4C",x"3B",x"AF",
		x"08",x"3C",x"4B",x"B0",x"07",x"3C",x"4B",x"AD",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"47",x"27",x"08",x"4C",x"2F",x"A7",
		x"08",x"4C",x"3B",x"25",x"08",x"4C",x"00",x"70",x"08",x"44",x"3B",x"23",x"07",x"3C",x"4B",x"2A",
		x"08",x"3C",x"4B",x"2B",x"08",x"4C",x"2B",x"AA",x"08",x"3C",x"2B",x"AB",x"08",x"4C",x"00",x"70",
		x"0A",x"44",x"00",x"70",x"08",x"44",x"4B",x"2C",x"08",x"4C",x"3B",x"2E",x"08",x"4C",x"3B",x"2F",
		x"08",x"3C",x"2B",x"30",x"07",x"3C",x"2B",x"2D",x"08",x"4C",x"00",x"70",x"08",x"44",x"00",x"70",
		x"08",x"44",x"00",x"70",x"08",x"44",x"00",x"70",x"0A",x"44",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",
		x"FE",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"01",x"00",x"01",x"01",x"02",x"02",x"02",x"02",x"03",
		x"03",x"03",x"7F",x"1E",x"4E",x"BB",x"4C",x"D8",x"4E",x"59",x"4E",x"7F",x"BB",x"4D",x"7F",x"47",
		x"27",x"08",x"50",x"2D",x"26",x"08",x"50",x"3B",x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",
		x"24",x"07",x"40",x"4B",x"28",x"08",x"40",x"00",x"70",x"08",x"48",x"30",x"29",x"08",x"44",x"00",
		x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"49",x"A6",x"08",x"50",x"2F",x"A7",x"08",x"50",x"3B",
		x"25",x"08",x"50",x"00",x"70",x"08",x"48",x"3B",x"24",x"07",x"40",x"46",x"A9",x"08",x"44",x"00",
		x"70",x"08",x"48",x"2B",x"A8",x"08",x"40",x"00",x"70",x"08",x"48",x"00",x"70",x"0A",x"48",x"73",
		x"A7",x"88",x"60",x"8B",x"27",x"88",x"60",x"7F",x"25",x"88",x"60",x"00",x"70",x"88",x"68",x"7F",
		x"24",x"87",x"70",x"74",x"29",x"88",x"6C",x"00",x"70",x"88",x"68",x"8A",x"A9",x"88",x"6C",x"00",
		x"70",x"88",x"68",x"00",x"70",x"8A",x"68",x"05",x"AF",x"F0",x"50",x"F0",x"AA",x"05",x"AF",x"E8",
		x"50",x"E8",x"AA",x"05",x"AF",x"E0",x"50",x"E0",x"AA",x"05",x"AF",x"D8",x"50",x"D8",x"AA",x"05",
		x"B7",x"58",x"48",x"58",x"AA",x"01",x"04",x"01",x"03",x"04",x"01",x"02",x"03",x"04",x"01",x"02",
		x"01",x"03",x"04",x"01",x"02",x"01",x"03",x"01",x"04",x"7F",x"FF",x"00",x"FF",x"FF",x"FE",x"FE",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"00",x"E8",x"E5",x"E3",x"E2",
		x"E1",x"E0",x"DF",x"DE",x"DD",x"DD",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DE",x"DF",
		x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E7",x"E9",x"EB",x"ED",x"F0",x"AA",x"80",x"7B",x"78",x"76",
		x"74",x"73",x"72",x"71",x"70",x"70",x"6F",x"6F",x"6F",x"70",x"70",x"71",x"72",x"73",x"74",x"75",
		x"76",x"77",x"78",x"AA",x"EE",x"F0",x"DB",x"A0",x"E6",x"C8",x"D6",x"78",x"EB",x"F0",x"DB",x"A0",
		x"E6",x"C8",x"E6",x"C8",x"1B",x"C8",x"23",x"A0",x"2B",x"78",x"12",x"F0",x"1B",x"C8",x"23",x"A0",
		x"12",x"F0",x"1B",x"C8",x"02",x"97",x"38",x"68",x"38",x"02",x"9F",x"54",x"10",x"54",x"02",x"DF",
		x"58",x"A0",x"55",x"02",x"EF",x"6D",x"20",x"79",x"02",x"DF",x"9A",x"10",x"8E",x"02",x"EF",x"AF",
		x"20",x"BB",x"02",x"DF",x"DC",x"10",x"D0",x"02",x"FF",x"F0",x"80",x"F7",x"02",x"7F",x"F8",x"00",
		x"F8",x"00",x"CB",x"57",x"CB",x"6F",x"00",x"CB",x"99",x"CB",x"B1",x"00",x"CB",x"DB",x"CB",x"F3",
		x"00",x"63",x"18",x"63",x"54",x"01",x"63",x"D5",x"63",x"F8",x"00",x"33",x"78",x"33",x"90",x"00",
		x"33",x"BA",x"33",x"D2",x"00",x"53",x"18",x"53",x"54",x"01",x"53",x"92",x"53",x"B8",x"00",x"5B",
		x"76",x"5B",x"92",x"00",x"73",x"B6",x"73",x"D6",x"00",x"83",x"95",x"83",x"B5",x"00",x"93",x"38",
		x"93",x"54",x"01",x"BB",x"70",x"BB",x"98",x"01",x"6B",x"54",x"6B",x"75",x"AA",x"06",x"8F",x"90",
		x"70",x"90",x"06",x"8F",x"98",x"70",x"98",x"06",x"8F",x"A0",x"70",x"A0",x"00",x"63",x"18",x"63",
		x"58",x"00",x"63",x"80",x"63",x"A8",x"00",x"63",x"D0",x"63",x"F8",x"00",x"53",x"18",x"53",x"58",
		x"00",x"53",x"A8",x"53",x"D0",x"00",x"9B",x"80",x"9B",x"A8",x"00",x"9B",x"D0",x"9B",x"F8",x"01",
		x"23",x"58",x"23",x"80",x"01",x"DB",x"58",x"DB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"A3",x"A8",x"A3",x"D0",x"00",x"2B",x"D0",x"2B",x"F8",x"00",x"D3",x"D0",
		x"D3",x"F8",x"00",x"93",x"38",x"93",x"58",x"02",x"97",x"38",x"68",x"38",x"03",x"EF",x"58",x"10",
		x"58",x"03",x"F7",x"80",x"88",x"80",x"03",x"77",x"80",x"08",x"80",x"02",x"A7",x"A8",x"50",x"A8",
		x"02",x"E7",x"A8",x"B8",x"A8",x"02",x"3F",x"A8",x"18",x"A8",x"03",x"EF",x"D0",x"10",x"D0",x"02",
		x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"63",x"18",x"63",x"58",x"00",x"63",x"88",x"63",x"D0",x"00",
		x"53",x"18",x"53",x"58",x"00",x"53",x"88",x"53",x"D0",x"00",x"E3",x"68",x"E3",x"90",x"00",x"E3",
		x"B8",x"E3",x"D0",x"00",x"CB",x"90",x"CB",x"B0",x"00",x"B3",x"58",x"B3",x"78",x"00",x"9B",x"80",
		x"9B",x"A0",x"00",x"93",x"38",x"93",x"58",x"00",x"23",x"88",x"23",x"C0",x"00",x"1B",x"C0",x"1B",
		x"E8",x"02",x"97",x"38",x"68",x"38",x"02",x"B7",x"58",x"10",x"58",x"02",x"EF",x"68",x"E0",x"68",
		x"02",x"D7",x"70",x"C8",x"70",x"02",x"BF",x"78",x"B0",x"78",x"02",x"A7",x"80",x"90",x"80",x"02",
		x"67",x"88",x"48",x"88",x"02",x"27",x"88",x"10",x"88",x"02",x"EF",x"90",x"C8",x"90",x"02",x"A7",
		x"A0",x"98",x"A0",x"02",x"BF",x"A8",x"B0",x"A8",x"02",x"D7",x"B0",x"C8",x"B0",x"02",x"EF",x"B8",
		x"E0",x"B8",x"02",x"27",x"C0",x"10",x"C0",x"02",x"EF",x"D0",x"D8",x"D0",x"02",x"67",x"D0",x"50",
		x"D0",x"02",x"CF",x"D8",x"C0",x"D8",x"02",x"B7",x"E0",x"A8",x"E0",x"02",x"9F",x"E8",x"88",x"E8",
		x"02",x"27",x"E8",x"10",x"E8",x"02",x"EF",x"F8",x"10",x"F8",x"AA",x"00",x"7B",x"80",x"7B",x"A8",
		x"00",x"7B",x"D0",x"7B",x"F8",x"00",x"33",x"58",x"33",x"80",x"00",x"53",x"58",x"53",x"80",x"00",
		x"AB",x"58",x"AB",x"80",x"00",x"CB",x"58",x"CB",x"80",x"00",x"2B",x"80",x"2B",x"A8",x"00",x"D3",
		x"80",x"D3",x"A8",x"00",x"23",x"A8",x"23",x"D0",x"00",x"5B",x"A8",x"5B",x"D0",x"00",x"A3",x"A8",
		x"A3",x"D0",x"00",x"DB",x"A8",x"DB",x"D0",x"00",x"1B",x"D0",x"1B",x"F8",x"00",x"E3",x"D0",x"E3",
		x"F8",x"05",x"B7",x"30",x"48",x"30",x"05",x"CF",x"58",x"30",x"58",x"05",x"D7",x"80",x"28",x"80",
		x"05",x"DF",x"A8",x"20",x"A8",x"05",x"E7",x"D0",x"18",x"D0",x"05",x"EF",x"F8",x"10",x"F8",x"AA",
		x"10",x"82",x"85",x"8B",x"10",x"85",x"80",x"8B",x"10",x"87",x"85",x"8B",x"81",x"80",x"80",x"8B",
		x"81",x"82",x"85",x"8B",x"81",x"85",x"80",x"8B",x"05",x"88",x"77",x"01",x"68",x"77",x"01",x"6C",
		x"77",x"03",x"49",x"77",x"05",x"08",x"77",x"01",x"E8",x"76",x"01",x"EC",x"76",x"05",x"C8",x"76",
		x"05",x"88",x"76",x"02",x"69",x"76",x"02",x"4A",x"76",x"05",x"28",x"76",x"05",x"E8",x"75",x"01",
		x"CA",x"75",x"03",x"A9",x"75",x"01",x"88",x"75",x"01",x"8C",x"75",x"05",x"48",x"75",x"01",x"28",
		x"75",x"01",x"2A",x"75",x"01",x"2C",x"75",x"01",x"08",x"75",x"01",x"0A",x"75",x"01",x"0C",x"75",
		x"03",x"C8",x"74",x"03",x"AA",x"74",x"03",x"88",x"74",x"05",x"2F",x"77",x"05",x"0F",x"77",x"02",
		x"F0",x"76",x"02",x"CF",x"76",x"02",x"D2",x"76",x"05",x"8F",x"76",x"05",x"6F",x"76",x"01",x"4F",
		x"76",x"01",x"53",x"76",x"05",x"2F",x"76",x"05",x"EF",x"75",x"02",x"D0",x"75",x"02",x"B1",x"75",
		x"05",x"8F",x"75",x"03",x"50",x"75",x"05",x"2F",x"75",x"01",x"0F",x"75",x"01",x"13",x"75",x"01",
		x"EF",x"74",x"01",x"F1",x"74",x"01",x"F3",x"74",x"02",x"D1",x"74",x"00",x"00",x"00",x"23",x"68",
		x"01",x"11",x"00",x"00",x"00",x"10",x"DB",x"68",x"01",x"40",x"00",x"00",x"08",x"01",x"01",x"01",
		x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"01",x"C0",x"FF",
		x"01",x"FF",x"FF",x"34",x"C3",x"39",x"00",x"67",x"80",x"69",x"1A",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"0B",x"4B",
		x"14",x"18",x"0B",x"4B",x"1E",x"18",x"0B",x"3B",x"14",x"18",x"0B",x"3B",x"3D",x"01",x"03",x"02",
		x"4D",x"01",x"04",x"01",x"27",x"70",x"01",x"E0",x"00",x"00",x"7F",x"40",x"01",x"78",x"02",x"00",
		x"27",x"49",x"0C",x"F0",x"7F",x"49",x"0C",x"88",x"1E",x"07",x"03",x"09",x"24",x"64",x"BB",x"C0",
		x"23",x"8D",x"7B",x"B4",x"1B",x"8C",x"7C",x"64",x"4B",x"0E",x"04",x"02",x"23",x"46",x"03",x"68",
		x"DB",x"46",x"03",x"68",x"17",x"50",x"00",x"5C",x"E7",x"D0",x"00",x"5C",x"8C",x"50",x"00",x"84",
		x"73",x"D0",x"00",x"84",x"17",x"50",x"00",x"D4",x"E7",x"D0",x"00",x"D4",x"53",x"73",x"0A",x"A0",
		x"8B",x"74",x"0A",x"F0",x"DB",x"75",x"0A",x"A0",x"5B",x"73",x"0A",x"C8",x"E3",x"74",x"0A",x"60",
		x"1B",x"75",x"0A",x"80",x"DB",x"73",x"0A",x"C8",x"93",x"74",x"0A",x"F0",x"33",x"75",x"0A",x"50",
		x"44",x"03",x"08",x"04",x"37",x"F4",x"37",x"C0",x"37",x"8C",x"77",x"70",x"77",x"A4",x"77",x"D8",
		x"11",x"01",x"00",x"06",x"7B",x"1F",x"D2",x"28",x"1E",x"1E",x"03",x"06",x"7D",x"1F",x"D2",x"28",
		x"1E",x"1E",x"05",x"06",x"7F",x"C3",x"28",x"1E",x"3A",x"27",x"62",x"E5",x"EF",x"00",x"00",x"99",
		x"3E",x"B0",x"28",x"E0",x"28",x"01",x"29",x"00",x"00",x"E1",x"AF",x"32",x"60",x"60",x"06",x"0A",
		x"11",x"20",x"00",x"DD",x"21",x"00",x"67",x"CD",x"C3",x"3E",x"06",x"05",x"DD",x"21",x"00",x"64",
		x"CD",x"C3",x"3E",x"3A",x"60",x"60",x"A7",x"C8",x"FE",x"01",x"C8",x"FE",x"03",x"3E",x"03",x"D8",
		x"3E",x"07",x"C9",x"DD",x"CB",x"00",x"46",x"CA",x"FA",x"3E",x"79",x"DD",x"96",x"05",x"D2",x"D3",
		x"3E",x"ED",x"44",x"3C",x"95",x"DA",x"DE",x"3E",x"DD",x"96",x"0A",x"D2",x"FA",x"3E",x"FD",x"7E",
		x"03",x"DD",x"96",x"03",x"D2",x"E9",x"3E",x"ED",x"44",x"94",x"DA",x"F3",x"3E",x"DD",x"96",x"09",
		x"D2",x"FA",x"3E",x"3A",x"60",x"60",x"3C",x"32",x"60",x"60",x"DD",x"19",x"10",x"C5",x"C9",x"00",
		x"5C",x"76",x"49",x"4A",x"01",x"09",x"08",x"01",x"3F",x"7D",x"77",x"1E",x"19",x"1E",x"24",x"15",
		x"1E",x"14",x"1F",x"10",x"1F",x"16",x"10",x"11",x"1D",x"15",x"22",x"19",x"13",x"11",x"10",x"19",
		x"1E",x"13",x"2B",x"3F",x"21",x"AF",x"74",x"11",x"E0",x"FF",x"36",x"9F",x"19",x"36",x"9E",x"C9",
		x"50",x"52",x"4F",x"47",x"52",x"41",x"4D",x"2C",x"57",x"45",x"20",x"57",x"4F",x"55",x"4C",x"44",
		x"20",x"54",x"45",x"41",x"43",x"48",x"20",x"59",x"4F",x"55",x"2E",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"54",x"45",x"4C",x"2E",x"54",x"4F",x"4B",x"59",x"4F",x"2D",x"4A",x"41",x"50",x"41",x"4E",x"20",
		x"30",x"34",x"34",x"28",x"32",x"34",x"34",x"29",x"32",x"31",x"35",x"31",x"20",x"20",x"20",x"20",
		x"45",x"58",x"54",x"45",x"4E",x"54",x"49",x"4F",x"4E",x"20",x"33",x"30",x"34",x"20",x"20",x"20",
		x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"44",x"45",x"53",x"49",x"47",x"4E",x"20",x"20",x"20",
		x"49",x"4B",x"45",x"47",x"41",x"4D",x"49",x"20",x"43",x"4F",x"2E",x"20",x"4C",x"49",x"4D",x"2E",
		x"CD",x"A6",x"3F",x"C3",x"5F",x"0D",x"3E",x"02",x"F7",x"06",x"02",x"21",x"6C",x"77",x"36",x"10",
		x"23",x"23",x"36",x"C0",x"21",x"8C",x"74",x"10",x"F5",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"4D",x"69",x"36",x"03",x"2C",x"2C",x"C9",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"7F",x"7F",x"18",x"3C",x"76",x"63",x"41",x"00",x"00",x"7F",x"7F",x"49",x"49",x"49",x"41",
		x"00",x"1C",x"3E",x"63",x"41",x"49",x"79",x"79",x"00",x"7C",x"7E",x"13",x"11",x"13",x"7E",x"7C",
		x"00",x"7F",x"7F",x"0E",x"1C",x"0E",x"7F",x"7F",x"00",x"00",x"41",x"7F",x"7F",x"41",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"3F",x"3F",x"3F",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"05",x"1D",x"3D",x"3F",x"3E",x"3E",x"3F",x"3F",x"1E",x"1E",x"1C",x"09",x"01",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"03",x"07",x"07",x"1F",x"3C",x"1F",x"1F",x"1F",x"1F",x"3C",x"FF",x"FF",x"1C",x"00",x"00",
		x"00",x"10",x"30",x"20",x"40",x"60",x"70",x"70",x"60",x"40",x"70",x"30",x"18",x"1C",x"0C",x"00",
		x"00",x"03",x"04",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"01",x"03",x"1B",x"3C",x"1F",x"1F",x"1F",x"1F",x"3C",x"1B",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"FF",x"FF",x"FF",x"3E",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"3F",x"3E",x"3E",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"FF",x"FF",x"FF",x"3E",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3C",x"3F",x"3F",x"3E",x"3E",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"FF",x"FF",x"FF",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"01",x"01",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"05",x"01",
		x"01",x"03",x"07",x"1F",x"3F",x"3F",x"3E",x"3F",x"3F",x"3F",x"1F",x"1F",x"1D",x"09",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"67",x"7F",x"FF",x"FF",x"FF",x"FF",x"9E",x"1C",x"0D",x"09",x"03",x"06",x"04",
		x"01",x"01",x"21",x"6C",x"FE",x"FE",x"FE",x"FF",x"FF",x"BF",x"DE",x"66",x"20",x"00",x"00",x"00",
		x"00",x"00",x"27",x"77",x"DF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"5F",x"77",x"27",x"00",x"00",
		x"00",x"00",x"06",x"0E",x"1D",x"1B",x"1B",x"1B",x"1A",x"1A",x"1B",x"0A",x"03",x"03",x"03",x"01",
		x"00",x"00",x"03",x"04",x"08",x"0A",x"11",x"10",x"10",x"16",x"0E",x"08",x"04",x"03",x"00",x"00",
		x"02",x"0F",x"04",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"04",x"0F",x"02",
		x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",
		x"00",x"00",x"00",x"00",x"4F",x"7F",x"C0",x"40",x"40",x"C0",x"7F",x"4F",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"00",x"00",x"00",
		x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",
		x"02",x"0F",x"04",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"04",x"0F",x"02",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"03",x"03",x"03",x"01",x"00",x"00",x"00",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"00",x"1E",x"36",x"60",x"C0",x"CC",x"ED",x"F1",x"ED",x"CC",x"C0",x"60",x"36",x"1E",x"0E",x"00",
		x"00",x"1E",x"36",x"60",x"C0",x"CC",x"ED",x"F1",x"ED",x"CC",x"C0",x"60",x"36",x"1E",x"0E",x"00",
		x"FE",x"47",x"87",x"14",x"85",x"04",x"89",x"F0",x"F0",x"89",x"04",x"85",x"14",x"87",x"47",x"FE",
		x"00",x"01",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"87",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"00",x"00",x"00",
		x"01",x"0F",x"07",x"0F",x"07",x"23",x"13",x"09",x"51",x"31",x"11",x"01",x"01",x"03",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"11",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"03",x"03",x"01",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"03",x"01",x"01",
		x"00",x"00",x"00",x"00",x"C0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FC",x"F0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"0F",x"1F",x"3F",x"7F",
		x"F4",x"F9",x"FD",x"FE",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E6",x"E2",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F",x"1F",
		x"3C",x"78",x"78",x"FC",x"F7",x"E3",x"E1",x"C0",x"CC",x"4C",x"00",x"04",x"04",x"00",x"00",x"00",
		x"00",x"00",x"01",x"01",x"03",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"0C",x"08",
		x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",
		x"00",x"20",x"5C",x"7F",x"FF",x"7F",x"7F",x"1F",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",x"07",x"07",x"0B",x"00",x"00",x"00",x"00",
		x"FC",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"0E",x"00",x"00",
		x"00",x"1C",x"3E",x"7F",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"10",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"40",x"61",x"63",x"66",x"6C",x"7A",x"7A",x"6C",x"66",x"63",x"61",x"40",x"00",x"00",
		x"00",x"00",x"04",x"06",x"06",x"06",x"06",x"07",x"07",x"06",x"06",x"06",x"06",x"04",x"00",x"00",
		x"00",x"10",x"08",x"00",x"00",x"00",x"00",x"01",x"00",x"21",x"00",x"00",x"04",x"00",x"00",x"00",
		x"08",x"00",x"00",x"00",x"00",x"01",x"23",x"03",x"05",x"01",x"02",x"00",x"10",x"02",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"08",x"00",x"01",x"24",x"00",x"00",x"05",x"08",x"40",x"00",x"00",x"00",x"04",x"00",x"00",x"00",
		x"02",x"08",x"40",x"20",x"04",x"40",x"01",x"04",x"08",x"00",x"02",x"00",x"00",x"00",x"00",x"00",
		x"80",x"10",x"08",x"04",x"06",x"03",x"10",x"2F",x"03",x"01",x"01",x"0A",x"05",x"00",x"00",x"20",
		x"01",x"40",x"00",x"00",x"02",x"01",x"00",x"00",x"01",x"03",x"06",x"00",x"10",x"01",x"00",x"10",
		x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",
		x"F7",x"F7",x"F7",x"F7",x"FB",x"FD",x"CE",x"B6",x"B6",x"CE",x"FD",x"FB",x"F7",x"F7",x"F7",x"F7",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"F7",x"F7",x"F4",x"F4",x"F7",x"F4",x"F4",x"F7",x"F4",x"F5",x"F4",x"F7",x"FF",x"F7",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"01",x"02",x"0A",x"08",x"05",x"00",x"05",x"05",x"02",x"00",x"01",x"00",
		x"0F",x"0F",x"1F",x"1E",x"1E",x"3E",x"3C",x"3C",x"7C",x"78",x"79",x"FE",x"FE",x"70",x"30",x"10",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"06",x"07",x"06",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"06",x"07",x"06",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1F",x"1C",x"1C",x"1E",x"1F",x"0F",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1E",x"1E",x"1E",x"1E",x"1E",x"0E",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1F",x"1F",x"1E",x"1C",x"1C",x"0F",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"20",x"20",x"20",x"20",x"10",x"08",x"04",x"03",x"00",
		x"00",x"00",x"00",x"01",x"02",x"05",x"0A",x"0A",x"0A",x"0A",x"05",x"02",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"05",x"05",x"02",x"01",x"00",x"00",x"00",x"00",x"00",
		x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"00",x"00",x"00",x"00",x"00",x"20",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"00",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"20",x"47",x"1E",x"FE",x"FE",x"1E",x"47",x"20",x"30",x"18",x"0F",x"07",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"00",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1D",x"08",x"02",x"17",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",
		x"03",x"07",x"0F",x"3C",x"3D",x"3E",x"3F",x"3D",x"3D",x"3F",x"3E",x"3D",x"3C",x"0F",x"07",x"03",
		x"00",x"00",x"07",x"0F",x"1F",x"5F",x"E6",x"ED",x"7D",x"08",x"02",x"30",x"38",x"3C",x"3C",x"1C",
		x"20",x"50",x"88",x"88",x"88",x"88",x"88",x"56",x"26",x"0C",x"0C",x"0C",x"0C",x"00",x"00",x"00",
		x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"09",x"0A",x"0A",x"0A",x"0E",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"3F",x"3F",x"3F",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"05",x"1D",x"3D",x"3F",x"3E",x"3E",x"3F",x"3F",x"1E",x"1E",x"1C",x"09",x"01",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"03",x"07",x"07",x"1F",x"3C",x"1F",x"1F",x"1F",x"1F",x"3C",x"FF",x"FF",x"1C",x"00",x"00",
		x"00",x"10",x"30",x"20",x"40",x"60",x"70",x"70",x"60",x"40",x"70",x"30",x"18",x"1C",x"0C",x"00",
		x"00",x"03",x"04",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"01",x"03",x"1B",x"3C",x"1F",x"1F",x"1F",x"1F",x"3C",x"1B",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"FF",x"FF",x"FF",x"3E",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"3F",x"3E",x"3E",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3D",x"3F",x"FF",x"FF",x"FF",x"3E",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"3C",x"3F",x"3F",x"3E",x"3E",x"3F",x"1E",x"1E",x"1C",x"08",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"FF",x"FF",x"FF",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"04",x"00",
		x"00",x"01",x"01",x"02",x"0E",x"1E",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0E",x"05",x"01",
		x"01",x"03",x"07",x"1F",x"3F",x"3F",x"3E",x"3F",x"3F",x"3F",x"1F",x"1F",x"1D",x"09",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"67",x"7F",x"FF",x"FF",x"FF",x"FF",x"9E",x"1C",x"0D",x"09",x"03",x"06",x"04",
		x"01",x"01",x"21",x"6C",x"FE",x"FE",x"FE",x"FF",x"FF",x"BF",x"DE",x"66",x"20",x"00",x"00",x"00",
		x"00",x"00",x"27",x"77",x"DF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"5F",x"77",x"27",x"00",x"00",
		x"00",x"00",x"06",x"0E",x"1D",x"1B",x"1B",x"1B",x"1A",x"1A",x"1B",x"0A",x"03",x"03",x"03",x"01",
		x"00",x"00",x"03",x"04",x"08",x"0A",x"11",x"10",x"10",x"16",x"0E",x"08",x"04",x"03",x"00",x"00",
		x"02",x"0F",x"04",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"04",x"0F",x"02",
		x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",
		x"00",x"00",x"00",x"00",x"4F",x"7F",x"C0",x"40",x"40",x"C0",x"7F",x"4F",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"00",x"00",x"00",
		x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",
		x"02",x"0F",x"04",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"04",x"0F",x"02",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"03",x"03",x"03",x"01",x"00",x"00",x"00",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"1F",x"3F",x"7F",x"FF",x"FF",x"BF",x"9E",x"C1",x"E1",x"C6",x"8F",x"CF",x"E6",x"73",x"1F",x"00",
		x"00",x"1E",x"36",x"60",x"C0",x"CC",x"ED",x"F1",x"ED",x"CC",x"C0",x"60",x"36",x"1E",x"0E",x"00",
		x"00",x"1E",x"36",x"60",x"C0",x"CC",x"ED",x"F1",x"ED",x"CC",x"C0",x"60",x"36",x"1E",x"0E",x"00",
		x"FE",x"47",x"87",x"14",x"85",x"04",x"89",x"F0",x"F0",x"89",x"04",x"85",x"14",x"87",x"47",x"FE",
		x"00",x"01",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"87",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"00",x"00",x"00",
		x"01",x"0F",x"07",x"0F",x"07",x"23",x"13",x"09",x"51",x"31",x"11",x"01",x"01",x"03",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"11",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"03",x"03",x"01",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"03",x"01",x"01",
		x"00",x"00",x"00",x"00",x"C0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FC",x"F0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"0F",x"1F",x"3F",x"7F",
		x"F4",x"F9",x"FD",x"FE",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E6",x"E2",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F",x"1F",
		x"3C",x"78",x"78",x"FC",x"F7",x"E3",x"E1",x"C0",x"CC",x"4C",x"00",x"04",x"04",x"00",x"00",x"00",
		x"00",x"00",x"01",x"01",x"03",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"0C",x"08",
		x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",
		x"00",x"20",x"5C",x"7F",x"FF",x"7F",x"7F",x"1F",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",x"07",x"07",x"0B",x"00",x"00",x"00",x"00",
		x"FC",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"0E",x"00",x"00",
		x"00",x"1C",x"3E",x"7F",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"10",x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"40",x"61",x"63",x"66",x"6C",x"7A",x"7A",x"6C",x"66",x"63",x"61",x"40",x"00",x"00",
		x"00",x"00",x"04",x"06",x"06",x"06",x"06",x"07",x"07",x"06",x"06",x"06",x"06",x"04",x"00",x"00",
		x"00",x"10",x"08",x"00",x"00",x"00",x"00",x"01",x"00",x"21",x"00",x"00",x"04",x"00",x"00",x"00",
		x"08",x"00",x"00",x"00",x"00",x"01",x"23",x"03",x"05",x"01",x"02",x"00",x"10",x"02",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"08",x"00",x"01",x"24",x"00",x"00",x"05",x"08",x"40",x"00",x"00",x"00",x"04",x"00",x"00",x"00",
		x"02",x"08",x"40",x"20",x"04",x"40",x"01",x"04",x"08",x"00",x"02",x"00",x"00",x"00",x"00",x"00",
		x"80",x"10",x"08",x"04",x"06",x"03",x"10",x"2F",x"03",x"01",x"01",x"0A",x"05",x"00",x"00",x"20",
		x"01",x"40",x"00",x"00",x"02",x"01",x"00",x"00",x"01",x"03",x"06",x"00",x"10",x"01",x"00",x"10",
		x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",x"08",x"08",x"09",x"0B",x"0A",x"0B",x"09",x"08",
		x"F7",x"F7",x"F7",x"F7",x"FB",x"FD",x"CE",x"B6",x"B6",x"CE",x"FD",x"FB",x"F7",x"F7",x"F7",x"F7",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"F7",x"F7",x"F4",x"F4",x"F7",x"F4",x"F4",x"F7",x"F4",x"F5",x"F4",x"F7",x"FF",x"F7",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"01",x"02",x"0A",x"08",x"05",x"00",x"05",x"05",x"02",x"00",x"01",x"00",
		x"0F",x"0F",x"1F",x"1E",x"1E",x"3E",x"3C",x"3C",x"7C",x"78",x"79",x"FE",x"FE",x"70",x"30",x"10",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"06",x"07",x"06",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"06",x"07",x"06",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1F",x"1C",x"1C",x"1E",x"1F",x"0F",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1E",x"1E",x"1E",x"1E",x"1E",x"0E",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"1F",x"1F",x"1F",x"1E",x"1C",x"1C",x"0F",x"0F",x"07",x"03",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"20",x"20",x"20",x"20",x"10",x"08",x"04",x"03",x"00",
		x"00",x"00",x"00",x"01",x"02",x"05",x"0A",x"0A",x"0A",x"0A",x"05",x"02",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"05",x"05",x"02",x"01",x"00",x"00",x"00",x"00",x"00",
		x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"00",x"00",x"00",x"00",x"00",x"20",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"00",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"20",x"47",x"1E",x"FE",x"FE",x"1E",x"47",x"20",x"30",x"18",x"0F",x"07",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"00",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1D",x"08",x"02",x"17",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",
		x"03",x"07",x"0F",x"3C",x"3D",x"3E",x"3F",x"3D",x"3D",x"3F",x"3E",x"3D",x"3C",x"0F",x"07",x"03",
		x"00",x"00",x"07",x"0F",x"1F",x"5F",x"E6",x"ED",x"7D",x"08",x"02",x"30",x"38",x"3C",x"3C",x"1C",
		x"20",x"50",x"88",x"88",x"88",x"88",x"88",x"56",x"26",x"0C",x"0C",x"0C",x"0C",x"00",x"00",x"00",
		x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"09",x"0A",x"0A",x"0A",x"0E",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00",
		x"00",x"00",x"00",x"E3",x"F3",x"FB",x"B9",x"10",x"43",x"83",x"83",x"01",x"00",x"00",x"00",x"00",
		x"E0",x"E6",x"C7",x"87",x"C1",x"C0",x"00",x"40",x"00",x"80",x"80",x"C0",x"DC",x"FC",x"C0",x"00",
		x"1E",x"1C",x"20",x"60",x"C0",x"C0",x"E0",x"E3",x"E3",x"63",x"61",x"E0",x"40",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"07",x"07",x"87",x"83",x"0B",x"08",x"08",x"08",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"06",x"0F",x"0F",x"0F",x"37",x"33",x"30",x"20",x"00",x"00",x"00",x"00",
		x"C0",x"C0",x"00",x"00",x"0C",x"0E",x"0E",x"06",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"60",x"E0",x"E0",x"81",x"01",x"01",x"81",x"C1",x"C1",x"81",x"01",x"01",x"81",x"E0",x"E0",x"60",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"03",x"C3",x"C3",x"C1",x"80",x"43",x"03",x"83",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"C3",x"E3",x"E3",x"C1",x"C0",x"C3",x"C3",x"C3",x"C1",x"E0",x"E0",x"E0",x"C0",
		x"00",x"06",x"07",x"03",x"C1",x"C0",x"C0",x"00",x"40",x"00",x"00",x"00",x"1C",x"3C",x"00",x"00",
		x"00",x"06",x"07",x"03",x"C1",x"E0",x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FC",x"FC",x"E0",x"C0",
		x"1E",x"1C",x"00",x"00",x"C0",x"C0",x"E0",x"E3",x"C3",x"A3",x"81",x"00",x"00",x"00",x"00",x"00",
		x"1E",x"1C",x"00",x"00",x"C0",x"C0",x"E0",x"E3",x"E3",x"63",x"E1",x"60",x"60",x"E0",x"E0",x"C0",
		x"84",x"8C",x"D8",x"9C",x"C8",x"E0",x"E0",x"00",x"20",x"80",x"C0",x"40",x"40",x"C0",x"CC",x"9C",
		x"C1",x"E5",x"42",x"82",x"C1",x"C0",x"80",x"41",x"03",x"87",x"8E",x"8D",x"83",x"C6",x"CC",x"C0",
		x"00",x"20",x"70",x"58",x"7B",x"7F",x"1F",x"2F",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"08",x"A8",x"B8",x"B0",x"38",x"60",x"40",x"C0",x"80",x"D0",x"F0",x"E0",x"40",x"00",
		x"80",x"40",x"E0",x"F0",x"E0",x"C0",x"40",x"40",x"40",x"68",x"78",x"F8",x"D0",x"40",x"00",x"00",
		x"00",x"40",x"40",x"68",x"38",x"20",x"B8",x"A0",x"A0",x"B8",x"B0",x"38",x"68",x"40",x"40",x"00",
		x"40",x"C0",x"DC",x"FF",x"FF",x"C7",x"02",x"00",x"00",x"00",x"00",x"E0",x"F0",x"F0",x"60",x"00",
		x"00",x"00",x"C0",x"20",x"10",x"10",x"08",x"88",x"48",x"08",x"10",x"10",x"20",x"C0",x"00",x"00",
		x"40",x"F0",x"20",x"20",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"20",x"20",x"F0",x"40",
		x"A0",x"F0",x"D0",x"D8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"D8",x"D0",x"F0",x"A0",
		x"00",x"00",x"00",x"00",x"F2",x"FE",x"03",x"02",x"02",x"03",x"FF",x"F2",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"C0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0",x"C0",x"00",x"00",x"00",
		x"A0",x"F0",x"D0",x"D8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"D8",x"D0",x"F0",x"A0",
		x"40",x"F0",x"20",x"20",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"20",x"20",x"F0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"02",x"08",x"04",x"02",x"F8",x"FC",x"FC",x"FC",x"FC",x"FC",x"FA",x"02",x"0A",x"14",x"02",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"1F",x"27",x"47",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"47",x"27",x"1F",x"1F",
		x"6F",x"F7",x"F7",x"73",x"7B",x"7B",x"7B",x"73",x"7B",x"7B",x"7B",x"73",x"F7",x"F7",x"67",x"0F",
		x"00",x"00",x"C0",x"C0",x"40",x"C0",x"C0",x"40",x"C0",x"40",x"C0",x"40",x"C0",x"C0",x"00",x"00",
		x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"F8",x"F8",x"F8",x"F4",x"F0",x"F0",x"28",x"00",x"00",x"00",
		x"00",x"01",x"02",x"E4",x"F8",x"FA",x"FC",x"FC",x"FC",x"F8",x"FA",x"FC",x"F8",x"F8",x"30",x"20",
		x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",
		x"00",x"05",x"02",x"07",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FC",x"F8",x"F0",
		x"00",x"00",x"00",x"00",x"03",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"60",x"B0",x"40",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"78",x"00",x"CC",x"F8",x"FE",x"FD",x"FC",x"F9",x"F8",x"F8",x"F8",
		x"FC",x"F8",x"FC",x"FC",x"32",x"84",x"C3",x"F0",x"F8",x"F0",x"F0",x"A0",x"04",x"02",x"00",x"00",
		x"F8",x"F8",x"F8",x"F0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E6",x"FC",x"78",x"F8",x"FC",
		x"00",x"01",x"07",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"3F",x"9F",x"CF",x"E3",x"C1",x"80",x"08",x"10",x"20",x"20",x"20",x"20",x"20",x"00",
		x"60",x"F0",x"F8",x"FC",x"FC",x"FE",x"FC",x"EC",x"CE",x"CE",x"C0",x"C0",x"E0",x"E0",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0B",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"FF",x"FE",x"FC",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F8",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"18",x"30",x"F6",x"F7",x"F7",x"F3",x"FB",x"F9",x"FC",x"E4",x"C2",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"90",x"30",x"70",x"F0",x"F0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"49",x"2A",x"08",x"7E",x"08",x"2A",x"49",x"80",x"00",x"02",x"09",x"80",x"08",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"81",x"C3",x"E3",x"33",x"1B",x"AF",x"AF",x"1B",x"33",x"E3",x"C3",x"81",x"00",x"00",
		x"20",x"70",x"71",x"53",x"DB",x"8B",x"8B",x"FF",x"FF",x"8B",x"8B",x"DB",x"53",x"71",x"70",x"20",
		x"00",x"00",x"00",x"00",x"00",x"78",x"FC",x"CC",x"FC",x"FC",x"CC",x"78",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"78",x"FC",x"FE",x"CE",x"FE",x"FE",x"CC",x"FC",x"78",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"18",x"38",x"9F",x"37",x"25",x"09",x"5E",x"17",x"0E",x"10",x"21",x"0F",x"13",x"04",x"00",
		x"00",x"00",x"00",x"07",x"13",x"03",x"38",x"7F",x"07",x"00",x"02",x"43",x"07",x"06",x"10",x"00",
		x"20",x"04",x"02",x"0B",x"37",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"13",x"21",x"42",x"00",
		x"00",x"00",x"03",x"03",x"7F",x"FF",x"7F",x"7F",x"FF",x"FF",x"7F",x"7F",x"8D",x"00",x"22",x"00",
		x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",
		x"FE",x"FF",x"FF",x"83",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"83",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"DF",x"5F",x"5F",x"5F",x"DF",x"5F",x"5F",x"DF",x"5F",x"5F",x"5F",x"DF",x"FF",x"DF",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"60",x"70",x"70",x"70",x"70",x"F0",x"70",x"70",x"70",x"F0",x"70",x"70",x"F0",x"70",x"70",x"E0",
		x"00",x"00",x"20",x"70",x"10",x"00",x"00",x"20",x"70",x"A8",x"F4",x"52",x"7A",x"34",x"00",x"00",
		x"00",x"20",x"10",x"08",x"0C",x"DE",x"FE",x"FE",x"FE",x"7C",x"F8",x"78",x"F0",x"80",x"00",x"00",
		x"00",x"00",x"10",x"08",x"08",x"FC",x"FC",x"FE",x"FE",x"7E",x"FE",x"7E",x"FC",x"98",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"78",x"38",x"38",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"78",x"78",x"78",x"78",x"78",x"70",x"70",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"F8",x"38",x"38",x"78",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C0",x"20",x"10",x"08",x"04",x"04",x"04",x"04",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",
		x"00",x"00",x"00",x"80",x"40",x"A0",x"50",x"50",x"50",x"50",x"A0",x"40",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"A0",x"A0",x"40",x"80",x"00",x"00",x"00",x"00",x"00",
		x"82",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"9A",x"00",x"00",x"00",x"00",x"00",x"84",x"82",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"04",x"02",x"84",x"54",x"12",x"12",x"12",x"12",x"14",x"14",x"14",x"12",x"02",x"02",x"04",x"00",
		x"00",x"00",x"00",x"00",x"DE",x"2E",x"76",x"6A",x"6A",x"6A",x"76",x"2E",x"DE",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"80",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FC",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"F4",x"E0",x"4A",x"1C",x"B8",x"F0",x"F0",x"E0",x"C0",x"00",
		x"38",x"BC",x"9C",x"CC",x"80",x"40",x"00",x"80",x"80",x"00",x"46",x"86",x"CE",x"8C",x"8C",x"00",
		x"00",x"00",x"F0",x"F8",x"FC",x"FE",x"33",x"DF",x"DE",x"88",x"20",x"03",x"07",x"0F",x"0E",x"0C",
		x"00",x"00",x"1F",x"7F",x"FF",x"7F",x"3F",x"2F",x"5E",x"0F",x"47",x"07",x"07",x"0F",x"07",x"03",
		x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"40",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",
		x"00",x"00",x"00",x"E3",x"F3",x"FB",x"B9",x"10",x"43",x"83",x"83",x"01",x"00",x"00",x"00",x"00",
		x"E0",x"E6",x"C7",x"87",x"C1",x"C0",x"00",x"40",x"00",x"80",x"80",x"C0",x"DC",x"FC",x"C0",x"00",
		x"1E",x"1C",x"20",x"60",x"C0",x"C0",x"E0",x"E3",x"E3",x"63",x"61",x"E0",x"40",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"07",x"07",x"87",x"83",x"0B",x"08",x"08",x"08",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"06",x"0F",x"0F",x"0F",x"37",x"33",x"30",x"20",x"00",x"00",x"00",x"00",
		x"C0",x"C0",x"00",x"00",x"0C",x"0E",x"0E",x"06",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"00",
		x"60",x"E0",x"E0",x"81",x"01",x"01",x"81",x"C1",x"C1",x"81",x"01",x"01",x"81",x"E0",x"E0",x"60",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"03",x"C3",x"C3",x"C1",x"80",x"43",x"03",x"83",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"C3",x"E3",x"E3",x"C1",x"C0",x"C3",x"C3",x"C3",x"C1",x"E0",x"E0",x"E0",x"C0",
		x"00",x"06",x"07",x"03",x"C1",x"C0",x"C0",x"00",x"40",x"00",x"00",x"00",x"1C",x"3C",x"00",x"00",
		x"00",x"06",x"07",x"03",x"C1",x"E0",x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FC",x"FC",x"E0",x"C0",
		x"1E",x"1C",x"00",x"00",x"C0",x"C0",x"E0",x"E3",x"C3",x"A3",x"81",x"00",x"00",x"00",x"00",x"00",
		x"1E",x"1C",x"00",x"00",x"C0",x"C0",x"E0",x"E3",x"E3",x"63",x"E1",x"60",x"60",x"E0",x"E0",x"C0",
		x"84",x"8C",x"D8",x"9C",x"C8",x"E0",x"E0",x"00",x"20",x"80",x"C0",x"40",x"40",x"C0",x"CC",x"9C",
		x"C1",x"E5",x"42",x"82",x"C1",x"C0",x"80",x"41",x"03",x"87",x"8E",x"8D",x"83",x"C6",x"CC",x"C0",
		x"00",x"20",x"70",x"58",x"7B",x"7F",x"1F",x"2F",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"08",x"A8",x"B8",x"B0",x"38",x"60",x"40",x"C0",x"80",x"D0",x"F0",x"E0",x"40",x"00",
		x"80",x"40",x"E0",x"F0",x"E0",x"C0",x"40",x"40",x"40",x"68",x"78",x"F8",x"D0",x"40",x"00",x"00",
		x"00",x"40",x"40",x"68",x"38",x"20",x"B8",x"A0",x"A0",x"B8",x"B0",x"38",x"68",x"40",x"40",x"00",
		x"40",x"C0",x"DC",x"FF",x"FF",x"C7",x"02",x"00",x"00",x"00",x"00",x"E0",x"F0",x"F0",x"60",x"00",
		x"00",x"00",x"C0",x"20",x"10",x"10",x"08",x"88",x"48",x"08",x"10",x"10",x"20",x"C0",x"00",x"00",
		x"40",x"F0",x"20",x"20",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"20",x"20",x"F0",x"40",
		x"A0",x"F0",x"D0",x"D8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"D8",x"D0",x"F0",x"A0",
		x"00",x"00",x"00",x"00",x"F2",x"FE",x"03",x"02",x"02",x"03",x"FF",x"F2",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"C0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0",x"C0",x"00",x"00",x"00",
		x"A0",x"F0",x"D0",x"D8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"D8",x"D0",x"F0",x"A0",
		x"40",x"F0",x"20",x"20",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"20",x"20",x"F0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"02",x"08",x"04",x"02",x"F8",x"FC",x"FC",x"FC",x"FC",x"FC",x"FA",x"02",x"0A",x"14",x"02",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"33",x"39",x"78",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"3D",x"19",x"03",
		x"1F",x"27",x"47",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"43",x"47",x"27",x"1F",x"1F",
		x"6F",x"F7",x"F7",x"73",x"7B",x"7B",x"7B",x"73",x"7B",x"7B",x"7B",x"73",x"F7",x"F7",x"67",x"0F",
		x"00",x"00",x"C0",x"C0",x"40",x"C0",x"C0",x"40",x"C0",x"40",x"C0",x"40",x"C0",x"C0",x"00",x"00",
		x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"F8",x"F8",x"F8",x"F4",x"F0",x"F0",x"28",x"00",x"00",x"00",
		x"00",x"01",x"02",x"E4",x"F8",x"FA",x"FC",x"FC",x"FC",x"F8",x"FA",x"FC",x"F8",x"F8",x"30",x"20",
		x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",
		x"00",x"05",x"02",x"07",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FC",x"F8",x"F0",
		x"00",x"00",x"00",x"00",x"03",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"60",x"B0",x"40",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"78",x"00",x"CC",x"F8",x"FE",x"FD",x"FC",x"F9",x"F8",x"F8",x"F8",
		x"FC",x"F8",x"FC",x"FC",x"32",x"84",x"C3",x"F0",x"F8",x"F0",x"F0",x"A0",x"04",x"02",x"00",x"00",
		x"F8",x"F8",x"F8",x"F0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E6",x"FC",x"78",x"F8",x"FC",
		x"00",x"01",x"07",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"3F",x"9F",x"CF",x"E3",x"C1",x"80",x"08",x"10",x"20",x"20",x"20",x"20",x"20",x"00",
		x"60",x"F0",x"F8",x"FC",x"FC",x"FE",x"FC",x"EC",x"CE",x"CE",x"C0",x"C0",x"E0",x"E0",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0B",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"FF",x"FE",x"FC",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F8",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"18",x"30",x"F6",x"F7",x"F7",x"F3",x"FB",x"F9",x"FC",x"E4",x"C2",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"90",x"30",x"70",x"F0",x"F0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"49",x"2A",x"08",x"7E",x"08",x"2A",x"49",x"80",x"00",x"02",x"09",x"80",x"08",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"81",x"C3",x"E3",x"33",x"1B",x"AF",x"AF",x"1B",x"33",x"E3",x"C3",x"81",x"00",x"00",
		x"20",x"70",x"71",x"53",x"DB",x"8B",x"8B",x"FF",x"FF",x"8B",x"8B",x"DB",x"53",x"71",x"70",x"20",
		x"00",x"00",x"00",x"00",x"00",x"78",x"FC",x"CC",x"FC",x"FC",x"CC",x"78",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"78",x"FC",x"FE",x"CE",x"FE",x"FE",x"CC",x"FC",x"78",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"18",x"38",x"9F",x"37",x"25",x"09",x"5E",x"17",x"0E",x"10",x"21",x"0F",x"13",x"04",x"00",
		x"00",x"00",x"00",x"07",x"13",x"03",x"38",x"7F",x"07",x"00",x"02",x"43",x"07",x"06",x"10",x"00",
		x"20",x"04",x"02",x"0B",x"37",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"13",x"21",x"42",x"00",
		x"00",x"00",x"03",x"03",x"7F",x"FF",x"7F",x"7F",x"FF",x"FF",x"7F",x"7F",x"8D",x"00",x"22",x"00",
		x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",x"60",x"E0",x"A0",x"20",x"20",x"20",x"A0",x"E0",
		x"FE",x"FF",x"FF",x"83",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"BB",x"83",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"DF",x"5F",x"5F",x"5F",x"DF",x"5F",x"5F",x"DF",x"5F",x"5F",x"5F",x"DF",x"FF",x"DF",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"60",x"70",x"70",x"70",x"70",x"F0",x"70",x"70",x"70",x"F0",x"70",x"70",x"F0",x"70",x"70",x"E0",
		x"00",x"00",x"20",x"70",x"10",x"00",x"00",x"20",x"70",x"A8",x"F4",x"52",x"7A",x"34",x"00",x"00",
		x"00",x"20",x"10",x"08",x"0C",x"DE",x"FE",x"FE",x"FE",x"7C",x"F8",x"78",x"F0",x"80",x"00",x"00",
		x"00",x"00",x"10",x"08",x"08",x"FC",x"FC",x"FE",x"FE",x"7E",x"FE",x"7E",x"FC",x"98",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"78",x"38",x"38",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"78",x"78",x"78",x"78",x"78",x"70",x"70",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"F8",x"F8",x"F8",x"38",x"38",x"78",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C0",x"20",x"10",x"08",x"04",x"04",x"04",x"04",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",
		x"00",x"00",x"00",x"80",x"40",x"A0",x"50",x"50",x"50",x"50",x"A0",x"40",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"A0",x"A0",x"40",x"80",x"00",x"00",x"00",x"00",x"00",
		x"82",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"9A",x"00",x"00",x"00",x"00",x"00",x"84",x"82",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"04",x"02",x"84",x"54",x"12",x"12",x"12",x"12",x"14",x"14",x"14",x"12",x"02",x"02",x"04",x"00",
		x"00",x"00",x"00",x"00",x"DE",x"2E",x"76",x"6A",x"6A",x"6A",x"76",x"2E",x"DE",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"02",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"80",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FC",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"F4",x"E0",x"4A",x"1C",x"B8",x"F0",x"F0",x"E0",x"C0",x"00",
		x"38",x"BC",x"9C",x"CC",x"80",x"40",x"00",x"80",x"80",x"00",x"46",x"86",x"CE",x"8C",x"8C",x"00",
		x"00",x"00",x"F0",x"F8",x"FC",x"FE",x"33",x"DF",x"DE",x"88",x"20",x"03",x"07",x"0F",x"0E",x"0C",
		x"00",x"00",x"1F",x"7F",x"FF",x"7F",x"3F",x"2F",x"5E",x"0F",x"47",x"07",x"07",x"0F",x"07",x"03",
		x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"40",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"05",x"1D",x"65",x"E1",x"F9",x"D9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"03",x"07",x"07",x"1F",x"7B",x"7B",x"7B",x"7B",x"7B",x"7B",x"3F",x"3F",x"1C",x"00",x"00",
		x"00",x"07",x"1F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"7F",x"7F",x"3F",x"1F",x"03",x"00",x"00",
		x"00",x"03",x"07",x"07",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"07",x"03",
		x"00",x"00",x"01",x"03",x"1B",x"7B",x"7B",x"7B",x"7B",x"7B",x"7B",x"1B",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E3",x"1F",x"1F",x"1F",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E7",x"1F",x"1F",x"1F",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"64",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"71",x"1F",x"1F",x"1F",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"01",x"03",x"07",x"1F",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4D",x"45",x"05",x"01",x"00",x"00",
		x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"40",x"6C",x"6F",x"7F",x"FF",x"DF",x"DF",x"DF",x"9F",x"1F",x"0F",x"0F",x"07",x"06",x"04",
		x"01",x"01",x"3B",x"7F",x"FF",x"BF",x"BF",x"BF",x"BF",x"BF",x"DF",x"67",x"31",x"10",x"10",x"00",
		x"10",x"10",x"3F",x"77",x"DF",x"BF",x"BF",x"BF",x"BF",x"BF",x"FF",x"5F",x"77",x"3F",x"10",x"10",
		x"00",x"01",x"07",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"06",x"06",x"03",x"01",
		x"00",x"00",x"03",x"07",x"0F",x"0D",x"1E",x"1F",x"1F",x"19",x"09",x"0F",x"07",x"03",x"00",x"00",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"00",x"00",x"00",x"1F",x"3F",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF",x"3F",x"1F",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"0C",x"1B",x"1A",x"19",x"18",x"0C",x"0F",x"07",x"03",x"00",x"00",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"1E",x"3F",x"3F",x"3F",x"7D",x"7F",x"3E",x"1E",x"3F",x"7D",x"3F",x"1F",x"0C",x"00",x"0F",
		x"00",x"1E",x"3F",x"3F",x"3F",x"6F",x"7F",x"3E",x"1E",x"3F",x"7F",x"3F",x"1B",x"0C",x"00",x"0F",
		x"00",x"1E",x"3B",x"3F",x"3F",x"7F",x"7F",x"3E",x"1E",x"3F",x"77",x"3F",x"1F",x"0C",x"00",x"0F",
		x"0F",x"01",x"09",x"1F",x"3F",x"3F",x"1A",x"0E",x"1A",x"3F",x"3F",x"1F",x"09",x"01",x"01",x"0F",
		x"0F",x"01",x"09",x"1F",x"3F",x"3F",x"1A",x"0E",x"1A",x"3F",x"3F",x"1F",x"09",x"01",x"01",x"0F",
		x"38",x"FC",x"FF",x"EF",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF",x"FF",x"EF",x"FF",x"FC",x"38",
		x"00",x"00",x"09",x"00",x"00",x"08",x"08",x"08",x"08",x"04",x"04",x"03",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"08",x"00",x"00",x"48",x"B4",x"00",x"00",x"00",x"00",
		x"00",x"00",x"38",x"3C",x"7C",x"7F",x"FF",x"FC",x"FC",x"FC",x"78",x"20",x"00",x"00",x"06",x"0E",
		x"00",x"00",x"00",x"00",x"00",x"EE",x"60",x"00",x"10",x"08",x"08",x"04",x"02",x"02",x"01",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"06",x"04",x"04",x"01",x"06",x"0E",
		x"00",x"00",x"00",x"00",x"C0",x"78",x"00",x"00",x"00",x"00",x"00",x"17",x"E7",x"87",x"06",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"40",
		x"0F",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"03",x"87",x"C7",x"7F",x"3F",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"04",x"08",x"09",x"09",x"08",x"10",x"10",x"10",
		x"03",x"07",x"07",x"03",x"08",x"1C",x"1E",x"3F",x"3F",x"3B",x"1F",x"03",x"03",x"03",x"01",x"00",
		x"00",x"00",x"01",x"01",x"02",x"02",x"02",x"04",x"04",x"04",x"08",x"08",x"08",x"08",x"08",x"08",
		x"00",x"80",x"C0",x"40",x"61",x"3A",x"0E",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"0A",x"32",x"41",x"40",x"80",x"00",x"00",
		x"60",x"F0",x"A0",x"80",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"0E",x"08",x"00",x"00",
		x"0C",x"0C",x"06",x"06",x"06",x"04",x"08",x"10",x"20",x"00",x"80",x"60",x"18",x"0C",x"00",x"00",
		x"00",x"18",x"20",x"40",x"80",x"00",x"00",x"21",x"11",x"09",x"04",x"04",x"06",x"06",x"06",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"01",x"03",x"06",x"0C",x"15",x"15",x"0C",x"06",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"44",x"02",x"01",x"05",x"43",x"0F",x"16",x"03",x"0E",x"5B",x"21",x"00",x"00",x"00",x"00",
		x"00",x"00",x"28",x"87",x"33",x"1E",x"0C",x"44",x"32",x"1E",x"0D",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"12",x"01",x"00",x"22",x"00",x"02",x"40",x"10",x"02",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"00",x"20",x"00",x"43",x"10",x"00",x"00",x"40",x"21",x"02",x"00",x"00",x"00",x"00",
		x"80",x"0A",x"75",x"1A",x"09",x"04",x"2F",x"50",x"9C",x"0E",x"06",x"35",x"4A",x"07",x"00",x"20",
		x"08",x"80",x"00",x"00",x"09",x"86",x"40",x"01",x"02",x"14",x"09",x"00",x"01",x"A6",x"43",x"00",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",
		x"0D",x"2D",x"0D",x"2F",x"07",x"03",x"31",x"79",x"79",x"31",x"03",x"07",x"2F",x"0D",x"2D",x"0D",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"7F",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"03",x"01",x"06",x"0D",x"05",x"07",x"02",x"07",x"02",x"02",x"01",x"01",x"00",x"00",
		x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"7F",x"7F",x"7E",x"F9",x"F8",x"70",x"30",x"10",
		x"02",x"00",x"05",x"02",x"01",x"03",x"06",x"04",x"09",x"09",x"09",x"09",x"0C",x"06",x"03",x"00",
		x"00",x"00",x"01",x"00",x"01",x"03",x"06",x"04",x"09",x"09",x"09",x"09",x"0D",x"06",x"03",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"30",x"30",x"30",x"30",x"18",x"0C",x"07",x"03",x"00",
		x"00",x"00",x"00",x"01",x"03",x"06",x"0C",x"0C",x"0C",x"0C",x"06",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"06",x"06",x"03",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"20",x"10",x"08",x"04",x"00",x"00",x"00",x"38",x"00",x"00",x"04",x"08",x"10",x"20",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"7F",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"7F",x"00",
		x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"00",x"00",x"00",
		x"07",x"0F",x"1E",x"3F",x"3F",x"7F",x"7E",x"7E",x"7F",x"7E",x"7F",x"3F",x"3F",x"1E",x"0F",x"07",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"00",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1D",x"08",x"02",x"17",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",
		x"00",x"01",x"0D",x"1C",x"61",x"C9",x"ED",x"C7",x"C7",x"ED",x"C9",x"61",x"9C",x"0D",x"01",x"00",
		x"03",x"07",x"05",x"08",x"1B",x"19",x"05",x"3F",x"3F",x"0F",x"05",x"37",x"3F",x"3F",x"3E",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"0C",x"0E",x"0F",x"0F",x"07",x"03",x"00",
		x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"09",x"0A",x"0A",x"0A",x"0E",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"05",x"1D",x"65",x"E1",x"F9",x"D9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"03",x"07",x"07",x"1F",x"7B",x"7B",x"7B",x"7B",x"7B",x"7B",x"3F",x"3F",x"1C",x"00",x"00",
		x"00",x"07",x"1F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"7F",x"7F",x"3F",x"1F",x"03",x"00",x"00",
		x"00",x"03",x"07",x"07",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"07",x"03",
		x"00",x"00",x"01",x"03",x"1B",x"7B",x"7B",x"7B",x"7B",x"7B",x"7B",x"1B",x"03",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E3",x"1F",x"1F",x"1F",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"65",x"E7",x"1F",x"1F",x"1F",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"64",x"E1",x"F9",x"E9",x"C1",x"55",x"4C",x"44",x"04",x"00",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"71",x"1F",x"1F",x"1F",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"00",x"00",x"00",x"02",x"0E",x"32",x"70",x"7C",x"74",x"60",x"2A",x"26",x"22",x"02",x"00",x"00",
		x"01",x"03",x"07",x"1F",x"65",x"E1",x"F9",x"E9",x"C1",x"55",x"4D",x"45",x"05",x"01",x"00",x"00",
		x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"40",x"6C",x"6F",x"7F",x"FF",x"DF",x"DF",x"DF",x"9F",x"1F",x"0F",x"0F",x"07",x"06",x"04",
		x"01",x"01",x"3B",x"7F",x"FF",x"BF",x"BF",x"BF",x"BF",x"BF",x"DF",x"67",x"31",x"10",x"10",x"00",
		x"10",x"10",x"3F",x"77",x"DF",x"BF",x"BF",x"BF",x"BF",x"BF",x"FF",x"5F",x"77",x"3F",x"10",x"10",
		x"00",x"01",x"07",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"06",x"06",x"03",x"01",
		x"00",x"00",x"03",x"07",x"0F",x"0D",x"1E",x"1F",x"1F",x"19",x"09",x"0F",x"07",x"03",x"00",x"00",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"00",x"00",x"00",x"1F",x"3F",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF",x"3F",x"1F",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"0C",x"1B",x"1A",x"19",x"18",x"0C",x"0F",x"07",x"03",x"00",x"00",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"1E",x"3F",x"3F",x"3F",x"7D",x"7F",x"3E",x"1E",x"3F",x"7D",x"3F",x"1F",x"0C",x"00",x"0F",
		x"00",x"1E",x"3F",x"3F",x"3F",x"6F",x"7F",x"3E",x"1E",x"3F",x"7F",x"3F",x"1B",x"0C",x"00",x"0F",
		x"00",x"1E",x"3B",x"3F",x"3F",x"7F",x"7F",x"3E",x"1E",x"3F",x"77",x"3F",x"1F",x"0C",x"00",x"0F",
		x"0F",x"01",x"09",x"1F",x"3F",x"3F",x"1A",x"0E",x"1A",x"3F",x"3F",x"1F",x"09",x"01",x"01",x"0F",
		x"0F",x"01",x"09",x"1F",x"3F",x"3F",x"1A",x"0E",x"1A",x"3F",x"3F",x"1F",x"09",x"01",x"01",x"0F",
		x"38",x"FC",x"FF",x"EF",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF",x"FF",x"EF",x"FF",x"FC",x"38",
		x"00",x"00",x"09",x"00",x"00",x"08",x"08",x"08",x"08",x"04",x"04",x"03",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"08",x"00",x"00",x"48",x"B4",x"00",x"00",x"00",x"00",
		x"00",x"00",x"38",x"3C",x"7C",x"7F",x"FF",x"FC",x"FC",x"FC",x"78",x"20",x"00",x"00",x"06",x"0E",
		x"00",x"00",x"00",x"00",x"00",x"EE",x"60",x"00",x"10",x"08",x"08",x"04",x"02",x"02",x"01",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"06",x"04",x"04",x"01",x"06",x"0E",
		x"00",x"00",x"00",x"00",x"C0",x"78",x"00",x"00",x"00",x"00",x"00",x"17",x"E7",x"87",x"06",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"40",
		x"0F",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"03",x"87",x"C7",x"7F",x"3F",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"04",x"08",x"09",x"09",x"08",x"10",x"10",x"10",
		x"03",x"07",x"07",x"03",x"08",x"1C",x"1E",x"3F",x"3F",x"3B",x"1F",x"03",x"03",x"03",x"01",x"00",
		x"00",x"00",x"01",x"01",x"02",x"02",x"02",x"04",x"04",x"04",x"08",x"08",x"08",x"08",x"08",x"08",
		x"00",x"80",x"C0",x"40",x"61",x"3A",x"0E",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"0A",x"32",x"41",x"40",x"80",x"00",x"00",
		x"60",x"F0",x"A0",x"80",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"0E",x"08",x"00",x"00",
		x"0C",x"0C",x"06",x"06",x"06",x"04",x"08",x"10",x"20",x"00",x"80",x"60",x"18",x"0C",x"00",x"00",
		x"00",x"18",x"20",x"40",x"80",x"00",x"00",x"21",x"11",x"09",x"04",x"04",x"06",x"06",x"06",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"01",x"03",x"06",x"0C",x"15",x"15",x"0C",x"06",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"44",x"02",x"01",x"05",x"43",x"0F",x"16",x"03",x"0E",x"5B",x"21",x"00",x"00",x"00",x"00",
		x"00",x"00",x"28",x"87",x"33",x"1E",x"0C",x"44",x"32",x"1E",x"0D",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"12",x"01",x"00",x"22",x"00",x"02",x"40",x"10",x"02",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"00",x"20",x"00",x"43",x"10",x"00",x"00",x"40",x"21",x"02",x"00",x"00",x"00",x"00",
		x"80",x"0A",x"75",x"1A",x"09",x"04",x"2F",x"50",x"9C",x"0E",x"06",x"35",x"4A",x"07",x"00",x"20",
		x"08",x"80",x"00",x"00",x"09",x"86",x"40",x"01",x"02",x"14",x"09",x"00",x"01",x"A6",x"43",x"00",
		x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",
		x"0D",x"2D",x"0D",x"2F",x"07",x"03",x"31",x"79",x"79",x"31",x"03",x"07",x"2F",x"0D",x"2D",x"0D",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"7F",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"03",x"01",x"06",x"0D",x"05",x"07",x"02",x"07",x"02",x"02",x"01",x"01",x"00",x"00",
		x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"7F",x"7F",x"7E",x"F9",x"F8",x"70",x"30",x"10",
		x"02",x"00",x"05",x"02",x"01",x"03",x"06",x"04",x"09",x"09",x"09",x"09",x"0C",x"06",x"03",x"00",
		x"00",x"00",x"01",x"00",x"01",x"03",x"06",x"04",x"09",x"09",x"09",x"09",x"0D",x"06",x"03",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"30",x"30",x"30",x"30",x"18",x"0C",x"07",x"03",x"00",
		x"00",x"00",x"00",x"01",x"03",x"06",x"0C",x"0C",x"0C",x"0C",x"06",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"06",x"06",x"03",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"20",x"10",x"08",x"04",x"00",x"00",x"00",x"38",x"00",x"00",x"04",x"08",x"10",x"20",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"7F",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"7F",x"00",
		x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"02",x"02",x"02",x"01",x"00",x"00",x"00",x"00",
		x"07",x"0F",x"1E",x"3F",x"3F",x"7F",x"7E",x"7E",x"7F",x"7E",x"7F",x"3F",x"3F",x"1E",x"0F",x"07",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"00",
		x"0F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1D",x"08",x"02",x"17",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",
		x"00",x"01",x"0D",x"1C",x"61",x"C9",x"ED",x"C7",x"C7",x"ED",x"C9",x"61",x"9C",x"0D",x"01",x"00",
		x"03",x"07",x"05",x"08",x"1B",x"19",x"05",x"3F",x"3F",x"0F",x"05",x"37",x"3F",x"3F",x"3E",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"0C",x"0E",x"0F",x"0F",x"07",x"03",x"00",
		x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"08",x"08",x"04",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"08",x"0D",x"0B",x"09",x"08",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"09",x"0A",x"0A",x"0A",x"0E",x"00",
		x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08",x"07",x"00",x"06",x"09",x"09",x"09",x"06",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"E7",x"E5",x"E8",x"BF",x"FF",x"FF",x"39",x"00",x"00",x"00",x"00",
		x"00",x"06",x"8F",x"9F",x"FD",x"FC",x"F8",x"B8",x"F8",x"FC",x"FC",x"BC",x"5C",x"3C",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"FF",x"1D",x"18",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"F0",x"FE",x"FF",x"FF",x"FF",x"F7",x"FB",x"F8",x"F8",x"F8",x"60",x"00",x"00",
		x"00",x"80",x"C0",x"F0",x"FE",x"FF",x"FF",x"BF",x"FF",x"F3",x"F0",x"E0",x"80",x"00",x"00",x"00",
		x"80",x"80",x"F0",x"F8",x"FC",x"FE",x"FE",x"DE",x"44",x"C0",x"C0",x"C0",x"80",x"80",x"00",x"00",
		x"00",x"C0",x"C0",x"FD",x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FF",x"FF",x"FD",x"C0",x"C0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"FF",x"FF",x"FD",x"F8",x"BF",x"FF",x"FF",x"39",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FD",x"F8",x"FF",x"FF",x"FF",x"F9",x"C0",x"00",x"00",x"00",
		x"00",x"06",x"0F",x"1F",x"FD",x"FC",x"F8",x"F8",x"B8",x"FC",x"7C",x"1C",x"1C",x"3C",x"00",x"00",
		x"00",x"06",x"0F",x"1F",x"FD",x"FC",x"F8",x"F8",x"F8",x"FC",x"FC",x"DC",x"1C",x"1C",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"DF",x"FD",x"38",x"00",x"00",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"FF",x"FD",x"78",x"00",x"00",x"00",x"00",
		x"04",x"0C",x"18",x"9C",x"CE",x"FF",x"FF",x"FE",x"DC",x"FC",x"FC",x"7C",x"4C",x"CC",x"4C",x"1C",
		x"80",x"80",x"00",x"F8",x"FC",x"FE",x"FE",x"BF",x"FF",x"FF",x"FE",x"9F",x"0F",x"06",x"0C",x"00",
		x"00",x"80",x"80",x"A0",x"83",x"81",x"E1",x"D3",x"FF",x"6F",x"0E",x"0E",x"1F",x"36",x"25",x"00",
		x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"80",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"80",x"80",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"40",x"00",x"00",
		x"00",x"40",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"40",x"00",
		x"60",x"E0",x"E0",x"E0",x"F0",x"E0",x"C0",x"C0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"78",x"B8",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"00",x"00",x"00",x"F8",x"FC",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FC",x"F8",x"00",x"00",x"00",
		x"00",x"00",x"C0",x"E0",x"70",x"B0",x"58",x"B8",x"B8",x"38",x"70",x"F0",x"E0",x"C0",x"00",x"00",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"00",x"80",x"8F",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",
		x"40",x"42",x"48",x"44",x"42",x"00",x"00",x"00",x"00",x"00",x"78",x"02",x"42",x"0A",x"14",x"02",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"E0",x"D8",x"B8",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"B8",x"D8",x"E0",x"E0",
		x"D0",x"F8",x"D8",x"8C",x"DC",x"FC",x"DC",x"8C",x"DC",x"FC",x"DC",x"8C",x"D8",x"F8",x"D8",x"F0",
		x"00",x"00",x"40",x"80",x"80",x"C0",x"00",x"80",x"C0",x"80",x"C0",x"80",x"80",x"40",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"08",x"0C",x"0C",x"14",x"1C",x"1C",x"0C",
		x"01",x"03",x"07",x"E3",x"07",x"05",x"03",x"03",x"03",x"07",x"05",x"03",x"06",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"40",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
		x"0E",x"1A",x"1D",x"18",x"00",x"10",x"30",x"30",x"60",x"40",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"3C",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",x"01",x"03",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"E0",x"70",x"B0",x"F8",x"18",x"00",
		x"00",x"00",x"00",x"00",x"00",x"78",x"FE",x"33",x"07",x"81",x"83",x"03",x"03",x"01",x"00",x"00",
		x"03",x"07",x"03",x"03",x"05",x"07",x"07",x"03",x"00",x"0C",x"0E",x"5E",x"FF",x"FF",x"CF",x"C6",
		x"00",x"00",x"00",x"00",x"00",x"60",x"E0",x"E0",x"E0",x"E0",x"C0",x"C1",x"83",x"87",x"07",x"03",
		x"00",x"01",x"07",x"3C",x"C0",x"00",x"00",x"00",x"00",x"00",x"FC",x"07",x"01",x"00",x"00",x"00",
		x"00",x"00",x"C0",x"60",x"30",x"1C",x"3E",x"7E",x"F6",x"EE",x"DC",x"DC",x"DC",x"D8",x"D0",x"60",
		x"40",x"80",x"00",x"00",x"00",x"42",x"33",x"07",x"07",x"07",x"07",x"07",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"40",x"60",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"0C",x"0E",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"10",x"70",x"70",x"F0",x"F0",x"F0",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"80",x"40",x"E0",x"30",x"18",x"54",x"54",x"18",x"30",x"E0",x"40",x"80",x"00",x"00",
		x"20",x"50",x"70",x"50",x"D8",x"88",x"88",x"04",x"04",x"88",x"88",x"D8",x"50",x"70",x"50",x"20",
		x"00",x"00",x"00",x"78",x"FE",x"86",x"03",x"73",x"7B",x"3B",x"33",x"86",x"FE",x"3C",x"00",x"00",
		x"00",x"80",x"78",x"FC",x"86",x"03",x"71",x"F9",x"F9",x"79",x"7B",x"32",x"86",x"FC",x"38",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"14",x"64",x"EB",x"03",x"94",x"A7",x"6F",x"35",x"05",x"2A",x"30",x"0C",x"02",x"00",
		x"00",x"80",x"F6",x"38",x"0F",x"3D",x"CF",x"84",x"5B",x"07",x"01",x"8F",x"7C",x"38",x"08",x"00",
		x"0C",x"13",x"3D",x"F4",x"C9",x"07",x"1C",x"18",x"70",x"9E",x"23",x"04",x"EC",x"9E",x"25",x"CC",
		x"00",x"0D",x"04",x"FE",x"83",x"0E",x"BC",x"BC",x"78",x"9C",x"8F",x"87",x"7B",x"9D",x"01",x"44",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"00",x"54",x"00",x"7C",x"7C",x"5C",x"4C",x"64",x"54",x"6C",x"74",x"7C",x"7C",x"00",x"54",x"00",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"FF",x"F7",x"FF",x"F7",x"F7",x"FF",x"F7",x"F7",x"FF",x"F7",x"F7",x"FF",x"01",x"FE",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E0",x"F0",x"F0",x"F0",x"F0",x"70",x"F0",x"F0",x"F0",x"70",x"F0",x"F0",x"70",x"F0",x"F0",x"60",
		x"00",x"30",x"58",x"08",x"A0",x"C0",x"F8",x"DE",x"8F",x"57",x"0B",x"2D",x"04",x"08",x"00",x"00",
		x"70",x"DA",x"EC",x"36",x"D3",x"21",x"01",x"81",x"C1",x"E3",x"E6",x"C6",x"0E",x"7C",x"BC",x"00",
		x"20",x"F0",x"68",x"34",x"F6",x"02",x"03",x"E1",x"F1",x"F1",x"F1",x"E1",x"83",x"66",x"BE",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",
		x"00",x"00",x"00",x"80",x"C0",x"60",x"30",x"30",x"30",x"30",x"60",x"C0",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"60",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"84",x"88",x"90",x"20",x"00",x"00",x"00",x"1C",x"00",x"00",x"20",x"90",x"88",x"84",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"FE",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"FE",x"00",
		x"04",x"0E",x"8C",x"CC",x"EE",x"EE",x"EE",x"EE",x"EC",x"EC",x"6C",x"0E",x"0E",x"0E",x"04",x"00",
		x"00",x"00",x"00",x"00",x"DE",x"3E",x"7E",x"7E",x"7E",x"7E",x"7E",x"3E",x"DE",x"00",x"00",x"00",
		x"80",x"00",x"00",x"00",x"80",x"00",x"04",x"02",x"FC",x"00",x"00",x"80",x"00",x"00",x"00",x"80",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FC",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"F4",x"E0",x"4A",x"1C",x"B8",x"F0",x"F0",x"E0",x"C0",x"00",
		x"38",x"BC",x"9C",x"DC",x"FC",x"BC",x"F8",x"F8",x"F8",x"FC",x"BE",x"FE",x"DE",x"8C",x"8C",x"00",
		x"E0",x"F0",x"50",x"08",x"6C",x"CC",x"A0",x"FE",x"FE",x"F8",x"D0",x"FB",x"FF",x"FF",x"3E",x"0C",
		x"5E",x"3F",x"07",x"05",x"09",x"7B",x"01",x"3D",x"7F",x"7F",x"BF",x"FF",x"FF",x"F0",x"F8",x"70",
		x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"40",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"E7",x"E5",x"E8",x"BF",x"FF",x"FF",x"39",x"00",x"00",x"00",x"00",
		x"00",x"06",x"8F",x"9F",x"FD",x"FC",x"F8",x"B8",x"F8",x"FC",x"FC",x"BC",x"5C",x"3C",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"FF",x"1D",x"18",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"F0",x"FE",x"FF",x"FF",x"FF",x"F7",x"FB",x"F8",x"F8",x"F8",x"60",x"00",x"00",
		x"00",x"80",x"C0",x"F0",x"FE",x"FF",x"FF",x"BF",x"FF",x"F3",x"F0",x"E0",x"80",x"00",x"00",x"00",
		x"80",x"80",x"F0",x"F8",x"FC",x"FE",x"FE",x"DE",x"44",x"C0",x"C0",x"C0",x"80",x"80",x"00",x"00",
		x"00",x"C0",x"C0",x"FD",x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FF",x"FF",x"FD",x"C0",x"C0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"FF",x"FF",x"FD",x"F8",x"BF",x"FF",x"FF",x"39",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FD",x"F8",x"FF",x"FF",x"FF",x"F9",x"C0",x"00",x"00",x"00",
		x"00",x"06",x"0F",x"1F",x"FD",x"FC",x"F8",x"F8",x"B8",x"FC",x"7C",x"1C",x"1C",x"3C",x"00",x"00",
		x"00",x"06",x"0F",x"1F",x"FD",x"FC",x"F8",x"F8",x"F8",x"FC",x"FC",x"DC",x"1C",x"1C",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"DF",x"FD",x"38",x"00",x"00",x"00",x"00",
		x"1E",x"1C",x"1C",x"1C",x"FC",x"FC",x"F8",x"FB",x"FF",x"FF",x"FD",x"78",x"00",x"00",x"00",x"00",
		x"04",x"0C",x"18",x"9C",x"CE",x"FF",x"FF",x"FE",x"DC",x"FC",x"FC",x"7C",x"4C",x"CC",x"4C",x"1C",
		x"80",x"80",x"00",x"F8",x"FC",x"FE",x"FE",x"BF",x"FF",x"FF",x"FE",x"9F",x"0F",x"06",x"0C",x"00",
		x"00",x"80",x"80",x"A0",x"83",x"81",x"E1",x"D3",x"FF",x"6F",x"0E",x"0E",x"1F",x"36",x"25",x"00",
		x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"80",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"80",x"80",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"40",x"00",x"00",
		x"00",x"40",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"40",x"00",
		x"60",x"E0",x"E0",x"E0",x"F0",x"E0",x"C0",x"C0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"78",x"B8",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"00",x"00",x"00",x"F8",x"FC",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FC",x"F8",x"00",x"00",x"00",
		x"00",x"00",x"C0",x"E0",x"70",x"B0",x"58",x"B8",x"B8",x"38",x"70",x"F0",x"E0",x"C0",x"00",x"00",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"E0",x"00",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"00",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"00",x"80",x"8F",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",
		x"40",x"42",x"48",x"44",x"42",x"00",x"00",x"00",x"00",x"00",x"78",x"02",x"42",x"0A",x"14",x"02",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"CC",x"E6",x"EF",x"C3",x"E7",x"E7",x"E7",x"C3",x"F7",x"F7",x"E7",x"C3",x"E7",x"F6",x"E6",x"FC",
		x"E0",x"D8",x"B8",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"B8",x"D8",x"E0",x"E0",
		x"D0",x"F8",x"D8",x"8C",x"DC",x"FC",x"DC",x"8C",x"DC",x"FC",x"DC",x"8C",x"D8",x"F8",x"D8",x"F0",
		x"00",x"00",x"40",x"80",x"80",x"C0",x"00",x"80",x"C0",x"80",x"C0",x"80",x"80",x"40",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"08",x"0C",x"0C",x"14",x"1C",x"1C",x"0C",
		x"01",x"03",x"07",x"E3",x"07",x"05",x"03",x"03",x"03",x"07",x"05",x"03",x"06",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"40",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
		x"0E",x"1A",x"1D",x"18",x"00",x"10",x"30",x"30",x"60",x"40",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"3C",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",x"01",x"03",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"E0",x"70",x"B0",x"F8",x"18",x"00",
		x"00",x"00",x"00",x"00",x"00",x"78",x"FE",x"33",x"07",x"81",x"83",x"03",x"03",x"01",x"00",x"00",
		x"03",x"07",x"03",x"03",x"05",x"07",x"07",x"03",x"00",x"0C",x"0E",x"5E",x"FF",x"FF",x"CF",x"C6",
		x"00",x"00",x"00",x"00",x"00",x"60",x"E0",x"E0",x"E0",x"E0",x"C0",x"C1",x"83",x"87",x"07",x"03",
		x"00",x"01",x"07",x"3C",x"C0",x"00",x"00",x"00",x"00",x"00",x"FC",x"07",x"01",x"00",x"00",x"00",
		x"00",x"00",x"C0",x"60",x"30",x"1C",x"3E",x"7E",x"F6",x"EE",x"DC",x"DC",x"DC",x"D8",x"D0",x"60",
		x"40",x"80",x"00",x"00",x"00",x"42",x"33",x"07",x"07",x"07",x"07",x"07",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"40",x"60",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"0C",x"0E",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"10",x"70",x"70",x"F0",x"F0",x"F0",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"80",x"40",x"E0",x"30",x"18",x"54",x"54",x"18",x"30",x"E0",x"40",x"80",x"00",x"00",
		x"20",x"50",x"70",x"50",x"D8",x"88",x"88",x"04",x"04",x"88",x"88",x"D8",x"50",x"70",x"50",x"20",
		x"00",x"00",x"00",x"78",x"FE",x"86",x"03",x"73",x"7B",x"3B",x"33",x"86",x"FE",x"3C",x"00",x"00",
		x"00",x"80",x"78",x"FC",x"86",x"03",x"71",x"F9",x"F9",x"79",x"7B",x"32",x"86",x"FC",x"38",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"14",x"64",x"EB",x"03",x"94",x"A7",x"6F",x"35",x"05",x"2A",x"30",x"0C",x"02",x"00",
		x"00",x"80",x"F6",x"38",x"0F",x"3D",x"CF",x"84",x"5B",x"07",x"01",x"8F",x"7C",x"38",x"08",x"00",
		x"0C",x"13",x"3D",x"F4",x"C9",x"07",x"1C",x"18",x"70",x"9E",x"23",x"04",x"EC",x"9E",x"25",x"CC",
		x"00",x"0D",x"04",x"FE",x"83",x"0E",x"BC",x"BC",x"78",x"9C",x"8F",x"87",x"7B",x"9D",x"01",x"44",
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"00",x"54",x"00",x"7C",x"7C",x"5C",x"4C",x"64",x"54",x"6C",x"74",x"7C",x"7C",x"00",x"54",x"00",
		x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"FF",x"F7",x"FF",x"F7",x"F7",x"FF",x"F7",x"F7",x"FF",x"F7",x"F7",x"FF",x"01",x"FE",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E0",x"F0",x"F0",x"F0",x"F0",x"70",x"F0",x"F0",x"F0",x"70",x"F0",x"F0",x"70",x"F0",x"F0",x"60",
		x"00",x"30",x"58",x"08",x"A0",x"C0",x"F8",x"DE",x"8F",x"57",x"0B",x"2D",x"04",x"08",x"00",x"00",
		x"70",x"DA",x"EC",x"36",x"D3",x"21",x"01",x"81",x"C1",x"E3",x"E6",x"C6",x"0E",x"7C",x"BC",x"00",
		x"20",x"F0",x"68",x"34",x"F6",x"02",x"03",x"E1",x"F1",x"F1",x"F1",x"E1",x"83",x"66",x"BE",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",
		x"00",x"00",x"00",x"80",x"C0",x"60",x"30",x"30",x"30",x"30",x"60",x"C0",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"60",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"84",x"88",x"90",x"20",x"00",x"00",x"00",x"1C",x"00",x"00",x"20",x"90",x"88",x"84",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"FE",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"FE",x"00",
		x"04",x"0E",x"8C",x"CC",x"EE",x"EE",x"EE",x"EE",x"EC",x"EC",x"6C",x"0E",x"0E",x"0E",x"04",x"00",
		x"00",x"00",x"00",x"00",x"DE",x"3E",x"7E",x"7E",x"7E",x"7E",x"7E",x"3E",x"DE",x"00",x"00",x"00",
		x"80",x"00",x"00",x"00",x"80",x"00",x"04",x"02",x"FC",x"00",x"00",x"80",x"00",x"00",x"00",x"80",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FC",x"F8",x"F0",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"F4",x"E0",x"4A",x"1C",x"B8",x"F0",x"F0",x"E0",x"C0",x"00",
		x"38",x"BC",x"9C",x"DC",x"FC",x"BC",x"F8",x"F8",x"F8",x"FC",x"BE",x"FE",x"DE",x"8C",x"8C",x"00",
		x"E0",x"F0",x"50",x"08",x"6C",x"CC",x"A0",x"FE",x"FE",x"F8",x"D0",x"FB",x"FF",x"FF",x"3E",x"0C",
		x"5E",x"3F",x"07",x"05",x"09",x"7B",x"01",x"3D",x"7F",x"7F",x"BF",x"FF",x"FF",x"F0",x"F8",x"70",
		x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"20",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"40",x"00",
		x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20",x"20",x"C0",x"00",
		x"55",x"04",x"52",x"C5",x"A5",x"8A",x"40",x"8A",x"80",x"B9",x"02",x"BA",x"40",x"BB",x"40",x"FA",
		x"77",x"77",x"53",x"3F",x"6A",x"AA",x"AB",x"34",x"00",x"FB",x"97",x"67",x"6B",x"AB",x"34",x"00",
		x"E9",x"0F",x"FA",x"47",x"00",x"53",x"0F",x"37",x"17",x"6A",x"07",x"AA",x"AB",x"03",x"D8",x"E6",
		x"3C",x"34",x"00",x"FB",x"97",x"67",x"6B",x"AB",x"34",x"00",x"04",x"22",x"D5",x"23",x"2B",x"34",
		x"81",x"14",x"45",x"04",x"52",x"80",x"37",x"B4",x"33",x"C6",x"51",x"53",x"F0",x"96",x"51",x"04",
		x"45",x"83",x"05",x"85",x"A5",x"B8",x"20",x"B0",x"00",x"D5",x"27",x"AE",x"AF",x"C5",x"8A",x"80",
		x"14",x"73",x"26",x"74",x"A5",x"0A",x"37",x"B2",x"A8",x"27",x"AE",x"AF",x"A9",x"B4",x"35",x"14",
		x"73",x"04",x"62",x"93",x"B8",x"20",x"F0",x"03",x"05",x"C6",x"69",x"F0",x"03",x"09",x"C6",x"69",
		x"B8",x"08",x"A5",x"B5",x"D4",x"1A",x"D4",x"38",x"8A",x"80",x"C6",x"62",x"B9",x"03",x"34",x"3F",
		x"B4",x"35",x"E9",x"8E",x"B9",x"04",x"B4",x"35",x"E9",x"96",x"FA",x"03",x"F9",x"A9",x"C6",x"86",
		x"9A",x"7F",x"B4",x"35",x"E9",x"A2",x"04",x"86",x"BB",x"20",x"34",x"15",x"FB",x"77",x"77",x"53",
		x"3F",x"6B",x"AB",x"26",x"74",x"E6",x"AA",x"34",x"15",x"FB",x"77",x"77",x"53",x"3F",x"6B",x"AB",
		x"26",x"74",x"E6",x"B7",x"04",x"62",x"BA",x"08",x"B9",x"FF",x"8A",x"80",x"A5",x"B5",x"FA",x"AB",
		x"34",x"31",x"34",x"31",x"FA",x"97",x"67",x"6A",x"F6",x"62",x"AB",x"34",x"31",x"34",x"31",x"34",
		x"31",x"FA",x"AB",x"34",x"31",x"34",x"31",x"FA",x"97",x"67",x"97",x"67",x"6A",x"AA",x"04",x"CE",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"B8",x"03",x"34",x"23",x"E8",x"02",x"B8",x"03",x"34",x"0D",x"E8",x"08",x"83",x"27",x"AE",x"AF",
		x"D5",x"AE",x"AF",x"C4",x"7B",x"FB",x"47",x"E7",x"53",x"1F",x"AF",x"FB",x"47",x"E7",x"53",x"E0",
		x"AE",x"A4",x"35",x"FB",x"77",x"77",x"AE",x"53",x"3F",x"AF",x"FE",x"53",x"C0",x"AE",x"D5",x"C4",
		x"7B",x"FB",x"77",x"77",x"AE",x"53",x"3F",x"AF",x"FE",x"53",x"C0",x"AE",x"D5",x"A4",x"35",x"FE",
		x"6F",x"E6",x"44",x"1F",x"6F",x"E6",x"48",x"1F",x"AE",x"83",x"AB",x"D5",x"FB",x"1B",x"C5",x"B4",
		x"33",x"C6",x"9E",x"F2",x"9F",x"A8",x"D4",x"1A",x"D4",x"38",x"D4",x"4B",x"C6",x"4B",x"B9",x"03",
		x"8A",x"80",x"34",x"3F",x"D5",x"34",x"3F",x"D4",x"7B",x"E9",x"62",x"B9",x"04",x"D5",x"D4",x"7B",
		x"E9",x"6D",x"FA",x"03",x"F9",x"A9",x"C6",x"58",x"9A",x"7F",x"D5",x"D4",x"7B",x"E9",x"7A",x"24",
		x"58",x"AB",x"D5",x"FB",x"1B",x"C5",x"B4",x"33",x"C6",x"9E",x"F2",x"9F",x"A8",x"D4",x"1A",x"D4",
		x"38",x"D4",x"4B",x"C6",x"82",x"FA",x"A9",x"D5",x"D4",x"7B",x"E9",x"97",x"24",x"8F",x"83",x"BE",
		x"80",x"A4",x"A2",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"03",x"06",x"09",x"0C",x"0F",x"12",x"15",x"18",x"1B",x"1E",x"21",x"24",x"27",x"2A",x"2D",
		x"30",x"33",x"36",x"39",x"3C",x"3F",x"42",x"45",x"48",x"4B",x"4E",x"51",x"54",x"57",x"5A",x"5D",
		x"60",x"5D",x"5A",x"57",x"54",x"51",x"4E",x"4B",x"48",x"45",x"42",x"3F",x"3C",x"39",x"36",x"33",
		x"30",x"2D",x"2A",x"27",x"24",x"21",x"1E",x"1B",x"18",x"15",x"12",x"0F",x"0C",x"09",x"06",x"03",
		x"FC",x"6E",x"AC",x"FD",x"7F",x"AD",x"77",x"77",x"53",x"3F",x"A3",x"A8",x"C5",x"FC",x"6E",x"AC",
		x"FD",x"7F",x"AD",x"77",x"77",x"43",x"C0",x"A3",x"D5",x"68",x"39",x"16",x"5F",x"44",x"40",x"C5",
		x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"05",x"0A",x"0F",x"14",x"19",x"1E",x"23",x"28",x"2D",x"32",x"37",x"3C",x"41",x"46",x"4B",
		x"50",x"55",x"5A",x"5F",x"64",x"69",x"6E",x"73",x"78",x"7D",x"82",x"87",x"8C",x"91",x"96",x"9B",
		x"9F",x"9B",x"96",x"91",x"8C",x"87",x"82",x"7D",x"78",x"73",x"6E",x"69",x"64",x"5F",x"5A",x"55",
		x"50",x"4B",x"46",x"41",x"3C",x"37",x"32",x"2D",x"28",x"23",x"1E",x"19",x"14",x"0F",x"0A",x"05",
		x"00",x"2A",x"80",x"1C",x"84",x"0E",x"88",x"8A",x"88",x"00",x"16",x"84",x"0B",x"84",x"84",x"00",
		x"00",x"18",x"84",x"0C",x"80",x"80",x"00",x"10",x"B8",x"B4",x"B0",x"00",x"12",x"90",x"09",x"90",
		x"90",x"12",x"90",x"90",x"94",x"90",x"94",x"90",x"94",x"09",x"94",x"94",x"12",x"94",x"94",x"98",
		x"94",x"98",x"94",x"00",x"00",x"09",x"B0",x"B2",x"B4",x"12",x"BA",x"B6",x"00",x"0E",x"A4",x"1C",
		x"E8",x"90",x"D8",x"88",x"38",x"E0",x"80",x"00",x"60",x"CA",x"82",x"20",x"CC",x"84",x"40",x"D0",
		x"86",x"CA",x"82",x"08",x"DA",x"89",x"D9",x"89",x"DA",x"89",x"D9",x"89",x"DA",x"89",x"D9",x"89",
		x"DA",x"89",x"D9",x"89",x"08",x"DA",x"89",x"D9",x"89",x"DA",x"89",x"D9",x"89",x"DA",x"89",x"D9",
		x"89",x"DA",x"89",x"D9",x"89",x"7F",x"DA",x"8A",x"00",x"00",x"24",x"88",x"82",x"88",x"82",x"12",
		x"D8",x"88",x"D6",x"88",x"D8",x"82",x"D6",x"82",x"D6",x"88",x"88",x"D6",x"82",x"82",x"24",x"DA",
		x"87",x"D9",x"83",x"DA",x"87",x"D7",x"83",x"09",x"D8",x"88",x"D7",x"88",x"D8",x"88",x"D7",x"88",
		x"D8",x"82",x"D7",x"82",x"D8",x"82",x"D7",x"82",x"48",x"D8",x"88",x"00",x"00",x"00",x"20",x"E8",
		x"88",x"82",x"E2",x"88",x"10",x"82",x"A4",x"20",x"DC",x"88",x"82",x"84",x"18",x"E0",x"87",x"08",
		x"A2",x"20",x"E4",x"88",x"E7",x"82",x"E8",x"88",x"EA",x"82",x"20",x"EA",x"88",x"EC",x"82",x"88",
		x"82",x"EC",x"88",x"82",x"F0",x"90",x"88",x"EC",x"88",x"82",x"10",x"84",x"AA",x"E8",x"8C",x"AA",
		x"20",x"E7",x"92",x"8A",x"10",x"84",x"A4",x"E2",x"8C",x"A4",x"00",x"1B",x"E2",x"88",x"09",x"A4",
		x"12",x"82",x"A8",x"12",x"88",x"A4",x"E2",x"82",x"A4",x"12",x"E0",x"80",x"09",x"82",x"83",x"86",
		x"88",x"8A",x"8C",x"24",x"D0",x"88",x"00",x"20",x"80",x"DC",x"98",x"E0",x"9A",x"E2",x"9C",x"20",
		x"90",x"E4",x"88",x"10",x"E3",x"90",x"A4",x"20",x"88",x"DA",x"8A",x"EA",x"84",x"10",x"E8",x"8A",
		x"A4",x"20",x"84",x"E2",x"82",x"E2",x"87",x"16",x"E8",x"88",x"0A",x"A3",x"10",x"E4",x"82",x"A0",
		x"15",x"C8",x"80",x"2B",x"CA",x"83",x"40",x"CB",x"80",x"00",x"10",x"E8",x"A4",x"E8",x"A4",x"E6",
		x"A2",x"E6",x"A2",x"E4",x"A0",x"E4",x"A0",x"E2",x"9C",x"E2",x"9C",x"10",x"E0",x"90",x"A0",x"E4",
		x"88",x"A0",x"E4",x"80",x"A0",x"E4",x"88",x"A8",x"20",x"EA",x"96",x"E8",x"90",x"40",x"F0",x"80",
		x"00",x"10",x"E8",x"A4",x"E8",x"A4",x"E6",x"A2",x"E6",x"A2",x"E4",x"A0",x"E4",x"A0",x"E2",x"9C",
		x"E2",x"9C",x"20",x"E0",x"90",x"10",x"88",x"08",x"A0",x"A2",x"20",x"E4",x"90",x"E0",x"88",x"20",
		x"E2",x"92",x"10",x"8A",x"08",x"A2",x"A4",x"20",x"E6",x"92",x"E2",x"8A",x"20",x"E8",x"88",x"10",
		x"82",x"A8",x"EA",x"88",x"A8",x"E6",x"82",x"A4",x"E8",x"80",x"2B",x"83",x"40",x"80",x"00",x"0A",
		x"E8",x"A4",x"EA",x"A6",x"14",x"EC",x"A8",x"28",x"E8",x"A4",x"0A",x"E8",x"A4",x"EA",x"A6",x"14",
		x"EC",x"A8",x"28",x"E8",x"A4",x"00",x"0A",x"E0",x"98",x"E0",x"98",x"3C",x"E0",x"98",x"12",x"88",
		x"84",x"88",x"84",x"88",x"84",x"88",x"84",x"88",x"84",x"88",x"84",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"A3",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"20",x"10",x"05",x"06",x"12",x"40",x"16",x"01",x"02",x"00",x"04",x"14",x"FA",x"1E",x"2D",
		x"10",x"00",x"13",x"00",x"11",x"00",x"14",x"83",x"FE",x"85",x"FE",x"85",x"FE",x"00",x"15",x"00",
		x"0A",x"00",x"95",x"FE",x"85",x"FE",x"85",x"FE",x"00",x"00",x"00",x"09",x"00",x"FE",x"84",x"FE",
		x"83",x"FE",x"00",x"A3",x"83",x"D5",x"B8",x"20",x"80",x"37",x"53",x"0F",x"20",x"37",x"17",x"60",
		x"96",x"64",x"B6",x"BD",x"46",x"BA",x"F0",x"A3",x"C6",x"5D",x"F2",x"5F",x"34",x"3F",x"E9",x"5D",
		x"FF",x"96",x"56",x"FE",x"C6",x"75",x"FA",x"03",x"F8",x"A9",x"27",x"AE",x"AF",x"C4",x"7B",x"27",
		x"AE",x"AF",x"C4",x"7B",x"F0",x"A3",x"C6",x"5F",x"F2",x"8C",x"92",x"7D",x"B2",x"81",x"D2",x"E5",
		x"8A",x"80",x"A8",x"D4",x"1A",x"D4",x"38",x"C6",x"64",x"B9",x"08",x"C4",x"7B",x"34",x"4A",x"04",
		x"52",x"34",x"81",x"04",x"52",x"C5",x"BE",x"80",x"F4",x"06",x"04",x"52",x"76",x"91",x"C5",x"04",
		x"74",x"B0",x"08",x"A4",x"46",x"D5",x"FB",x"1B",x"C5",x"A3",x"C6",x"9E",x"96",x"A2",x"14",x"45",
		x"04",x"52",x"D2",x"B6",x"97",x"F7",x"97",x"F7",x"A9",x"23",x"80",x"62",x"16",x"AE",x"16",x"B2",
		x"A4",x"AE",x"E9",x"A9",x"A4",x"95",x"F4",x"06",x"A4",x"95",x"95",x"BB",x"F0",x"FB",x"E7",x"E7",
		x"47",x"53",x"03",x"96",x"C6",x"17",x"37",x"17",x"6B",x"AB",x"03",x"E0",x"F6",x"D7",x"85",x"27",
		x"AE",x"AF",x"B8",x"20",x"A0",x"C4",x"7B",x"FB",x"47",x"E7",x"53",x"1F",x"AF",x"FB",x"47",x"E7",
		x"53",x"E0",x"AE",x"C4",x"7B",x"B0",x"04",x"C5",x"F9",x"F2",x"ED",x"04",x"C6",x"D5",x"A4",x"46",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"28",x"00",x"2A",x"61",x"2C",x"E6",x"2F",x"91",x"32",x"66",x"FF",x"FF",x"35",x"65",x"38",x"92",
		x"3B",x"EF",x"3F",x"75",x"43",x"46",x"47",x"46",x"4B",x"83",x"BB",x"00",x"B9",x"30",x"B1",x"FF",
		x"D4",x"27",x"96",x"20",x"E8",x"20",x"83",x"B9",x"30",x"FB",x"96",x"2D",x"11",x"F1",x"96",x"34",
		x"FB",x"1B",x"E3",x"83",x"FB",x"1B",x"84",x"F8",x"D4",x"27",x"C6",x"5C",x"F2",x"46",x"AA",x"D4",
		x"27",x"F2",x"46",x"A9",x"D4",x"27",x"A8",x"D4",x"5D",x"F8",x"83",x"D2",x"54",x"D5",x"BE",x"00",
		x"BF",x"00",x"C5",x"83",x"D4",x"27",x"D5",x"A8",x"D4",x"5D",x"C5",x"F8",x"83",x"F8",x"53",x"0F",
		x"E7",x"AC",x"A3",x"AF",x"FC",x"17",x"A3",x"AE",x"F8",x"53",x"30",x"47",x"AC",x"FF",x"97",x"67",
		x"AF",x"FE",x"67",x"AE",x"1C",x"FC",x"03",x"FC",x"96",x"6D",x"83",x"42",x"03",x"80",x"62",x"76",
		x"A2",x"FC",x"6E",x"AC",x"FD",x"7F",x"AD",x"77",x"77",x"43",x"C0",x"A3",x"A8",x"C5",x"FC",x"6E",
		x"AC",x"FD",x"7F",x"AD",x"77",x"77",x"43",x"C0",x"A3",x"D5",x"68",x"39",x"16",x"A0",x"C4",x"81",
		x"C5",x"83",x"44",x"40",x"A3",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"03",x"06",x"09",x"0C",x"0F",x"12",x"15",x"18",x"1B",x"1E",x"21",x"24",x"27",x"2A",x"2D",
		x"30",x"33",x"36",x"39",x"3C",x"3F",x"42",x"45",x"48",x"4B",x"4E",x"51",x"54",x"57",x"5A",x"5D",
		x"60",x"5D",x"5A",x"57",x"54",x"51",x"4E",x"4B",x"48",x"45",x"42",x"3F",x"3C",x"39",x"36",x"33",
		x"30",x"2D",x"2A",x"27",x"24",x"21",x"1E",x"1B",x"18",x"15",x"12",x"0F",x"0C",x"09",x"06",x"03",
		x"02",x"04",x"06",x"0C",x"14",x"FF",x"A8",x"A3",x"28",x"17",x"A3",x"A9",x"12",x"24",x"C9",x"F4",
		x"24",x"9A",x"7F",x"B8",x"00",x"B9",x"FF",x"F4",x"24",x"9A",x"7F",x"B8",x"00",x"B9",x"FF",x"F4",
		x"24",x"8A",x"80",x"83",x"BF",x"00",x"9A",x"BF",x"A5",x"23",x"B0",x"48",x"3A",x"BA",x"08",x"81",
		x"E9",x"3B",x"AB",x"C8",x"F8",x"F2",x"BA",x"43",x"B0",x"3A",x"FB",x"77",x"AB",x"F2",x"78",x"76",
		x"5B",x"1F",x"FF",x"A3",x"F2",x"4A",x"37",x"17",x"E4",x"4E",x"CF",x"00",x"23",x"EC",x"6E",x"AE",
		x"F6",x"59",x"27",x"AE",x"39",x"EA",x"AC",x"E4",x"2D",x"E4",x"54",x"A5",x"CF",x"FF",x"F2",x"62",
		x"E4",x"64",x"27",x"AF",x"A3",x"37",x"17",x"6E",x"F6",x"71",x"27",x"AE",x"39",x"EA",x"AC",x"E4",
		x"2D",x"00",x"AE",x"39",x"EA",x"AC",x"E4",x"2D",x"76",x"93",x"B5",x"CF",x"FF",x"F2",x"81",x"E4",
		x"83",x"27",x"AF",x"A3",x"6E",x"AE",x"E6",x"90",x"23",x"FF",x"AE",x"39",x"EA",x"AC",x"E4",x"2D",
		x"00",x"E4",x"8B",x"1F",x"FF",x"A3",x"F2",x"9C",x"00",x"00",x"E4",x"9F",x"CF",x"FF",x"A3",x"6E",
		x"E6",x"AA",x"23",x"FF",x"AE",x"39",x"EA",x"AC",x"E4",x"2D",x"E4",x"A4",x"FB",x"C6",x"B4",x"00",
		x"00",x"00",x"E4",x"3B",x"81",x"C6",x"BA",x"FB",x"E4",x"3B",x"8A",x"40",x"A5",x"83",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"FF",x"05",x"FF",x"02",x"00",
		x"C0",x"F0",x"F0",x"F8",x"38",x"7C",x"3C",x"7A",x"38",x"D1",x"E1",x"E1",x"E1",x"E0",x"E2",x"F0",
		x"F1",x"D1",x"DC",x"4E",x"9E",x"0F",x"0F",x"1E",x"1E",x"0E",x"1E",x"1E",x"1A",x"58",x"E1",x"E1",
		x"C0",x"F0",x"F0",x"F8",x"38",x"7C",x"3C",x"7A",x"38",x"D1",x"E1",x"E1",x"E1",x"E0",x"E2",x"F0",
		x"F1",x"D1",x"DC",x"4E",x"9E",x"0F",x"0F",x"1E",x"1E",x"0E",x"1E",x"1E",x"1A",x"58",x"E1",x"E1",
		x"C0",x"F0",x"F0",x"F8",x"38",x"7C",x"3C",x"7A",x"38",x"D1",x"E1",x"E1",x"E1",x"E0",x"E2",x"F0",
		x"F1",x"D1",x"DC",x"4E",x"9E",x"0F",x"0F",x"1E",x"1E",x"0E",x"1E",x"1E",x"1A",x"58",x"E1",x"E1",
		x"C0",x"F0",x"F0",x"F8",x"38",x"7C",x"3C",x"7A",x"38",x"D1",x"E1",x"E1",x"E1",x"E0",x"E2",x"F0",
		x"F1",x"D1",x"DC",x"4E",x"9E",x"0F",x"0F",x"1E",x"1E",x"0E",x"1E",x"1E",x"1A",x"58",x"E1",x"E1",
		x"1E",x"0E",x"3E",x"8F",x"27",x"0C",x"DC",x"38",x"7C",x"78",x"38",x"EC",x"6C",x"7C",x"78",x"70",
		x"CC",x"78",x"78",x"70",x"F8",x"78",x"78",x"78",x"78",x"66",x"B8",x"E4",x"E1",x"E0",x"E6",x"63",
		x"1E",x"0E",x"3E",x"8F",x"27",x"0C",x"DC",x"38",x"7C",x"78",x"38",x"EC",x"6C",x"7C",x"78",x"70",
		x"CC",x"78",x"78",x"70",x"F8",x"78",x"78",x"78",x"78",x"66",x"B8",x"E4",x"E1",x"E0",x"E6",x"63",
		x"1E",x"0E",x"3E",x"8F",x"27",x"0C",x"DC",x"38",x"7C",x"78",x"38",x"EC",x"6C",x"7C",x"78",x"70",
		x"CC",x"78",x"78",x"70",x"F8",x"78",x"78",x"78",x"78",x"66",x"B8",x"E4",x"E1",x"E0",x"E6",x"63",
		x"1E",x"0E",x"3E",x"8F",x"27",x"0C",x"DC",x"38",x"7C",x"78",x"38",x"EC",x"6C",x"7C",x"78",x"70",
		x"CC",x"78",x"78",x"70",x"F8",x"78",x"78",x"78",x"78",x"66",x"B8",x"E4",x"E1",x"E0",x"E6",x"63",
		x"1E",x"47",x"13",x"93",x"C6",x"E5",x"70",x"73",x"3C",x"1C",x"67",x"1F",x"19",x"E0",x"E2",x"78",
		x"CC",x"3E",x"39",x"1E",x"0E",x"63",x"8B",x"91",x"F0",x"E3",x"38",x"EC",x"73",x"1C",x"4E",x"33",
		x"1E",x"47",x"13",x"93",x"C6",x"E5",x"70",x"73",x"3C",x"1C",x"67",x"1F",x"19",x"E0",x"E2",x"78",
		x"CC",x"3E",x"39",x"1E",x"0E",x"63",x"8B",x"91",x"F0",x"E3",x"38",x"EC",x"73",x"1C",x"4E",x"33",
		x"1E",x"47",x"13",x"93",x"C6",x"E5",x"70",x"73",x"3C",x"1C",x"67",x"1F",x"19",x"E0",x"E2",x"78",
		x"CC",x"3E",x"39",x"1E",x"0E",x"63",x"8B",x"91",x"F0",x"E3",x"38",x"EC",x"73",x"1C",x"4E",x"33",
		x"1E",x"47",x"13",x"93",x"C6",x"E5",x"70",x"73",x"3C",x"1C",x"67",x"1F",x"19",x"E0",x"E2",x"78",
		x"CC",x"3E",x"39",x"1E",x"0E",x"63",x"8B",x"91",x"F0",x"E3",x"38",x"EC",x"73",x"1C",x"4E",x"33",
		x"E4",x"E2",x"E4",x"E4",x"D3",x"53",x"55",x"8D",x"53",x"33",x"33",x"34",x"D5",x"4D",x"55",x"35",
		x"8D",x"4D",x"55",x"4D",x"33",x"35",x"4D",x"33",x"34",x"D5",x"55",x"4D",x"94",x"CD",x"33",x"33",
		x"E4",x"E2",x"E4",x"E4",x"D3",x"53",x"55",x"8D",x"53",x"33",x"33",x"34",x"D5",x"4D",x"55",x"35",
		x"8D",x"4D",x"55",x"4D",x"33",x"35",x"4D",x"33",x"34",x"D5",x"55",x"4D",x"94",x"CD",x"33",x"33",
		x"E4",x"E2",x"E4",x"E4",x"D3",x"53",x"55",x"8D",x"53",x"33",x"33",x"34",x"D5",x"4D",x"55",x"35",
		x"8D",x"4D",x"55",x"4D",x"33",x"35",x"4D",x"33",x"34",x"D5",x"55",x"4D",x"94",x"CD",x"33",x"33",
		x"E4",x"E2",x"E4",x"E4",x"D3",x"53",x"55",x"8D",x"53",x"33",x"33",x"34",x"D5",x"4D",x"55",x"35",
		x"8D",x"4D",x"55",x"4D",x"33",x"35",x"4D",x"33",x"34",x"D5",x"55",x"4D",x"94",x"CD",x"33",x"33",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"55",x"55",x"55",x"56",x"66",x"66",x"66",x"66",x"66",
		x"66",x"55",x"65",x"55",x"56",x"66",x"66",x"66",x"59",x"99",x"99",x"99",x"95",x"55",x"55",x"66",
		x"65",x"66",x"66",x"66",x"66",x"59",x"59",x"59",x"59",x"59",x"59",x"59",x"96",x"56",x"59",x"59",
		x"66",x"56",x"66",x"66",x"66",x"66",x"55",x"55",x"95",x"56",x"59",x"99",x"99",x"99",x"95",x"99",
		x"99",x"99",x"99",x"99",x"99",x"59",x"59",x"99",x"96",x"66",x"56",x"55",x"99",x"99",x"A6",x"96",
		x"56",x"59",x"56",x"66",x"66",x"66",x"99",x"96",x"66",x"59",x"96",x"95",x"95",x"4D",x"93",x"66",
		x"65",x"99",x"66",x"59",x"59",x"39",x"39",x"56",x"59",x"5A",x"56",x"5A",x"5A",x"69",x"5A",x"59",
		x"64",x"E4",x"CD",x"4C",x"E4",x"E6",x"66",x"69",x"6A",x"66",x"A6",x"63",x"4D",x"4B",x"4D",x"59",
		x"59",x"9A",x"56",x"36",x"36",x"36",x"97",x"27",x"25",x"8E",x"8D",x"8A",x"CD",x"4D",x"4C",x"D6",
		x"65",x"A6",x"A6",x"66",x"64",x"D5",x"35",x"36",x"56",x"CE",x"4D",x"4A",x"6A",x"9B",x"26",x"26",
		x"36",x"DD",x"CC",x"88",x"89",x"22",x"CB",x"DD",x"DD",x"CA",x"92",x"46",x"65",x"95",x"65",x"96",
		x"65",x"95",x"95",x"4C",x"D3",x"4D",x"59",x"56",x"66",x"66",x"66",x"66",x"56",x"35",x"55",x"59",
		x"99",x"99",x"99",x"66",x"59",x"99",x"99",x"96",x"59",x"96",x"66",x"66",x"66",x"56",x"56",x"66",
		x"59",x"99",x"96",x"66",x"53",x"55",x"9A",x"65",x"99",x"94",x"D9",x"99",x"55",x"99",x"99",x"59",
		x"99",x"55",x"99",x"99",x"55",x"66",x"65",x"95",x"99",x"99",x"59",x"99",x"8D",x"99",x"99",x"56",
		x"65",x"96",x"59",x"59",x"95",x"66",x"66",x"59",x"66",x"65",x"55",x"9A",x"4D",x"56",x"64",x"D3",
		x"00",x"66",x"4E",x"56",x"99",x"53",x"9A",x"4E",x"4D",x"A9",x"54",x"DD",x"33",x"1D",x"C9",x"93",
		x"3D",x"49",x"25",x"E4",x"92",x"5E",x"48",x"95",x"E4",x"89",x"DD",x"44",x"BB",x"31",x"25",x"E4",
		x"46",x"5E",x"44",x"65",x"E4",x"45",x"5D",x"84",x"55",x"D8",x"45",x"67",x"61",x"16",x"76",x"12",
		x"6A",x"E1",x"4C",x"CF",x"21",x"A9",x"7A",x"1B",x"27",x"61",x"6C",x"9E",x"8D",x"98",x"E8",x"DC",
		x"C1",x"47",x"EC",x"09",x"FD",x"81",x"1F",x"E2",x"01",x"FF",x"02",x"1F",x"E0",x"C1",x"FE",x"0C",
		x"1F",x"C0",x"A0",x"FF",x"07",x"07",x"F0",x"70",x"7F",x"07",x"07",x"F0",x"70",x"7F",x"23",x"83",
		x"F0",x"38",x"3F",x"83",x"C3",x"F2",x"1C",x"3F",x"21",x"E0",x"FC",x"8E",x"0F",x"C0",x"F0",x"7F",
		x"07",x"83",x"F0",x"3C",x"3F",x"03",x"C3",x"F8",x"1E",x"1F",x"80",x"F0",x"FE",x"07",x"87",x"E0",
		x"78",x"3F",x"03",x"E1",x"F8",x"1E",x"0F",x"C0",x"F0",x"FC",x"07",x"8F",x"E0",x"3C",x"3F",x"03",
		x"C3",x"F8",x"1E",x"0F",x"C0",x"F8",x"7C",x"27",x"C3",x"E0",x"1E",x"3F",x"80",x"F0",x"FC",x"07",
		x"87",x"F0",x"3C",x"3F",x"01",x"E1",x"FC",x"0F",x"0F",x"C0",x"7C",x"3E",x"0B",x"E1",x"F0",x"0F",
		x"1F",x"80",x"F8",x"7C",x"13",x"C3",x"F0",x"1F",x"1F",x"80",x"78",x"FC",x"13",x"C3",x"F0",x"1E",
		x"0F",x"C0",x"F8",x"FC",x"07",x"C3",x"F0",x"1E",x"1F",x"84",x"F0",x"7C",x"27",x"C3",x"E0",x"1E",
		x"3F",x"01",x"F0",x"FC",x"0F",x"87",x"E0",x"3C",x"3F",x"01",x"E1",x"F8",x"1F",x"0F",x"C0",x"F8",
		x"7C",x"13",x"C3",x"F0",x"1E",x"1F",x"81",x"F0",x"FC",x"07",x"87",x"F0",x"1E",x"1F",x"09",x"F0",
		x"F8",x"07",x"8F",x"E0",x"78",x"3F",x"03",x"E1",x"F0",x"1E",x"1F",x"88",x"F0",x"FC",x"07",x"87",
		x"00",x"E2",x"38",x"3F",x"03",x"E1",x"F8",x"1E",x"1F",x"80",x"F0",x"FE",x"07",x"87",x"E1",x"38",
		x"1F",x"83",x"E1",x"F8",x"1E",x"0F",x"C0",x"F0",x"FC",x"0D",x"87",x"F0",x"78",x"3F",x"07",x"83",
		x"F0",x"3C",x"3F",x"03",x"C1",x"F8",x"9C",x"1F",x"81",x"E0",x"FC",x"1E",x"0F",x"C4",x"F0",x"FC",
		x"0F",x"07",x"C0",x"F8",x"7E",x"07",x"07",x"E2",x"78",x"7E",x"07",x"87",x"E0",x"3C",x"3F",x"03",
		x"C3",x"F0",x"3C",x"3F",x"03",x"C3",x"F0",x"3C",x"3F",x"03",x"C3",x"F0",x"2C",x"3F",x"22",x"C3",
		x"E2",x"2C",x"3F",x"06",x"C3",x"E2",x"3C",x"3F",x"21",x"C3",x"E4",x"78",x"3E",x"05",x"C7",x"E0",
		x"78",x"7E",x"05",x"87",x"E4",x"38",x"7E",x"0B",x"0F",x"C8",x"70",x"FC",x"87",x"1F",x"81",x"61",
		x"F9",x"0E",x"1F",x"83",x"C1",x"F2",x"3C",x"3E",x"23",x"87",x"E4",x"38",x"7C",x"87",x"0F",x"98",
		x"71",x"F9",x"0E",x"1F",x"81",x"C3",x"F0",x"5C",x"3E",x"21",x"87",x"E6",x"38",x"7C",x"47",x"0F",
		x"88",x"71",x"F9",x"0E",x"1F",x"11",x"C3",x"E6",x"1C",x"7C",x"87",x"0F",x"98",x"E1",x"F1",x"0E",
		x"3E",x"23",x"87",x"C8",x"38",x"FC",x"47",x"8F",x"80",x"E3",x"E2",x"1E",x"3E",x"23",x"87",x"8C",
		x"71",x"F0",x"C7",x"1E",x"31",x"C3",x"C7",x"1C",x"78",x"E1",x"8F",x"1C",x"71",x"E3",x"C6",x"1C",
		x"71",x"C7",x"87",x"18",x"F1",x"C7",x"1E",x"1C",x"63",x"C7",x"9C",x"70",x"79",x"8E",x"1E",x"75",
		x"C1",x"C7",x"3C",x"38",x"C7",x"87",x"1A",x"F0",x"E3",x"1E",x"1E",x"27",x"83",x"8D",x"78",x"38",
		x"AF",x"0E",x"33",x"E0",x"E2",x"7C",x"38",x"7F",x"07",x"07",x"E0",x"E0",x"FC",x"3C",x"1F",x"87",
		x"07",x"E0",x"71",x"FC",x"1C",x"1F",x"81",x"8B",x"F0",x"70",x"FE",x"0E",x"0F",x"C1",x"C3",x"F8",
		x"0F",x"38",x"3F",x"07",x"0F",x"C1",x"C1",x"FC",x"1C",x"3F",x"07",x"0F",x"E0",x"71",x"BC",x"1C",
		x"1F",x"83",x"87",x"E2",x"61",x"FC",x"0E",x"3F",x"03",x"87",x"E0",x"61",x"FC",x"5C",x"3B",x"13",
		x"86",x"E2",x"71",x"9C",x"4E",x"1F",x"19",x"8E",x"70",x"38",x"FC",x"27",x"39",x"C0",x"E3",x"71",
		x"B8",x"EE",x"07",x"1B",x"8D",x"C6",x"71",x"38",x"CC",x"66",x"3B",x"8C",x"C7",x"71",x"B8",x"CC",
		x"27",x"39",x"C0",x"E7",x"71",x"B8",x"CC",x"63",x"39",x"88",x"E7",x"71",x"19",x"CC",x"67",x"3B",
		x"88",x"C6",x"72",x"39",x"9C",x"C6",x"73",x"19",x"CC",x"62",x"73",x"B8",x"9C",x"6E",x"27",x"1D",
		x"88",x"CE",x"63",x"39",x"9C",x"8E",x"76",x"31",x"1B",x"C4",x"4E",x"73",x"13",x"9D",x"88",x"E7",
		x"62",x"3B",x"99",x"8E",x"C4",x"83",x"FB",x"01",x"FC",x"88",x"EE",x"62",x"3B",x"D8",x"1D",x"E6",
		x"07",x"79",x"83",x"BC",x"C0",x"EF",x"B0",x"37",x"9C",x"0D",x"E7",x"03",x"7B",x"80",x"DF",x"60",
		x"37",x"DC",x"04",x"FE",x"03",x"7B",x"C0",x"6F",x"78",x"0D",x"EE",x"07",x"77",x"81",x"CE",x"C6",
		x"3B",x"3C",x"13",x"BB",x"03",x"5D",x"86",x"37",x"26",x"65",x"D8",x"CB",x"24",x"E6",x"38",x"CE",
		x"67",x"64",x"D3",x"32",x"64",x"FB",x"26",x"61",x"BB",x"24",x"ED",x"99",x"99",x"39",x"16",x"72",
		x"4E",x"33",x"32",x"73",x"96",x"66",x"66",x"33",x"66",x"36",x"66",x"39",x"A6",x"71",x"98",x"9C",
		x"DD",x"91",x"99",x"99",x"B1",x"4C",x"E3",x"33",x"33",x"38",x"CC",x"CB",x"31",x"CC",x"E6",x"64",
		x"59",x"93",x"33",x"99",x"8B",x"33",x"8C",x"CB",x"1C",x"CC",x"C9",x"9C",x"CC",x"C9",x"9D",x"8C",
		x"66",x"CD",x"33",x"8C",x"E9",x"99",x"93",x"99",x"99",x"99",x"33",x"98",x"E6",x"66",x"2C",x"E0",
		x"00",x"00",x"00",x"AB",x"35",x"4C",x"65",x"9A",x"D9",x"8C",x"A6",x"B6",x"69",x"24",x"CD",x"B6",
		x"65",x"29",x"AD",x"B2",x"62",x"4C",x"DD",x"98",x"C9",x"9B",x"5B",x"32",x"8C",x"6D",x"B9",x"A4",
		x"99",x"B7",x"64",x"44",x"57",x"76",x"C9",x"25",x"77",x"6A",x"28",x"99",x"EE",x"D4",x"44",x"B5",
		x"D9",x"88",x"46",x"EB",x"99",x"89",x"99",x"EE",x"53",x"19",x"9C",x"F6",x"22",x"26",x"D9",x"98",
		x"C4",x"6E",x"F6",x"93",x"33",x"39",x"C8",x"85",x"76",x"79",x"26",x"31",x"76",x"C4",x"C6",x"76",
		x"7A",x"22",x"25",x"B3",x"91",x"85",x"CD",x"E9",x"14",x"CC",x"E6",x"64",x"67",x"37",x"A6",x"32",
		x"73",x"B3",x"42",x"9D",x"9B",x"33",x"19",x"99",x"C9",x"86",x"EE",x"B3",x"31",x"93",x"99",x"98",
		x"CE",x"CC",x"C6",x"66",x"67",x"32",x"33",x"BB",x"94",x"CC",x"99",x"CC",x"C4",x"F6",x"EA",x"66",
		x"62",x"76",x"31",x"4F",x"B4",x"4B",x"13",x"33",x"B0",x"9D",x"B9",x"13",x"66",x"33",x"63",x"3B",
		x"39",x"0D",x"60",x"B6",x"66",x"27",x"E9",x"33",x"31",x"B3",x"91",x"9C",x"E1",x"33",x"A4",x"F9",
		x"4C",x"6E",x"33",x"91",x"9D",x"98",x"EC",x"E5",x"36",x"27",x"33",x"19",x"B8",x"33",x"49",x"D8",
		x"C6",x"EE",x"98",x"9C",x"4E",x"62",x"67",x"8C",x"C8",x"D9",x"C4",x"EE",x"33",x"13",x"93",x"89",
		x"9E",x"61",x"9E",x"CD",x"66",x"71",x"46",x"76",x"63",x"33",x"C8",x"4F",x"26",x"53",x"3C",x"C1",
		x"E4",x"EC",x"67",x"D0",x"7C",x"1B",x"99",x"E1",x"1E",x"0D",x"C6",x"7C",x"0F",x"86",x"C3",x"F8",
		x"0F",x"07",x"C2",x"FC",x"0F",x"0D",x"C3",x"F0",x"1E",x"1B",x"8F",x"C0",x"E4",x"2E",x"37",x"83",
		x"B1",x"B8",x"DC",x"0B",x"85",x"C2",x"F0",x"3C",x"3E",x"17",x"81",x"E1",x"71",x"F8",x"1E",x"1B",
		x"0F",x"8D",x"C1",x"E1",x"B8",x"DC",x"1E",x"1B",x"8D",x"C1",x"E1",x"B8",x"D8",x"2E",x"33",x"1F",
		x"83",x"63",x"E3",x"30",x"D8",x"EE",x"37",x"07",x"8D",x"C6",x"E0",x"71",x"38",x"F8",x"4C",x"2F",
		x"33",x"83",x"8D",x"8E",x"E2",x"72",x"71",x"BC",x"1C",x"9C",x"6E",x"0E",x"67",x"1B",x"83",x"39",
		x"CD",x"C1",x"CC",x"E2",x"70",x"F2",x"63",x"B8",x"73",x"38",x"D8",x"39",x"9C",x"CE",x"1E",x"CC",
		x"67",x"1C",x"67",x"1B",x"86",x"37",x"19",x"C7",x"19",x"CC",x"C3",x"8C",x"E3",x"70",x"E6",x"71",
		x"B8",x"71",x"39",x"CC",x"1C",x"CE",x"67",x"0E",x"27",x"1B",x"87",x"19",x"8E",x"E1",x"C4",x"E3",
		x"78",x"78",x"3C",x"DC",x"1E",x"66",x"3B",x"83",x"9D",x"8C",x"E0",x"F0",x"F1",x"B8",x"38",x"DE",
		x"36",x"0F",x"0B",x"86",x"E1",x"F0",x"78",x"DC",x"1E",x"17",x"19",x"C1",x"E2",x"71",x"BC",x"1E",
		x"27",x"9B",x"C0",x"F0",x"78",x"FC",x"0F",x"07",x"89",x"E2",x"70",x"9C",x"7E",x"07",x"89",x"C6",
		x"F0",x"3C",x"4E",x"37",x"C0",x"E3",x"71",x"9E",x"43",x"89",x"E3",x"70",x"5C",x"27",x"0B",x"E1",
		x"98",x"9E",x"37",x"82",x"71",x"38",x"DF",x"04",x"E6",x"61",x"3E",x"33",x"0D",x"C3",x"78",x"53",
		x"13",x"8E",x"F1",x"1C",x"93",x"1D",x"E0",x"B1",x"46",x"7B",x"89",x"32",x"8D",x"3B",x"84",x"94",
		x"C5",x"9C",x"E2",x"4C",x"67",x"AE",x"72",x"22",x"4E",x"6F",x"9A",x"14",x"62",x"CF",x"7B",x"21",
		x"42",x"36",x"EF",x"64",x"98",x"C6",x"6E",x"F6",x"98",x"C2",x"2C",x"EF",x"34",x"91",x"11",x"5B",
		x"7A",x"D1",x"24",x"49",x"B6",x"E7",x"24",x"92",x"46",x"DD",x"DA",x"49",x"32",x"4A",x"CF",x"59",
		x"25",x"2A",x"56",x"77",x"35",x"14",x"AA",x"99",x"B7",x"35",x"25",x"2A",x"65",x"AD",x"B5",x"30",
		x"0F",x"0C",x"00",x"0F",x"0F",x"0B",x"0F",x"00",x"0F",x"0A",x"0F",x"0D",x"0F",x"0C",x"0F",x"03",
		x"0F",x"03",x"0B",x"0F",x"0F",x"00",x"0D",x"03",x"0F",x"0F",x"0C",x"00",x"0F",x"0F",x"0A",x"00",
		x"0F",x"0F",x"0A",x"03",x"0F",x"00",x"03",x"05",x"0F",x"0D",x"00",x"05",x"0F",x"0C",x"03",x"0A",
		x"0F",x"00",x"00",x"0C",x"0F",x"0F",x"0B",x"03",x"0F",x"0E",x"0A",x"0C",x"0F",x"0B",x"0F",x"0F",
		x"0F",x"0C",x"00",x"0F",x"0F",x"0B",x"0F",x"00",x"0F",x"0A",x"0F",x"0D",x"0F",x"03",x"0A",x"00",
		x"0F",x"03",x"0A",x"00",x"0F",x"03",x"0A",x"00",x"0F",x"03",x"0A",x"00",x"0F",x"0F",x"0A",x"00",
		x"0F",x"0F",x"0A",x"03",x"0F",x"00",x"03",x"05",x"0F",x"0D",x"00",x"05",x"0F",x"0C",x"03",x"0A",
		x"0F",x"00",x"00",x"0C",x"0F",x"0F",x"0B",x"03",x"0F",x"0E",x"0A",x"0C",x"0F",x"0B",x"0F",x"0F",
		x"0F",x"0C",x"00",x"0F",x"0F",x"0B",x"0F",x"00",x"0F",x"0A",x"0F",x"0D",x"0F",x"0A",x"0F",x"00",
		x"0F",x"0A",x"0F",x"00",x"0F",x"0A",x"0F",x"00",x"0F",x"0A",x"0F",x"00",x"0F",x"0F",x"0A",x"00",
		x"0F",x"0F",x"0A",x"03",x"0F",x"00",x"03",x"05",x"0F",x"0D",x"00",x"05",x"0F",x"0C",x"03",x"0A",
		x"0F",x"00",x"00",x"0C",x"0F",x"0F",x"0B",x"03",x"0F",x"0E",x"0A",x"0C",x"0F",x"0B",x"0F",x"0F",
		x"0F",x"0C",x"00",x"0F",x"0F",x"0B",x"0F",x"00",x"0F",x"0A",x"0F",x"0D",x"0F",x"0C",x"00",x"0B",
		x"0F",x"0C",x"00",x"0B",x"0F",x"0C",x"00",x"0B",x"0F",x"0C",x"00",x"0B",x"0F",x"0F",x"0A",x"00",
		x"0F",x"0F",x"0A",x"03",x"0F",x"00",x"03",x"05",x"0F",x"0D",x"00",x"05",x"0F",x"0C",x"03",x"0A",
		x"0F",x"00",x"00",x"0C",x"0F",x"0F",x"0B",x"03",x"0F",x"0E",x"0A",x"0C",x"0F",x"0B",x"0F",x"0F",
		x"0F",x"06",x"0E",x"01",x"0F",x"00",x"01",x"00",x"0F",x"00",x"01",x"0F",x"0F",x"0F",x"01",x"0E",
		x"0F",x"01",x"00",x"01",x"0F",x"00",x"01",x"00",x"0F",x"01",x"0F",x"0E",x"0F",x"05",x"00",x"00",
		x"0F",x"05",x"00",x"01",x"0F",x"00",x"01",x"01",x"0F",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"00",
		x"0F",x"00",x"0E",x"0F",x"0F",x"01",x"00",x"01",x"0F",x"02",x"00",x"0F",x"0F",x"00",x"01",x"0F",
		x"0F",x"06",x"0E",x"01",x"0F",x"00",x"01",x"00",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"00",x"00",
		x"0F",x"01",x"00",x"00",x"0F",x"01",x"00",x"00",x"0F",x"01",x"00",x"00",x"0F",x"05",x"00",x"00",
		x"0F",x"05",x"00",x"01",x"0F",x"00",x"01",x"01",x"0F",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"00",
		x"0F",x"00",x"0E",x"0F",x"0F",x"01",x"00",x"01",x"0F",x"02",x"00",x"0F",x"0F",x"00",x"01",x"0F",
		x"0F",x"06",x"0E",x"01",x"0F",x"00",x"01",x"00",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"07",x"0E",
		x"0F",x"01",x"07",x"0E",x"0F",x"01",x"07",x"0E",x"0F",x"01",x"07",x"0E",x"0F",x"05",x"00",x"00",
		x"0F",x"05",x"00",x"01",x"0F",x"00",x"01",x"01",x"0F",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"00",
		x"0F",x"00",x"0E",x"0F",x"0F",x"01",x"00",x"01",x"0F",x"02",x"00",x"0F",x"0F",x"00",x"01",x"0F",
		x"0F",x"06",x"0E",x"01",x"0F",x"00",x"01",x"00",x"0F",x"00",x"01",x"0F",x"0F",x"0F",x"0E",x"00",
		x"0F",x"0F",x"0E",x"00",x"0F",x"0F",x"0E",x"00",x"0F",x"0F",x"0E",x"00",x"0F",x"05",x"00",x"00",
		x"0F",x"05",x"00",x"01",x"0F",x"00",x"01",x"01",x"0F",x"0F",x"00",x"01",x"0F",x"0F",x"01",x"00",
		x"0F",x"00",x"0E",x"0F",x"0F",x"01",x"00",x"01",x"0F",x"02",x"00",x"0F",x"0F",x"00",x"01",x"0F",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"01",x"01",x"02",x"06",x"06",x"04",x"06",x"06",x"06",x"06",x"03",x"06",x"03",x"04",x"03",
		x"06",x"06",x"06",x"06",x"04",x"03",x"04",x"05",x"04",x"06",x"05",x"03",x"05",x"03",x"06",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",
		x"7F",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7C",x"7A",x"6D",x"4D",x"37",x"34",x"40",
		x"52",x"7F",x"AD",x"BD",x"C2",x"BF",x"B7",x"B0",x"A7",x"9E",x"8F",x"6A",x"4D",x"41",x"46",x"52",
		x"77",x"A5",x"B9",x"BD",x"B9",x"B1",x"A8",x"A1",x"98",x"8F",x"76",x"53",x"3E",x"3B",x"41",x"58",
		x"87",x"A7",x"B1",x"B1",x"AD",x"A5",x"9E",x"96",x"8D",x"86",x"6B",x"4C",x"3B",x"3A",x"43",x"5B",
		x"87",x"A4",x"AD",x"AD",x"A7",x"A1",x"99",x"93",x"8C",x"84",x"6E",x"50",x"3E",x"3B",x"41",x"55",
		x"80",x"9F",x"A8",x"AB",x"A5",x"9F",x"99",x"93",x"8D",x"87",x"7C",x"5F",x"47",x"3E",x"41",x"4C",
		x"6A",x"92",x"A4",x"AA",x"A7",x"A2",x"9C",x"95",x"90",x"8A",x"84",x"76",x"59",x"46",x"41",x"47",
		x"55",x"77",x"98",x"A4",x"A8",x"A5",x"9F",x"99",x"93",x"8F",x"89",x"84",x"76",x"5B",x"49",x"46",
		x"4A",x"58",x"79",x"98",x"A4",x"A7",x"A4",x"9F",x"99",x"93",x"8F",x"89",x"84",x"79",x"61",x"4F",
		x"49",x"4C",x"56",x"71",x"92",x"A1",x"A4",x"A2",x"9E",x"98",x"93",x"8F",x"8A",x"86",x"7F",x"6A",
		x"56",x"4C",x"4D",x"55",x"68",x"89",x"9B",x"A2",x"A2",x"9F",x"99",x"95",x"90",x"8C",x"87",x"83",
		x"76",x"61",x"52",x"4F",x"53",x"5E",x"7A",x"93",x"9E",x"A2",x"9F",x"9B",x"96",x"92",x"8D",x"89",
		x"84",x"80",x"6E",x"5B",x"52",x"52",x"58",x"67",x"84",x"98",x"9F",x"9F",x"9C",x"98",x"93",x"90",
		x"8C",x"87",x"83",x"7D",x"6B",x"5B",x"53",x"55",x"5B",x"6D",x"87",x"98",x"9C",x"9C",x"99",x"95",
		x"90",x"8D",x"89",x"86",x"83",x"7C",x"6B",x"5C",x"56",x"58",x"5E",x"6E",x"89",x"96",x"9B",x"9B",
		x"99",x"95",x"90",x"8C",x"89",x"86",x"83",x"7D",x"6E",x"5F",x"59",x"59",x"5F",x"6D",x"84",x"93",
		x"99",x"9B",x"98",x"93",x"90",x"8C",x"89",x"86",x"83",x"7F",x"71",x"64",x"5C",x"5B",x"5F",x"6B",
		x"81",x"90",x"98",x"98",x"96",x"93",x"8F",x"8C",x"89",x"86",x"83",x"80",x"77",x"68",x"5F",x"5E",
		x"61",x"68",x"7C",x"8D",x"95",x"98",x"96",x"93",x"90",x"8C",x"89",x"86",x"84",x"81",x"7C",x"6D",
		x"62",x"5F",x"61",x"65",x"74",x"87",x"92",x"96",x"95",x"92",x"8F",x"8C",x"89",x"87",x"84",x"81",
		x"7F",x"76",x"68",x"62",x"62",x"65",x"6D",x"80",x"8D",x"93",x"95",x"92",x"90",x"8D",x"8A",x"87",
		x"86",x"83",x"80",x"7C",x"70",x"65",x"62",x"64",x"68",x"76",x"87",x"90",x"93",x"92",x"90",x"8D",
		x"8A",x"89",x"86",x"83",x"81",x"7F",x"77",x"6B",x"64",x"64",x"67",x"6D",x"7D",x"8C",x"90",x"93",
		x"92",x"8F",x"8C",x"8A",x"87",x"84",x"83",x"81",x"7D",x"73",x"6A",x"65",x"67",x"6A",x"73",x"83",
		x"8D",x"90",x"90",x"8F",x"8D",x"8A",x"87",x"86",x"84",x"81",x"80",x"7A",x"70",x"68",x"67",x"68",
		x"6D",x"77",x"86",x"8D",x"90",x"8F",x"8D",x"8C",x"89",x"87",x"84",x"83",x"80",x"7F",x"79",x"6E",
		x"6A",x"68",x"6B",x"70",x"7D",x"89",x"8D",x"8F",x"8F",x"8C",x"8A",x"87",x"86",x"84",x"83",x"81",
		x"7F",x"77",x"6E",x"6A",x"6A",x"6D",x"73",x"80",x"8A",x"8D",x"8F",x"8D",x"8C",x"89",x"87",x"84",
		x"83",x"81",x"80",x"7D",x"76",x"6E",x"6B",x"6B",x"6E",x"76",x"81",x"8A",x"8D",x"8D",x"8C",x"8A",
		x"87",x"86",x"84",x"83",x"81",x"80",x"7D",x"74",x"6E",x"6D",x"6D",x"70",x"77",x"83",x"8A",x"8D",
		x"8D",x"8C",x"8A",x"87",x"86",x"84",x"83",x"81",x"80",x"7C",x"74",x"6E",x"6D",x"6E",x"71",x"79",
		x"84",x"8A",x"8C",x"8C",x"8A",x"89",x"87",x"84",x"83",x"81",x"81",x"80",x"7D",x"76",x"70",x"6E",
		x"6E",x"71",x"77",x"81",x"89",x"8C",x"8C",x"8A",x"89",x"87",x"86",x"84",x"83",x"81",x"80",x"80",
		x"7F",x"7C",x"76",x"70",x"6E",x"6E",x"71",x"77",x"81",x"89",x"8A",x"8A",x"8A",x"87",x"86",x"86",
		x"84",x"83",x"81",x"81",x"81",x"80",x"80",x"86",x"92",x"96",x"96",x"93",x"8D",x"81",x"73",x"6A",
		x"65",x"65",x"67",x"6A",x"6D",x"6E",x"71",x"74",x"77",x"79",x"7C",x"7F",x"89",x"93",x"98",x"98",
		x"95",x"8F",x"80",x"73",x"6B",x"68",x"6A",x"6D",x"70",x"73",x"76",x"79",x"7A",x"7D",x"7F",x"81",
		x"8A",x"96",x"9B",x"9B",x"98",x"92",x"84",x"76",x"6E",x"6B",x"6D",x"6E",x"71",x"74",x"77",x"79",
		x"7C",x"7D",x"80",x"83",x"8F",x"99",x"9C",x"9B",x"96",x"8F",x"7F",x"73",x"6D",x"6B",x"6D",x"6E",
		x"73",x"74",x"77",x"7A",x"7C",x"7F",x"81",x"89",x"95",x"9B",x"9B",x"98",x"93",x"84",x"76",x"6E",
		x"6B",x"6D",x"6E",x"71",x"74",x"77",x"7A",x"7C",x"7F",x"80",x"87",x"95",x"9B",x"9B",x"98",x"93",
		x"87",x"77",x"6E",x"6B",x"6D",x"6E",x"71",x"74",x"76",x"79",x"7C",x"7D",x"80",x"87",x"93",x"9B",
		x"9B",x"96",x"92",x"84",x"76",x"6E",x"6B",x"6D",x"6E",x"71",x"74",x"77",x"79",x"7C",x"7D",x"80",
		x"8A",x"96",x"9B",x"99",x"96",x"8F",x"80",x"73",x"6D",x"6B",x"6D",x"70",x"73",x"74",x"77",x"7A",
		x"7C",x"7F",x"83",x"8F",x"98",x"9B",x"98",x"93",x"8A",x"7A",x"70",x"6B",x"6B",x"6D",x"70",x"73",
		x"76",x"77",x"7A",x"7D",x"7F",x"89",x"95",x"99",x"99",x"96",x"8F",x"81",x"73",x"6D",x"6B",x"6D",
		x"70",x"73",x"74",x"77",x"79",x"7C",x"7F",x"84",x"90",x"98",x"99",x"96",x"92",x"86",x"77",x"6E",
		x"6B",x"6D",x"6E",x"71",x"74",x"77",x"79",x"7C",x"7F",x"81",x"8D",x"96",x"99",x"98",x"93",x"8A",
		x"7C",x"71",x"6D",x"6D",x"6E",x"71",x"74",x"76",x"79",x"7A",x"7D",x"80",x"8A",x"95",x"98",x"96",
		x"93",x"8D",x"7F",x"73",x"6E",x"6D",x"6E",x"71",x"74",x"76",x"79",x"7A",x"7D",x"7F",x"87",x"92",
		x"96",x"98",x"95",x"8F",x"81",x"74",x"6E",x"6D",x"6E",x"71",x"74",x"76",x"79",x"7A",x"7D",x"7F",
		x"86",x"90",x"96",x"96",x"93",x"8F",x"83",x"76",x"70",x"6E",x"6E",x"71",x"74",x"76",x"79",x"7A",
		x"7D",x"7F",x"84",x"8F",x"95",x"95",x"93",x"8F",x"83",x"77",x"71",x"70",x"70",x"71",x"74",x"76",
		x"79",x"7A",x"7D",x"7F",x"83",x"8D",x"92",x"93",x"92",x"8F",x"84",x"79",x"73",x"70",x"71",x"73",
		x"76",x"77",x"79",x"7A",x"7C",x"7F",x"83",x"8C",x"92",x"93",x"92",x"8F",x"84",x"7A",x"74",x"71",
		x"71",x"73",x"76",x"77",x"79",x"7A",x"7D",x"7F",x"81",x"8A",x"90",x"92",x"90",x"8D",x"86",x"7A",
		x"74",x"71",x"73",x"74",x"76",x"77",x"7A",x"7A",x"7C",x"7F",x"81",x"89",x"8F",x"90",x"8F",x"8C",
		x"86",x"7C",x"76",x"73",x"73",x"74",x"76",x"79",x"79",x"7A",x"7D",x"7F",x"80",x"87",x"8D",x"8F",
		x"8D",x"8C",x"86",x"7C",x"77",x"74",x"74",x"76",x"77",x"79",x"7A",x"7C",x"7D",x"7D",x"80",x"86",
		x"8C",x"8D",x"8D",x"8C",x"86",x"7F",x"77",x"76",x"74",x"76",x"77",x"79",x"7A",x"7C",x"7C",x"7D",
		x"80",x"84",x"8A",x"8D",x"8C",x"8A",x"86",x"7F",x"79",x"76",x"76",x"76",x"77",x"79",x"7A",x"7C",
		x"7D",x"7F",x"7F",x"83",x"8A",x"8C",x"8C",x"8A",x"87",x"7F",x"79",x"76",x"76",x"77",x"77",x"79",
		x"7A",x"7C",x"7D",x"7F",x"7F",x"84",x"89",x"8A",x"8C",x"8A",x"87",x"80",x"7A",x"77",x"77",x"77",
		x"79",x"7A",x"7A",x"7C",x"7D",x"7F",x"7F",x"83",x"87",x"8A",x"8A",x"89",x"87",x"80",x"7A",x"79",
		x"77",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7F",x"7F",x"81",x"86",x"89",x"89",x"89",x"86",x"80",
		x"7C",x"79",x"77",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7D",x"7F",x"81",x"86",x"89",x"89",x"89",
		x"87",x"81",x"7C",x"79",x"79",x"79",x"7A",x"7A",x"7C",x"7D",x"7D",x"7F",x"7F",x"81",x"86",x"87",
		x"89",x"87",x"86",x"81",x"7C",x"79",x"79",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7F",x"7F",x"81",
		x"86",x"87",x"87",x"87",x"84",x"80",x"7C",x"7A",x"79",x"7A",x"7A",x"7C",x"7C",x"7D",x"7D",x"7F",
		x"83",x"86",x"87",x"86",x"86",x"83",x"7D",x"7A",x"79",x"7A",x"7A",x"7C",x"7C",x"7D",x"7D",x"7F",
		x"83",x"86",x"86",x"86",x"84",x"81",x"7D",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7D",x"7F",x"81",
		x"84",x"86",x"86",x"84",x"83",x"7F",x"7C",x"7A",x"7A",x"7A",x"7C",x"7D",x"7D",x"7F",x"81",x"84",
		x"86",x"84",x"83",x"81",x"7D",x"7A",x"7A",x"7A",x"7A",x"7C",x"7D",x"7D",x"80",x"83",x"84",x"84",
		x"84",x"83",x"7F",x"7C",x"7A",x"7A",x"7C",x"7C",x"7D",x"7D",x"80",x"83",x"84",x"84",x"84",x"83",
		x"7F",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7F",x"80",x"83",x"84",x"84",x"84",x"81",x"7F",x"7C",
		x"7C",x"7C",x"7C",x"7D",x"7D",x"7F",x"81",x"83",x"84",x"84",x"83",x"80",x"7D",x"7C",x"7C",x"7C",
		x"7C",x"7D",x"7F",x"80",x"83",x"84",x"84",x"83",x"81",x"7F",x"7D",x"7C",x"7C",x"7D",x"7D",x"7F",
		x"80",x"81",x"83",x"83",x"83",x"81",x"7F",x"7D",x"7C",x"7C",x"7C",x"7D",x"7D",x"80",x"81",x"83",
		x"83",x"83",x"81",x"7F",x"7D",x"7C",x"7C",x"7C",x"7D",x"7D",x"80",x"81",x"81",x"83",x"83",x"81",
		x"7F",x"7D",x"7C",x"7C",x"7C",x"7D",x"7F",x"80",x"83",x"83",x"83",x"83",x"81",x"7F",x"7D",x"7C",
		x"7C",x"7D",x"7D",x"7F",x"80",x"81",x"83",x"83",x"81",x"80",x"7D",x"7C",x"7C",x"7C",x"7D",x"7D",
		x"80",x"81",x"81",x"83",x"81",x"81",x"7F",x"7D",x"7C",x"7D",x"7D",x"7D",x"7F",x"80",x"81",x"83",
		x"83",x"81",x"80",x"7F",x"7D",x"7D",x"7C",x"7D",x"7D",x"7F",x"80",x"81",x"83",x"81",x"81",x"7F",
		x"7D",x"7D",x"7C",x"7D",x"7D",x"7F",x"80",x"81",x"81",x"81",x"81",x"80",x"7F",x"7D",x"7D",x"7D",
		x"7D",x"7F",x"80",x"81",x"81",x"81",x"81",x"81",x"7F",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"80",
		x"81",x"81",x"81",x"81",x"80",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"80",x"81",x"81",x"81",x"81",
		x"80",x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"80",x"81",x"81",x"81",x"80",x"7F",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7F",x"80",x"81",x"81",x"81",x"81",x"80",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",
		x"80",x"81",x"81",x"81",x"81",x"80",x"7F",x"7D",x"7D",x"7F",x"7F",x"7F",x"80",x"81",x"81",x"81",
		x"81",x"80",x"7F",x"7D",x"7D",x"7D",x"7D",x"7F",x"80",x"80",x"81",x"81",x"81",x"80",x"7F",x"7D",
		x"7D",x"7D",x"7D",x"7F",x"80",x"81",x"81",x"81",x"81",x"80",x"7F",x"7D",x"7D",x"7D",x"7D",x"7F",
		x"7F",x"80",x"81",x"81",x"81",x"80",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7F",x"80",x"80",x"81",
		x"81",x"80",x"80",x"7F",x"7D",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"81",x"81",x"80",x"80",x"7F",
		x"7D",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"81",x"81",x"80",x"80",x"7F",x"7D",x"7D",x"7D",x"7D",
		x"7F",x"80",x"80",x"81",x"81",x"80",x"80",x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"80",
		x"81",x"81",x"80",x"7F",x"7F",x"7D",x"7F",x"7F",x"7F",x"80",x"80",x"81",x"81",x"80",x"80",x"7F",
		x"7F",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"80",x"80",x"81",x"80",x"7F",x"7D",x"7D",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"81",x"80",x"80",x"80",x"7F",x"7D",x"7D",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"81",x"80",x"80",x"80",
		x"7F",x"7D",x"7F",x"7D",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"81",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7F",x"7F",x"7F",x"7D",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",
		x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",
		x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",x"7A",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"80",x"7E",x"7E",x"7E",x"7E",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",
		x"7A",x"7A",x"7A",x"7C",x"7E",x"80",x"82",x"84",x"86",x"84",x"84",x"82",x"82",x"7C",x"7A",x"78",
		x"76",x"76",x"76",x"76",x"78",x"78",x"7A",x"7C",x"7C",x"7E",x"84",x"88",x"8C",x"8E",x"8C",x"8C",
		x"8A",x"88",x"80",x"7A",x"74",x"72",x"72",x"72",x"72",x"74",x"76",x"78",x"78",x"7A",x"7C",x"80",
		x"88",x"8E",x"94",x"96",x"96",x"94",x"92",x"8E",x"84",x"7A",x"72",x"6E",x"6C",x"6C",x"6E",x"6E",
		x"70",x"72",x"76",x"78",x"7A",x"7C",x"82",x"8A",x"92",x"98",x"9A",x"9C",x"9C",x"9A",x"94",x"88",
		x"7A",x"70",x"6C",x"68",x"68",x"6A",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7C",x"7E",x"84",x"8E",
		x"94",x"9A",x"9C",x"9E",x"9E",x"9C",x"96",x"84",x"76",x"6E",x"68",x"64",x"66",x"66",x"6A",x"6C",
		x"70",x"72",x"76",x"78",x"7C",x"7E",x"82",x"88",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"94",
		x"84",x"76",x"6C",x"66",x"64",x"64",x"66",x"68",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7E",x"80",
		x"84",x"8A",x"92",x"98",x"9E",x"A0",x"A0",x"A0",x"9C",x"8E",x"7C",x"70",x"68",x"64",x"64",x"64",
		x"66",x"68",x"6C",x"6E",x"72",x"74",x"78",x"7A",x"7E",x"80",x"82",x"86",x"8E",x"96",x"9C",x"9E",
		x"A0",x"A0",x"A0",x"9A",x"8A",x"78",x"6E",x"68",x"64",x"62",x"64",x"66",x"6A",x"6C",x"6E",x"72",
		x"74",x"78",x"7A",x"7E",x"80",x"82",x"84",x"8C",x"94",x"9A",x"9C",x"A0",x"A0",x"A0",x"9E",x"94",
		x"80",x"74",x"6A",x"64",x"62",x"64",x"66",x"68",x"6A",x"6E",x"70",x"72",x"76",x"78",x"7A",x"7C",
		x"7E",x"80",x"82",x"86",x"8E",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9C",x"8C",x"7C",x"70",x"68",
		x"64",x"62",x"64",x"66",x"68",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7C",x"7E",x"80",x"82",x"82",
		x"84",x"88",x"90",x"98",x"9C",x"A0",x"A0",x"A2",x"A0",x"98",x"88",x"78",x"6C",x"66",x"62",x"62",
		x"64",x"66",x"68",x"6C",x"6E",x"70",x"74",x"76",x"78",x"7C",x"7C",x"7E",x"80",x"82",x"84",x"86",
		x"8E",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"80",x"72",x"68",x"64",x"62",x"62",x"64",
		x"66",x"68",x"6C",x"70",x"72",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"82",x"84",x"86",x"88",
		x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"A0",x"9A",x"8A",x"7A",x"6C",x"64",x"62",x"60",x"62",x"64",
		x"66",x"6A",x"6C",x"70",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"82",x"84",x"86",x"86",
		x"8C",x"92",x"98",x"9C",x"A0",x"A2",x"A0",x"A0",x"98",x"86",x"74",x"6A",x"64",x"60",x"60",x"62",
		x"64",x"66",x"6A",x"6C",x"70",x"74",x"76",x"7A",x"7C",x"7E",x"7E",x"80",x"82",x"84",x"84",x"86",
		x"86",x"88",x"8E",x"96",x"9A",x"9E",x"A0",x"A2",x"A0",x"9C",x"92",x"7E",x"70",x"68",x"62",x"60",
		x"60",x"62",x"64",x"68",x"6C",x"70",x"72",x"74",x"78",x"7A",x"7C",x"7E",x"80",x"80",x"82",x"82",
		x"84",x"84",x"86",x"86",x"8A",x"92",x"98",x"9C",x"9E",x"A0",x"A0",x"9E",x"9A",x"8C",x"7A",x"6E",
		x"66",x"62",x"60",x"62",x"64",x"66",x"68",x"6C",x"70",x"72",x"74",x"78",x"7A",x"7C",x"7E",x"80",
		x"82",x"82",x"82",x"84",x"84",x"84",x"86",x"86",x"8C",x"94",x"9A",x"9E",x"9E",x"A0",x"A0",x"9E",
		x"98",x"86",x"74",x"68",x"62",x"60",x"60",x"62",x"64",x"66",x"6A",x"6E",x"70",x"74",x"76",x"78",
		x"7A",x"7C",x"7E",x"80",x"80",x"80",x"82",x"84",x"84",x"86",x"86",x"8C",x"94",x"98",x"9C",x"9E",
		x"A0",x"A0",x"9E",x"9A",x"8A",x"78",x"6C",x"64",x"60",x"60",x"60",x"62",x"66",x"68",x"6C",x"6E",
		x"72",x"74",x"78",x"7A",x"7C",x"7E",x"7E",x"80",x"82",x"82",x"84",x"84",x"84",x"88",x"90",x"98",
		x"9C",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"7E",x"70",x"66",x"62",x"60",x"60",x"62",x"64",x"68",
		x"6C",x"6E",x"70",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"82",x"84",x"84",x"86",x"8C",
		x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"A0",x"9A",x"88",x"78",x"6C",x"64",x"60",x"60",x"62",x"64",
		x"66",x"6A",x"6E",x"70",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"82",x"84",x"86",x"88",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"A0",x"98",x"86",x"76",x"6A",x"64",x"60",x"60",x"62",
		x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"7A",x"7C",x"7E",x"7E",x"80",x"82",x"82",x"84",x"86",
		x"88",x"90",x"96",x"9C",x"9E",x"A2",x"A2",x"A0",x"9E",x"92",x"80",x"70",x"68",x"62",x"60",x"62",
		x"62",x"64",x"68",x"6C",x"6E",x"72",x"74",x"76",x"7A",x"7C",x"7E",x"80",x"82",x"84",x"84",x"86",
		x"8A",x"90",x"96",x"9C",x"A0",x"A0",x"A2",x"A0",x"9E",x"90",x"7E",x"70",x"68",x"64",x"62",x"62",
		x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"80",x"82",x"84",x"86",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"96",x"84",x"74",x"6A",x"64",x"60",x"60",x"62",
		x"64",x"68",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7C",x"7E",x"80",x"82",x"82",x"84",x"88",x"90",
		x"96",x"9C",x"A0",x"A2",x"A2",x"A0",x"9E",x"92",x"7E",x"70",x"66",x"62",x"60",x"60",x"62",x"66",
		x"68",x"6C",x"70",x"72",x"76",x"78",x"7A",x"7E",x"7E",x"82",x"82",x"88",x"90",x"98",x"9C",x"A0",
		x"A2",x"A2",x"A0",x"9C",x"8C",x"7A",x"6E",x"66",x"62",x"60",x"62",x"64",x"68",x"6A",x"6E",x"70",
		x"74",x"76",x"7A",x"7C",x"7E",x"82",x"84",x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"94",
		x"80",x"72",x"68",x"64",x"62",x"62",x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"7A",x"7C",x"7E",
		x"82",x"88",x"90",x"98",x"9C",x"A0",x"A2",x"A2",x"A0",x"9C",x"8A",x"78",x"6C",x"66",x"64",x"62",
		x"64",x"66",x"68",x"6C",x"6E",x"72",x"74",x"78",x"7A",x"7E",x"82",x"8A",x"94",x"98",x"9E",x"A0",
		x"A2",x"A2",x"9E",x"94",x"80",x"72",x"6A",x"64",x"62",x"64",x"64",x"68",x"6A",x"6E",x"72",x"74",
		x"78",x"7C",x"7E",x"84",x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"9C",x"8E",x"7C",x"6E",x"66",
		x"64",x"62",x"62",x"64",x"68",x"6C",x"6E",x"72",x"76",x"78",x"7C",x"80",x"8A",x"92",x"98",x"9C",
		x"A0",x"A0",x"A0",x"9C",x"90",x"7C",x"6E",x"68",x"62",x"62",x"64",x"66",x"68",x"6C",x"6E",x"72",
		x"76",x"7A",x"7E",x"84",x"8E",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"98",x"86",x"76",x"6C",x"64",
		x"62",x"62",x"64",x"66",x"6A",x"6E",x"70",x"74",x"78",x"7C",x"82",x"8C",x"94",x"9A",x"9E",x"A0",
		x"A0",x"A0",x"98",x"86",x"76",x"6C",x"66",x"64",x"62",x"64",x"68",x"6A",x"6E",x"72",x"76",x"78",
		x"7E",x"86",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"90",x"7E",x"70",x"68",x"64",x"64",x"64",
		x"66",x"68",x"6C",x"70",x"74",x"78",x"7C",x"84",x"8E",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"92",
		x"80",x"72",x"68",x"64",x"64",x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"7C",x"86",x"90",x"96",
		x"9C",x"9E",x"A0",x"A0",x"9E",x"8E",x"7C",x"6E",x"66",x"64",x"62",x"64",x"66",x"68",x"6C",x"70",
		x"74",x"7A",x"82",x"8E",x"96",x"9A",x"9E",x"A0",x"A0",x"9E",x"94",x"82",x"74",x"6A",x"66",x"64",
		x"64",x"66",x"68",x"6C",x"70",x"74",x"78",x"80",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9E",x"96",
		x"84",x"74",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"78",x"80",x"8A",x"92",x"98",
		x"9C",x"A0",x"A0",x"9E",x"94",x"80",x"72",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",
		x"7A",x"84",x"8E",x"94",x"9A",x"9E",x"9E",x"9E",x"9C",x"8C",x"7C",x"6E",x"66",x"64",x"64",x"64",
		x"68",x"6C",x"6E",x"72",x"76",x"80",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9E",x"92",x"80",x"72",
		x"6A",x"66",x"64",x"66",x"68",x"6A",x"6E",x"72",x"76",x"7E",x"88",x"90",x"98",x"9A",x"9E",x"9E",
		x"9E",x"96",x"84",x"74",x"6C",x"66",x"64",x"64",x"66",x"6A",x"6C",x"70",x"74",x"7C",x"86",x"90",
		x"96",x"9C",x"9E",x"9E",x"9E",x"96",x"84",x"74",x"6A",x"66",x"64",x"64",x"66",x"6A",x"6C",x"70",
		x"76",x"7E",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9E",x"94",x"80",x"72",x"6A",x"66",x"64",x"66",
		x"68",x"6A",x"6E",x"72",x"78",x"82",x"8C",x"92",x"9A",x"9E",x"9E",x"9E",x"9C",x"8C",x"7A",x"6E",
		x"66",x"62",x"62",x"64",x"68",x"6C",x"70",x"74",x"7C",x"88",x"90",x"98",x"9C",x"9E",x"9E",x"9E",
		x"96",x"84",x"74",x"6A",x"66",x"64",x"66",x"66",x"6A",x"6E",x"72",x"78",x"82",x"8C",x"94",x"98",
		x"9C",x"9E",x"9E",x"9A",x"8A",x"78",x"6E",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"80",
		x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9C",x"8E",x"7C",x"70",x"68",x"64",x"64",x"66",x"68",x"6C",
		x"6E",x"74",x"7C",x"88",x"90",x"96",x"9A",x"9E",x"9E",x"9C",x"90",x"7E",x"72",x"68",x"66",x"64",
		x"66",x"68",x"6C",x"6E",x"72",x"7C",x"86",x"90",x"96",x"9A",x"9C",x"9E",x"9C",x"92",x"7E",x"72",
		x"68",x"64",x"64",x"64",x"68",x"6A",x"6E",x"74",x"7E",x"88",x"90",x"96",x"9A",x"9E",x"9E",x"9C",
		x"90",x"7C",x"70",x"6A",x"66",x"64",x"66",x"68",x"6C",x"6E",x"74",x"7E",x"8A",x"92",x"96",x"9C",
		x"9E",x"9E",x"9C",x"8E",x"7C",x"70",x"68",x"64",x"64",x"66",x"68",x"6C",x"70",x"76",x"80",x"8A",
		x"92",x"98",x"9C",x"9E",x"9E",x"9A",x"88",x"78",x"6E",x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",
		x"7A",x"86",x"8E",x"94",x"9A",x"9C",x"9E",x"9E",x"96",x"84",x"74",x"6A",x"66",x"64",x"64",x"66",
		x"68",x"6C",x"72",x"7C",x"88",x"90",x"96",x"9A",x"9E",x"9E",x"9C",x"90",x"7E",x"70",x"68",x"66",
		x"64",x"66",x"68",x"6C",x"70",x"78",x"82",x"8C",x"94",x"98",x"9C",x"9E",x"9E",x"9A",x"88",x"78",
		x"6C",x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",x"7C",x"86",x"90",x"96",x"9A",x"9E",x"9E",x"9C",
		x"90",x"7E",x"70",x"68",x"64",x"64",x"64",x"68",x"6C",x"6E",x"76",x"82",x"8A",x"94",x"98",x"9C",
		x"9E",x"9E",x"98",x"86",x"74",x"6A",x"66",x"62",x"64",x"66",x"6A",x"6C",x"72",x"7E",x"88",x"90",
		x"96",x"9C",x"9E",x"9E",x"9A",x"8C",x"7A",x"70",x"68",x"64",x"64",x"66",x"68",x"6C",x"72",x"7A",
		x"86",x"8E",x"94",x"9A",x"9E",x"9E",x"9C",x"92",x"7E",x"72",x"68",x"64",x"64",x"66",x"68",x"6C",
		x"6E",x"76",x"82",x"8C",x"94",x"98",x"9C",x"9E",x"9E",x"96",x"82",x"74",x"6C",x"66",x"64",x"66",
		x"68",x"6A",x"6E",x"72",x"7C",x"86",x"90",x"96",x"9A",x"9E",x"9E",x"9E",x"92",x"80",x"72",x"6A",
		x"66",x"64",x"66",x"68",x"6A",x"6E",x"72",x"7A",x"86",x"8E",x"96",x"9A",x"9E",x"A0",x"9E",x"94",
		x"82",x"74",x"6C",x"66",x"64",x"66",x"68",x"6A",x"6E",x"72",x"78",x"80",x"8A",x"94",x"98",x"9C",
		x"9E",x"A0",x"9C",x"8C",x"7A",x"6E",x"68",x"64",x"64",x"64",x"68",x"6C",x"6E",x"72",x"7A",x"82",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"9C",x"8C",x"7A",x"6E",x"68",x"64",x"64",x"66",x"68",x"6C",
		x"70",x"74",x"78",x"80",x"8A",x"92",x"9A",x"9C",x"9E",x"9E",x"9C",x"92",x"7E",x"72",x"68",x"64",
		x"64",x"66",x"68",x"6A",x"6E",x"70",x"74",x"7A",x"84",x"8E",x"94",x"9A",x"9E",x"9E",x"9E",x"9C",
		x"8C",x"7A",x"6E",x"68",x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"76",x"7A",x"84",x"8E",x"96",
		x"9A",x"9E",x"A0",x"9E",x"9C",x"8C",x"7C",x"6E",x"68",x"66",x"64",x"66",x"68",x"6A",x"6E",x"72",
		x"76",x"78",x"80",x"8A",x"92",x"9A",x"9C",x"A0",x"A0",x"A0",x"96",x"82",x"74",x"6A",x"66",x"64",
		x"64",x"66",x"68",x"6C",x"70",x"72",x"76",x"7C",x"84",x"8E",x"94",x"9A",x"9E",x"A0",x"A0",x"9E",
		x"92",x"80",x"72",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"76",x"7A",x"82",x"8E",
		x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"94",x"82",x"74",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",
		x"70",x"72",x"76",x"7A",x"7E",x"88",x"92",x"98",x"9E",x"A0",x"A0",x"A0",x"9C",x"8C",x"7A",x"6E",
		x"68",x"64",x"64",x"66",x"66",x"6A",x"6C",x"70",x"72",x"78",x"7A",x"80",x"88",x"92",x"9A",x"9C",
		x"A0",x"A0",x"A0",x"9C",x"8A",x"7A",x"6E",x"68",x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"74",
		x"78",x"7C",x"80",x"88",x"92",x"98",x"9C",x"A0",x"A0",x"A0",x"9E",x"90",x"7C",x"70",x"68",x"64",
		x"64",x"64",x"66",x"68",x"6C",x"6E",x"72",x"76",x"78",x"7E",x"84",x"8E",x"96",x"9A",x"9E",x"A0",
		x"A0",x"9E",x"96",x"84",x"74",x"6C",x"66",x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"74",x"78",
		x"7C",x"80",x"88",x"90",x"98",x"9C",x"9E",x"A0",x"A0",x"A0",x"94",x"80",x"72",x"6A",x"64",x"64",
		x"64",x"66",x"68",x"6C",x"6E",x"72",x"74",x"78",x"7C",x"7E",x"88",x"90",x"98",x"9C",x"9E",x"A0",
		x"A0",x"9E",x"94",x"82",x"72",x"6A",x"64",x"62",x"64",x"64",x"68",x"6A",x"6E",x"70",x"74",x"78",
		x"7A",x"7E",x"84",x"8E",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"9A",x"8A",x"78",x"6C",x"66",x"64",
		x"62",x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"7A",x"7C",x"80",x"88",x"90",x"98",x"9C",x"A0",
		x"A2",x"A0",x"A0",x"96",x"84",x"74",x"6A",x"64",x"62",x"64",x"64",x"68",x"6A",x"6E",x"70",x"74",
		x"78",x"7A",x"7E",x"82",x"8A",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"7E",x"70",x"68",
		x"62",x"62",x"64",x"64",x"68",x"6C",x"6E",x"72",x"76",x"7A",x"7C",x"80",x"84",x"8C",x"94",x"9A",
		x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"7E",x"72",x"6A",x"64",x"62",x"64",x"66",x"68",x"6A",x"6E",
		x"70",x"74",x"78",x"7A",x"7E",x"80",x"88",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"96",x"84",
		x"74",x"6A",x"64",x"62",x"62",x"64",x"66",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7C",x"7E",x"84",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A2",x"9E",x"8E",x"7C",x"70",x"68",x"64",x"62",x"64",x"64",
		x"68",x"6A",x"6E",x"72",x"74",x"78",x"7A",x"7E",x"80",x"88",x"90",x"96",x"9C",x"A0",x"A2",x"A2",
		x"A2",x"98",x"86",x"76",x"6A",x"66",x"62",x"62",x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"78",
		x"7C",x"7E",x"82",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A2",x"A0",x"96",x"82",x"74",x"6A",x"64",
		x"62",x"62",x"64",x"68",x"6A",x"6E",x"70",x"74",x"76",x"78",x"7C",x"7E",x"82",x"8A",x"92",x"9A",
		x"9E",x"A0",x"A2",x"A0",x"9E",x"94",x"80",x"72",x"6A",x"64",x"62",x"64",x"64",x"68",x"6A",x"6E",
		x"70",x"74",x"76",x"7A",x"7C",x"7E",x"82",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A2",x"A0",x"96",
		x"82",x"74",x"6A",x"64",x"62",x"62",x"62",x"66",x"6A",x"6C",x"70",x"74",x"76",x"7A",x"7C",x"80",
		x"82",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A0",x"A0",x"9A",x"88",x"78",x"6C",x"66",x"62",x"62",
		x"64",x"66",x"6A",x"6C",x"70",x"72",x"76",x"78",x"7C",x"7E",x"80",x"84",x"8C",x"94",x"9A",x"9E",
		x"A0",x"A2",x"A0",x"9C",x"8E",x"7C",x"70",x"66",x"62",x"62",x"62",x"64",x"66",x"6A",x"6E",x"70",
		x"74",x"76",x"7A",x"7C",x"80",x"82",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A2",x"A0",x"98",x"86",
		x"76",x"6A",x"64",x"62",x"62",x"64",x"66",x"6A",x"6C",x"6E",x"72",x"74",x"78",x"7C",x"7E",x"80",
		x"84",x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"80",x"72",x"68",x"64",x"62",x"62",
		x"64",x"66",x"6A",x"6E",x"70",x"74",x"76",x"78",x"7C",x"7E",x"80",x"86",x"8E",x"96",x"9A",x"9E",
		x"A0",x"A2",x"A2",x"9C",x"8C",x"7C",x"6E",x"66",x"64",x"62",x"64",x"64",x"68",x"6A",x"6E",x"70",
		x"74",x"78",x"7A",x"7E",x"80",x"82",x"88",x"92",x"98",x"9C",x"A0",x"A2",x"A0",x"A0",x"9A",x"88",
		x"78",x"6C",x"64",x"62",x"60",x"62",x"64",x"68",x"6A",x"6E",x"72",x"76",x"78",x"7C",x"80",x"82",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",x"80",x"70",x"68",x"62",x"62",x"62",x"64",
		x"66",x"6A",x"6E",x"72",x"74",x"78",x"7C",x"7E",x"84",x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",
		x"9E",x"90",x"7C",x"70",x"68",x"64",x"62",x"62",x"66",x"68",x"6C",x"6E",x"72",x"74",x"78",x"7C",
		x"80",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A0",x"9E",x"90",x"7E",x"70",x"68",x"64",x"62",x"62",
		x"64",x"68",x"6A",x"6E",x"72",x"74",x"78",x"7C",x"82",x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",
		x"9A",x"88",x"78",x"6C",x"66",x"64",x"62",x"66",x"68",x"6A",x"6E",x"70",x"74",x"78",x"7A",x"82",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"9A",x"86",x"76",x"6C",x"66",x"62",x"62",x"64",x"66",
		x"6A",x"6E",x"70",x"74",x"78",x"7E",x"86",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"92",x"7E",
		x"70",x"68",x"64",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"76",x"7C",x"86",x"8E",x"96",x"9C",
		x"9E",x"A0",x"A0",x"9E",x"92",x"80",x"72",x"6A",x"64",x"62",x"64",x"66",x"68",x"6C",x"70",x"74",
		x"76",x"7C",x"86",x"90",x"96",x"9C",x"A0",x"A0",x"A0",x"9E",x"90",x"7C",x"70",x"68",x"64",x"64",
		x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"80",x"8C",x"94",x"9A",x"9C",x"A0",x"A0",x"A0",x"96",
		x"84",x"74",x"6C",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"78",x"7E",x"8A",x"92",x"98",
		x"9C",x"A0",x"A0",x"A0",x"98",x"88",x"76",x"6C",x"66",x"64",x"64",x"66",x"68",x"6C",x"6E",x"72",
		x"76",x"80",x"8A",x"92",x"98",x"9C",x"9E",x"A0",x"9E",x"96",x"84",x"76",x"6A",x"64",x"62",x"62",
		x"66",x"68",x"6C",x"70",x"72",x"78",x"82",x"8C",x"94",x"98",x"9C",x"9E",x"9E",x"9E",x"92",x"80",
		x"72",x"68",x"64",x"64",x"64",x"66",x"6A",x"6E",x"70",x"74",x"7C",x"86",x"90",x"96",x"9A",x"9E",
		x"9E",x"A0",x"98",x"86",x"76",x"6C",x"66",x"64",x"64",x"66",x"6A",x"6C",x"70",x"74",x"7A",x"84",
		x"8E",x"94",x"9A",x"9E",x"9E",x"9E",x"9A",x"8A",x"7A",x"6E",x"66",x"64",x"64",x"66",x"68",x"6C",
		x"6E",x"72",x"78",x"82",x"8C",x"94",x"9A",x"9C",x"A0",x"A0",x"9C",x"8A",x"7A",x"6E",x"66",x"64",
		x"64",x"66",x"68",x"6C",x"6E",x"74",x"7A",x"86",x"8E",x"96",x"9A",x"9E",x"A0",x"A0",x"9A",x"88",
		x"78",x"6C",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"7C",x"88",x"90",x"98",x"9C",x"9E",
		x"A0",x"9E",x"94",x"82",x"74",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"76",x"82",x"8C",
		x"94",x"9A",x"9E",x"A0",x"A0",x"9A",x"8A",x"7A",x"6E",x"68",x"64",x"64",x"66",x"68",x"6C",x"70",
		x"74",x"7E",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9C",x"92",x"7E",x"70",x"68",x"64",x"64",x"64",
		x"68",x"6A",x"6E",x"72",x"7A",x"86",x"8E",x"96",x"9A",x"9E",x"A0",x"9E",x"96",x"84",x"74",x"6A",
		x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",x"7A",x"84",x"8C",x"94",x"9A",x"9C",x"9E",x"9E",x"98",
		x"86",x"76",x"6C",x"66",x"64",x"64",x"66",x"6A",x"6C",x"70",x"78",x"82",x"8C",x"94",x"9A",x"9C",
		x"9E",x"9E",x"98",x"86",x"76",x"6C",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"78",x"84",x"8E",
		x"96",x"9A",x"9E",x"9E",x"9E",x"96",x"84",x"74",x"6A",x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",
		x"7C",x"86",x"8E",x"96",x"9A",x"9E",x"9E",x"9E",x"94",x"80",x"72",x"6A",x"64",x"64",x"64",x"68",
		x"6A",x"6E",x"74",x"7E",x"88",x"90",x"96",x"9A",x"9E",x"9E",x"9C",x"8E",x"7C",x"6E",x"68",x"64",
		x"64",x"66",x"68",x"6C",x"70",x"76",x"82",x"8C",x"94",x"98",x"9C",x"9E",x"9E",x"98",x"88",x"76",
		x"6C",x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",x"7C",x"86",x"90",x"96",x"9A",x"9E",x"9E",x"9C",
		x"90",x"7E",x"70",x"68",x"64",x"62",x"64",x"68",x"6C",x"70",x"78",x"82",x"8C",x"94",x"9A",x"9E",
		x"9E",x"9E",x"98",x"88",x"78",x"6C",x"66",x"64",x"64",x"66",x"6A",x"6E",x"72",x"7C",x"86",x"90",
		x"96",x"9A",x"9E",x"9E",x"9E",x"90",x"7C",x"70",x"68",x"64",x"64",x"64",x"68",x"6A",x"70",x"78",
		x"84",x"8C",x"94",x"9A",x"9C",x"9E",x"9E",x"96",x"84",x"74",x"6A",x"66",x"64",x"64",x"68",x"6A",
		x"6E",x"74",x"7E",x"8A",x"90",x"98",x"9C",x"9E",x"9E",x"9A",x"8A",x"7A",x"6E",x"66",x"64",x"64",
		x"66",x"68",x"6C",x"70",x"7C",x"86",x"90",x"96",x"9A",x"9E",x"9E",x"9C",x"90",x"7C",x"70",x"68",
		x"64",x"64",x"66",x"68",x"6C",x"70",x"78",x"84",x"8C",x"94",x"9A",x"9C",x"9E",x"9E",x"92",x"80",
		x"72",x"6A",x"64",x"64",x"64",x"68",x"6A",x"6E",x"76",x"82",x"8C",x"94",x"98",x"9C",x"9E",x"9E",
		x"96",x"82",x"74",x"6A",x"64",x"64",x"64",x"68",x"6A",x"6E",x"76",x"80",x"8A",x"92",x"98",x"9C",
		x"9E",x"9E",x"98",x"84",x"76",x"6C",x"66",x"64",x"64",x"66",x"6A",x"6E",x"76",x"80",x"8A",x"92",
		x"98",x"9C",x"9E",x"9E",x"98",x"86",x"76",x"6C",x"66",x"64",x"66",x"68",x"6A",x"6E",x"76",x"80",
		x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"98",x"86",x"76",x"6A",x"66",x"64",x"64",x"68",x"6A",x"6E",
		x"74",x"80",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"98",x"86",x"76",x"6C",x"66",x"64",x"66",x"68",
		x"6C",x"6E",x"74",x"7C",x"88",x"90",x"96",x"9C",x"9E",x"9E",x"9C",x"90",x"7C",x"70",x"68",x"64",
		x"64",x"66",x"68",x"6C",x"70",x"74",x"7E",x"8A",x"92",x"98",x"9C",x"9E",x"A0",x"9C",x"8A",x"7A",
		x"6E",x"68",x"66",x"64",x"66",x"68",x"6C",x"70",x"74",x"7E",x"88",x"90",x"98",x"9C",x"9E",x"A0",
		x"9E",x"90",x"7E",x"72",x"68",x"66",x"64",x"66",x"68",x"6A",x"6E",x"72",x"78",x"80",x"8A",x"94",
		x"98",x"9C",x"9E",x"9E",x"9C",x"8E",x"7C",x"70",x"68",x"64",x"64",x"66",x"68",x"6C",x"6E",x"72",
		x"78",x"80",x"8A",x"94",x"98",x"9E",x"A0",x"A0",x"9E",x"90",x"7E",x"70",x"68",x"64",x"64",x"64",
		x"68",x"6A",x"6E",x"72",x"74",x"7C",x"86",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9A",x"86",x"76",
		x"6C",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"72",x"78",x"7E",x"88",x"92",x"98",x"9C",x"A0",
		x"A0",x"A0",x"96",x"84",x"74",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"78",x"7E",
		x"88",x"90",x"98",x"9C",x"A0",x"A0",x"A0",x"9A",x"88",x"76",x"6C",x"66",x"62",x"62",x"64",x"68",
		x"6C",x"70",x"72",x"76",x"7A",x"82",x"8C",x"94",x"9A",x"A0",x"A0",x"A0",x"A0",x"96",x"84",x"74",
		x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"6E",x"72",x"76",x"7A",x"82",x"8C",x"94",x"9A",x"9E",
		x"A0",x"A0",x"A0",x"96",x"82",x"74",x"6A",x"64",x"64",x"64",x"66",x"68",x"6C",x"70",x"72",x"76",
		x"7A",x"7E",x"88",x"90",x"98",x"9C",x"A0",x"A2",x"A2",x"9C",x"8C",x"7A",x"6E",x"66",x"64",x"62",
		x"64",x"68",x"6A",x"6E",x"70",x"74",x"78",x"7C",x"82",x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",
		x"98",x"84",x"76",x"6C",x"66",x"64",x"62",x"64",x"68",x"6A",x"6E",x"72",x"74",x"78",x"7C",x"82",
		x"8C",x"94",x"9A",x"9E",x"A0",x"A0",x"A0",x"9A",x"8A",x"78",x"6C",x"66",x"64",x"62",x"64",x"66",
		x"6A",x"6C",x"70",x"74",x"76",x"7A",x"80",x"88",x"90",x"98",x"9E",x"A0",x"A2",x"A0",x"9E",x"90",
		x"7E",x"70",x"68",x"64",x"62",x"64",x"66",x"6A",x"6C",x"6E",x"72",x"76",x"78",x"7C",x"82",x"8A",
		x"94",x"9A",x"9E",x"A0",x"A2",x"A2",x"9C",x"8C",x"7A",x"6E",x"66",x"64",x"64",x"64",x"66",x"6A",
		x"6C",x"70",x"74",x"76",x"7A",x"7C",x"82",x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9C",x"8A",
		x"78",x"6C",x"66",x"64",x"62",x"64",x"66",x"6A",x"6C",x"70",x"74",x"76",x"7A",x"7E",x"82",x"8A",
		x"92",x"9A",x"9E",x"A2",x"A2",x"A2",x"9E",x"90",x"7E",x"70",x"68",x"64",x"62",x"64",x"64",x"68",
		x"6A",x"6E",x"72",x"76",x"7A",x"7C",x"7E",x"86",x"8E",x"96",x"9C",x"9E",x"A2",x"A2",x"A0",x"98",
		x"86",x"76",x"6C",x"66",x"62",x"62",x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"7A",x"7E",x"80",
		x"88",x"92",x"98",x"9E",x"A0",x"A2",x"A2",x"A0",x"94",x"80",x"72",x"68",x"64",x"62",x"62",x"64",
		x"68",x"6A",x"6E",x"70",x"74",x"78",x"7A",x"7E",x"82",x"8A",x"92",x"98",x"9E",x"A0",x"A2",x"A2",
		x"9E",x"92",x"80",x"72",x"68",x"64",x"62",x"62",x"64",x"68",x"6A",x"6E",x"70",x"74",x"78",x"7A",
		x"7E",x"80",x"88",x"90",x"98",x"9E",x"A0",x"A2",x"A2",x"A0",x"96",x"84",x"74",x"6A",x"64",x"62",
		x"62",x"64",x"68",x"6A",x"6C",x"70",x"74",x"76",x"7A",x"7C",x"80",x"86",x"8E",x"96",x"9C",x"9E",
		x"A2",x"A2",x"A0",x"9A",x"88",x"78",x"6C",x"66",x"62",x"62",x"64",x"66",x"6A",x"6C",x"70",x"72",
		x"76",x"7A",x"7C",x"7E",x"82",x"8A",x"94",x"9A",x"9E",x"A0",x"A2",x"A2",x"9E",x"92",x"7E",x"70",
		x"66",x"62",x"60",x"62",x"64",x"66",x"6A",x"6E",x"72",x"74",x"78",x"7C",x"7E",x"80",x"86",x"8E",
		x"96",x"9C",x"A0",x"A2",x"A2",x"A0",x"9C",x"8C",x"7C",x"70",x"68",x"64",x"64",x"64",x"66",x"68",
		x"6C",x"6E",x"70",x"74",x"78",x"7A",x"7E",x"80",x"86",x"8E",x"96",x"9C",x"A0",x"A2",x"A2",x"A0",
		x"9C",x"8A",x"78",x"6C",x"66",x"62",x"62",x"64",x"66",x"68",x"6C",x"6E",x"72",x"76",x"78",x"7C",
		x"7E",x"80",x"86",x"90",x"96",x"9C",x"A0",x"A2",x"A2",x"A0",x"9A",x"8A",x"78",x"6C",x"66",x"64",
		x"62",x"64",x"66",x"68",x"6C",x"6E",x"72",x"74",x"78",x"7A",x"7E",x"80",x"84",x"8E",x"94",x"9A",
		x"A0",x"A2",x"A2",x"A2",x"9C",x"8C",x"7A",x"6E",x"66",x"62",x"62",x"62",x"64",x"68",x"6A",x"6E",
		x"70",x"74",x"76",x"7A",x"7E",x"80",x"84",x"8C",x"94",x"9A",x"9E",x"A0",x"A2",x"A0",x"9E",x"92",
		x"80",x"72",x"68",x"64",x"62",x"62",x"64",x"66",x"6A",x"6E",x"70",x"74",x"76",x"7A",x"7C",x"7E",
		x"82",x"88",x"90",x"98",x"9C",x"A0",x"A2",x"A2",x"A0",x"9A",x"88",x"76",x"6C",x"64",x"62",x"62",
		x"64",x"66",x"68",x"6C",x"6E",x"72",x"76",x"78",x"7C",x"7E",x"80",x"84",x"8C",x"94",x"9A",x"9E",
		x"A0",x"A2",x"A0",x"9E",x"90",x"7E",x"70",x"68",x"62",x"62",x"64",x"64",x"68",x"6C",x"6E",x"72",
		x"74",x"76",x"7A",x"7C",x"80",x"82",x"86",x"8E",x"96",x"9C",x"A0",x"A2",x"A2",x"A0",x"9C",x"8C",
		x"7A",x"6E",x"66",x"64",x"62",x"64",x"66",x"68",x"6C",x"6E",x"72",x"74",x"76",x"7A",x"7C",x"7E",
		x"82",x"88",x"90",x"98",x"9C",x"A0",x"A2",x"A0",x"A0",x"98",x"88",x"78",x"6C",x"66",x"62",x"62",
		x"64",x"66",x"68",x"6C",x"6E",x"72",x"76",x"78",x"7A",x"7E",x"82",x"88",x"92",x"98",x"9C",x"A0",
		x"A2",x"A0",x"9E",x"96",x"84",x"74",x"6A",x"64",x"62",x"62",x"64",x"66",x"68",x"6C",x"70",x"72",
		x"76",x"7A",x"7C",x"80",x"88",x"90",x"98",x"9C",x"A0",x"A2",x"A0",x"9E",x"96",x"84",x"74",x"6A",
		x"64",x"62",x"62",x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"7A",x"7E",x"84",x"8C",x"94",x"9A",
		x"9E",x"A0",x"A0",x"9E",x"9A",x"88",x"78",x"6C",x"66",x"64",x"64",x"64",x"66",x"6A",x"6C",x"70",
		x"72",x"76",x"7A",x"7E",x"86",x"90",x"96",x"9C",x"9E",x"A0",x"A0",x"9E",x"96",x"84",x"74",x"6C",
		x"66",x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"74",x"78",x"7C",x"82",x"8C",x"94",x"9A",x"9E",
		x"A0",x"A0",x"A0",x"98",x"86",x"76",x"6C",x"66",x"62",x"62",x"64",x"68",x"6A",x"6E",x"72",x"76",
		x"78",x"7E",x"86",x"90",x"98",x"9C",x"A0",x"A0",x"A0",x"9C",x"92",x"80",x"72",x"6A",x"66",x"64",
		x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"7A",x"82",x"8C",x"94",x"9A",x"9E",x"A0",x"9E",x"9C",
		x"94",x"82",x"74",x"6A",x"66",x"64",x"64",x"66",x"68",x"6C",x"70",x"74",x"76",x"7C",x"84",x"8E",
		x"96",x"9C",x"9E",x"A0",x"9E",x"9C",x"90",x"7E",x"72",x"68",x"66",x"64",x"64",x"68",x"6A",x"6E",
		x"70",x"74",x"78",x"7E",x"88",x"92",x"98",x"9C",x"9E",x"A0",x"9E",x"98",x"88",x"78",x"6C",x"66",
		x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"76",x"7C",x"86",x"90",x"96",x"9A",x"9E",x"9E",x"9C",
		x"98",x"8A",x"7A",x"6E",x"68",x"64",x"64",x"66",x"68",x"6A",x"6E",x"72",x"76",x"7C",x"86",x"90",
		x"96",x"9C",x"9E",x"9E",x"9E",x"98",x"88",x"78",x"6E",x"68",x"64",x"64",x"66",x"6A",x"6C",x"70",
		x"74",x"78",x"80",x"8A",x"92",x"98",x"9C",x"9E",x"9E",x"9C",x"92",x"80",x"74",x"6C",x"66",x"66",
		x"66",x"68",x"6A",x"6E",x"72",x"74",x"7A",x"86",x"8E",x"94",x"9A",x"9C",x"9C",x"9A",x"96",x"88",
		x"78",x"6E",x"68",x"66",x"66",x"68",x"6A",x"6C",x"70",x"74",x"78",x"82",x"8C",x"94",x"9A",x"9C",
		x"9E",x"9C",x"98",x"8C",x"7A",x"70",x"6A",x"66",x"64",x"66",x"6A",x"6C",x"70",x"74",x"78",x"82",
		x"8C",x"94",x"9A",x"9C",x"9E",x"9C",x"98",x"8A",x"7C",x"70",x"6A",x"66",x"66",x"66",x"68",x"6C",
		x"70",x"74",x"7A",x"84",x"8C",x"94",x"9A",x"9C",x"9E",x"9C",x"96",x"88",x"78",x"6E",x"68",x"66",
		x"66",x"68",x"6A",x"6E",x"70",x"74",x"7C",x"86",x"90",x"96",x"9A",x"9C",x"9C",x"9A",x"92",x"82",
		x"74",x"6C",x"68",x"66",x"66",x"68",x"6C",x"6E",x"72",x"78",x"82",x"8C",x"94",x"98",x"9C",x"9C",
		x"9C",x"96",x"8A",x"7A",x"70",x"6A",x"66",x"66",x"68",x"6A",x"6E",x"70",x"74",x"7C",x"88",x"90",
		x"96",x"9A",x"9C",x"9C",x"98",x"90",x"7E",x"72",x"6A",x"66",x"66",x"66",x"6A",x"6C",x"70",x"74",
		x"7A",x"84",x"8E",x"94",x"98",x"9C",x"9C",x"9A",x"92",x"84",x"76",x"6C",x"68",x"66",x"66",x"68",
		x"6C",x"6E",x"72",x"78",x"82",x"8C",x"94",x"98",x"9A",x"9C",x"9A",x"94",x"86",x"78",x"6E",x"68",
		x"68",x"68",x"6A",x"6C",x"6E",x"72",x"78",x"82",x"8C",x"94",x"98",x"9A",x"9A",x"9A",x"94",x"86",
		x"78",x"6E",x"68",x"66",x"66",x"68",x"6C",x"6E",x"72",x"7A",x"84",x"8C",x"94",x"98",x"9A",x"9A",
		x"98",x"92",x"82",x"76",x"6C",x"68",x"68",x"68",x"6A",x"6E",x"70",x"74",x"7C",x"86",x"8E",x"96",
		x"9A",x"9C",x"9A",x"98",x"90",x"80",x"74",x"6C",x"68",x"66",x"66",x"6A",x"6C",x"70",x"74",x"7E",
		x"88",x"90",x"96",x"9A",x"9A",x"98",x"96",x"8C",x"7C",x"72",x"6A",x"68",x"68",x"68",x"6A",x"6E",
		x"70",x"76",x"80",x"8A",x"92",x"98",x"9A",x"9A",x"98",x"94",x"88",x"78",x"70",x"6A",x"68",x"68",
		x"68",x"6C",x"70",x"72",x"7A",x"84",x"8E",x"94",x"98",x"9A",x"9A",x"96",x"90",x"82",x"74",x"6E",
		x"68",x"68",x"68",x"6A",x"6C",x"70",x"74",x"7E",x"88",x"90",x"96",x"9A",x"9A",x"98",x"94",x"8A",
		x"7A",x"70",x"6A",x"68",x"66",x"6A",x"6C",x"6E",x"72",x"7A",x"84",x"8C",x"94",x"98",x"9A",x"98",
		x"96",x"8E",x"80",x"74",x"6C",x"68",x"68",x"68",x"6A",x"6E",x"70",x"76",x"80",x"8A",x"92",x"96",
		x"9A",x"9A",x"98",x"92",x"84",x"76",x"6E",x"68",x"68",x"68",x"6A",x"6C",x"70",x"74",x"7E",x"88",
		x"90",x"96",x"98",x"9A",x"98",x"94",x"8A",x"7A",x"70",x"6A",x"68",x"68",x"68",x"6C",x"6E",x"72",
		x"7A",x"86",x"8E",x"94",x"98",x"9A",x"98",x"96",x"8C",x"7E",x"72",x"6C",x"68",x"68",x"6A",x"6C",
		x"6E",x"70",x"78",x"84",x"8C",x"92",x"96",x"98",x"98",x"96",x"90",x"80",x"74",x"6E",x"6A",x"68",
		x"6A",x"6C",x"6E",x"72",x"78",x"82",x"8C",x"92",x"96",x"98",x"98",x"96",x"90",x"82",x"76",x"6E",
		x"6A",x"68",x"6A",x"6C",x"6E",x"70",x"76",x"80",x"8A",x"92",x"96",x"98",x"98",x"96",x"90",x"82",
		x"76",x"6E",x"6A",x"68",x"6A",x"6C",x"6E",x"72",x"78",x"82",x"8C",x"92",x"96",x"98",x"98",x"96",
		x"90",x"80",x"76",x"6E",x"6A",x"6A",x"6A",x"6C",x"6E",x"72",x"78",x"82",x"8A",x"92",x"96",x"98",
		x"98",x"96",x"90",x"82",x"76",x"6E",x"6A",x"6A",x"6A",x"6C",x"6E",x"72",x"76",x"82",x"8C",x"92",
		x"96",x"98",x"96",x"94",x"8C",x"7E",x"74",x"6C",x"6A",x"6A",x"6A",x"6C",x"6E",x"72",x"78",x"80",
		x"8A",x"92",x"96",x"98",x"98",x"96",x"90",x"84",x"76",x"6E",x"6A",x"6A",x"6A",x"6C",x"6E",x"70",
		x"74",x"7A",x"84",x"8C",x"94",x"98",x"9A",x"98",x"96",x"90",x"82",x"76",x"6E",x"6A",x"6A",x"6A",
		x"6C",x"6E",x"72",x"74",x"78",x"82",x"8C",x"92",x"96",x"98",x"98",x"96",x"90",x"84",x"78",x"70",
		x"6C",x"6A",x"6A",x"6C",x"6E",x"70",x"74",x"76",x"7E",x"88",x"90",x"94",x"98",x"98",x"96",x"94",
		x"8C",x"7E",x"74",x"6C",x"6A",x"68",x"6A",x"6C",x"6E",x"70",x"74",x"78",x"7E",x"88",x"92",x"98",
		x"9A",x"9A",x"98",x"96",x"8C",x"80",x"74",x"6E",x"6C",x"6A",x"6A",x"6C",x"6E",x"72",x"74",x"78",
		x"7C",x"86",x"8E",x"94",x"98",x"9A",x"98",x"96",x"90",x"84",x"78",x"70",x"6C",x"6A",x"6A",x"6A",
		x"6C",x"6E",x"72",x"74",x"78",x"7C",x"86",x"8E",x"96",x"98",x"9A",x"98",x"96",x"90",x"84",x"76",
		x"70",x"6A",x"6A",x"6A",x"6C",x"6E",x"70",x"72",x"76",x"78",x"7C",x"86",x"8E",x"94",x"98",x"9A",
		x"98",x"96",x"90",x"86",x"7A",x"72",x"6C",x"6A",x"6A",x"6C",x"6E",x"70",x"72",x"74",x"78",x"7A",
		x"80",x"8A",x"90",x"96",x"9A",x"9A",x"98",x"94",x"8E",x"82",x"76",x"70",x"6C",x"6A",x"6A",x"6C",
		x"6E",x"70",x"72",x"76",x"78",x"7A",x"80",x"8A",x"92",x"96",x"9A",x"98",x"98",x"94",x"8E",x"80",
		x"76",x"6E",x"6A",x"6A",x"6A",x"6C",x"6E",x"70",x"72",x"76",x"78",x"7A",x"7E",x"88",x"90",x"96",
		x"98",x"9A",x"98",x"96",x"90",x"86",x"7A",x"70",x"6C",x"6A",x"68",x"6A",x"6C",x"6E",x"72",x"74",
		x"78",x"7A",x"7C",x"82",x"8C",x"92",x"96",x"9A",x"9A",x"96",x"94",x"8E",x"82",x"76",x"70",x"6C",
		x"6A",x"6A",x"6C",x"6E",x"70",x"72",x"74",x"76",x"7A",x"7C",x"80",x"8A",x"92",x"96",x"98",x"98",
		x"98",x"94",x"90",x"84",x"78",x"72",x"6C",x"6C",x"6A",x"6C",x"6E",x"70",x"72",x"76",x"78",x"7A",
		x"7C",x"80",x"88",x"90",x"96",x"98",x"98",x"98",x"96",x"92",x"88",x"7C",x"72",x"6E",x"6C",x"6A",
		x"6C",x"6C",x"6E",x"72",x"74",x"76",x"78",x"7C",x"7E",x"82",x"8A",x"92",x"96",x"98",x"98",x"96",
		x"94",x"8E",x"84",x"78",x"72",x"6C",x"6C",x"6A",x"6C",x"6E",x"70",x"72",x"74",x"76",x"7A",x"7C",
		x"7E",x"82",x"8C",x"92",x"96",x"9A",x"98",x"96",x"94",x"8E",x"84",x"78",x"70",x"6C",x"6A",x"6A",
		x"6C",x"6E",x"70",x"72",x"74",x"76",x"7A",x"7C",x"7E",x"82",x"8A",x"92",x"96",x"98",x"98",x"96",
		x"94",x"90",x"86",x"7A",x"72",x"6E",x"6C",x"6A",x"6C",x"6C",x"6E",x"72",x"74",x"76",x"78",x"7C",
		x"7E",x"80",x"86",x"8E",x"94",x"98",x"98",x"98",x"94",x"92",x"8A",x"7E",x"74",x"6E",x"6C",x"6A",
		x"6C",x"6C",x"6E",x"70",x"72",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"88",x"90",x"94",x"98",x"98",
		x"96",x"94",x"90",x"88",x"7C",x"74",x"6E",x"6C",x"6C",x"6C",x"6E",x"70",x"72",x"74",x"76",x"78",
		x"7A",x"7C",x"7E",x"82",x"8A",x"90",x"96",x"98",x"98",x"96",x"92",x"8E",x"86",x"7A",x"72",x"6E",
		x"6A",x"6A",x"6C",x"6C",x"6E",x"72",x"74",x"76",x"7A",x"7C",x"7E",x"80",x"82",x"88",x"90",x"94",
		x"98",x"98",x"96",x"94",x"90",x"88",x"7E",x"74",x"70",x"6E",x"6C",x"6C",x"6E",x"70",x"72",x"74",
		x"76",x"78",x"7A",x"7C",x"7E",x"80",x"84",x"8C",x"92",x"96",x"96",x"96",x"94",x"90",x"8C",x"82",
		x"78",x"70",x"6E",x"6C",x"6C",x"6E",x"6E",x"70",x"72",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"80",
		x"88",x"90",x"94",x"96",x"96",x"96",x"94",x"90",x"88",x"7E",x"74",x"70",x"6C",x"6C",x"6C",x"6E",
		x"70",x"72",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"84",x"8A",x"90",x"96",x"96",x"96",x"94",
		x"92",x"8E",x"84",x"7A",x"74",x"70",x"6E",x"6C",x"6C",x"6E",x"70",x"72",x"74",x"76",x"78",x"7A",
		x"7C",x"7E",x"80",x"84",x"8C",x"92",x"96",x"96",x"94",x"94",x"90",x"8C",x"82",x"78",x"72",x"6E",
		x"6E",x"6C",x"6E",x"70",x"70",x"72",x"74",x"78",x"78",x"7C",x"7C",x"7E",x"80",x"84",x"8C",x"92",
		x"96",x"96",x"96",x"94",x"90",x"8C",x"82",x"78",x"72",x"6E",x"6E",x"6E",x"6E",x"70",x"70",x"72",
		x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"84",x"8A",x"92",x"94",x"96",x"96",x"94",x"90",x"8C",
		x"84",x"7A",x"72",x"6E",x"6C",x"6C",x"6E",x"6E",x"70",x"72",x"74",x"78",x"7A",x"7C",x"7E",x"7E",
		x"80",x"84",x"8A",x"90",x"94",x"96",x"96",x"94",x"90",x"8E",x"86",x"7C",x"76",x"70",x"6E",x"6E",
		x"6E",x"70",x"72",x"72",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"86",x"8E",x"92",x"94",
		x"94",x"94",x"90",x"8E",x"8A",x"80",x"78",x"72",x"70",x"6E",x"6E",x"70",x"70",x"72",x"74",x"76",
		x"78",x"7A",x"7C",x"7E",x"80",x"80",x"82",x"88",x"8E",x"92",x"94",x"94",x"92",x"90",x"8C",x"86",
		x"7C",x"76",x"72",x"6E",x"6E",x"6E",x"70",x"72",x"72",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",
		x"80",x"84",x"8C",x"90",x"94",x"94",x"94",x"92",x"8E",x"8A",x"82",x"7A",x"74",x"70",x"6E",x"6E",
		x"6E",x"70",x"72",x"74",x"76",x"78",x"7A",x"7C",x"7C",x"7E",x"80",x"82",x"86",x"8C",x"92",x"94",
		x"94",x"92",x"90",x"8E",x"88",x"80",x"78",x"72",x"70",x"6E",x"6E",x"70",x"70",x"72",x"74",x"76",
		x"78",x"7A",x"7C",x"7E",x"7E",x"80",x"86",x"8C",x"90",x"94",x"92",x"92",x"90",x"8C",x"88",x"7E",
		x"78",x"72",x"70",x"70",x"6E",x"70",x"72",x"72",x"74",x"78",x"78",x"7A",x"7C",x"7E",x"80",x"86",
		x"8C",x"90",x"92",x"92",x"92",x"8E",x"8C",x"86",x"7E",x"76",x"72",x"6E",x"6E",x"70",x"70",x"72",
		x"74",x"76",x"78",x"7A",x"7C",x"7E",x"80",x"82",x"8A",x"90",x"92",x"92",x"92",x"90",x"8C",x"8A",
		x"82",x"7A",x"74",x"72",x"70",x"70",x"70",x"72",x"74",x"76",x"78",x"7A",x"7A",x"7C",x"7E",x"84",
		x"8A",x"90",x"92",x"92",x"90",x"8E",x"8C",x"88",x"80",x"78",x"74",x"72",x"70",x"70",x"72",x"72",
		x"74",x"76",x"78",x"7A",x"7A",x"7E",x"82",x"88",x"8E",x"90",x"92",x"90",x"8E",x"8C",x"88",x"82",
		x"7A",x"74",x"72",x"70",x"70",x"72",x"72",x"74",x"76",x"78",x"7A",x"7C",x"7E",x"82",x"8A",x"8E",
		x"90",x"90",x"90",x"8E",x"8A",x"86",x"7E",x"78",x"74",x"72",x"70",x"72",x"72",x"74",x"76",x"78",
		x"7A",x"7C",x"7C",x"80",x"88",x"8C",x"90",x"90",x"8E",x"8E",x"8C",x"88",x"80",x"7A",x"74",x"72",
		x"70",x"70",x"72",x"74",x"76",x"76",x"78",x"7A",x"7C",x"82",x"88",x"8C",x"90",x"90",x"8E",x"8C",
		x"8A",x"86",x"80",x"78",x"74",x"72",x"70",x"72",x"72",x"74",x"74",x"76",x"7A",x"7A",x"7E",x"84",
		x"8A",x"8E",x"90",x"90",x"8E",x"8C",x"88",x"82",x"7C",x"76",x"74",x"72",x"72",x"72",x"74",x"76",
		x"76",x"78",x"7A",x"7C",x"82",x"88",x"8E",x"8E",x"8E",x"8E",x"8C",x"8A",x"84",x"7C",x"76",x"72",
		x"72",x"72",x"72",x"74",x"76",x"78",x"7A",x"7A",x"7C",x"84",x"88",x"8C",x"8E",x"8E",x"8E",x"8A",
		x"8A",x"84",x"7C",x"78",x"74",x"72",x"72",x"72",x"74",x"76",x"76",x"7A",x"7A",x"7E",x"84",x"8A",
		x"8C",x"8E",x"8C",x"8C",x"8A",x"86",x"80",x"7A",x"76",x"74",x"72",x"74",x"74",x"76",x"76",x"78",
		x"7A",x"7C",x"80",x"88",x"8C",x"8E",x"8E",x"8C",x"8A",x"88",x"84",x"7C",x"78",x"74",x"74",x"72",
		x"74",x"74",x"76",x"78",x"7A",x"7C",x"80",x"86",x"8A",x"8C",x"8E",x"8C",x"8C",x"88",x"86",x"80",
		x"78",x"76",x"74",x"72",x"72",x"74",x"76",x"76",x"78",x"7A",x"7E",x"86",x"8A",x"8C",x"8C",x"8C",
		x"8A",x"88",x"86",x"80",x"7A",x"76",x"74",x"74",x"74",x"74",x"76",x"78",x"7A",x"7C",x"80",x"86",
		x"8A",x"8C",x"8C",x"8C",x"8A",x"88",x"84",x"7E",x"7A",x"76",x"74",x"74",x"74",x"74",x"76",x"78",
		x"7A",x"7A",x"80",x"86",x"8A",x"8C",x"8C",x"8C",x"8A",x"88",x"82",x"7C",x"78",x"74",x"74",x"74",
		x"74",x"76",x"76",x"78",x"7A",x"7E",x"84",x"88",x"8A",x"8C",x"8C",x"8A",x"88",x"86",x"80",x"7A",
		x"76",x"74",x"74",x"74",x"76",x"76",x"78",x"7A",x"7C",x"82",x"86",x"8A",x"8A",x"8A",x"8A",x"88",
		x"86",x"80",x"7A",x"76",x"76",x"74",x"74",x"76",x"76",x"78",x"78",x"7A",x"80",x"86",x"8A",x"8C",
		x"8C",x"8A",x"88",x"86",x"82",x"7C",x"78",x"76",x"74",x"74",x"76",x"76",x"78",x"78",x"7A",x"80",
		x"86",x"88",x"8A",x"8C",x"8A",x"8A",x"86",x"84",x"7E",x"78",x"76",x"74",x"74",x"76",x"76",x"78",
		x"7A",x"7A",x"7E",x"84",x"88",x"8A",x"8A",x"8A",x"8A",x"88",x"84",x"7E",x"78",x"76",x"74",x"76",
		x"76",x"76",x"78",x"7A",x"7C",x"80",x"86",x"88",x"8A",x"8A",x"8A",x"88",x"86",x"82",x"7C",x"78",
		x"76",x"76",x"74",x"76",x"78",x"78",x"7A",x"7C",x"82",x"86",x"88",x"8A",x"8A",x"88",x"88",x"84",
		x"82",x"7C",x"78",x"76",x"76",x"76",x"76",x"78",x"78",x"7A",x"7C",x"82",x"86",x"88",x"8A",x"8A",
		x"88",x"86",x"84",x"80",x"7A",x"78",x"76",x"76",x"76",x"76",x"78",x"7A",x"7A",x"7E",x"84",x"88",
		x"8A",x"88",x"88",x"88",x"86",x"82",x"7E",x"7A",x"76",x"76",x"76",x"76",x"78",x"78",x"7A",x"7C",
		x"82",x"86",x"88",x"8A",x"8A",x"88",x"86",x"84",x"80",x"7C",x"78",x"76",x"76",x"76",x"76",x"78",
		x"7A",x"7A",x"7E",x"84",x"86",x"88",x"8A",x"88",x"86",x"86",x"82",x"7E",x"7A",x"76",x"76",x"76",
		x"76",x"78",x"78",x"78",x"7C",x"82",x"86",x"88",x"8A",x"88",x"88",x"86",x"84",x"80",x"7C",x"78",
		x"76",x"76",x"78",x"78",x"78",x"7A",x"7C",x"80",x"84",x"88",x"88",x"88",x"88",x"86",x"84",x"82",
		x"7C",x"78",x"76",x"76",x"76",x"78",x"78",x"7A",x"7C",x"80",x"84",x"86",x"88",x"88",x"88",x"86",
		x"84",x"80",x"7C",x"7A",x"76",x"76",x"76",x"76",x"78",x"7A",x"7A",x"7E",x"84",x"86",x"88",x"88",
		x"88",x"86",x"84",x"82",x"7E",x"7A",x"78",x"76",x"76",x"78",x"78",x"7A",x"7A",x"7E",x"84",x"86",
		x"88",x"88",x"88",x"88",x"86",x"82",x"7E",x"7A",x"78",x"78",x"76",x"78",x"78",x"7A",x"7A",x"7E",
		x"82",x"86",x"88",x"88",x"88",x"86",x"86",x"82",x"7E",x"7C",x"78",x"78",x"78",x"76",x"78",x"7A",
		x"7A",x"7E",x"82",x"86",x"86",x"88",x"88",x"86",x"86",x"82",x"7E",x"7A",x"78",x"78",x"78",x"78",
		x"78",x"7A",x"7A",x"7C",x"82",x"84",x"86",x"88",x"86",x"86",x"84",x"82",x"7E",x"7A",x"78",x"78",
		x"78",x"78",x"78",x"78",x"7A",x"7E",x"82",x"86",x"88",x"88",x"88",x"86",x"86",x"82",x"7E",x"7C",
		x"7A",x"78",x"78",x"78",x"78",x"7A",x"7A",x"7E",x"82",x"84",x"86",x"86",x"86",x"86",x"84",x"82",
		x"7E",x"7A",x"78",x"76",x"76",x"76",x"78",x"78",x"7A",x"7C",x"82",x"86",x"88",x"88",x"88",x"88",
		x"86",x"84",x"80",x"7C",x"7A",x"78",x"78",x"78",x"7A",x"7A",x"7A",x"7C",x"7E",x"82",x"86",x"86",
		x"88",x"88",x"86",x"84",x"82",x"7E",x"7A",x"78",x"78",x"78",x"78",x"78",x"7A",x"7A",x"7C",x"7E",
		x"82",x"84",x"86",x"86",x"86",x"86",x"84",x"82",x"7E",x"7C",x"7A",x"78",x"78",x"78",x"7A",x"7A",
		x"7A",x"7C",x"7E",x"80",x"84",x"86",x"88",x"88",x"86",x"86",x"84",x"82",x"7E",x"7A",x"7A",x"78",
		x"78",x"78",x"7A",x"7A",x"7A",x"7C",x"7C",x"80",x"84",x"86",x"88",x"88",x"86",x"84",x"84",x"82",
		x"7E",x"7C",x"7A",x"78",x"78",x"78",x"7A",x"7A",x"7A",x"7C",x"7C",x"7E",x"82",x"84",x"86",x"86",
		x"86",x"86",x"84",x"82",x"80",x"7C",x"7A",x"7A",x"78",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7C",
		x"7E",x"82",x"84",x"86",x"88",x"86",x"86",x"86",x"84",x"80",x"7C",x"7A",x"78",x"78",x"78",x"7A",
		x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"82",x"84",x"86",x"86",x"86",x"86",x"84",x"82",x"80",x"7C",
		x"7A",x"7A",x"78",x"78",x"7A",x"7A",x"7A",x"7A",x"7C",x"7E",x"7E",x"80",x"82",x"86",x"86",x"86",
		x"86",x"86",x"84",x"82",x"7E",x"7C",x"7A",x"78",x"78",x"78",x"78",x"78",x"7A",x"7A",x"7C",x"7E",
		x"7E",x"80",x"84",x"86",x"88",x"88",x"88",x"86",x"84",x"82",x"80",x"7C",x"7A",x"7A",x"7A",x"7A",
		x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"82",x"84",x"86",x"86",x"86",x"84",x"84",x"82",
		x"80",x"7E",x"7A",x"78",x"78",x"78",x"7A",x"7A",x"7A",x"7C",x"7C",x"7E",x"7E",x"7E",x"80",x"84",
		x"86",x"86",x"86",x"86",x"84",x"84",x"82",x"80",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",
		x"7C",x"7C",x"7E",x"7E",x"7E",x"80",x"84",x"86",x"86",x"86",x"86",x"84",x"84",x"82",x"80",x"7C",
		x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"80",x"82",x"84",x"86",
		x"86",x"86",x"84",x"84",x"82",x"80",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"80",x"82",x"86",x"86",x"86",x"86",x"84",x"84",x"82",x"7E",x"7C",x"7A",
		x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"80",x"84",x"84",x"86",
		x"86",x"84",x"84",x"82",x"82",x"7E",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",
		x"7E",x"7E",x"7E",x"80",x"82",x"84",x"86",x"86",x"84",x"84",x"82",x"82",x"82",x"7E",x"7C",x"7A",
		x"7A",x"78",x"7A",x"7A",x"7A",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"82",x"84",x"84",
		x"84",x"84",x"84",x"82",x"82",x"80",x"7E",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",
		x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"84",x"84",x"84",x"84",x"82",x"82",x"82",x"7E",x"7C",
		x"7C",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"80",x"7E",x"7E",x"82",x"84",
		x"84",x"84",x"84",x"84",x"84",x"82",x"80",x"7E",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"82",x"84",x"84",x"84",x"84",x"84",x"84",x"82",x"80",
		x"7E",x"7C",x"7C",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"82",x"84",x"84",x"84",x"84",x"82",x"82",x"80",x"7E",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"80",x"82",x"84",x"84",x"84",x"84",x"84",
		x"82",x"82",x"80",x"7E",x"7C",x"7C",x"7C",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"80",x"80",x"82",x"84",x"84",x"84",x"84",x"82",x"82",x"80",x"7E",x"7C",x"7A",x"7A",
		x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",x"84",x"84",
		x"84",x"84",x"84",x"82",x"82",x"80",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"82",x"84",x"82",x"82",x"82",x"82",x"80",
		x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"80",x"82",x"82",x"84",x"82",x"82",x"82",x"82",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"7E",x"80",x"80",x"82",x"82",x"84",x"84",
		x"82",x"82",x"82",x"80",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"80",x"7E",x"80",x"80",x"82",x"84",x"84",x"84",x"82",x"82",x"80",x"80",x"7E",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",x"82",x"84",x"84",x"82",
		x"82",x"82",x"80",x"80",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"7E",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"80",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7E",x"7C",x"7E",x"7E",x"7E",x"80",x"7E",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"80",
		x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"82",
		x"80",x"80",x"7E",x"7E",x"7E",x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",
		x"80",x"80",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",x"82",x"82",x"82",x"80",x"80",x"80",
		x"7E",x"7E",x"7C",x"7C",x"7C",x"7C",x"7C",x"7E",x"7E",x"7C",x"7E",x"7E",x"7E",x"80",x"80",x"82",
		x"82",x"82",x"82",x"82",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"7E",x"7E",x"7E",x"7C",
		x"7C",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",x"82",x"82",x"82",x"82",
		x"80",x"7E",x"7E",x"7E",x"7E",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",
		x"82",x"82",x"82",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7E",x"7C",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"82",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7C",x"7E",
		x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"82",x"82",x"80",x"80",x"80",
		x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",
		x"82",x"82",x"82",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"80",x"80",x"80",x"82",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7C",x"7C",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"82",x"82",x"80",x"80",x"80",x"80",x"80",x"7E",x"7C",x"7C",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"80",x"80",x"80",x"82",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",
		x"82",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7C",x"7E",x"7E",
		x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7C",x"7C",x"7E",x"7C",
		x"7C",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"7E",x"7C",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",
		x"7E",x"7E",x"7C",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"7E",x"7E",x"7C",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"82",x"80",x"80",
		x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7E",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7E",x"7E",x"7E",x"7E",x"7E",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"7F",x"80",x"80",x"7F",x"7F",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",
		x"80",x"7F",x"80",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"7F",
		x"7F",x"7F",x"7F",x"80",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"80",x"7F",x"7F",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",
		x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"81",x"81",x"83",x"83",x"84",x"84",x"84",
		x"84",x"84",x"84",x"84",x"83",x"83",x"83",x"83",x"81",x"81",x"81",x"80",x"80",x"80",x"7F",x"7F",
		x"7D",x"7D",x"7D",x"7D",x"7C",x"7C",x"79",x"77",x"76",x"74",x"73",x"73",x"74",x"74",x"76",x"77",
		x"77",x"7A",x"7A",x"7D",x"7F",x"80",x"81",x"81",x"83",x"84",x"86",x"87",x"87",x"87",x"89",x"89",
		x"89",x"89",x"89",x"87",x"87",x"87",x"87",x"87",x"86",x"86",x"86",x"84",x"84",x"84",x"83",x"83",
		x"81",x"81",x"81",x"81",x"80",x"80",x"80",x"80",x"83",x"87",x"8A",x"8C",x"8D",x"8D",x"8C",x"8A",
		x"87",x"84",x"83",x"80",x"7D",x"7A",x"77",x"74",x"73",x"71",x"70",x"6E",x"6D",x"6D",x"6B",x"6B",
		x"6B",x"6B",x"6D",x"6D",x"6D",x"6E",x"70",x"70",x"70",x"6E",x"6B",x"6A",x"68",x"68",x"68",x"6A",
		x"6B",x"6E",x"71",x"74",x"77",x"7A",x"7F",x"81",x"84",x"89",x"8A",x"8D",x"90",x"93",x"95",x"96",
		x"98",x"99",x"9B",x"9B",x"9B",x"9B",x"99",x"99",x"99",x"98",x"96",x"96",x"95",x"93",x"92",x"93",
		x"96",x"9B",x"9F",x"A1",x"A1",x"A1",x"9E",x"99",x"95",x"8F",x"89",x"84",x"7F",x"79",x"73",x"6E",
		x"6A",x"67",x"62",x"61",x"5E",x"5C",x"5B",x"59",x"59",x"59",x"59",x"5B",x"5B",x"5C",x"5E",x"5F",
		x"62",x"64",x"67",x"68",x"6B",x"6E",x"70",x"73",x"76",x"77",x"7A",x"7C",x"7D",x"80",x"81",x"83",
		x"84",x"86",x"87",x"89",x"89",x"8A",x"8A",x"8C",x"8C",x"8D",x"8D",x"8D",x"8D",x"8D",x"8D",x"8C",
		x"8C",x"8C",x"89",x"84",x"81",x"7D",x"7A",x"79",x"79",x"77",x"79",x"79",x"7A",x"7C",x"7D",x"7F",
		x"80",x"81",x"84",x"86",x"87",x"89",x"8A",x"8A",x"8C",x"8D",x"8D",x"8F",x"8F",x"8F",x"8F",x"8F",
		x"8F",x"8F",x"8F",x"8D",x"8D",x"8D",x"8C",x"8A",x"8A",x"89",x"89",x"87",x"87",x"87",x"86",x"86",
		x"86",x"87",x"8F",x"96",x"9C",x"A2",x"A4",x"A4",x"9F",x"9B",x"96",x"8F",x"89",x"81",x"7A",x"74",
		x"6E",x"68",x"62",x"5E",x"59",x"56",x"55",x"52",x"50",x"50",x"50",x"50",x"50",x"52",x"53",x"55",
		x"56",x"59",x"5B",x"59",x"58",x"58",x"58",x"59",x"5C",x"5F",x"62",x"67",x"6B",x"70",x"74",x"79",
		x"7F",x"83",x"87",x"8A",x"8F",x"92",x"96",x"99",x"9C",x"9E",x"A1",x"A2",x"A4",x"A5",x"AA",x"B3",
		x"BA",x"C0",x"C3",x"C5",x"C3",x"C0",x"BC",x"B6",x"B0",x"A8",x"A1",x"99",x"92",x"8A",x"84",x"7D",
		x"79",x"73",x"6E",x"6A",x"67",x"64",x"61",x"5F",x"5E",x"5C",x"5C",x"5C",x"5C",x"5C",x"5E",x"5F",
		x"5F",x"61",x"62",x"64",x"67",x"68",x"6A",x"6D",x"6E",x"71",x"73",x"76",x"77",x"79",x"7A",x"7C",
		x"7D",x"7F",x"80",x"7D",x"7A",x"79",x"77",x"77",x"77",x"77",x"79",x"7A",x"7C",x"7F",x"80",x"83",
		x"86",x"87",x"8A",x"8C",x"8F",x"90",x"92",x"93",x"95",x"95",x"96",x"96",x"98",x"98",x"98",x"99",
		x"99",x"9E",x"A4",x"AA",x"B0",x"B3",x"B3",x"B1",x"AE",x"AA",x"A4",x"9E",x"96",x"90",x"89",x"83",
		x"7C",x"76",x"71",x"6B",x"67",x"64",x"61",x"5E",x"5B",x"59",x"58",x"58",x"58",x"58",x"58",x"58",
		x"59",x"5B",x"5C",x"5E",x"5F",x"5F",x"5E",x"5C",x"5C",x"5C",x"5E",x"61",x"62",x"65",x"6A",x"6D",
		x"71",x"74",x"79",x"7D",x"81",x"84",x"87",x"8C",x"8F",x"92",x"93",x"96",x"98",x"99",x"9B",x"9B",
		x"9C",x"9C",x"9C",x"9C",x"9C",x"9C",x"9B",x"99",x"99",x"98",x"96",x"95",x"95",x"93",x"92",x"90",
		x"90",x"95",x"9B",x"A2",x"A7",x"AA",x"AB",x"A8",x"A5",x"9F",x"98",x"92",x"8A",x"81",x"7C",x"74",
		x"6E",x"68",x"62",x"5E",x"5B",x"56",x"55",x"53",x"52",x"50",x"50",x"50",x"50",x"52",x"53",x"55",
		x"56",x"59",x"5B",x"5E",x"61",x"64",x"67",x"6A",x"6D",x"70",x"73",x"76",x"79",x"7C",x"7D",x"80",
		x"83",x"84",x"86",x"89",x"8A",x"8C",x"8C",x"8D",x"8F",x"90",x"90",x"92",x"92",x"92",x"92",x"92",
		x"90",x"90",x"8F",x"8D",x"89",x"84",x"81",x"7F",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7F",
		x"80",x"81",x"84",x"86",x"87",x"89",x"8A",x"8C",x"8D",x"8D",x"8F",x"8F",x"90",x"90",x"90",x"90",
		x"90",x"90",x"8F",x"8F",x"8D",x"8D",x"8C",x"8C",x"8A",x"8A",x"89",x"87",x"86",x"84",x"84",x"83",
		x"81",x"81",x"80",x"80",x"7F",x"7F",x"7D",x"7C",x"7C",x"7C",x"7A",x"7A",x"79",x"79",x"79",x"79",
		x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"76",x"76",x"76",x"76",x"77",x"77",x"77",x"77",x"77",
		x"77",x"77",x"77",x"77",x"77",x"77",x"79",x"79",x"79",x"7A",x"7C",x"7D",x"84",x"90",x"9B",x"A2",
		x"A7",x"A7",x"A5",x"A1",x"9B",x"95",x"8D",x"86",x"7F",x"79",x"71",x"6D",x"67",x"62",x"5F",x"5C",
		x"59",x"58",x"56",x"56",x"56",x"56",x"56",x"58",x"59",x"5B",x"5E",x"5F",x"62",x"65",x"68",x"6B",
		x"6E",x"71",x"74",x"77",x"7A",x"7D",x"80",x"81",x"81",x"80",x"7F",x"7D",x"7D",x"7F",x"80",x"81",
		x"83",x"86",x"89",x"8A",x"8D",x"90",x"93",x"95",x"98",x"99",x"9B",x"9C",x"9E",x"9F",x"9F",x"9F",
		x"9F",x"9F",x"9F",x"9F",x"9E",x"9E",x"9E",x"9C",x"9B",x"99",x"99",x"98",x"9B",x"A2",x"A8",x"AE",
		x"B0",x"B0",x"AD",x"AA",x"A4",x"9E",x"96",x"8F",x"87",x"80",x"79",x"71",x"6B",x"67",x"61",x"5C",
		x"59",x"56",x"53",x"52",x"50",x"50",x"50",x"50",x"50",x"52",x"53",x"56",x"58",x"59",x"5C",x"5F",
		x"61",x"64",x"67",x"6A",x"6D",x"6E",x"71",x"74",x"77",x"79",x"7A",x"7A",x"79",x"76",x"76",x"76",
		x"76",x"77",x"79",x"7C",x"7D",x"80",x"83",x"86",x"89",x"8A",x"8D",x"90",x"92",x"95",x"96",x"98",
		x"99",x"99",x"9B",x"9B",x"9C",x"9B",x"9B",x"9B",x"9B",x"99",x"99",x"98",x"98",x"96",x"95",x"93",
		x"92",x"90",x"8F",x"8D",x"8C",x"8A",x"89",x"87",x"86",x"84",x"84",x"83",x"84",x"89",x"90",x"98",
		x"9E",x"A1",x"A1",x"9F",x"9B",x"96",x"90",x"89",x"81",x"7C",x"74",x"6D",x"67",x"62",x"5C",x"58",
		x"55",x"52",x"4F",x"4D",x"4C",x"4A",x"47",x"43",x"41",x"40",x"40",x"41",x"44",x"49",x"4C",x"52",
		x"56",x"5C",x"62",x"68",x"6D",x"73",x"79",x"7D",x"83",x"87",x"8C",x"90",x"93",x"96",x"99",x"9C",
		x"9E",x"9F",x"A1",x"A2",x"A4",x"A4",x"A4",x"A4",x"A4",x"A4",x"A2",x"A2",x"A1",x"A1",x"A1",x"A5",
		x"AE",x"B4",x"BA",x"BC",x"BA",x"B7",x"B1",x"AB",x"A4",x"9C",x"93",x"8C",x"83",x"7C",x"76",x"6E",
		x"68",x"62",x"5F",x"5B",x"58",x"55",x"53",x"52",x"52",x"52",x"52",x"52",x"53",x"55",x"56",x"58",
		x"59",x"5B",x"5E",x"5C",x"5B",x"5B",x"5B",x"5C",x"5F",x"62",x"65",x"68",x"6D",x"71",x"76",x"7A",
		x"7F",x"83",x"87",x"8C",x"8F",x"92",x"95",x"98",x"9B",x"9C",x"9E",x"9F",x"A1",x"A1",x"A2",x"A2",
		x"A2",x"A2",x"A2",x"A4",x"AA",x"B1",x"B7",x"BC",x"BC",x"BC",x"B9",x"B3",x"AD",x"A7",x"9F",x"98",
		x"8F",x"87",x"80",x"79",x"73",x"6D",x"68",x"64",x"5F",x"5C",x"59",x"56",x"55",x"55",x"53",x"55",
		x"55",x"55",x"56",x"58",x"5B",x"5C",x"5E",x"61",x"62",x"65",x"68",x"6A",x"6B",x"6B",x"6A",x"68",
		x"68",x"6A",x"6A",x"6D",x"6E",x"71",x"76",x"79",x"7C",x"80",x"83",x"86",x"8A",x"8D",x"90",x"92",
		x"95",x"96",x"98",x"9B",x"9B",x"9C",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9C",x"9B",x"99",x"98",
		x"98",x"96",x"95",x"93",x"92",x"90",x"8F",x"8C",x"8A",x"89",x"87",x"86",x"84",x"84",x"86",x"8D",
		x"95",x"9C",x"A2",x"A4",x"A2",x"9F",x"99",x"93",x"8C",x"84",x"7F",x"77",x"70",x"68",x"64",x"5E",
		x"59",x"55",x"52",x"4F",x"4D",x"4C",x"4A",x"4A",x"4C",x"4C",x"4D",x"50",x"52",x"55",x"56",x"58",
		x"56",x"56",x"56",x"56",x"59",x"5C",x"61",x"65",x"6A",x"6E",x"74",x"79",x"7F",x"83",x"87",x"8C",
		x"90",x"95",x"98",x"9B",x"9E",x"A1",x"A4",x"A5",x"A7",x"A8",x"AB",x"B0",x"B9",x"C0",x"C5",x"C8",
		x"C8",x"C5",x"C0",x"BC",x"B6",x"AE",x"A7",x"9E",x"96",x"8F",x"87",x"81",x"7C",x"74",x"70",x"6B",
		x"67",x"62",x"5F",x"5E",x"5B",x"59",x"59",x"59",x"59",x"59",x"5B",x"5B",x"5C",x"5E",x"5F",x"61",
		x"64",x"65",x"67",x"68",x"68",x"67",x"65",x"65",x"65",x"65",x"68",x"6A",x"6D",x"70",x"73",x"77",
		x"7A",x"7F",x"81",x"86",x"89",x"8D",x"8F",x"92",x"95",x"96",x"99",x"9B",x"9C",x"9C",x"9E",x"9E",
		x"9E",x"9E",x"9E",x"9C",x"9C",x"9B",x"99",x"99",x"98",x"96",x"93",x"92",x"90",x"8F",x"8D",x"8C",
		x"89",x"87",x"86",x"84",x"83",x"81",x"81",x"81",x"83",x"8A",x"93",x"9B",x"9F",x"A1",x"A1",x"9C",
		x"98",x"92",x"8A",x"84",x"7C",x"76",x"6E",x"68",x"62",x"5C",x"58",x"55",x"52",x"4F",x"4D",x"4D",
		x"4C",x"4C",x"4D",x"4D",x"4F",x"50",x"53",x"55",x"58",x"5B",x"5F",x"62",x"65",x"6A",x"6D",x"70",
		x"74",x"77",x"7A",x"7D",x"80",x"83",x"84",x"87",x"89",x"8A",x"8D",x"8F",x"8F",x"90",x"92",x"92",
		x"93",x"93",x"92",x"8D",x"89",x"86",x"84",x"83",x"81",x"83",x"83",x"83",x"84",x"86",x"87",x"89",
		x"8A",x"8C",x"8D",x"8F",x"90",x"90",x"92",x"92",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",
		x"92",x"90",x"90",x"8F",x"8D",x"8D",x"8C",x"8A",x"89",x"89",x"87",x"86",x"84",x"83",x"83",x"81",
		x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"81",x"89",x"92",x"99",x"9E",x"A1",x"9F",x"9C",x"98",x"93",
		x"8C",x"86",x"7F",x"77",x"71",x"6B",x"65",x"61",x"5C",x"58",x"55",x"53",x"50",x"4F",x"4F",x"4F",
		x"4F",x"50",x"52",x"53",x"55",x"58",x"59",x"5C",x"5F",x"62",x"65",x"68",x"6B",x"6E",x"70",x"73",
		x"73",x"71",x"70",x"70",x"71",x"73",x"74",x"77",x"7A",x"7F",x"81",x"84",x"89",x"8C",x"8F",x"93",
		x"96",x"98",x"9B",x"9C",x"9E",x"A1",x"A1",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A1",
		x"A1",x"A5",x"AB",x"B3",x"B9",x"BA",x"BA",x"B7",x"B3",x"AD",x"A5",x"9F",x"96",x"8F",x"87",x"80",
		x"79",x"71",x"6B",x"65",x"61",x"5E",x"59",x"56",x"55",x"53",x"52",x"50",x"50",x"50",x"52",x"50",
		x"4F",x"4C",x"4A",x"4A",x"4C",x"4F",x"52",x"55",x"59",x"5E",x"62",x"68",x"6D",x"71",x"77",x"7C",
		x"80",x"84",x"87",x"8C",x"8F",x"92",x"95",x"98",x"99",x"9B",x"9C",x"9E",x"9E",x"9F",x"9F",x"9F",
		x"9F",x"9F",x"9E",x"9E",x"9E",x"9C",x"9F",x"A7",x"AE",x"B4",x"B6",x"B7",x"B6",x"B1",x"AB",x"A5",
		x"9E",x"96",x"8D",x"86",x"7F",x"77",x"70",x"6A",x"65",x"5F",x"5B",x"58",x"55",x"53",x"52",x"50",
		x"50",x"50",x"52",x"52",x"53",x"55",x"56",x"59",x"5C",x"5E",x"61",x"64",x"67",x"6A",x"6D",x"70",
		x"73",x"76",x"77",x"7A",x"7C",x"7D",x"7C",x"7A",x"79",x"79",x"79",x"7A",x"7C",x"7D",x"7F",x"81",
		x"84",x"87",x"89",x"8C",x"8F",x"90",x"93",x"95",x"98",x"99",x"99",x"9B",x"9C",x"9C",x"9C",x"9C",
		x"9C",x"9C",x"9B",x"9B",x"99",x"99",x"98",x"98",x"96",x"98",x"9E",x"A5",x"AB",x"AE",x"B0",x"AE",
		x"AB",x"A7",x"A1",x"99",x"92",x"8A",x"81",x"7C",x"74",x"6D",x"67",x"62",x"5E",x"59",x"56",x"53",
		x"52",x"50",x"4F",x"4F",x"4F",x"4F",x"50",x"52",x"53",x"56",x"58",x"5B",x"5E",x"61",x"64",x"67",
		x"6A",x"6D",x"70",x"73",x"76",x"77",x"7A",x"7D",x"7F",x"81",x"83",x"84",x"87",x"87",x"89",x"8A",
		x"8C",x"8A",x"87",x"84",x"81",x"80",x"80",x"80",x"80",x"81",x"83",x"84",x"86",x"87",x"89",x"8A",
		x"8D",x"8F",x"90",x"92",x"93",x"93",x"95",x"95",x"96",x"96",x"96",x"96",x"95",x"95",x"95",x"93",
		x"93",x"92",x"92",x"92",x"90",x"8F",x"8F",x"8F",x"92",x"99",x"A1",x"A5",x"A7",x"A7",x"A5",x"A1",
		x"9C",x"96",x"8F",x"87",x"81",x"7A",x"74",x"6D",x"67",x"62",x"5E",x"5B",x"56",x"53",x"52",x"50",
		x"50",x"50",x"50",x"52",x"52",x"53",x"55",x"58",x"59",x"5C",x"5F",x"62",x"64",x"67",x"6A",x"6D",
		x"70",x"73",x"76",x"79",x"7A",x"7D",x"80",x"81",x"83",x"84",x"86",x"87",x"89",x"8A",x"8C",x"8A",
		x"87",x"84",x"81",x"80",x"7F",x"7F",x"7F",x"80",x"81",x"83",x"84",x"86",x"87",x"8A",x"8C",x"8D",
		x"8F",x"90",x"92",x"93",x"95",x"95",x"96",x"96",x"96",x"96",x"96",x"96",x"96",x"96",x"96",x"95",
		x"95",x"95",x"95",x"96",x"9E",x"A4",x"AA",x"AD",x"AD",x"AB",x"A8",x"A2",x"9C",x"96",x"8F",x"87",
		x"80",x"7A",x"73",x"6D",x"67",x"62",x"5E",x"5B",x"58",x"55",x"53",x"52",x"52",x"52",x"52",x"52",
		x"53",x"55",x"56",x"59",x"5B",x"5E",x"5F",x"62",x"65",x"68",x"6A",x"6D",x"70",x"73",x"74",x"77",
		x"79",x"7A",x"7A",x"79",x"77",x"76",x"74",x"76",x"77",x"79",x"7A",x"7C",x"7F",x"81",x"84",x"87",
		x"8A",x"8D",x"90",x"92",x"95",x"96",x"98",x"99",x"9B",x"9C",x"9C",x"9E",x"9E",x"9E",x"9E",x"9C",
		x"9C",x"9C",x"9B",x"9B",x"99",x"98",x"96",x"95",x"93",x"92",x"90",x"8F",x"8D",x"8C",x"8A",x"89",
		x"86",x"86",x"84",x"84",x"89",x"8F",x"95",x"99",x"9B",x"99",x"96",x"93",x"8D",x"87",x"81",x"7C",
		x"76",x"70",x"6A",x"65",x"5F",x"5C",x"59",x"56",x"53",x"52",x"50",x"50",x"50",x"50",x"52",x"53",
		x"55",x"58",x"59",x"5C",x"5F",x"61",x"64",x"67",x"6A",x"6B",x"6D",x"6B",x"6B",x"6A",x"6B",x"6B",
		x"6E",x"70",x"73",x"77",x"7A",x"7D",x"81",x"84",x"89",x"8C",x"90",x"93",x"96",x"99",x"9B",x"9E",
		x"9F",x"A1",x"A1",x"A2",x"A2",x"A4",x"A4",x"A4",x"A4",x"A4",x"A2",x"A1",x"9F",x"9E",x"9C",x"9B",
		x"99",x"98",x"96",x"95",x"93",x"92",x"92",x"96",x"9C",x"A1",x"A2",x"A2",x"A1",x"9E",x"98",x"92",
		x"8C",x"86",x"7F",x"79",x"71",x"6B",x"67",x"61",x"5E",x"59",x"56",x"53",x"52",x"50",x"4F",x"4D",
		x"4A",x"46",x"43",x"43",x"43",x"46",x"49",x"4C",x"50",x"55",x"59",x"5F",x"65",x"6A",x"70",x"76",
		x"7A",x"80",x"84",x"89",x"8D",x"90",x"95",x"98",x"9B",x"9C",x"9E",x"9F",x"A1",x"A2",x"A2",x"A4",
		x"A4",x"A4",x"A4",x"A7",x"AE",x"B4",x"B7",x"B9",x"B7",x"B4",x"B0",x"AB",x"A4",x"9E",x"96",x"8F",
		x"87",x"80",x"79",x"73",x"6D",x"68",x"64",x"61",x"5E",x"5B",x"59",x"58",x"58",x"56",x"56",x"58",
		x"59",x"59",x"5B",x"5E",x"5F",x"62",x"64",x"67",x"68",x"6B",x"6E",x"70",x"73",x"76",x"79",x"7A",
		x"7D",x"7F",x"80",x"83",x"84",x"84",x"86",x"86",x"83",x"80",x"7D",x"7D",x"7C",x"7C",x"7D",x"7D",
		x"7F",x"80",x"83",x"84",x"86",x"89",x"8A",x"8D",x"8F",x"90",x"92",x"93",x"95",x"96",x"96",x"96",
		x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"99",x"9E",x"A5",x"AA",x"AD",x"AD",x"AA",x"A7",
		x"A2",x"9C",x"96",x"8F",x"89",x"81",x"7C",x"76",x"70",x"6A",x"65",x"61",x"5E",x"5B",x"58",x"56",
		x"56",x"55",x"55",x"55",x"55",x"56",x"58",x"59",x"5B",x"5E",x"5F",x"62",x"64",x"67",x"6A",x"6B",
		x"6E",x"71",x"73",x"76",x"77",x"7A",x"7C",x"7C",x"79",x"77",x"76",x"76",x"76",x"77",x"79",x"7A",
		x"7D",x"7F",x"81",x"84",x"87",x"8A",x"8C",x"8F",x"92",x"93",x"96",x"98",x"99",x"9B",x"9C",x"9C",
		x"9E",x"9E",x"9E",x"9E",x"9E",x"9C",x"9C",x"9B",x"9B",x"99",x"99",x"9E",x"A4",x"A8",x"AA",x"AA",
		x"A8",x"A5",x"A1",x"9B",x"93",x"8D",x"87",x"80",x"7A",x"74",x"6E",x"68",x"64",x"5F",x"5C",x"59",
		x"58",x"56",x"55",x"55",x"55",x"55",x"56",x"56",x"58",x"59",x"5B",x"5C",x"5F",x"61",x"64",x"67",
		x"6A",x"6B",x"6E",x"71",x"73",x"76",x"79",x"7A",x"7C",x"7D",x"7C",x"79",x"77",x"77",x"77",x"77",
		x"79",x"7A",x"7C",x"7F",x"80",x"83",x"86",x"89",x"8C",x"8F",x"90",x"93",x"95",x"98",x"98",x"9B",
		x"9C",x"9C",x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"9C",x"9C",x"9B",x"99",x"98",x"96",x"95",x"93",
		x"90",x"8F",x"8D",x"8C",x"8A",x"8A",x"8F",x"95",x"98",x"99",x"99",x"98",x"93",x"90",x"8A",x"84",
		x"80",x"7A",x"74",x"70",x"6A",x"65",x"61",x"5E",x"5C",x"59",x"58",x"56",x"56",x"55",x"55",x"55",
		x"56",x"55",x"52",x"50",x"4F",x"4F",x"50",x"53",x"56",x"5B",x"5F",x"64",x"68",x"6E",x"73",x"79",
		x"7D",x"81",x"86",x"8C",x"8F",x"93",x"96",x"99",x"9C",x"9F",x"A1",x"A2",x"A4",x"A5",x"A7",x"AA",
		x"B0",x"B4",x"B9",x"BA",x"BA",x"B7",x"B4",x"AE",x"A8",x"A2",x"9C",x"95",x"8D",x"87",x"81",x"7C",
		x"76",x"71",x"6D",x"68",x"65",x"62",x"61",x"5F",x"5E",x"5C",x"5C",x"5C",x"5C",x"5E",x"5F",x"61",
		x"61",x"62",x"64",x"67",x"68",x"6A",x"6D",x"6E",x"70",x"71",x"73",x"74",x"71",x"70",x"6E",x"6E",
		x"6E",x"70",x"71",x"74",x"77",x"7A",x"7D",x"81",x"84",x"87",x"8C",x"8F",x"90",x"93",x"96",x"98",
		x"9B",x"9C",x"9E",x"9F",x"9F",x"A1",x"A2",x"A8",x"AE",x"B3",x"B4",x"B6",x"B4",x"B0",x"AB",x"A7",
		x"A1",x"9B",x"93",x"8D",x"87",x"81",x"7A",x"76",x"71",x"6D",x"68",x"65",x"62",x"5F",x"5E",x"5C",
		x"5C",x"5B",x"5B",x"5B",x"5C",x"5C",x"5E",x"5F",x"61",x"62",x"64",x"67",x"68",x"6A",x"6D",x"6E",
		x"71",x"73",x"74",x"76",x"77",x"77",x"74",x"73",x"71",x"71",x"71",x"73",x"74",x"76",x"79",x"7C",
		x"7F",x"81",x"84",x"87",x"8A",x"8D",x"90",x"93",x"95",x"98",x"99",x"9C",x"9C",x"9E",x"9E",x"9E",
		x"9E",x"9E",x"9E",x"9C",x"9B",x"99",x"98",x"96",x"95",x"93",x"92",x"8F",x"8D",x"8C",x"8A",x"87",
		x"86",x"83",x"81",x"80",x"7F",x"7D",x"7C",x"79",x"79",x"77",x"76",x"76",x"76",x"76",x"77",x"7C",
		x"81",x"86",x"89",x"89",x"89",x"87",x"84",x"81",x"7F",x"7A",x"77",x"73",x"70",x"6D",x"6A",x"67",
		x"64",x"62",x"61",x"61",x"61",x"5F",x"61",x"61",x"61",x"62",x"64",x"65",x"67",x"6A",x"6B",x"6D",
		x"70",x"73",x"74",x"76",x"79",x"7A",x"7C",x"7F",x"80",x"81",x"83",x"84",x"86",x"87",x"89",x"89",
		x"8A",x"8A",x"8C",x"8C",x"8C",x"8D",x"8D",x"8F",x"8F",x"8F",x"8D",x"8D",x"8D",x"8D",x"8C",x"8C",
		x"8A",x"86",x"81",x"7D",x"7A",x"79",x"77",x"77",x"77",x"77",x"79",x"7A",x"7C",x"7F",x"81",x"83",
		x"86",x"87",x"8A",x"8C",x"8D",x"90",x"92",x"92",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"92",
		x"90",x"90",x"8F",x"8D",x"8C",x"8A",x"89",x"87",x"86",x"84",x"83",x"81",x"80",x"7F",x"7D",x"7C",
		x"7A",x"79",x"79",x"77",x"77",x"76",x"76",x"77",x"7C",x"80",x"84",x"87",x"89",x"89",x"87",x"84",
		x"81",x"7F",x"7A",x"77",x"73",x"70",x"6D",x"6A",x"67",x"65",x"64",x"62",x"61",x"61",x"61",x"61",
		x"61",x"61",x"62",x"64",x"65",x"67",x"68",x"6A",x"6D",x"70",x"71",x"73",x"76",x"79",x"7A",x"7C",
		x"7F",x"80",x"81",x"83",x"84",x"86",x"87",x"89",x"89",x"89",x"86",x"81",x"80",x"7F",x"7D",x"7D",
		x"7D",x"7F",x"80",x"81",x"84",x"86",x"89",x"8C",x"8D",x"90",x"92",x"95",x"96",x"98",x"99",x"99",
		x"9B",x"9B",x"9B",x"9B",x"99",x"99",x"98",x"96",x"95",x"93",x"93",x"90",x"8F",x"8D",x"8A",x"89",
		x"87",x"86",x"84",x"83",x"81",x"80",x"7F",x"7D",x"7F",x"83",x"86",x"89",x"8A",x"8A",x"89",x"86",
		x"83",x"80",x"7C",x"79",x"74",x"71",x"6E",x"6A",x"67",x"65",x"62",x"61",x"5F",x"5F",x"5F",x"5F",
		x"5F",x"5F",x"61",x"61",x"62",x"64",x"67",x"68",x"6A",x"6B",x"6D",x"70",x"71",x"73",x"74",x"74",
		x"71",x"71",x"70",x"70",x"70",x"73",x"74",x"77",x"7A",x"7D",x"81",x"84",x"87",x"8C",x"8F",x"92",
		x"95",x"98",x"99",x"9B",x"9E",x"9E",x"9F",x"9F",x"9F",x"9F",x"9F",x"9E",x"9E",x"9C",x"9B",x"99",
		x"98",x"96",x"93",x"92",x"90",x"8D",x"8C",x"89",x"87",x"86",x"84",x"83",x"80",x"80",x"7D",x"7C",
		x"7C",x"7A",x"79",x"77",x"77",x"76",x"76",x"74",x"74",x"74",x"74",x"74",x"74",x"74",x"77",x"7C",
		x"81",x"84",x"87",x"89",x"87",x"87",x"84",x"83",x"80",x"7D",x"7A",x"76",x"73",x"71",x"6E",x"6D",
		x"6B",x"6A",x"68",x"68",x"67",x"67",x"67",x"67",x"68",x"68",x"65",x"62",x"5F",x"5E",x"5F",x"5F",
		x"62",x"64",x"68",x"6B",x"70",x"74",x"79",x"7D",x"81",x"86",x"8A",x"8D",x"90",x"95",x"96",x"99",
		x"9B",x"9C",x"9E",x"9F",x"9F",x"9F",x"9F",x"A1",x"A2",x"A5",x"AA",x"AB",x"AB",x"AB",x"A8",x"A5",
		x"A1",x"9C",x"96",x"92",x"8C",x"87",x"81",x"7D",x"79",x"76",x"73",x"70",x"6D",x"6A",x"68",x"67",
		x"65",x"65",x"65",x"64",x"65",x"65",x"65",x"67",x"67",x"68",x"6A",x"6B",x"6D",x"6E",x"70",x"71",
		x"73",x"74",x"76",x"77",x"76",x"74",x"71",x"70",x"70",x"70",x"71",x"73",x"74",x"77",x"7A",x"7D",
		x"80",x"83",x"86",x"89",x"8C",x"8F",x"92",x"93",x"95",x"96",x"98",x"99",x"99",x"99",x"99",x"98",
		x"98",x"96",x"96",x"95",x"93",x"92",x"90",x"8F",x"8D",x"8C",x"8A",x"89",x"86",x"84",x"84",x"83",
		x"81",x"84",x"87",x"8A",x"8C",x"8C",x"8C",x"8A",x"87",x"84",x"80",x"7D",x"79",x"76",x"73",x"70",
		x"6D",x"6A",x"68",x"67",x"65",x"64",x"64",x"64",x"64",x"64",x"64",x"65",x"65",x"67",x"68",x"6A",
		x"6B",x"6D",x"6E",x"70",x"71",x"70",x"6D",x"6B",x"6A",x"6B",x"6D",x"6E",x"71",x"74",x"77",x"7C",
		x"7F",x"81",x"86",x"89",x"8C",x"8F",x"92",x"95",x"96",x"98",x"99",x"9B",x"9C",x"9C",x"9C",x"9C",
		x"9C",x"9B",x"99",x"99",x"98",x"96",x"96",x"95",x"93",x"95",x"98",x"99",x"99",x"99",x"98",x"96",
		x"93",x"8F",x"8C",x"87",x"83",x"7F",x"7A",x"77",x"73",x"70",x"6D",x"6A",x"68",x"65",x"65",x"64",
		x"64",x"62",x"62",x"62",x"64",x"64",x"65",x"67",x"67",x"68",x"6A",x"6D",x"6E",x"70",x"71",x"73",
		x"74",x"76",x"76",x"74",x"73",x"71",x"70",x"70",x"71",x"73",x"76",x"79",x"7C",x"7F",x"81",x"84",
		x"87",x"8C",x"8D",x"90",x"93",x"95",x"96",x"98",x"99",x"99",x"99",x"99",x"99",x"99",x"98",x"98",
		x"96",x"95",x"93",x"92",x"90",x"8F",x"8D",x"8C",x"89",x"87",x"86",x"84",x"83",x"81",x"80",x"7F",
		x"7F",x"7D",x"7C",x"7A",x"7A",x"79",x"79",x"77",x"77",x"77",x"76",x"76",x"76",x"76",x"76",x"76",
		x"76",x"76",x"76",x"76",x"77",x"7A",x"7F",x"83",x"86",x"87",x"89",x"89",x"87",x"86",x"84",x"81",
		x"80",x"7D",x"7C",x"79",x"77",x"74",x"73",x"71",x"70",x"70",x"6E",x"6E",x"6E",x"6E",x"6E",x"70",
		x"70",x"70",x"71",x"73",x"73",x"74",x"74",x"76",x"77",x"79",x"7A",x"7C",x"7D",x"7D",x"7F",x"80",
		x"80",x"81",x"83",x"83",x"83",x"84",x"84",x"86",x"86",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"89",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"86",x"86",x"84",x"80",x"7C",x"79",x"77",x"76",
		x"76",x"76",x"77",x"79",x"7A",x"7D",x"7F",x"80",x"83",x"86",x"87",x"89",x"8A",x"8C",x"8D",x"8F",
		x"8F",x"90",x"90",x"90",x"90",x"8F",x"8F",x"8F",x"8D",x"8C",x"8C",x"8A",x"89",x"87",x"86",x"86",
		x"83",x"83",x"81",x"80",x"7F",x"7D",x"7D",x"7C",x"7A",x"7A",x"79",x"79",x"77",x"76",x"76",x"76",
		x"76",x"76",x"74",x"74",x"76",x"76",x"76",x"79",x"7C",x"80",x"83",x"84",x"84",x"84",x"84",x"83",
		x"80",x"7F",x"7D",x"7A",x"79",x"77",x"74",x"73",x"71",x"70",x"70",x"6E",x"6E",x"6E",x"6E",x"6E",
		x"6E",x"6E",x"70",x"70",x"71",x"73",x"74",x"76",x"77",x"77",x"79",x"7A",x"7C",x"7D",x"7D",x"7F",
		x"7F",x"7D",x"7A",x"79",x"77",x"77",x"79",x"7A",x"7C",x"7F",x"80",x"83",x"86",x"89",x"8C",x"8D",
		x"8F",x"92",x"93",x"95",x"95",x"96",x"96",x"96",x"96",x"96",x"96",x"95",x"95",x"93",x"92",x"92",
		x"90",x"8F",x"8C",x"8A",x"89",x"87",x"86",x"86",x"84",x"83",x"81",x"80",x"80",x"81",x"84",x"86",
		x"87",x"87",x"87",x"86",x"83",x"81",x"7F",x"7C",x"79",x"76",x"73",x"71",x"6E",x"6D",x"6B",x"6A",
		x"6A",x"68",x"68",x"68",x"67",x"68",x"68",x"68",x"6A",x"6B",x"6D",x"6E",x"70",x"71",x"73",x"74",
		x"76",x"77",x"77",x"7A",x"7A",x"7C",x"7D",x"7F",x"7F",x"7D",x"7A",x"79",x"79",x"79",x"79",x"7A",
		x"7C",x"7F",x"80",x"83",x"86",x"87",x"8A",x"8C",x"8F",x"90",x"92",x"92",x"93",x"95",x"95",x"95",
		x"95",x"95",x"95",x"93",x"93",x"92",x"90",x"90",x"8F",x"8D",x"8C",x"8A",x"89",x"87",x"86",x"86",
		x"84",x"83",x"81",x"81",x"81",x"83",x"86",x"87",x"89",x"89",x"87",x"86",x"83",x"81",x"7F",x"7C",
		x"79",x"77",x"74",x"73",x"70",x"6E",x"6D",x"6B",x"6B",x"6A",x"6A",x"6A",x"6A",x"6A",x"6A",x"6A",
		x"6B",x"6D",x"6D",x"6E",x"70",x"70",x"71",x"73",x"74",x"76",x"77",x"79",x"79",x"7A",x"79",x"76",
		x"74",x"74",x"74",x"76",x"77",x"7A",x"7D",x"7F",x"81",x"84",x"87",x"89",x"8C",x"8F",x"90",x"92",
		x"93",x"93",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"93",x"92",x"92",x"90",x"8F",x"8D",x"8C",
		x"8A",x"89",x"89",x"87",x"86",x"84",x"83",x"81",x"80",x"80",x"7F",x"7F",x"7D",x"7C",x"7C",x"7D",
		x"7F",x"81",x"83",x"83",x"83",x"83",x"81",x"80",x"7F",x"7C",x"7A",x"79",x"76",x"74",x"73",x"71",
		x"70",x"70",x"70",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"70",x"70",x"70",x"70",x"6E",x"6D",
		x"6B",x"6B",x"6D",x"6E",x"70",x"73",x"76",x"77",x"7A",x"7D",x"80",x"83",x"86",x"87",x"8A",x"8C",
		x"8D",x"8F",x"90",x"92",x"92",x"92",x"93",x"92",x"92",x"92",x"92",x"90",x"90",x"8F",x"8F",x"8D",
		x"8C",x"8A",x"8A",x"89",x"87",x"86",x"84",x"84",x"83",x"81",x"81",x"80",x"80",x"7F",x"7F",x"80",
		x"80",x"81",x"83",x"83",x"83",x"81",x"80",x"80",x"7F",x"7D",x"7C",x"7A",x"79",x"77",x"76",x"74",
		x"73",x"73",x"73",x"71",x"71",x"71",x"71",x"71",x"71",x"73",x"73",x"74",x"74",x"76",x"76",x"76",
		x"76",x"74",x"73",x"73",x"73",x"73",x"74",x"76",x"77",x"79",x"7A",x"7D",x"7F",x"81",x"83",x"84",
		x"87",x"89",x"8A",x"8C",x"8D",x"8D",x"8F",x"8F",x"8F",x"8F",x"8F",x"8F",x"8F",x"8D",x"8D",x"8D",
		x"8C",x"8C",x"8A",x"89",x"87",x"87",x"86",x"86",x"84",x"83",x"81",x"81",x"80",x"80",x"7F",x"7F",
		x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7D",
		x"80",x"83",x"84",x"86",x"86",x"86",x"84",x"84",x"83",x"80",x"7F",x"7D",x"7C",x"7A",x"79",x"77",
		x"76",x"76",x"74",x"74",x"74",x"74",x"73",x"73",x"73",x"73",x"74",x"74",x"74",x"76",x"76",x"77",
		x"77",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7D",x"7D",x"7C",x"7A",x"79",x"77",x"77",x"79",x"7A",
		x"7A",x"7D",x"7F",x"81",x"83",x"84",x"87",x"89",x"8A",x"8C",x"8D",x"8F",x"8F",x"8F",x"90",x"90",
		x"90",x"90",x"8F",x"8F",x"8F",x"8D",x"8D",x"8C",x"8C",x"8A",x"89",x"89",x"87",x"86",x"86",x"84",
		x"84",x"83",x"84",x"86",x"87",x"87",x"87",x"87",x"86",x"84",x"83",x"81",x"7F",x"7D",x"7A",x"79",
		x"76",x"74",x"73",x"71",x"71",x"70",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"70",
		x"6E",x"6D",x"6B",x"6B",x"6B",x"6B",x"6D",x"70",x"71",x"74",x"77",x"79",x"7C",x"7F",x"81",x"83",
		x"86",x"87",x"89",x"8A",x"8C",x"8D",x"8F",x"8F",x"90",x"90",x"90",x"90",x"90",x"8F",x"8F",x"8D",
		x"8D",x"8D",x"8C",x"8C",x"8A",x"89",x"89",x"8A",x"8C",x"8D",x"8D",x"8D",x"8C",x"8A",x"89",x"87",
		x"84",x"83",x"80",x"7D",x"7C",x"79",x"77",x"76",x"74",x"73",x"71",x"71",x"70",x"70",x"70",x"70",
		x"70",x"70",x"70",x"70",x"71",x"71",x"73",x"74",x"74",x"76",x"76",x"77",x"79",x"79",x"7A",x"7A",
		x"7A",x"79",x"77",x"76",x"76",x"76",x"77",x"79",x"7A",x"7D",x"7F",x"80",x"83",x"84",x"86",x"89",
		x"8A",x"8A",x"8C",x"8D",x"8D",x"8D",x"8F",x"8F",x"8F",x"8F",x"8F",x"8F",x"8D",x"8D",x"8D",x"8C",
		x"8C",x"8A",x"89",x"89",x"89",x"8A",x"8C",x"8C",x"8C",x"8C",x"8A",x"89",x"86",x"84",x"83",x"80",
		x"7D",x"7C",x"79",x"77",x"76",x"74",x"73",x"71",x"71",x"70",x"70",x"6E",x"6E",x"6E",x"6E",x"70",
		x"70",x"71",x"71",x"73",x"73",x"74",x"74",x"76",x"77",x"79",x"79",x"7A",x"7A",x"7C",x"7C",x"7D",
		x"7F",x"7F",x"7F",x"7F",x"7D",x"7C",x"7A",x"7A",x"7A",x"7A",x"7C",x"7D",x"7F",x"80",x"81",x"83",
		x"84",x"86",x"87",x"89",x"8A",x"8A",x"8A",x"8C",x"8C",x"8D",x"8D",x"8D",x"8C",x"8C",x"8C",x"8A",
		x"8A",x"8A",x"89",x"89",x"87",x"86",x"86",x"84",x"83",x"83",x"81",x"81",x"80",x"80",x"7F",x"7F",
		x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7F",x"80",x"81",x"83",x"81",x"81",x"81",
		x"80",x"7F",x"7D",x"7D",x"7C",x"7A",x"79",x"77",x"76",x"76",x"74",x"74",x"74",x"74",x"74",x"74",
		x"74",x"74",x"74",x"76",x"76",x"76",x"77",x"77",x"79",x"79",x"7A",x"7A",x"7C",x"7C",x"7D",x"7D",
		x"7F",x"7F",x"80",x"80",x"7F",x"7D",x"7C",x"7A",x"7A",x"7A",x"7C",x"7C",x"7D",x"7F",x"80",x"81",
		x"83",x"84",x"86",x"87",x"89",x"89",x"8A",x"8A",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
		x"8A",x"8A",x"89",x"89",x"87",x"87",x"86",x"86",x"84",x"84",x"83",x"83",x"81",x"81",x"80",x"80",
		x"7F",x"7F",x"7F",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",
		x"7C",x"7D",x"7F",x"81",x"81",x"83",x"83",x"81",x"81",x"80",x"80",x"7F",x"7D",x"7D",x"7C",x"7A",
		x"7A",x"79",x"77",x"77",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"77",x"77",x"77",
		x"79",x"79",x"79",x"7A",x"7A",x"7C",x"7C",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"80",x"81",x"81",
		x"83",x"83",x"83",x"83",x"83",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
		x"83",x"83",x"83",x"83",x"80",x"7F",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7F",x"7F",x"80",
		x"81",x"83",x"83",x"84",x"86",x"86",x"86",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"86",
		x"86",x"84",x"84",x"84",x"83",x"83",x"81",x"81",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7D",x"7D",
		x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",
		x"7C",x"7D",x"80",x"81",x"81",x"83",x"83",x"81",x"81",x"80",x"80",x"7F",x"7F",x"7D",x"7C",x"7C",
		x"7A",x"79",x"79",x"79",x"77",x"77",x"77",x"77",x"77",x"77",x"79",x"79",x"79",x"79",x"7A",x"7A",
		x"7A",x"7A",x"7A",x"79",x"77",x"77",x"77",x"79",x"79",x"7A",x"7C",x"7D",x"7F",x"80",x"81",x"83",
		x"84",x"86",x"87",x"89",x"89",x"8A",x"8A",x"8A",x"8A",x"8A",x"8A",x"8A",x"8A",x"8A",x"8A",x"89",
		x"89",x"89",x"89",x"87",x"86",x"86",x"86",x"84",x"84",x"86",x"86",x"87",x"87",x"87",x"86",x"84",
		x"83",x"83",x"80",x"7F",x"7D",x"7C",x"7A",x"79",x"79",x"77",x"76",x"76",x"74",x"74",x"74",x"74",
		x"74",x"74",x"74",x"74",x"74",x"74",x"76",x"77",x"77",x"79",x"79",x"79",x"7A",x"7A",x"7C",x"7C",
		x"7C",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7F",
		x"7F",x"80",x"81",x"81",x"83",x"84",x"86",x"86",x"87",x"87",x"89",x"89",x"89",x"89",x"89",x"89",
		x"89",x"89",x"89",x"89",x"8A",x"8C",x"8C",x"8C",x"8A",x"8A",x"89",x"87",x"86",x"84",x"83",x"81",
		x"80",x"7F",x"7D",x"7C",x"7A",x"79",x"79",x"77",x"77",x"76",x"76",x"76",x"76",x"76",x"76",x"76",
		x"76",x"76",x"76",x"77",x"77",x"77",x"77",x"79",x"79",x"7A",x"7A",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7A",x"7A",x"79",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7F",x"80",x"81",x"83",x"83",x"84",x"84",
		x"86",x"86",x"87",x"87",x"87",x"89",x"89",x"89",x"89",x"87",x"87",x"87",x"87",x"86",x"86",x"86",
		x"86",x"84",x"84",x"83",x"83",x"83",x"81",x"81",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7D",x"7F",x"80",x"80",x"81",x"81",x"83",x"81",x"81",x"81",x"80",x"80",x"7F",x"7F",x"7D",
		x"7D",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",
		x"7A",x"7A",x"79",x"79",x"77",x"79",x"79",x"79",x"7A",x"7C",x"7C",x"7D",x"7F",x"80",x"81",x"83",
		x"83",x"84",x"84",x"86",x"86",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"89",x"89",x"8A",x"89",x"89",x"89",x"87",x"86",x"84",x"83",x"81",x"80",x"80",x"7F",x"7D",x"7C",
		x"7C",x"7A",x"7A",x"79",x"79",x"79",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"79",x"79",x"79",
		x"79",x"79",x"7A",x"79",x"79",x"77",x"77",x"77",x"79",x"79",x"7A",x"7A",x"7C",x"7D",x"7F",x"80",
		x"80",x"81",x"83",x"83",x"84",x"84",x"86",x"86",x"86",x"86",x"87",x"87",x"87",x"86",x"86",x"86",
		x"86",x"86",x"86",x"84",x"84",x"84",x"83",x"83",x"83",x"81",x"81",x"81",x"80",x"80",x"80",x"80",
		x"80",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"81",x"81",x"81",x"81",x"81",x"80",x"80",x"7F",x"7F",
		x"7D",x"7D",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"79",x"79",x"79",x"79",x"79",x"79",x"79",x"79",
		x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7D",x"7D",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7F",x"7F",x"80",x"80",x"81",x"83",x"83",x"84",x"84",x"84",
		x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"86",x"84",x"84",x"84",x"83",
		x"83",x"83",x"81",x"81",x"81",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"7F",x"7F",x"7F",x"7D",x"7D",x"7C",x"7C",x"7C",x"7A",x"7A",x"7A",x"7A",x"7C",x"7A",x"7A",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"80",
		x"80",x"80",x"81",x"81",x"83",x"83",x"83",x"83",x"83",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
		x"84",x"84",x"84",x"83",x"83",x"83",x"83",x"83",x"81",x"81",x"81",x"81",x"80",x"80",x"80",x"80",
		x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"80",x"7F",x"7F",x"7F",x"7F",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"80",x"80",x"80",x"81",x"81",x"83",x"83",x"83",x"83",x"84",
		x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"83",x"83",x"83",x"83",x"83",x"83",x"84",
		x"84",x"83",x"83",x"83",x"81",x"81",x"81",x"80",x"80",x"7F",x"7F",x"7D",x"7D",x"7D",x"7C",x"7C",
		x"7C",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7A",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7A",x"7A",x"7C",x"7C",x"7C",x"7D",x"7D",x"7F",x"7F",x"7F",x"80",x"80",
		x"81",x"81",x"81",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",
		x"83",x"83",x"83",x"81",x"81",x"81",x"81",x"81",x"81",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",
		x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",
		x"80",x"81",x"81",x"81",x"81",x"83",x"81",x"83",x"83",x"83",x"83",x"81",x"83",x"83",x"83",x"83",
		x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"81",x"81",x"81",x"80",x"80",x"80",x"7F",x"7F",x"7F",
		x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"81",
		x"81",x"81",x"81",x"81",x"81",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"81",x"81",
		x"81",x"81",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",
		x"7D",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"81",x"81",
		x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"80",x"81",x"81",x"81",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",
		x"80",x"80",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",x"81",
		x"81",x"81",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7F",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",
		x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"81",x"81",x"81",x"81",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7D",x"7F",x"7D",x"7D",x"7D",
		x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"81",x"81",x"81",
		x"81",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7D",x"7F",x"7D",x"7F",x"7D",x"7D",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"80",x"7F",x"7F",x"7F",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
		x"7F",x"7F",x"80",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"80",x"7F",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"82",
		x"7C",x"7C",x"80",x"87",x"87",x"7C",x"80",x"8B",x"82",x"7C",x"82",x"87",x"82",x"77",x"69",x"7C",
		x"90",x"B1",x"DB",x"D7",x"B6",x"95",x"6E",x"7C",x"95",x"BA",x"DB",x"BF",x"9E",x"82",x"A3",x"B1",
		x"9E",x"B6",x"B6",x"A7",x"87",x"87",x"A7",x"C8",x"BF",x"90",x"7C",x"82",x"82",x"82",x"80",x"7C",
		x"82",x"82",x"80",x"7C",x"82",x"87",x"99",x"99",x"82",x"69",x"43",x"56",x"7C",x"99",x"B6",x"95",
		x"77",x"51",x"43",x"69",x"82",x"A7",x"AC",x"82",x"69",x"43",x"51",x"77",x"90",x"B1",x"99",x"77",
		x"56",x"3F",x"64",x"80",x"A3",x"AC",x"87",x"69",x"48",x"27",x"31",x"51",x"72",x"90",x"80",x"60",
		x"43",x"60",x"82",x"A3",x"B6",x"8B",x"72",x"4D",x"48",x"72",x"8B",x"B1",x"9E",x"80",x"60",x"43",
		x"5B",x"80",x"95",x"72",x"64",x"87",x"90",x"69",x"6E",x"8B",x"AC",x"D2",x"BF",x"9E",x"80",x"90",
		x"B1",x"D2",x"E5",x"C4",x"A7",x"80",x"7C",x"95",x"BA",x"BA",x"90",x"72",x"51",x"35",x"43",x"64",
		x"82",x"69",x"51",x"69",x"51",x"4D",x"5B",x"7C",x"82",x"5B",x"60",x"64",x"4D",x"31",x"3F",x"64",
		x"7C",x"6E",x"48",x"31",x"51",x"77",x"90",x"B6",x"BA",x"99",x"7C",x"56",x"5B",x"80",x"9E",x"90",
		x"69",x"4D",x"2C",x"14",x"31",x"51",x"77",x"82",x"69",x"43",x"3F",x"69",x"82",x"A7",x"9E",x"77",
		x"5B",x"69",x"60",x"4D",x"60",x"6E",x"5B",x"51",x"64",x"7C",x"A7",x"A3",x"87",x"64",x"69",x"8B",
		x"80",x"82",x"99",x"87",x"7C",x"4D",x"3F",x"5B",x"80",x"87",x"80",x"87",x"7C",x"69",x"4D",x"2C",
		x"31",x"60",x"77",x"6E",x"43",x"2C",x"48",x"69",x"8B",x"B1",x"BA",x"9E",x"77",x"51",x"51",x"77",
		x"99",x"90",x"6E",x"80",x"A3",x"BA",x"A3",x"8B",x"A7",x"B6",x"99",x"87",x"AC",x"B1",x"90",x"69",
		x"6E",x"8B",x"AC",x"D7",x"EE",x"E0",x"B6",x"8B",x"77",x"99",x"B6",x"DB",x"E0",x"BA",x"95",x"95",
		x"B6",x"AC",x"B1",x"C4",x"BA",x"9E",x"87",x"95",x"C4",x"D2",x"B6",x"8B",x"87",x"8B",x"87",x"8B",
		x"80",x"82",x"87",x"87",x"80",x"82",x"87",x"95",x"A3",x"90",x"80",x"51",x"48",x"69",x"87",x"B1",
		x"AC",x"8B",x"6E",x"43",x"56",x"72",x"99",x"B6",x"99",x"80",x"51",x"43",x"64",x"80",x"AC",x"AC",
		x"8B",x"6E",x"43",x"4D",x"6E",x"90",x"B1",x"99",x"80",x"5B",x"31",x"22",x"3F",x"64",x"87",x"90",
		x"72",x"48",x"4D",x"6E",x"8B",x"B6",x"A3",x"82",x"60",x"3F",x"5B",x"77",x"A3",x"B1",x"90",x"77",
		x"48",x"48",x"69",x"87",x"87",x"64",x"6E",x"8B",x"80",x"60",x"77",x"95",x"BF",x"CD",x"B6",x"87",
		x"7C",x"99",x"B6",x"E5",x"DB",x"BA",x"95",x"72",x"80",x"9E",x"BA",x"A7",x"82",x"69",x"3A",x"2C",
		x"4D",x"6E",x"7C",x"56",x"5B",x"60",x"43",x"4D",x"60",x"80",x"6E",x"51",x"64",x"5B",x"3F",x"2C",
		x"48",x"77",x"7C",x"60",x"3A",x"3A",x"5B",x"7C",x"9E",x"C4",x"AC",x"90",x"69",x"4D",x"64",x"87",
		x"99",x"80",x"60",x"3A",x"14",x"14",x"3A",x"64",x"82",x"7C",x"51",x"35",x"4D",x"69",x"95",x"A7",
		x"8B",x"69",x"5B",x"69",x"51",x"51",x"69",x"69",x"51",x"56",x"6E",x"8B",x"AC",x"95",x"6E",x"5B",
		x"77",x"82",x"77",x"8B",x"90",x"80",x"64",x"3F",x"43",x"6E",x"87",x"80",x"80",x"80",x"6E",x"60",
		x"35",x"27",x"3F",x"69",x"72",x"56",x"31",x"31",x"56",x"77",x"95",x"B6",x"A7",x"87",x"69",x"4D",
		x"64",x"82",x"99",x"77",x"6E",x"87",x"AC",x"B1",x"8B",x"8B",x"AC",x"A7",x"82",x"90",x"AC",x"9E",
		x"7C",x"60",x"7C",x"9E",x"BA",x"E0",x"E9",x"C4",x"A3",x"80",x"80",x"A3",x"BF",x"E0",x"CD",x"AC",
		x"8B",x"A7",x"BA",x"A7",x"BA",x"BF",x"B1",x"90",x"87",x"AC",x"CD",x"C8",x"A3",x"80",x"8B",x"87",
		x"87",x"87",x"80",x"82",x"87",x"82",x"80",x"82",x"87",x"99",x"9E",x"8B",x"69",x"48",x"51",x"77",
		x"99",x"B6",x"A3",x"7C",x"56",x"43",x"60",x"82",x"A7",x"B1",x"90",x"69",x"48",x"48",x"6E",x"90",
		x"B1",x"A3",x"7C",x"56",x"3F",x"56",x"7C",x"A3",x"AC",x"90",x"69",x"4D",x"27",x"27",x"51",x"6E",
		x"90",x"80",x"60",x"43",x"5B",x"80",x"9E",x"B6",x"8B",x"72",x"4D",x"43",x"6E",x"87",x"AC",x"A3",
		x"80",x"60",x"3F",x"56",x"7C",x"90",x"7C",x"64",x"82",x"90",x"6E",x"69",x"87",x"A3",x"C4",x"BA",
		x"95",x"77",x"82",x"A7",x"BF",x"C4",x"A3",x"82",x"60",x"4D",x"6E",x"90",x"99",x"7C",x"51",x"35",
		x"10",x"19",x"43",x"64",x"56",x"3A",x"48",x"3A",x"2C",x"3F",x"5B",x"6E",x"48",x"48",x"4D",x"3A",
		x"1E",x"22",x"48",x"69",x"60",x"35",x"1E",x"31",x"5B",x"7C",x"9E",x"B1",x"8B",x"6E",x"48",x"43",
		x"6E",x"8B",x"87",x"64",x"3F",x"22",x"01",x"1E",x"43",x"64",x"7C",x"60",x"3A",x"31",x"51",x"77",
		x"99",x"99",x"77",x"51",x"60",x"60",x"48",x"56",x"64",x"5B",x"4D",x"5B",x"72",x"95",x"9E",x"82",
		x"60",x"5B",x"82",x"7C",x"7C",x"90",x"87",x"77",x"56",x"3F",x"51",x"77",x"87",x"80",x"82",x"7C",
		x"6E",x"4D",x"2C",x"2C",x"51",x"77",x"6E",x"4D",x"31",x"3F",x"64",x"80",x"AC",x"BF",x"9E",x"82",
		x"56",x"51",x"72",x"90",x"95",x"72",x"77",x"99",x"BF",x"A7",x"87",x"A3",x"BA",x"99",x"8B",x"AC",
		x"B1",x"95",x"69",x"6E",x"8B",x"AC",x"D7",x"EE",x"E5",x"BA",x"90",x"7C",x"90",x"B6",x"DB",x"E5",
		x"C8",x"99",x"95",x"BA",x"B6",x"B1",x"C4",x"C4",x"A7",x"87",x"99",x"BA",x"D2",x"BF",x"95",x"82",
		x"90",x"8B",x"90",x"87",x"87",x"8B",x"8B",x"82",x"87",x"8B",x"95",x"A3",x"99",x"82",x"64",x"4D",
		x"6E",x"87",x"AC",x"B6",x"90",x"77",x"51",x"56",x"77",x"95",x"B6",x"A3",x"82",x"64",x"48",x"64",
		x"82",x"A3",x"B1",x"90",x"77",x"51",x"4D",x"72",x"8B",x"B1",x"A7",x"82",x"69",x"3F",x"22",x"3F",
		x"5B",x"87",x"95",x"7C",x"56",x"4D",x"72",x"8B",x"B1",x"AC",x"87",x"69",x"48",x"5B",x"7C",x"99",
		x"B6",x"99",x"7C",x"56",x"4D",x"69",x"8B",x"90",x"69",x"6E",x"90",x"87",x"64",x"77",x"90",x"BA",
		x"C4",x"AC",x"87",x"77",x"90",x"B1",x"C4",x"B6",x"95",x"77",x"56",x"5B",x"7C",x"99",x"8B",x"64",
		x"4D",x"27",x"14",x"2C",x"51",x"64",x"3F",x"3A",x"4D",x"31",x"35",x"43",x"6E",x"60",x"3F",x"4D",
		x"4D",x"31",x"19",x"31",x"5B",x"69",x"51",x"2C",x"22",x"4D",x"6E",x"8B",x"B6",x"A3",x"87",x"60",
		x"43",x"5B",x"7C",x"90",x"7C",x"5B",x"3A",x"10",x"10",x"31",x"51",x"80",x"77",x"56",x"35",x"43",
		x"64",x"87",x"9E",x"8B",x"69",x"56",x"64",x"51",x"4D",x"60",x"69",x"51",x"51",x"69",x"8B",x"A7",
		x"9E",x"77",x"5B",x"72",x"8B",x"7C",x"8B",x"95",x"87",x"69",x"43",x"43",x"64",x"8B",x"82",x"82",
		x"82",x"77",x"69",x"43",x"2C",x"43",x"69",x"7C",x"60",x"3A",x"35",x"51",x"7C",x"99",x"BF",x"B6",
		x"90",x"72",x"51",x"64",x"8B",x"9E",x"90",x"9E",x"B6",x"D7",x"E9",x"BF",x"9E",x"7C",x"7C",x"9E",
		x"BA",x"E0",x"D2",x"A7",x"8B",x"99",x"C4",x"DB",x"BA",x"A7",x"B1",x"AC",x"B6",x"B6",x"B1",x"B1",
		x"A7",x"A7",x"B1",x"B6",x"C8",x"BF",x"A3",x"82",x"69",x"87",x"A7",x"C8",x"D7",x"B1",x"90",x"6E",
		x"6E",x"90",x"AC",x"D2",x"C4",x"95",x"80",x"8B",x"B6",x"D2",x"CD",x"C8",x"A7",x"87",x"64",x"5B",
		x"82",x"9E",x"C4",x"BA",x"90",x"77",x"56",x"69",x"90",x"A3",x"8B",x"69",x"43",x"35",x"56",x"7C",
		x"9E",x"9E",x"80",x"56",x"3A",x"43",x"69",x"8B",x"AC",x"C4",x"A7",x"87",x"69",x"56",x"7C",x"7C",
		x"77",x"7C",x"72",x"60",x"60",x"77",x"6E",x"72",x"82",x"8B",x"82",x"69",x"5B",x"64",x"56",x"3F",
		x"35",x"56",x"7C",x"7C",x"77",x"77",x"69",x"5B",x"60",x"7C",x"90",x"7C",x"56",x"35",x"22",x"4D",
		x"69",x"8B",x"90",x"6E",x"4D",x"2C",x"35",x"3A",x"3A",x"48",x"56",x"51",x"35",x"22",x"43",x"69",
		x"82",x"A7",x"AC",x"8B",x"72",x"4D",x"51",x"77",x"95",x"B1",x"9E",x"80",x"60",x"48",x"64",x"82",
		x"A3",x"B1",x"90",x"72",x"51",x"51",x"72",x"90",x"B1",x"A3",x"82",x"64",x"4D",x"60",x"82",x"95",
		x"87",x"8B",x"82",x"80",x"8B",x"99",x"9E",x"87",x"69",x"72",x"95",x"AC",x"A3",x"A7",x"A3",x"95",
		x"77",x"69",x"82",x"AC",x"B1",x"90",x"72",x"48",x"51",x"72",x"95",x"B6",x"A3",x"82",x"60",x"3A",
		x"27",x"43",x"69",x"8B",x"95",x"7C",x"51",x"51",x"72",x"90",x"BA",x"D7",x"CD",x"A3",x"80",x"60",
		x"43",x"64",x"82",x"A7",x"B6",x"8B",x"72",x"4D",x"4D",x"77",x"90",x"B6",x"A7",x"80",x"64",x"43",
		x"60",x"82",x"9E",x"BF",x"DB",x"CD",x"B1",x"82",x"87",x"A7",x"C8",x"D2",x"BA",x"9E",x"77",x"5B",
		x"72",x"8B",x"BA",x"C8",x"A7",x"82",x"7C",x"99",x"BA",x"BF",x"90",x"9E",x"99",x"99",x"A7",x"9E",
		x"9E",x"99",x"95",x"99",x"9E",x"B1",x"B6",x"A3",x"87",x"60",x"64",x"82",x"A3",x"B6",x"9E",x"82",
		x"5B",x"3F",x"5B",x"77",x"A3",x"AC",x"90",x"6E",x"64",x"82",x"A3",x"B1",x"AC",x"9E",x"80",x"5B",
		x"3A",x"51",x"6E",x"99",x"AC",x"8B",x"72",x"43",x"3F",x"60",x"80",x"82",x"64",x"43",x"22",x"31",
		x"51",x"72",x"90",x"7C",x"5B",x"3A",x"27",x"43",x"69",x"82",x"B1",x"AC",x"8B",x"6E",x"43",x"51",
		x"72",x"69",x"6E",x"69",x"5B",x"4D",x"60",x"69",x"64",x"6E",x"7C",x"82",x"72",x"51",x"56",x"5B",
		x"43",x"27",x"35",x"5B",x"72",x"6E",x"6E",x"6E",x"56",x"51",x"60",x"80",x"87",x"64",x"48",x"27",
		x"2C",x"51",x"72",x"90",x"80",x"60",x"3A",x"2C",x"35",x"31",x"3A",x"51",x"56",x"48",x"2C",x"2C",
		x"51",x"6E",x"90",x"B6",x"9E",x"82",x"5B",x"43",x"60",x"7C",x"A7",x"B1",x"90",x"77",x"48",x"4D",
		x"6E",x"8B",x"B6",x"A7",x"82",x"5B",x"43",x"5B",x"82",x"A7",x"B6",x"95",x"72",x"4D",x"4D",x"6E",
		x"95",x"87",x"8B",x"87",x"80",x"82",x"90",x"9E",x"95",x"7C",x"64",x"82",x"AC",x"AC",x"A3",x"A7",
		x"99",x"8B",x"6E",x"77",x"95",x"B6",x"A3",x"80",x"60",x"43",x"64",x"82",x"A7",x"B6",x"90",x"72",
		x"51",x"31",x"35",x"56",x"77",x"95",x"87",x"69",x"4D",x"64",x"87",x"A3",x"C8",x"D7",x"B6",x"95",
		x"77",x"4D",x"51",x"72",x"90",x"BA",x"A7",x"87",x"64",x"43",x"64",x"80",x"A7",x"B6",x"95",x"7C",
		x"4D",x"4D",x"6E",x"90",x"B6",x"D2",x"DB",x"C8",x"9E",x"82",x"95",x"BF",x"D7",x"CD",x"B6",x"8B",
		x"69",x"60",x"80",x"A7",x"C8",x"C4",x"9E",x"77",x"87",x"A7",x"C4",x"AC",x"95",x"A3",x"99",x"A3",
		x"A3",x"A3",x"A3",x"99",x"99",x"9E",x"A7",x"BA",x"B6",x"99",x"77",x"60",x"72",x"95",x"B6",x"B1",
		x"99",x"72",x"4D",x"48",x"69",x"8B",x"B1",x"AC",x"82",x"64",x"72",x"90",x"B1",x"B1",x"AC",x"95",
		x"72",x"4D",x"3F",x"60",x"82",x"A7",x"A7",x"87",x"60",x"3F",x"48",x"72",x"90",x"7C",x"60",x"35",
		x"22",x"3F",x"69",x"8B",x"90",x"72",x"48",x"2C",x"31",x"56",x"7C",x"99",x"BA",x"A3",x"7C",x"60",
		x"43",x"6E",x"72",x"69",x"72",x"64",x"56",x"51",x"69",x"69",x"69",x"77",x"82",x"80",x"64",x"51",
		x"5B",x"56",x"35",x"27",x"4D",x"72",x"72",x"6E",x"72",x"64",x"56",x"56",x"72",x"8B",x"80",x"56",
		x"31",x"1E",x"3A",x"64",x"87",x"90",x"72",x"4D",x"2C",x"31",x"35",x"35",x"43",x"56",x"51",x"35",
		x"22",x"35",x"64",x"82",x"A3",x"B6",x"8B",x"72",x"4D",x"4D",x"77",x"90",x"B6",x"A7",x"80",x"64",
		x"43",x"60",x"82",x"A3",x"B6",x"95",x"77",x"51",x"48",x"72",x"8B",x"B6",x"AC",x"82",x"69",x"48",
		x"5B",x"82",x"95",x"87",x"8B",x"82",x"82",x"87",x"99",x"9E",x"8B",x"72",x"72",x"90",x"B1",x"A7",
		x"A7",x"A3",x"99",x"80",x"69",x"82",x"A3",x"B6",x"95",x"77",x"51",x"51",x"72",x"90",x"B1",x"A7",
		x"87",x"69",x"43",x"27",x"43",x"60",x"8B",x"99",x"80",x"60",x"51",x"77",x"90",x"B6",x"DB",x"CD",
		x"AC",x"87",x"64",x"48",x"5B",x"82",x"A7",x"BA",x"9E",x"77",x"51",x"4D",x"6E",x"90",x"B6",x"AC",
		x"82",x"69",x"48",x"60",x"82",x"9E",x"BF",x"DB",x"D7",x"BA",x"95",x"8B",x"A7",x"CD",x"D7",x"BF",
		x"A3",x"80",x"64",x"72",x"90",x"B1",x"C8",x"B1",x"8B",x"7C",x"99",x"BF",x"C4",x"9E",x"9E",x"9E",
		x"99",x"A7",x"A3",x"A3",x"9E",x"99",x"99",x"A3",x"AC",x"BA",x"A7",x"90",x"6E",x"64",x"82",x"A3",
		x"B6",x"A7",x"87",x"69",x"48",x"5B",x"7C",x"99",x"B1",x"99",x"77",x"64",x"82",x"A7",x"B6",x"B1",
		x"A3",x"82",x"64",x"43",x"51",x"72",x"90",x"AC",x"95",x"77",x"51",x"43",x"60",x"82",x"8B",x"69",
		x"4D",x"27",x"2C",x"56",x"72",x"95",x"82",x"60",x"3F",x"22",x"43",x"69",x"82",x"A7",x"B1",x"90",
		x"77",x"51",x"51",x"77",x"6E",x"6E",x"6E",x"60",x"4D",x"60",x"6E",x"64",x"6E",x"80",x"82",x"77",
		x"5B",x"56",x"60",x"48",x"31",x"35",x"5B",x"77",x"72",x"72",x"6E",x"60",x"56",x"60",x"7C",x"8B",
		x"69",x"4D",x"27",x"27",x"51",x"6E",x"90",x"82",x"64",x"43",x"27",x"35",x"35",x"3A",x"4D",x"56",
		x"4D",x"2C",x"27",x"4D",x"6E",x"8B",x"AC",x"A7",x"82",x"69",x"48",x"60",x"7C",x"A3",x"B6",x"95",
		x"7C",x"4D",x"4D",x"6E",x"8B",x"B6",x"A7",x"8B",x"69",x"43",x"5B",x"7C",x"A3",x"BA",x"99",x"80",
		x"51",x"4D",x"69",x"8B",x"8B",x"8B",x"8B",x"82",x"82",x"90",x"9E",x"99",x"7C",x"69",x"7C",x"A7",
		x"B1",x"A3",x"AC",x"9E",x"90",x"72",x"72",x"95",x"B6",x"AC",x"87",x"64",x"48",x"60",x"80",x"A7",
		x"B6",x"9E",x"77",x"56",x"35",x"31",x"5B",x"77",x"99",x"90",x"69",x"51",x"5B",x"82",x"A3",x"C8",
		x"DB",x"BF",x"99",x"7C",x"56",x"51",x"72",x"90",x"B1",x"AC",x"8B",x"6E",x"4D",x"48",x"48",x"43",
		x"48",x"51",x"5B",x"51",x"4D",x"5B",x"5B",x"51",x"56",x"60",x"60",x"56",x"43",x"4D",x"60",x"82",
		x"A7",x"BA",x"A3",x"80",x"5B",x"4D",x"6E",x"90",x"B6",x"B6",x"90",x"6E",x"77",x"99",x"8B",x"95",
		x"A3",x"99",x"7C",x"6E",x"82",x"A7",x"B1",x"95",x"72",x"6E",x"77",x"77",x"7C",x"6E",x"72",x"7C",
		x"77",x"72",x"77",x"7C",x"87",x"95",x"82",x"6E",x"48",x"43",x"69",x"82",x"A7",x"A3",x"80",x"60",
		x"43",x"56",x"77",x"95",x"AC",x"90",x"77",x"51",x"48",x"69",x"87",x"B1",x"A7",x"87",x"64",x"3F",
		x"56",x"77",x"9E",x"B6",x"99",x"7C",x"56",x"31",x"27",x"48",x"72",x"95",x"90",x"72",x"4D",x"5B",
		x"7C",x"9E",x"BF",x"A3",x"87",x"5B",x"4D",x"6E",x"87",x"B6",x"B6",x"95",x"77",x"4D",x"5B",x"77",
		x"99",x"8B",x"6E",x"80",x"99",x"82",x"6E",x"87",x"AC",x"D2",x"D7",x"BA",x"8B",x"90",x"AC",x"CD",
		x"F7",x"E0",x"C4",x"99",x"7C",x"90",x"B6",x"C8",x"AC",x"8B",x"6E",x"43",x"43",x"64",x"82",x"82",
		x"60",x"6E",x"69",x"56",x"60",x"77",x"90",x"77",x"64",x"77",x"64",x"48",x"3F",x"60",x"87",x"82",
		x"64",x"48",x"4D",x"72",x"8B",x"B6",x"D2",x"B6",x"99",x"6E",x"60",x"7C",x"9E",x"A7",x"87",x"69",
		x"48",x"1E",x"2C",x"4D",x"77",x"95",x"80",x"60",x"48",x"64",x"80",x"A3",x"B1",x"95",x"72",x"6E",
		x"77",x"60",x"64",x"77",x"72",x"60",x"69",x"80",x"A3",x"B6",x"A3",x"77",x"69",x"8B",x"90",x"87",
		x"9E",x"9E",x"8B",x"69",x"4D",x"51",x"7C",x"99",x"87",x"90",x"87",x"7C",x"69",x"43",x"35",x"56",
		x"7C",x"80",x"5B",x"3A",x"3F",x"64",x"8B",x"A7",x"C4",x"AC",x"8B",x"6E",x"5B",x"77",x"99",x"A7",
		x"7C",x"80",x"99",x"BF",x"BA",x"90",x"9E",x"BF",x"AC",x"8B",x"A7",x"BA",x"A3",x"80",x"6E",x"90",
		x"B1",x"CD",x"EE",x"EE",x"C8",x"A7",x"87",x"90",x"B1",x"D2",x"EE",x"D2",x"B1",x"95",x"BA",x"C4",
		x"B1",x"C8",x"C8",x"B6",x"95",x"95",x"BF",x"D7",x"CD",x"A3",x"87",x"95",x"8B",x"90",x"8B",x"87",
		x"8B",x"90",x"87",x"87",x"8B",x"95",x"A7",x"A3",x"8B",x"6E",x"51",x"60",x"82",x"AC",x"BF",x"A3",
		x"80",x"56",x"4D",x"6E",x"90",x"B6",x"B1",x"90",x"69",x"4D",x"56",x"7C",x"A3",x"BA",x"A3",x"7C",
		x"56",x"48",x"64",x"8B",x"B1",x"B1",x"90",x"69",x"4D",x"27",x"35",x"60",x"7C",x"99",x"82",x"60",
		x"4D",x"64",x"87",x"AC",x"B6",x"95",x"72",x"4D",x"51",x"72",x"99",x"B6",x"A7",x"82",x"5B",x"48",
		x"5B",x"87",x"99",x"77",x"69",x"8B",x"90",x"6E",x"6E",x"90",x"B1",x"C8",x"BA",x"90",x"77",x"82",
		x"AC",x"C8",x"BF",x"A7",x"80",x"5B",x"51",x"72",x"99",x"95",x"77",x"56",x"2C",x"14",x"1E",x"4D",
		x"69",x"4D",x"3A",x"4D",x"35",x"31",x"43",x"64",x"69",x"48",x"4D",x"4D",x"3A",x"1E",x"2C",x"56",
		x"6E",x"5B",x"31",x"22",x"3A",x"69",x"82",x"A7",x"B1",x"87",x"6E",x"48",x"51",x"77",x"90",x"87",
		x"60",x"3F",x"1E",x"06",x"2C",x"4D",x"72",x"80",x"5B",x"3A",x"35",x"5B",x"82",x"9E",x"95",x"72",
		x"51",x"64",x"5B",x"4D",x"5B",x"69",x"5B",x"51",x"64",x"7C",x"9E",x"9E",x"80",x"5B",x"69",x"8B",
		x"7C",x"82",x"95",x"87",x"77",x"51",x"3F",x"5B",x"82",x"87",x"80",x"82",x"7C",x"6E",x"48",x"2C",
		x"31",x"60",x"7C",x"69",x"48",x"31",x"4D",x"6E",x"8B",x"B6",x"BA",x"99",x"7C",x"51",x"5B",x"7C",
		x"99",x"90",x"72",x"80",x"A7",x"BF",x"A3",x"8B",x"AC",x"BA",x"95",x"8B",x"B6",x"B1",x"90",x"72",
		x"72",x"95",x"B1",x"DB",x"F7",x"DB",x"BA",x"90",x"80",x"99",x"B6",x"E5",x"E5",x"C4",x"9E",x"99",
		x"C4",x"B6",x"B6",x"C8",x"BF",x"A7",x"8B",x"9E",x"C4",x"D7",x"BA",x"8B",x"87",x"90",x"8B",x"90",
		x"87",x"87",x"8B",x"8B",x"82",x"87",x"8B",x"99",x"A7",x"99",x"80",x"60",x"4D",x"72",x"90",x"B1",
		x"B1",x"8B",x"72",x"4D",x"60",x"80",x"9E",x"B6",x"9E",x"80",x"5B",x"4D",x"6E",x"87",x"AC",x"B1",
		x"8B",x"72",x"4D",x"56",x"77",x"95",x"B1",x"9E",x"7C",x"60",x"35",x"27",x"48",x"64",x"90",x"90",
		x"77",x"51",x"51",x"77",x"95",x"B6",x"A3",x"82",x"64",x"48",x"64",x"82",x"A3",x"B1",x"90",x"77",
		x"51",x"51",x"6E",x"90",x"8B",x"64",x"77",x"95",x"80",x"64",x"80",x"99",x"BF",x"C4",x"A7",x"82",
		x"7C",x"95",x"B6",x"C4",x"AC",x"90",x"72",x"51",x"60",x"82",x"9E",x"82",x"60",x"43",x"1E",x"14",
		x"31",x"5B",x"64",x"3A",x"43",x"48",x"31",x"3A",x"4D",x"72",x"56",x"3F",x"51",x"48",x"27",x"19",
		x"3A",x"60",x"69",x"48",x"27",x"27",x"51",x"72",x"90",x"B1",x"9E",x"80",x"60",x"48",x"60",x"82",
		x"95",x"72",x"51",x"35",x"14",x"14",x"35",x"56",x"7C",x"72",x"51",x"31",x"48",x"6E",x"8B",x"A3",
		x"87",x"60",x"5B",x"69",x"4D",x"51",x"64",x"69",x"4D",x"5B",x"69",x"8B",x"AC",x"95",x"77",x"5B",
		x"7C",x"87",x"77",x"90",x"90",x"82",x"69",x"3F",x"48",x"69",x"87",x"82",x"82",x"82",x"72",x"64",
		x"3A",x"31",x"48",x"72",x"7C",x"56",x"35",x"35",x"5B",x"82",x"9E",x"C4",x"AC",x"87",x"6E",x"4D",
		x"6E",x"90",x"A3",x"80",x"77",x"90",x"B6",x"BA",x"90",x"99",x"BA",x"AC",x"87",x"9E",x"BA",x"A3",
		x"7C",x"6E",x"80",x"A7",x"C8",x"E9",x"F3",x"C8",x"A7",x"82",x"87",x"B1",x"C8",x"EE",x"D7",x"AC",
		x"95",x"AC",x"BF",x"B1",x"C4",x"C8",x"B6",x"95",x"90",x"B1",x"D7",x"CD",x"A7",x"8B",x"90",x"8B",
		x"90",x"8B",x"87",x"8B",x"90",x"87",x"82",x"8B",x"90",x"A7",x"A3",x"90",x"77",x"4D",x"60",x"7C",
		x"A3",x"BF",x"A3",x"87",x"5B",x"4D",x"6E",x"87",x"B6",x"B6",x"95",x"77",x"48",x"56",x"77",x"99",
		x"BA",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B1",x"95",x"77",x"4D",x"2C",x"31",x"56",x"7C",
		x"99",x"8B",x"64",x"48",x"64",x"80",x"A7",x"BA",x"99",x"7C",x"4D",x"51",x"6E",x"8B",x"BA",x"A7",
		x"8B",x"64",x"43",x"5B",x"7C",x"95",x"7C",x"69",x"82",x"90",x"72",x"69",x"87",x"B1",x"C8",x"BF",
		x"99",x"72",x"82",x"A3",x"C4",x"BF",x"A7",x"87",x"60",x"51",x"6E",x"95",x"99",x"77",x"56",x"31",
		x"14",x"1E",x"48",x"69",x"51",x"35",x"48",x"3A",x"31",x"3F",x"64",x"6E",x"48",x"48",x"4D",x"3F",
		x"1E",x"27",x"56",x"6E",x"64",x"3A",x"22",x"3A",x"60",x"82",x"A7",x"B1",x"95",x"6E",x"4D",x"4D",
		x"6E",x"95",x"87",x"69",x"48",x"1E",x"0B",x"1E",x"48",x"72",x"80",x"69",x"3A",x"35",x"5B",x"77",
		x"A3",x"99",x"7C",x"5B",x"64",x"60",x"4D",x"5B",x"6E",x"60",x"51",x"64",x"7C",x"9E",x"A7",x"82",
		x"64",x"64",x"82",x"80",x"80",x"95",x"8B",x"77",x"56",x"3F",x"56",x"80",x"8B",x"80",x"87",x"7C",
		x"72",x"51",x"2C",x"35",x"56",x"77",x"6E",x"4D",x"31",x"48",x"6E",x"87",x"AC",x"BF",x"9E",x"80",
		x"60",x"5B",x"7C",x"99",x"99",x"95",x"AC",x"C4",x"E5",x"CD",x"AC",x"8B",x"77",x"90",x"AC",x"D2",
		x"DB",x"BA",x"95",x"90",x"B6",x"D7",x"CD",x"A7",x"B6",x"AC",x"B1",x"B6",x"B1",x"B6",x"AC",x"A7",
		x"AC",x"B1",x"BF",x"C4",x"B1",x"95",x"72",x"7C",x"99",x"BA",x"D7",x"BF",x"9E",x"80",x"69",x"82",
		x"9E",x"C4",x"CD",x"AC",x"87",x"82",x"AC",x"C8",x"D2",x"CD",x"B6",x"95",x"6E",x"56",x"77",x"90",
		x"BA",x"C4",x"A3",x"82",x"56",x"60",x"80",x"9E",x"95",x"72",x"56",x"35",x"4D",x"6E",x"90",x"A3",
		x"87",x"69",x"43",x"3A",x"60",x"7C",x"9E",x"C4",x"B6",x"95",x"72",x"51",x"69",x"82",x"77",x"7C",
		x"77",x"64",x"5B",x"72",x"72",x"6E",x"7C",x"87",x"8B",x"77",x"56",x"64",x"64",x"43",x"31",x"43",
		x"6E",x"7C",x"72",x"77",x"72",x"5B",x"5B",x"6E",x"87",x"87",x"64",x"48",x"27",x"3A",x"5B",x"80",
		x"95",x"7C",x"60",x"3A",x"31",x"3A",x"35",x"43",x"56",x"56",x"43",x"2C",x"31",x"5B",x"77",x"9E",
		x"B6",x"99",x"80",x"51",x"48",x"69",x"82",x"B1",x"AC",x"8B",x"6E",x"43",x"56",x"72",x"99",x"B6",
		x"9E",x"82",x"56",x"43",x"64",x"80",x"AC",x"B1",x"90",x"72",x"48",x"51",x"72",x"90",x"87",x"8B",
		x"87",x"80",x"82",x"90",x"9E",x"90",x"72",x"69",x"82",x"AC",x"A7",x"A3",x"A7",x"95",x"87",x"64",
		x"77",x"9E",x"B6",x"9E",x"7C",x"56",x"43",x"64",x"87",x"AC",x"B1",x"90",x"69",x"4D",x"27",x"35",
		x"5B",x"7C",x"99",x"82",x"5B",x"48",x"69",x"8B",x"A7",x"CD",x"CD",x"AC",x"8B",x"6E",x"43",x"56",
		x"72",x"99",x"B6",x"9E",x"80",x"56",x"43",x"64",x"80",x"AC",x"B1",x"90",x"72",x"43",x"51",x"72",
		x"95",x"BA",x"D7",x"D7",x"BA",x"95",x"82",x"95",x"C4",x"D2",x"C8",x"A7",x"80",x"60",x"64",x"82",
		x"AC",x"C8",x"BA",x"90",x"72",x"8B",x"AC",x"C4",x"9E",x"95",x"9E",x"95",x"A3",x"9E",x"9E",x"9E",
		x"95",x"95",x"99",x"A7",x"B6",x"AC",x"90",x"6E",x"5B",x"72",x"99",x"B1",x"AC",x"8B",x"69",x"43",
		x"48",x"6E",x"95",x"AC",x"A3",x"7C",x"60",x"77",x"95",x"B1",x"AC",x"A7",x"8B",x"64",x"43",x"3F",
		x"64",x"87",x"A7",x"9E",x"7C",x"51",x"3A",x"4D",x"77",x"8B",x"72",x"56",x"27",x"22",x"43",x"64",
		x"90",x"87",x"69",x"48",x"22",x"35",x"56",x"7C",x"9E",x"B6",x"9E",x"77",x"51",x"43",x"69",x"6E",
		x"69",x"6E",x"60",x"4D",x"56",x"69",x"64",x"69",x"77",x"82",x"7C",x"5B",x"4D",x"5B",x"4D",x"2C",
		x"27",x"48",x"77",x"6E",x"6E",x"6E",x"60",x"51",x"56",x"77",x"8B",x"72",x"56",x"2C",x"1E",x"3F",
		x"60",x"8B",x"8B",x"69",x"43",x"27",x"31",x"35",x"35",x"48",x"56",x"4D",x"31",x"22",x"3F",x"69",
		x"87",x"A7",x"AC",x"82",x"69",x"43",x"51",x"7C",x"95",x"B6",x"99",x"7C",x"5B",x"43",x"64",x"82",
		x"A7",x"B1",x"8B",x"6E",x"48",x"4D",x"77",x"90",x"B6",x"A3",x"80",x"60",x"43",x"60",x"87",x"90",
		x"87",x"8B",x"80",x"80",x"87",x"9E",x"99",x"87",x"6E",x"77",x"99",x"B1",x"A7",x"A7",x"9E",x"95",
		x"77",x"69",x"87",x"A7",x"B1",x"8B",x"72",x"4D",x"56",x"77",x"95",x"B1",x"A3",x"80",x"64",x"3A",
		x"27",x"48",x"69",x"90",x"95",x"77",x"56",x"56",x"7C",x"95",x"BA",x"DB",x"C4",x"A3",x"80",x"5B",
		x"48",x"64",x"87",x"AC",x"B6",x"95",x"72",x"4D",x"51",x"72",x"99",x"B6",x"A7",x"82",x"60",x"48",
		x"60",x"82",x"A7",x"C4",x"DB",x"CD",x"B1",x"8B",x"87",x"B1",x"CD",x"D7",x"BF",x"99",x"7C",x"5B",
		x"77",x"95",x"BA",x"CD",x"A7",x"82",x"7C",x"99",x"BF",x"BF",x"95",x"9E",x"9E",x"9E",x"A7",x"A3",
		x"A3",x"9E",x"95",x"99",x"A3",x"B1",x"BA",x"A3",x"87",x"64",x"64",x"8B",x"A7",x"B6",x"A3",x"80",
		x"60",x"43",x"60",x"80",x"A3",x"AC",x"90",x"6E",x"64",x"8B",x"A7",x"B1",x"AC",x"99",x"7C",x"5B",
		x"3F",x"56",x"77",x"95",x"AC",x"8B",x"72",x"48",x"43",x"64",x"87",x"87",x"60",x"43",x"1E",x"31",
		x"5B",x"77",x"95",x"7C",x"5B",x"35",x"27",x"48",x"6E",x"87",x"AC",x"AC",x"87",x"6E",x"48",x"56",
		x"77",x"69",x"6E",x"69",x"5B",x"4D",x"64",x"69",x"64",x"6E",x"80",x"82",x"72",x"56",x"56",x"5B",
		x"43",x"2C",x"3A",x"64",x"77",x"6E",x"72",x"6E",x"5B",x"56",x"64",x"82",x"87",x"60",x"43",x"22",
		x"2C",x"56",x"72",x"95",x"7C",x"5B",x"3A",x"27",x"35",x"35",x"3F",x"4D",x"56",x"48",x"27",x"2C",
		x"56",x"72",x"95",x"B1",x"9E",x"80",x"60",x"48",x"64",x"82",x"A3",x"B1",x"90",x"72",x"4D",x"51",
		x"72",x"90",x"B1",x"A3",x"82",x"64",x"48",x"60",x"80",x"A3",x"B6",x"95",x"77",x"51",x"51",x"6E",
		x"90",x"90",x"8B",x"8B",x"80",x"82",x"95",x"9E",x"99",x"77",x"69",x"82",x"A7",x"AC",x"A7",x"AC",
		x"9E",x"8B",x"6E",x"72",x"95",x"BA",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",x"6E",
		x"51",x"2C",x"35",x"60",x"7C",x"9E",x"87",x"64",x"4D",x"64",x"8B",x"AC",x"CD",x"DB",x"B6",x"90",
		x"77",x"51",x"56",x"77",x"95",x"B6",x"A7",x"82",x"64",x"4D",x"64",x"82",x"A7",x"B6",x"95",x"77",
		x"51",x"51",x"72",x"90",x"B1",x"DB",x"DB",x"C8",x"9E",x"82",x"99",x"BA",x"D7",x"CD",x"B1",x"90",
		x"64",x"64",x"82",x"A3",x"CD",x"BF",x"9E",x"7C",x"8B",x"AC",x"C8",x"A7",x"95",x"A3",x"95",x"A7",
		x"A3",x"A3",x"A3",x"99",x"99",x"9E",x"A7",x"BA",x"B1",x"9E",x"77",x"5B",x"77",x"95",x"B1",x"B1",
		x"95",x"77",x"48",x"4D",x"69",x"8B",x"B1",x"A3",x"82",x"69",x"77",x"95",x"B1",x"B1",x"AC",x"90",
		x"72",x"48",x"3F",x"64",x"80",x"AC",x"A3",x"82",x"60",x"3A",x"51",x"72",x"8B",x"77",x"56",x"35",
		x"22",x"43",x"64",x"87",x"8B",x"6E",x"4D",x"2C",x"31",x"56",x"77",x"99",x"BA",x"9E",x"82",x"5B",
		x"43",x"69",x"72",x"6E",x"6E",x"69",x"56",x"56",x"69",x"69",x"69",x"77",x"82",x"82",x"60",x"4D",
		x"60",x"56",x"35",x"27",x"48",x"6E",x"72",x"6E",x"72",x"64",x"56",x"56",x"72",x"8B",x"77",x"5B",
		x"31",x"1E",x"43",x"60",x"8B",x"8B",x"72",x"51",x"27",x"35",x"35",x"35",x"48",x"56",x"56",x"35",
		x"22",x"3F",x"60",x"82",x"A7",x"B1",x"90",x"6E",x"4D",x"4D",x"72",x"95",x"B6",x"A7",x"82",x"5B",
		x"48",x"5B",x"82",x"A7",x"B6",x"99",x"72",x"51",x"4D",x"6E",x"95",x"B6",x"AC",x"87",x"60",x"48",
		x"56",x"82",x"95",x"87",x"90",x"82",x"82",x"87",x"99",x"9E",x"8B",x"6E",x"72",x"99",x"B1",x"A7",
		x"A7",x"A3",x"95",x"80",x"6E",x"82",x"A7",x"B6",x"90",x"77",x"4D",x"4D",x"77",x"90",x"B6",x"A7",
		x"82",x"64",x"43",x"2C",x"43",x"64",x"87",x"95",x"7C",x"56",x"51",x"7C",x"95",x"B6",x"D7",x"CD",
		x"A7",x"8B",x"64",x"48",x"64",x"80",x"A7",x"BA",x"99",x"7C",x"51",x"48",x"48",x"48",x"4D",x"4D",
		x"4D",x"51",x"51",x"51",x"51",x"56",x"56",x"56",x"56",x"5B",x"5B",x"5B",x"5B",x"5B",x"60",x"60",
		x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"64",x"69",x"69",x"69",x"69",x"69",x"69",x"6E",
		x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"77",
		x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"82",x"82",x"87",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",
		x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"7C",x"80",
		x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"80",x"80",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"7C",x"7C",
		x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"80",x"80",
		x"80",x"80",x"7C",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"77",x"72",
		x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"77",x"77",x"7C",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",
		x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"80",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",
		x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"82",x"80",x"77",
		x"80",x"82",x"80",x"77",x"80",x"82",x"7C",x"77",x"82",x"82",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"80",
		x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"72",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"7C",x"7C",
		x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",
		x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"80",x"82",
		x"80",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"77",x"80",
		x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"72",
		x"77",x"80",x"87",x"7C",x"77",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"82",x"80",x"77",x"7C",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"72",x"7C",x"7C",x"7C",x"7C",x"77",
		x"77",x"7C",x"7C",x"7C",x"7C",x"77",x"7C",x"80",x"77",x"77",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",
		x"80",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"7C",x"82",x"82",x"80",x"7C",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"82",
		x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"8B",x"82",x"8B",x"8B",x"8B",x"90",x"90",x"90",x"95",
		x"95",x"95",x"95",x"95",x"90",x"95",x"99",x"95",x"90",x"87",x"8B",x"87",x"80",x"7C",x"80",x"7C",
		x"72",x"72",x"72",x"6E",x"64",x"69",x"64",x"60",x"51",x"43",x"4D",x"48",x"51",x"56",x"51",x"51",
		x"51",x"51",x"56",x"64",x"60",x"64",x"69",x"69",x"6E",x"72",x"72",x"72",x"80",x"80",x"7C",x"82",
		x"8B",x"8B",x"87",x"90",x"99",x"95",x"95",x"99",x"99",x"90",x"95",x"99",x"95",x"8B",x"87",x"8B",
		x"82",x"7C",x"7C",x"80",x"77",x"77",x"77",x"6E",x"72",x"6E",x"69",x"6E",x"77",x"7C",x"72",x"6E",
		x"7C",x"7C",x"7C",x"80",x"87",x"87",x"7C",x"80",x"87",x"82",x"87",x"8B",x"87",x"82",x"82",x"80",
		x"7C",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"7C",x"80",x"82",x"82",x"82",x"80",x"87",
		x"87",x"87",x"87",x"87",x"87",x"82",x"80",x"87",x"82",x"87",x"8B",x"87",x"82",x"7C",x"82",x"87",
		x"80",x"7C",x"80",x"7C",x"77",x"77",x"7C",x"77",x"77",x"80",x"80",x"77",x"7C",x"77",x"72",x"77",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"72",x"72",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"72",
		x"77",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",
		x"80",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"80",x"80",x"80",x"80",x"77",x"7C",
		x"77",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"7C",
		x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"80",x"77",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",
		x"77",x"80",x"7C",x"77",x"77",x"77",x"77",x"77",x"7C",x"82",x"87",x"7C",x"7C",x"80",x"77",x"77",
		x"80",x"87",x"82",x"82",x"80",x"77",x"77",x"7C",x"87",x"95",x"7C",x"80",x"80",x"7C",x"82",x"80",
		x"82",x"87",x"87",x"80",x"77",x"80",x"82",x"80",x"87",x"87",x"82",x"7C",x"7C",x"7C",x"7C",x"80",
		x"80",x"82",x"80",x"7C",x"7C",x"77",x"72",x"77",x"80",x"82",x"7C",x"7C",x"7C",x"72",x"77",x"7C",
		x"82",x"80",x"77",x"7C",x"7C",x"72",x"77",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",
		x"80",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"72",x"7C",x"7C",x"7C",x"7C",x"77",x"77",
		x"77",x"77",x"80",x"7C",x"80",x"7C",x"80",x"7C",x"77",x"7C",x"80",x"7C",x"80",x"77",x"77",x"7C",
		x"82",x"82",x"7C",x"80",x"87",x"82",x"7C",x"80",x"87",x"82",x"82",x"82",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"82",x"80",x"82",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"82",
		x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"80",
		x"72",x"72",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"72",x"77",x"80",x"77",x"72",x"7C",x"80",x"7C",
		x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"7C",x"77",x"77",x"80",x"7C",x"80",x"82",x"80",x"77",x"72",
		x"7C",x"80",x"7C",x"82",x"82",x"7C",x"80",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",
		x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"80",x"82",x"80",
		x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"82",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",
		x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"77",
		x"72",x"7C",x"80",x"7C",x"80",x"82",x"80",x"77",x"77",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"7C",x"72",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"7C",x"80",x"7C",x"80",x"82",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"80",x"80",x"80",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"80",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",
		x"80",x"80",x"7C",x"7C",x"80",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"77",x"80",x"82",x"7C",x"7C",x"80",
		x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"77",x"7C",x"82",x"7C",
		x"77",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"77",x"7C",x"82",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",
		x"82",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",
		x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",
		x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",
		x"82",x"82",x"7C",x"7C",x"80",x"87",x"87",x"7C",x"80",x"87",x"82",x"7C",x"82",x"87",x"82",x"77",
		x"69",x"7C",x"95",x"B1",x"D7",x"D7",x"B1",x"95",x"72",x"7C",x"99",x"BF",x"DB",x"BF",x"9E",x"82",
		x"A7",x"AC",x"9E",x"B6",x"B6",x"A3",x"87",x"87",x"A7",x"C8",x"BA",x"8B",x"7C",x"82",x"82",x"82",
		x"80",x"7C",x"82",x"82",x"7C",x"7C",x"82",x"87",x"99",x"95",x"80",x"64",x"43",x"5B",x"80",x"99",
		x"B6",x"90",x"72",x"51",x"43",x"6E",x"87",x"AC",x"A7",x"82",x"64",x"43",x"51",x"7C",x"95",x"B6",
		x"95",x"77",x"51",x"3F",x"69",x"82",x"A7",x"AC",x"82",x"69",x"48",x"27",x"31",x"56",x"77",x"90",
		x"80",x"5B",x"43",x"64",x"82",x"A7",x"B1",x"8B",x"6E",x"48",x"4D",x"77",x"90",x"B6",x"9E",x"7C",
		x"60",x"43",x"60",x"82",x"95",x"77",x"69",x"87",x"90",x"6E",x"6E",x"8B",x"AC",x"CD",x"BF",x"99",
		x"7C",x"90",x"B6",x"D2",x"E9",x"BF",x"A3",x"7C",x"72",x"95",x"B6",x"B6",x"90",x"6E",x"4D",x"2C",
		x"3F",x"69",x"80",x"69",x"51",x"64",x"51",x"48",x"5B",x"7C",x"80",x"5B",x"60",x"60",x"4D",x"31",
		x"3F",x"64",x"80",x"6E",x"3F",x"31",x"48",x"77",x"90",x"B6",x"BF",x"95",x"7C",x"56",x"5B",x"80",
		x"99",x"90",x"6E",x"48",x"27",x"10",x"31",x"51",x"77",x"80",x"64",x"3F",x"3F",x"69",x"82",x"A7",
		x"99",x"72",x"5B",x"69",x"60",x"4D",x"60",x"6E",x"5B",x"51",x"64",x"7C",x"AC",x"A3",x"82",x"64",
		x"6E",x"8B",x"7C",x"82",x"95",x"87",x"7C",x"4D",x"3F",x"5B",x"80",x"82",x"80",x"82",x"77",x"69",
		x"48",x"27",x"35",x"64",x"77",x"6E",x"3F",x"2C",x"48",x"69",x"90",x"B6",x"BA",x"99",x"72",x"51",
		x"56",x"7C",x"9E",x"8B",x"6E",x"80",x"A7",x"BA",x"A3",x"8B",x"A7",x"B6",x"95",x"8B",x"AC",x"B1",
		x"8B",x"64",x"72",x"90",x"B1",x"DB",x"EE",x"DB",x"B1",x"8B",x"7C",x"95",x"BA",x"DB",x"E0",x"BF",
		x"95",x"95",x"BF",x"B1",x"B6",x"C4",x"BF",x"9E",x"87",x"99",x"BF",x"CD",x"B6",x"8B",x"82",x"8B",
		x"87",x"8B",x"82",x"82",x"87",x"87",x"80",x"82",x"87",x"95",x"A3",x"95",x"80",x"5B",x"4D",x"6E",
		x"87",x"AC",x"AC",x"8B",x"6E",x"4D",x"56",x"77",x"95",x"B1",x"99",x"7C",x"5B",x"48",x"64",x"82",
		x"A7",x"AC",x"87",x"6E",x"48",x"51",x"72",x"90",x"AC",x"9E",x"7C",x"60",x"35",x"22",x"43",x"60",
		x"8B",x"8B",x"72",x"4D",x"4D",x"72",x"90",x"B6",x"9E",x"82",x"5B",x"43",x"60",x"7C",x"A7",x"B1",
		x"90",x"72",x"43",x"4D",x"69",x"8B",x"82",x"64",x"72",x"90",x"7C",x"60",x"77",x"99",x"BF",x"BF",
		x"A3",x"77",x"77",x"90",x"B1",x"C4",x"AC",x"90",x"69",x"48",x"5B",x"80",x"95",x"82",x"60",x"43",
		x"14",x"10",x"31",x"51",x"5B",x"35",x"3F",x"43",x"2C",x"35",x"48",x"69",x"51",x"3F",x"4D",x"43",
		x"27",x"19",x"35",x"64",x"69",x"48",x"27",x"27",x"4D",x"6E",x"90",x"B1",x"99",x"80",x"56",x"3F",
		x"5B",x"80",x"8B",x"72",x"51",x"31",x"06",x"10",x"31",x"56",x"80",x"6E",x"4D",x"31",x"48",x"69",
		x"8B",x"9E",x"82",x"60",x"56",x"64",x"4D",x"4D",x"60",x"64",x"4D",x"56",x"69",x"90",x"A7",x"95",
		x"6E",x"56",x"77",x"87",x"7C",x"8B",x"90",x"82",x"60",x"3F",x"43",x"69",x"8B",x"80",x"82",x"80",
		x"72",x"60",x"3A",x"2C",x"43",x"6E",x"7C",x"56",x"35",x"35",x"56",x"80",x"99",x"BF",x"AC",x"87",
		x"6E",x"4D",x"69",x"8B",x"9E",x"80",x"77",x"90",x"B6",x"BA",x"90",x"95",x"B6",x"AC",x"87",x"99",
		x"B6",x"A3",x"7C",x"69",x"82",x"A7",x"C4",x"E5",x"EE",x"C8",x"A7",x"82",x"87",x"AC",x"C8",x"E9",
		x"D2",x"B1",x"90",x"B1",x"BF",x"AC",x"BF",x"C4",x"B6",x"95",x"8B",x"B6",x"D2",x"CD",x"A3",x"82",
		x"90",x"8B",x"8B",x"8B",x"82",x"8B",x"8B",x"87",x"82",x"8B",x"90",x"A3",x"A3",x"90",x"6E",x"4D",
		x"5B",x"80",x"A3",x"BA",x"A7",x"80",x"5B",x"4D",x"69",x"8B",x"B1",x"B6",x"90",x"6E",x"4D",x"51",
		x"77",x"9E",x"B6",x"A7",x"80",x"5B",x"48",x"60",x"82",x"AC",x"B1",x"95",x"6E",x"51",x"2C",x"31",
		x"5B",x"77",x"99",x"87",x"60",x"48",x"60",x"82",x"A7",x"B6",x"99",x"77",x"51",x"4D",x"6E",x"95",
		x"B6",x"AC",x"87",x"60",x"48",x"56",x"80",x"99",x"7C",x"64",x"87",x"95",x"72",x"69",x"8B",x"AC",
		x"C4",x"BA",x"90",x"77",x"80",x"A7",x"C4",x"BF",x"A7",x"82",x"5B",x"51",x"69",x"95",x"99",x"7C",
		x"5B",x"31",x"14",x"19",x"43",x"69",x"51",x"35",x"48",x"3A",x"31",x"3F",x"60",x"6E",x"48",x"48",
		x"51",x"3F",x"1E",x"22",x"51",x"6E",x"64",x"3A",x"22",x"3A",x"5B",x"80",x"A7",x"B1",x"8B",x"72",
		x"4D",x"4D",x"77",x"90",x"8B",x"64",x"43",x"22",x"06",x"27",x"48",x"6E",x"80",x"60",x"3A",x"35",
		x"56",x"80",x"9E",x"99",x"77",x"56",x"64",x"60",x"4D",x"5B",x"69",x"60",x"51",x"64",x"77",x"9E",
		x"A3",x"87",x"64",x"64",x"8B",x"80",x"80",x"95",x"8B",x"7C",x"56",x"43",x"56",x"80",x"8B",x"80",
		x"87",x"7C",x"72",x"4D",x"2C",x"31",x"5B",x"7C",x"6E",x"4D",x"31",x"48",x"6E",x"87",x"B1",x"BF",
		x"9E",x"82",x"56",x"5B",x"77",x"99",x"95",x"72",x"80",x"A3",x"C4",x"A7",x"8B",x"A7",x"BF",x"9E",
		x"8B",x"B1",x"B6",x"95",x"77",x"72",x"95",x"B1",x"D7",x"F7",x"E0",x"BF",x"99",x"80",x"99",x"B1",
		x"E0",x"E9",x"C8",x"A7",x"99",x"BF",x"B6",x"B6",x"CD",x"C4",x"AC",x"90",x"9E",x"C4",x"DB",x"BF",
		x"95",x"87",x"95",x"8B",x"90",x"87",x"87",x"90",x"8B",x"87",x"87",x"90",x"95",x"A7",x"9E",x"82",
		x"64",x"4D",x"72",x"8B",x"B1",x"BA",x"90",x"77",x"51",x"56",x"80",x"99",x"BA",x"A7",x"82",x"64",
		x"48",x"69",x"87",x"A7",x"BA",x"90",x"77",x"51",x"4D",x"77",x"90",x"B1",x"A7",x"82",x"69",x"3F",
		x"27",x"48",x"64",x"90",x"95",x"7C",x"5B",x"51",x"77",x"90",x"B6",x"AC",x"87",x"69",x"4D",x"60",
		x"80",x"9E",x"B6",x"99",x"7C",x"56",x"51",x"6E",x"90",x"90",x"69",x"72",x"95",x"87",x"64",x"7C",
		x"95",x"BF",x"C8",x"AC",x"87",x"7C",x"95",x"B6",x"C8",x"B6",x"95",x"77",x"56",x"60",x"80",x"9E",
		x"8B",x"64",x"4D",x"27",x"14",x"31",x"56",x"69",x"3F",x"3F",x"4D",x"31",x"3A",x"48",x"6E",x"60",
		x"3F",x"51",x"4D",x"2C",x"19",x"35",x"5B",x"6E",x"51",x"2C",x"27",x"51",x"6E",x"8B",x"B1",x"A3",
		x"82",x"64",x"48",x"5B",x"80",x"95",x"7C",x"56",x"3A",x"19",x"10",x"35",x"51",x"7C",x"77",x"56",
		x"31",x"43",x"69",x"87",x"A7",x"8B",x"64",x"56",x"69",x"51",x"4D",x"64",x"69",x"51",x"56",x"69",
		x"87",x"AC",x"99",x"7C",x"60",x"77",x"8B",x"7C",x"8B",x"95",x"87",x"72",x"43",x"43",x"64",x"87",
		x"82",x"82",x"82",x"77",x"64",x"43",x"27",x"43",x"6E",x"7C",x"64",x"3A",x"35",x"56",x"77",x"9E",
		x"BF",x"B6",x"95",x"6E",x"51",x"60",x"8B",x"A3",x"90",x"9E",x"B6",x"DB",x"E5",x"BA",x"9E",x"7C",
		x"7C",x"A3",x"BF",x"E0",x"CD",x"A3",x"8B",x"9E",x"C8",x"DB",x"B6",x"A7",x"B1",x"AC",x"BA",x"B6",
		x"B6",x"B1",x"A7",x"AC",x"B1",x"BA",x"CD",x"BF",x"A3",x"82",x"6E",x"8B",x"AC",x"CD",x"D7",x"AC",
		x"90",x"69",x"72",x"95",x"B1",x"D2",x"BF",x"95",x"80",x"90",x"BA",x"D2",x"CD",x"C8",x"A3",x"87",
		x"64",x"60",x"87",x"A3",x"C8",x"B6",x"90",x"72",x"56",x"6E",x"90",x"A3",x"8B",x"64",x"3F",x"35",
		x"5B",x"80",x"9E",x"9E",x"7C",x"56",x"3A",x"43",x"6E",x"8B",x"AC",x"C8",x"A7",x"82",x"64",x"51",
		x"80",x"7C",x"77",x"7C",x"6E",x"5B",x"60",x"72",x"6E",x"72",x"80",x"8B",x"82",x"69",x"5B",x"64",
		x"56",x"3A",x"31",x"5B",x"7C",x"77",x"72",x"77",x"69",x"5B",x"60",x"7C",x"90",x"80",x"56",x"31",
		x"27",x"43",x"6E",x"90",x"90",x"72",x"4D",x"2C",x"35",x"3A",x"3A",x"4D",x"5B",x"51",x"35",x"27",
		x"3F",x"69",x"87",x"AC",x"B1",x"87",x"6E",x"48",x"51",x"7C",x"95",x"B6",x"9E",x"7C",x"60",x"43",
		x"64",x"82",x"A7",x"B6",x"8B",x"72",x"4D",x"51",x"77",x"90",x"B1",x"9E",x"82",x"60",x"48",x"60",
		x"87",x"90",x"87",x"8B",x"80",x"80",x"8B",x"99",x"99",x"82",x"64",x"72",x"95",x"AC",x"A3",x"A7",
		x"9E",x"90",x"77",x"69",x"82",x"AC",x"AC",x"8B",x"6E",x"43",x"56",x"72",x"99",x"B6",x"9E",x"80",
		x"5B",x"35",x"27",x"43",x"6E",x"90",x"95",x"77",x"4D",x"56",x"77",x"95",x"BF",x"D7",x"C8",x"9E",
		x"7C",x"5B",x"43",x"69",x"87",x"A7",x"B6",x"8B",x"72",x"4D",x"51",x"77",x"90",x"B6",x"A3",x"80",
		x"60",x"43",x"64",x"82",x"A3",x"C4",x"DB",x"CD",x"B1",x"8B",x"8B",x"AC",x"CD",x"D2",x"BA",x"99",
		x"77",x"5B",x"72",x"90",x"B6",x"C4",x"A7",x"82",x"7C",x"9E",x"BF",x"BA",x"95",x"9E",x"99",x"99",
		x"A3",x"9E",x"9E",x"99",x"95",x"99",x"9E",x"AC",x"B6",x"9E",x"87",x"64",x"64",x"82",x"A3",x"B1",
		x"9E",x"80",x"5B",x"43",x"5B",x"7C",x"9E",x"AC",x"90",x"6E",x"64",x"87",x"A7",x"B1",x"AC",x"99",
		x"7C",x"5B",x"3F",x"51",x"72",x"90",x"A7",x"8B",x"6E",x"48",x"43",x"60",x"82",x"87",x"60",x"43",
		x"1E",x"2C",x"56",x"77",x"90",x"77",x"5B",x"35",x"27",x"48",x"69",x"87",x"B1",x"AC",x"8B",x"69",
		x"43",x"56",x"72",x"69",x"6E",x"69",x"5B",x"4D",x"60",x"69",x"60",x"6E",x"80",x"82",x"6E",x"4D",
		x"56",x"5B",x"3F",x"27",x"35",x"60",x"72",x"69",x"6E",x"69",x"56",x"51",x"60",x"80",x"82",x"60",
		x"43",x"22",x"31",x"51",x"72",x"90",x"7C",x"60",x"3A",x"2C",x"35",x"31",x"3A",x"51",x"56",x"43",
		x"27",x"2C",x"51",x"6E",x"95",x"B6",x"9E",x"80",x"56",x"43",x"64",x"80",x"AC",x"B1",x"90",x"72",
		x"48",x"51",x"6E",x"90",x"B6",x"A3",x"82",x"60",x"43",x"60",x"7C",x"A7",x"B6",x"95",x"77",x"4D",
		x"4D",x"6E",x"90",x"8B",x"8B",x"8B",x"80",x"82",x"90",x"9E",x"95",x"77",x"69",x"80",x"AC",x"AC",
		x"A3",x"AC",x"99",x"8B",x"69",x"77",x"99",x"B6",x"A7",x"80",x"5B",x"48",x"60",x"82",x"AC",x"B6",
		x"95",x"6E",x"51",x"2C",x"31",x"5B",x"7C",x"99",x"8B",x"64",x"4D",x"60",x"87",x"A7",x"C8",x"DB",
		x"B6",x"90",x"77",x"51",x"51",x"77",x"90",x"B1",x"A7",x"82",x"64",x"48",x"64",x"80",x"A3",x"B6",
		x"95",x"77",x"4D",x"51",x"72",x"90",x"BA",x"D7",x"DB",x"C4",x"99",x"82",x"95",x"BF",x"D7",x"CD",
		x"B1",x"87",x"64",x"60",x"82",x"A7",x"C8",x"BF",x"99",x"77",x"87",x"A7",x"C4",x"A7",x"95",x"A3",
		x"99",x"A7",x"A3",x"A3",x"9E",x"99",x"99",x"9E",x"A7",x"BA",x"B1",x"99",x"72",x"60",x"72",x"99",
		x"B6",x"B1",x"95",x"6E",x"4D",x"48",x"6E",x"90",x"B1",x"A7",x"80",x"60",x"77",x"95",x"B1",x"B1",
		x"AC",x"95",x"6E",x"48",x"3F",x"64",x"87",x"A7",x"A3",x"82",x"5B",x"3F",x"4D",x"77",x"90",x"77",
		x"5B",x"31",x"22",x"43",x"60",x"8B",x"8B",x"6E",x"4D",x"27",x"35",x"56",x"77",x"9E",x"B6",x"A3",
		x"7C",x"5B",x"43",x"69",x"72",x"69",x"72",x"64",x"51",x"51",x"69",x"69",x"69",x"77",x"82",x"80",
		x"60",x"51",x"60",x"51",x"35",x"2C",x"48",x"77",x"72",x"6E",x"72",x"64",x"56",x"56",x"72",x"8B",
		x"7C",x"5B",x"35",x"1E",x"3F",x"5B",x"8B",x"90",x"72",x"51",x"27",x"35",x"35",x"35",x"48",x"56",
		x"56",x"35",x"22",x"3A",x"60",x"82",x"A7",x"B1",x"95",x"6E",x"4D",x"4D",x"72",x"95",x"B6",x"A3",
		x"80",x"60",x"43",x"64",x"82",x"A3",x"B6",x"90",x"77",x"51",x"4D",x"77",x"90",x"B6",x"A7",x"82",
		x"64",x"48",x"5B",x"82",x"95",x"87",x"8B",x"82",x"82",x"87",x"9E",x"9E",x"8B",x"72",x"72",x"95",
		x"B1",x"A7",x"A7",x"A3",x"99",x"7C",x"69",x"82",x"A3",x"B6",x"90",x"77",x"51",x"51",x"77",x"90",
		x"B1",x"A7",x"82",x"69",x"3F",x"27",x"48",x"64",x"90",x"99",x"7C",x"5B",x"56",x"77",x"90",x"B6",
		x"DB",x"CD",x"A7",x"87",x"60",x"48",x"60",x"82",x"A7",x"B6",x"99",x"77",x"51",x"4D",x"72",x"95",
		x"B6",x"AC",x"87",x"64",x"48",x"5B",x"82",x"A3",x"C4",x"DB",x"D2",x"B6",x"90",x"87",x"AC",x"CD",
		x"D7",x"C4",x"9E",x"80",x"60",x"72",x"95",x"B6",x"CD",x"AC",x"87",x"7C",x"95",x"BF",x"C4",x"99",
		x"99",x"9E",x"9E",x"A7",x"A3",x"A3",x"9E",x"99",x"99",x"A3",x"AC",x"BA",x"A7",x"8B",x"69",x"60",
		x"87",x"A3",x"B6",x"A7",x"82",x"64",x"43",x"5B",x"7C",x"9E",x"B6",x"95",x"72",x"64",x"80",x"A7",
		x"B6",x"B1",x"A7",x"80",x"64",x"3F",x"4D",x"77",x"90",x"B1",x"95",x"77",x"51",x"43",x"60",x"82",
		x"8B",x"64",x"48",x"22",x"2C",x"56",x"77",x"95",x"80",x"5B",x"3F",x"22",x"48",x"69",x"87",x"A7",
		x"B1",x"90",x"72",x"4D",x"51",x"77",x"6E",x"6E",x"6E",x"60",x"4D",x"60",x"6E",x"64",x"6E",x"80",
		x"82",x"77",x"5B",x"56",x"5B",x"48",x"31",x"35",x"60",x"77",x"6E",x"72",x"6E",x"60",x"56",x"60",
		x"80",x"8B",x"64",x"48",x"27",x"27",x"56",x"6E",x"95",x"80",x"60",x"3F",x"27",x"35",x"35",x"3A",
		x"4D",x"56",x"48",x"2C",x"27",x"51",x"72",x"90",x"B1",x"A3",x"82",x"64",x"48",x"60",x"80",x"9E",
		x"B1",x"95",x"77",x"51",x"4D",x"72",x"8B",x"B1",x"A7",x"87",x"69",x"48",x"5B",x"80",x"9E",x"B6",
		x"99",x"7C",x"56",x"4D",x"69",x"90",x"90",x"8B",x"8B",x"80",x"82",x"90",x"9E",x"99",x"7C",x"69",
		x"80",x"A3",x"AC",x"A3",x"AC",x"9E",x"90",x"6E",x"72",x"90",x"B6",x"A7",x"87",x"64",x"43",x"60",
		x"7C",x"A7",x"B6",x"99",x"7C",x"56",x"31",x"31",x"51",x"7C",x"99",x"90",x"6E",x"4D",x"60",x"80",
		x"A3",x"CD",x"DB",x"C4",x"95",x"7C",x"56",x"4D",x"77",x"90",x"B6",x"AC",x"87",x"69",x"48",x"48",
		x"48",x"43",x"48",x"51",x"5B",x"51",x"4D",x"5B",x"5B",x"51",x"56",x"60",x"60",x"51",x"43",x"4D",
		x"60",x"87",x"AC",x"BF",x"A3",x"7C",x"56",x"51",x"72",x"95",x"BA",x"B6",x"90",x"6E",x"7C",x"99",
		x"8B",x"95",x"A3",x"99",x"7C",x"6E",x"87",x"AC",x"B1",x"95",x"72",x"72",x"77",x"77",x"77",x"6E",
		x"77",x"7C",x"77",x"72",x"77",x"7C",x"8B",x"95",x"82",x"6E",x"48",x"48",x"69",x"87",x"A7",x"9E",
		x"80",x"60",x"43",x"56",x"77",x"99",x"AC",x"90",x"72",x"51",x"48",x"69",x"87",x"AC",x"A7",x"82",
		x"64",x"48",x"56",x"77",x"99",x"B1",x"99",x"77",x"5B",x"31",x"2C",x"4D",x"6E",x"95",x"90",x"72",
		x"51",x"5B",x"80",x"99",x"BA",x"A3",x"82",x"60",x"4D",x"6E",x"8B",x"AC",x"B6",x"90",x"77",x"51",
		x"5B",x"7C",x"99",x"8B",x"69",x"82",x"9E",x"80",x"6E",x"8B",x"A3",x"D2",x"D7",x"B6",x"90",x"90",
		x"B1",x"CD",x"EE",x"E0",x"BF",x"99",x"80",x"90",x"B6",x"CD",x"AC",x"87",x"6E",x"48",x"43",x"64",
		x"87",x"82",x"5B",x"6E",x"69",x"56",x"60",x"77",x"90",x"72",x"64",x"72",x"60",x"43",x"3F",x"64",
		x"87",x"82",x"60",x"43",x"4D",x"77",x"8B",x"BA",x"CD",x"B1",x"95",x"69",x"60",x"7C",x"9E",x"A3",
		x"82",x"64",x"43",x"1E",x"31",x"51",x"77",x"95",x"80",x"60",x"48",x"64",x"82",x"A7",x"AC",x"90",
		x"6E",x"6E",x"77",x"5B",x"64",x"77",x"72",x"60",x"69",x"80",x"A7",x"B6",x"9E",x"77",x"69",x"8B",
		x"90",x"87",x"9E",x"9E",x"8B",x"64",x"4D",x"56",x"80",x"99",x"87",x"90",x"87",x"7C",x"64",x"3F",
		x"3A",x"56",x"7C",x"80",x"56",x"3A",x"43",x"69",x"8B",x"AC",x"C8",x"AC",x"8B",x"69",x"56",x"7C",
		x"99",x"A3",x"80",x"80",x"99",x"BF",x"BA",x"90",x"A3",x"BF",x"AC",x"8B",x"A7",x"BF",x"A3",x"7C",
		x"6E",x"87",x"B1",x"CD",x"F3",x"F3",x"C4",x"A7",x"82",x"90",x"B6",x"D2",x"EE",x"D2",x"AC",x"95",
		x"B6",x"BF",x"B1",x"C8",x"C8",x"B1",x"95",x"95",x"BA",x"DB",x"C8",x"A3",x"8B",x"95",x"8B",x"90",
		x"8B",x"87",x"8B",x"90",x"87",x"87",x"8B",x"95",x"A7",x"A3",x"90",x"6E",x"4D",x"64",x"80",x"A7",
		x"BF",x"9E",x"82",x"56",x"4D",x"72",x"95",x"B6",x"B1",x"8B",x"64",x"48",x"5B",x"80",x"A3",x"BA",
		x"9E",x"7C",x"56",x"48",x"69",x"8B",x"B1",x"B1",x"8B",x"64",x"48",x"27",x"3A",x"60",x"80",x"99",
		x"80",x"5B",x"48",x"69",x"8B",x"B1",x"B6",x"90",x"6E",x"4D",x"51",x"77",x"99",x"B6",x"A3",x"80",
		x"5B",x"48",x"60",x"87",x"95",x"72",x"69",x"90",x"90",x"69",x"72",x"95",x"B1",x"C8",x"B6",x"8B",
		x"77",x"87",x"B1",x"C8",x"BF",x"A3",x"7C",x"5B",x"56",x"77",x"9E",x"95",x"77",x"51",x"2C",x"14",
		x"22",x"4D",x"69",x"4D",x"3A",x"48",x"35",x"31",x"43",x"69",x"69",x"43",x"4D",x"4D",x"3A",x"1E",
		x"2C",x"5B",x"6E",x"60",x"31",x"22",x"3F",x"64",x"87",x"AC",x"AC",x"8B",x"69",x"48",x"4D",x"77",
		x"95",x"82",x"64",x"3F",x"19",x"0B",x"27",x"4D",x"77",x"7C",x"60",x"35",x"3A",x"5B",x"80",x"A3",
		x"90",x"72",x"56",x"64",x"5B",x"48",x"60",x"69",x"56",x"4D",x"64",x"7C",x"A3",x"A3",x"7C",x"5B",
		x"64",x"82",x"7C",x"82",x"95",x"87",x"72",x"4D",x"3F",x"60",x"82",x"87",x"80",x"82",x"77",x"6E",
		x"48",x"27",x"35",x"64",x"7C",x"64",x"43",x"31",x"4D",x"72",x"8B",x"BA",x"BA",x"99",x"7C",x"51",
		x"60",x"7C",x"99",x"8B",x"72",x"82",x"A7",x"BF",x"9E",x"8B",x"B1",x"BA",x"95",x"8B",x"B6",x"B1",
		x"8B",x"6E",x"77",x"99",x"B6",x"DB",x"F7",x"D7",x"BA",x"8B",x"80",x"9E",x"BA",x"E5",x"E5",x"BF",
		x"9E",x"9E",x"C4",x"B1",x"BA",x"C8",x"BF",x"A3",x"8B",x"A3",x"C8",x"D7",x"B6",x"8B",x"87",x"90",
		x"8B",x"90",x"87",x"87",x"8B",x"8B",x"82",x"87",x"8B",x"99",x"A7",x"95",x"80",x"5B",x"4D",x"77",
		x"90",x"B6",x"B1",x"87",x"6E",x"48",x"5B",x"82",x"9E",x"BA",x"9E",x"7C",x"5B",x"48",x"6E",x"8B",
		x"B1",x"B1",x"87",x"6E",x"48",x"56",x"7C",x"99",x"B6",x"9E",x"7C",x"60",x"3A",x"2C",x"48",x"69",
		x"8B",x"90",x"72",x"51",x"51",x"7C",x"95",x"BA",x"A3",x"80",x"64",x"43",x"64",x"82",x"A7",x"B6",
		x"90",x"77",x"4D",x"4D",x"72",x"90",x"8B",x"69",x"7C",x"95",x"82",x"69",x"80",x"9E",x"BA",x"BF",
		x"A3",x"80",x"77",x"99",x"BA",x"C4",x"B1",x"8B",x"6E",x"4D",x"60",x"87",x"9E",x"82",x"5B",x"43",
		x"1E",x"14",x"35",x"5B",x"60",x"35",x"43",x"43",x"31",x"3A",x"4D",x"72",x"51",x"3F",x"51",x"48",
		x"22",x"1E",x"3F",x"60",x"69",x"48",x"27",x"2C",x"56",x"72",x"95",x"B1",x"9E",x"7C",x"5B",x"48",
		x"60",x"82",x"90",x"72",x"51",x"31",x"10",x"14",x"3A",x"5B",x"7C",x"6E",x"4D",x"31",x"4D",x"6E",
		x"90",x"A3",x"82",x"60",x"5B",x"69",x"4D",x"51",x"64",x"64",x"4D",x"5B",x"69",x"90",x"AC",x"90",
		x"72",x"5B",x"80",x"87",x"7C",x"90",x"90",x"82",x"64",x"3F",x"48",x"6E",x"87",x"80",x"82",x"82",
		x"72",x"60",x"3A",x"27",x"4D",x"72",x"7C",x"5B",x"31",x"3A",x"5B",x"80",x"A3",x"BF",x"B1",x"8B",
		x"64",x"51",x"69",x"90",x"A3",x"80",x"77",x"95",x"BA",x"BA",x"95",x"99",x"BA",x"B1",x"8B",x"9E",
		x"BA",x"A7",x"7C",x"69",x"82",x"A3",x"C8",x"EE",x"F3",x"CD",x"A7",x"82",x"87",x"A7",x"D2",x"E9",
		x"DB",x"B1",x"90",x"B1",x"C4",x"B1",x"C4",x"C8",x"BA",x"95",x"90",x"B1",x"D2",x"CD",x"A7",x"87",
		x"90",x"90",x"90",x"8B",x"87",x"8B",x"90",x"8B",x"87",x"8B",x"90",x"A7",x"A3",x"90",x"72",x"4D",
		x"64",x"80",x"A7",x"BF",x"A3",x"82",x"5B",x"4D",x"6E",x"87",x"B6",x"B1",x"90",x"72",x"48",x"5B",
		x"77",x"99",x"BA",x"9E",x"82",x"5B",x"48",x"69",x"82",x"B1",x"B1",x"90",x"72",x"48",x"2C",x"31",
		x"56",x"80",x"99",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",x"7C",x"4D",x"51",x"72",x"90",
		x"BA",x"A7",x"87",x"64",x"43",x"60",x"80",x"95",x"77",x"69",x"87",x"90",x"6E",x"6E",x"8B",x"B1",
		x"C8",x"BA",x"95",x"72",x"87",x"A3",x"C4",x"BF",x"A3",x"87",x"5B",x"51",x"72",x"90",x"95",x"77",
		x"5B",x"35",x"10",x"22",x"43",x"64",x"51",x"35",x"4D",x"3A",x"31",x"43",x"60",x"6E",x"48",x"48",
		x"51",x"3A",x"1E",x"22",x"51",x"72",x"60",x"3A",x"27",x"3F",x"64",x"80",x"AC",x"B1",x"90",x"72",
		x"48",x"4D",x"6E",x"90",x"87",x"64",x"48",x"22",x"06",x"27",x"43",x"72",x"80",x"64",x"43",x"3A",
		x"5B",x"7C",x"9E",x"99",x"77",x"56",x"64",x"60",x"4D",x"5B",x"69",x"60",x"51",x"60",x"7C",x"A3",
		x"A7",x"87",x"60",x"64",x"87",x"82",x"82",x"99",x"8B",x"77",x"51",x"3F",x"5B",x"82",x"8B",x"80",
		x"87",x"7C",x"72",x"51",x"2C",x"35",x"5B",x"7C",x"6E",x"48",x"31",x"4D",x"72",x"8B",x"B1",x"BA",
		x"9E",x"80",x"5B",x"5B",x"7C",x"9E",x"95",x"95",x"AC",x"C8",x"E5",x"CD",x"AC",x"87",x"77",x"90",
		x"B1",x"D7",x"D7",x"B6",x"90",x"95",x"BA",x"D7",x"C8",x"A7",x"B6",x"AC",x"B1",x"B6",x"B1",x"B1",
		x"AC",x"A7",x"AC",x"B1",x"C4",x"C4",x"AC",x"90",x"72",x"7C",x"99",x"BA",x"D7",x"BF",x"99",x"7C",
		x"69",x"82",x"A3",x"C8",x"C8",x"A7",x"82",x"87",x"AC",x"C8",x"D2",x"CD",x"B6",x"90",x"72",x"5B",
		x"77",x"90",x"B6",x"BF",x"9E",x"82",x"60",x"60",x"80",x"9E",x"95",x"6E",x"51",x"31",x"4D",x"72",
		x"90",x"A7",x"82",x"64",x"43",x"3A",x"60",x"80",x"9E",x"BF",x"B6",x"90",x"77",x"56",x"6E",x"82",
		x"77",x"7C",x"72",x"64",x"5B",x"72",x"72",x"6E",x"7C",x"8B",x"8B",x"77",x"5B",x"64",x"60",x"48",
		x"31",x"43",x"6E",x"7C",x"72",x"77",x"6E",x"60",x"5B",x"6E",x"8B",x"87",x"60",x"43",x"22",x"3A",
		x"60",x"80",x"99",x"7C",x"5B",x"35",x"31",x"3A",x"35",x"43",x"56",x"56",x"43",x"27",x"35",x"5B",
		x"77",x"A3",x"B6",x"99",x"7C",x"51",x"48",x"69",x"87",x"B1",x"AC",x"8B",x"69",x"43",x"56",x"77",
		x"99",x"B6",x"99",x"80",x"56",x"48",x"69",x"82",x"B1",x"AC",x"90",x"6E",x"48",x"51",x"77",x"90",
		x"87",x"8B",x"87",x"80",x"82",x"95",x"9E",x"8B",x"72",x"69",x"87",x"B1",x"A7",x"A3",x"A7",x"95",
		x"87",x"64",x"7C",x"9E",x"B6",x"9E",x"77",x"51",x"48",x"64",x"8B",x"AC",x"AC",x"8B",x"64",x"48",
		x"27",x"35",x"60",x"80",x"99",x"80",x"5B",x"4D",x"64",x"8B",x"AC",x"CD",x"D2",x"A7",x"8B",x"69",
		x"4D",x"56",x"77",x"95",x"B1",x"99",x"7C",x"5B",x"48",x"69",x"82",x"A7",x"AC",x"8B",x"6E",x"4D",
		x"51",x"77",x"90",x"B6",x"D7",x"D2",x"BF",x"90",x"80",x"99",x"BA",x"D2",x"C4",x"A7",x"87",x"5B",
		x"64",x"82",x"A7",x"C8",x"B6",x"90",x"77",x"8B",x"AC",x"C4",x"9E",x"95",x"9E",x"95",x"A3",x"9E",
		x"9E",x"9E",x"95",x"95",x"99",x"A7",x"B6",x"A7",x"95",x"6E",x"5B",x"77",x"95",x"B1",x"A7",x"8B",
		x"6E",x"43",x"4D",x"6E",x"95",x"AC",x"9E",x"77",x"60",x"77",x"99",x"B1",x"AC",x"A7",x"87",x"64",
		x"3F",x"43",x"69",x"8B",x"A7",x"99",x"77",x"51",x"3A",x"4D",x"7C",x"8B",x"6E",x"51",x"22",x"22",
		x"43",x"64",x"90",x"82",x"69",x"43",x"22",x"3A",x"56",x"80",x"A3",x"B6",x"99",x"72",x"51",x"43",
		x"6E",x"6E",x"69",x"6E",x"60",x"4D",x"56",x"69",x"64",x"69",x"77",x"82",x"77",x"5B",x"4D",x"60",
		x"48",x"2C",x"27",x"4D",x"77",x"6E",x"6E",x"6E",x"60",x"51",x"56",x"77",x"8B",x"72",x"56",x"27",
		x"22",x"43",x"64",x"90",x"87",x"6E",x"48",x"22",x"35",x"31",x"35",x"48",x"56",x"51",x"2C",x"22",
		x"3F",x"64",x"87",x"AC",x"AC",x"87",x"64",x"43",x"51",x"77",x"99",x"B1",x"9E",x"7C",x"56",x"43",
		x"60",x"87",x"AC",x"B1",x"90",x"69",x"48",x"4D",x"72",x"95",x"B6",x"A3",x"80",x"5B",x"48",x"5B",
		x"87",x"90",x"82",x"90",x"80",x"82",x"87",x"99",x"99",x"82",x"69",x"72",x"9E",x"B1",x"A3",x"A7",
		x"9E",x"95",x"7C",x"6E",x"87",x"AC",x"B1",x"87",x"6E",x"48",x"56",x"7C",x"95",x"B6",x"9E",x"7C",
		x"60",x"35",x"27",x"4D",x"69",x"95",x"95",x"77",x"56",x"56",x"7C",x"95",x"BF",x"DB",x"C4",x"A3",
		x"80",x"56",x"48",x"64",x"8B",x"AC",x"B1",x"90",x"6E",x"4D",x"51",x"77",x"99",x"B6",x"A7",x"80",
		x"5B",x"48",x"60",x"87",x"A7",x"C8",x"DB",x"CD",x"B1",x"87",x"8B",x"B1",x"CD",x"D7",x"BA",x"95",
		x"77",x"5B",x"7C",x"99",x"BA",x"C8",x"A3",x"82",x"7C",x"99",x"C4",x"BA",x"95",x"9E",x"99",x"9E",
		x"A7",x"A3",x"A3",x"9E",x"95",x"9E",x"A3",x"B1",x"BA",x"9E",x"87",x"60",x"69",x"8B",x"A7",x"B6",
		x"9E",x"7C",x"5B",x"43",x"60",x"80",x"A3",x"B1",x"8B",x"6E",x"69",x"87",x"AC",x"B1",x"B1",x"9E",
		x"77",x"5B",x"3A",x"56",x"7C",x"99",x"B1",x"8B",x"6E",x"48",x"43",x"69",x"87",x"87",x"64",x"3F",
		x"22",x"31",x"56",x"80",x"95",x"80",x"5B",x"31",x"27",x"43",x"6E",x"8B",x"B1",x"B1",x"87",x"6E",
		x"43",x"56",x"77",x"69",x"72",x"69",x"5B",x"4D",x"60",x"69",x"64",x"6E",x"80",x"82",x"72",x"51",
		x"56",x"5B",x"43",x"27",x"3A",x"69",x"77",x"6E",x"6E",x"6E",x"5B",x"51",x"64",x"82",x"87",x"60",
		x"43",x"1E",x"31",x"5B",x"77",x"95",x"7C",x"5B",x"35",x"2C",x"35",x"35",x"3F",x"51",x"56",x"43",
		x"27",x"2C",x"5B",x"77",x"95",x"B1",x"9E",x"7C",x"5B",x"48",x"69",x"82",x"A7",x"AC",x"8B",x"72",
		x"4D",x"51",x"77",x"95",x"B1",x"A3",x"80",x"60",x"48",x"64",x"82",x"A3",x"B1",x"90",x"77",x"51",
		x"51",x"72",x"95",x"8B",x"8B",x"8B",x"80",x"87",x"95",x"9E",x"95",x"77",x"69",x"82",x"A7",x"AC",
		x"A7",x"AC",x"99",x"87",x"6E",x"77",x"99",x"BA",x"9E",x"82",x"5B",x"48",x"69",x"82",x"B1",x"B1",
		x"95",x"72",x"4D",x"2C",x"35",x"5B",x"80",x"99",x"8B",x"64",x"4D",x"69",x"87",x"AC",x"D2",x"D7",
		x"BA",x"90",x"72",x"4D",x"51",x"7C",x"95",x"BA",x"A7",x"82",x"64",x"48",x"69",x"87",x"A7",x"BA",
		x"90",x"77",x"51",x"51",x"77",x"95",x"B1",x"D7",x"DB",x"C4",x"A3",x"87",x"99",x"BF",x"D7",x"CD",
		x"AC",x"8B",x"69",x"64",x"87",x"A3",x"C8",x"BA",x"99",x"7C",x"8B",x"B1",x"C8",x"AC",x"99",x"A3",
		x"99",x"A3",x"A3",x"A3",x"A3",x"99",x"99",x"9E",x"A3",x"B6",x"AC",x"99",x"72",x"5B",x"77",x"95",
		x"B6",x"B1",x"90",x"72",x"48",x"4D",x"6E",x"8B",x"B6",x"A3",x"82",x"64",x"77",x"99",x"B1",x"B1",
		x"A7",x"90",x"72",x"43",x"43",x"64",x"82",x"AC",x"9E",x"82",x"5B",x"3A",x"51",x"72",x"8B",x"77",
		x"56",x"35",x"22",x"48",x"64",x"87",x"8B",x"6E",x"4D",x"2C",x"35",x"5B",x"77",x"9E",x"BA",x"9E",
		x"80",x"56",x"43",x"6E",x"72",x"6E",x"6E",x"64",x"56",x"56",x"6E",x"64",x"69",x"77",x"82",x"80",
		x"60",x"51",x"60",x"51",x"31",x"2C",x"4D",x"6E",x"72",x"6E",x"72",x"64",x"51",x"5B",x"72",x"87",
		x"77",x"56",x"35",x"22",x"43",x"60",x"87",x"8B",x"6E",x"51",x"2C",x"35",x"35",x"35",x"48",x"56",
		x"51",x"3A",x"27",x"3F",x"64",x"80",x"AC",x"B1",x"90",x"72",x"48",x"51",x"72",x"90",x"B6",x"A3",
		x"87",x"60",x"43",x"60",x"80",x"A7",x"B6",x"95",x"77",x"4D",x"4D",x"72",x"90",x"BA",x"A7",x"8B",
		x"64",x"48",x"5B",x"80",x"95",x"87",x"90",x"82",x"82",x"87",x"99",x"9E",x"87",x"6E",x"6E",x"95",
		x"B6",x"A3",x"AC",x"A3",x"95",x"80",x"69",x"87",x"AC",x"B6",x"8B",x"72",x"4D",x"51",x"7C",x"95",
		x"BA",x"A3",x"80",x"64",x"43",x"2C",x"48",x"69",x"8B",x"95",x"7C",x"56",x"51",x"7C",x"95",x"BA",
		x"D7",x"C8",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",x"77",x"4D",x"48",x"48",x"48",
		x"4D",x"4D",x"4D",x"51",x"51",x"51",x"51",x"56",x"56",x"56",x"56",x"5B",x"5B",x"5B",x"5B",x"5B",
		x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"64",x"69",x"69",x"69",x"69",x"69",
		x"69",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"6E",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",
		x"72",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"82",x"82",x"87",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",
		x"80",x"80",x"80",x"80",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"80",x"7C",x"7C",
		x"7C",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"7C",
		x"80",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",
		x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"80",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"80",x"80",x"7C",x"77",x"77",x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"7C",x"80",x"82",
		x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",
		x"7C",x"80",x"82",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",
		x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",
		x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"72",x"77",x"80",x"82",x"7C",x"77",x"82",x"82",x"7C",x"7C",
		x"82",x"82",x"77",x"7C",x"82",x"80",x"77",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",
		x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",
		x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",
		x"7C",x"77",x"72",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"7C",x"82",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"80",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"82",x"80",
		x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",
		x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",
		x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"80",x"80",x"77",x"7C",x"80",x"7C",x"77",x"7C",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"82",x"82",x"77",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"77",x"7C",x"7C",x"7C",x"7C",
		x"77",x"77",x"7C",x"7C",x"77",x"77",x"7C",x"7C",x"80",x"7C",x"7C",x"7C",x"80",x"7C",x"82",x"82",
		x"80",x"7C",x"7C",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"80",
		x"7C",x"80",x"87",x"87",x"87",x"8B",x"8B",x"8B",x"95",x"90",x"90",x"99",x"95",x"95",x"95",x"95",
		x"90",x"95",x"99",x"95",x"87",x"87",x"8B",x"82",x"7C",x"7C",x"80",x"77",x"6E",x"72",x"72",x"69",
		x"64",x"69",x"60",x"5B",x"48",x"48",x"4D",x"48",x"56",x"51",x"4D",x"51",x"51",x"51",x"5B",x"64",
		x"60",x"64",x"69",x"69",x"72",x"72",x"72",x"77",x"80",x"80",x"80",x"87",x"8B",x"87",x"8B",x"95",
		x"99",x"90",x"99",x"99",x"95",x"90",x"95",x"95",x"90",x"87",x"87",x"87",x"80",x"7C",x"80",x"7C",
		x"77",x"77",x"72",x"72",x"72",x"6E",x"69",x"72",x"7C",x"7C",x"6E",x"72",x"7C",x"7C",x"7C",x"82",
		x"87",x"82",x"7C",x"82",x"87",x"82",x"87",x"8B",x"82",x"82",x"82",x"80",x"80",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"80",x"7C",x"82",x"82",x"82",x"82",x"82",x"87",x"87",x"87",x"87",x"87",
		x"87",x"80",x"82",x"87",x"82",x"87",x"8B",x"87",x"80",x"7C",x"87",x"87",x"7C",x"80",x"80",x"77",
		x"7C",x"7C",x"7C",x"77",x"7C",x"80",x"7C",x"7C",x"7C",x"72",x"72",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"72",x"7C",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",
		x"80",x"80",x"82",x"80",x"77",x"80",x"82",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"77",x"72",x"77",x"7C",x"77",x"72",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"72",x"77",x"7C",x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"80",x"77",x"77",
		x"77",x"77",x"77",x"77",x"80",x"87",x"80",x"77",x"80",x"7C",x"77",x"7C",x"82",x"82",x"82",x"82",
		x"80",x"77",x"77",x"80",x"90",x"87",x"77",x"80",x"7C",x"80",x"82",x"80",x"87",x"87",x"82",x"7C",
		x"77",x"82",x"80",x"80",x"87",x"82",x"80",x"77",x"7C",x"7C",x"80",x"82",x"80",x"82",x"7C",x"7C",
		x"7C",x"77",x"72",x"7C",x"82",x"80",x"77",x"7C",x"7C",x"72",x"77",x"80",x"82",x"7C",x"77",x"7C",
		x"77",x"77",x"7C",x"82",x"82",x"77",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"82",x"7C",x"7C",
		x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"77",x"77",x"7C",x"7C",x"80",x"7C",x"77",x"77",x"77",x"7C",x"80",x"7C",
		x"7C",x"7C",x"80",x"77",x"77",x"80",x"80",x"80",x"7C",x"77",x"7C",x"80",x"87",x"80",x"7C",x"82",
		x"87",x"80",x"7C",x"82",x"82",x"82",x"82",x"82",x"82",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",
		x"80",x"82",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"82",x"80",x"7C",x"7C",x"82",x"80",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"77",x"6E",x"77",x"80",x"7C",
		x"80",x"82",x"80",x"72",x"72",x"7C",x"80",x"72",x"72",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"72",
		x"7C",x"80",x"77",x"72",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"72",x"77",x"80",x"7C",x"80",x"82",
		x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"80",x"82",x"80",x"82",x"80",x"7C",x"82",x"82",x"80",x"80",x"7C",x"7C",x"7C",
		x"80",x"82",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"82",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"82",x"7C",x"7C",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"77",x"72",x"80",x"7C",x"7C",
		x"82",x"80",x"7C",x"72",x"7C",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"82",x"80",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",
		x"80",x"7C",x"7C",x"7C",x"72",x"77",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"77",x"77",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",
		x"80",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",
		x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"7C",x"7C",x"80",x"82",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"82",x"80",x"7C",x"80",
		x"80",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",
		x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"80",x"82",
		x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",
		x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"77",x"7C",x"82",
		x"7C",x"77",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",
		x"77",x"7C",x"82",x"7C",x"77",x"80",x"80",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"80",x"80",x"77",
		x"7C",x"82",x"7C",x"77",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"82",x"7C",x"7C",
		x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",
		x"80",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"80",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",
		x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",x"7C",x"80",
		x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",
		x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",
		x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",x"80",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"82",x"80",x"7C",x"80",x"82",
		x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"77",x"7C",x"82",x"7C",
		x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",
		x"82",x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"82",x"80",x"7C",x"7C",x"82",
		x"80",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",
		x"7C",x"80",x"82",x"7C",x"7C",x"80",x"82",x"7C",x"7C",x"80",x"80",x"7C",x"7C",x"82",x"80",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"80",x"82",x"80",x"7C",x"80",
		x"82",x"8B",x"82",x"7C",x"87",x"87",x"80",x"80",x"87",x"87",x"80",x"6E",x"6E",x"87",x"A3",x"C4",
		x"E0",x"C8",x"A3",x"82",x"6E",x"8B",x"A7",x"CD",x"D2",x"B1",x"8B",x"8B",x"B6",x"A3",x"A7",x"B6",
		x"B1",x"95",x"80",x"95",x"BA",x"C8",x"B1",x"80",x"80",x"87",x"80",x"82",x"7C",x"80",x"82",x"82",
		x"7C",x"80",x"82",x"90",x"9E",x"90",x"77",x"51",x"43",x"64",x"87",x"AC",x"AC",x"87",x"64",x"43",
		x"4D",x"77",x"99",x"B1",x"9E",x"77",x"51",x"43",x"60",x"82",x"A7",x"AC",x"8B",x"64",x"43",x"4D",
		x"6E",x"95",x"B1",x"9E",x"7C",x"56",x"35",x"1E",x"43",x"64",x"87",x"8B",x"6E",x"4D",x"4D",x"77",
		x"90",x"B6",x"A3",x"7C",x"60",x"43",x"60",x"80",x"A3",x"B6",x"8B",x"72",x"4D",x"48",x"72",x"90",
		x"8B",x"69",x"77",x"90",x"80",x"64",x"7C",x"99",x"BF",x"CD",x"AC",x"87",x"80",x"A3",x"BF",x"E5",
		x"DB",x"B1",x"90",x"72",x"80",x"A7",x"BA",x"A7",x"80",x"60",x"3A",x"2C",x"51",x"77",x"7C",x"5B",
		x"5B",x"60",x"48",x"51",x"64",x"82",x"6E",x"5B",x"64",x"5B",x"3F",x"31",x"4D",x"72",x"7C",x"56",
		x"35",x"3A",x"5B",x"82",x"9E",x"C4",x"AC",x"87",x"69",x"4D",x"6E",x"90",x"9E",x"82",x"5B",x"3A",
		x"19",x"19",x"43",x"60",x"82",x"7C",x"51",x"3A",x"4D",x"72",x"95",x"A7",x"90",x"64",x"60",x"6E",
		x"56",x"56",x"69",x"6E",x"56",x"5B",x"6E",x"8B",x"AC",x"95",x"77",x"5B",x"80",x"8B",x"7C",x"8B",
		x"90",x"82",x"69",x"43",x"48",x"6E",x"8B",x"82",x"82",x"80",x"77",x"60",x"35",x"27",x"3F",x"72",
		x"77",x"5B",x"3A",x"35",x"5B",x"77",x"99",x"BF",x"AC",x"8B",x"69",x"4D",x"64",x"87",x"99",x"7C",
		x"72",x"8B",x"B6",x"B6",x"90",x"90",x"B6",x"AC",x"87",x"99",x"B6",x"A3",x"77",x"64",x"80",x"9E",
		x"C4",x"E5",x"EE",x"C8",x"9E",x"80",x"82",x"A3",x"C8",x"E5",x"D7",x"A7",x"8B",x"A7",x"BA",x"AC",
		x"BF",x"C4",x"B1",x"8B",x"8B",x"AC",x"CD",x"C8",x"9E",x"82",x"87",x"87",x"87",x"87",x"80",x"87",
		x"87",x"82",x"80",x"87",x"8B",x"9E",x"9E",x"8B",x"6E",x"4D",x"5B",x"7C",x"99",x"B6",x"9E",x"80",
		x"5B",x"48",x"69",x"82",x"A7",x"AC",x"8B",x"6E",x"4D",x"51",x"72",x"90",x"B1",x"9E",x"7C",x"5B",
		x"43",x"60",x"80",x"A3",x"AC",x"8B",x"6E",x"4D",x"22",x"2C",x"4D",x"72",x"95",x"82",x"64",x"48",
		x"60",x"80",x"9E",x"B1",x"90",x"72",x"51",x"4D",x"6E",x"87",x"AC",x"A3",x"82",x"64",x"43",x"56",
		x"7C",x"95",x"77",x"64",x"82",x"90",x"69",x"69",x"82",x"A3",x"C4",x"B6",x"95",x"77",x"80",x"A3",
		x"BF",x"BA",x"9E",x"82",x"5B",x"51",x"69",x"8B",x"95",x"72",x"51",x"35",x"10",x"1E",x"3F",x"64",
		x"4D",x"31",x"48",x"3A",x"31",x"3A",x"5B",x"6E",x"43",x"43",x"4D",x"3A",x"19",x"22",x"48",x"64",
		x"5B",x"35",x"1E",x"35",x"60",x"7C",x"A7",x"AC",x"8B",x"6E",x"43",x"48",x"6E",x"8B",x"82",x"60",
		x"48",x"1E",x"01",x"22",x"3F",x"6E",x"7C",x"60",x"3F",x"35",x"56",x"77",x"99",x"95",x"77",x"56",
		x"60",x"5B",x"48",x"56",x"64",x"5B",x"4D",x"5B",x"77",x"9E",x"A3",x"82",x"5B",x"60",x"82",x"80",
		x"80",x"95",x"87",x"77",x"4D",x"3A",x"51",x"80",x"87",x"7C",x"82",x"77",x"6E",x"51",x"2C",x"31",
		x"56",x"77",x"6E",x"43",x"2C",x"3F",x"69",x"8B",x"AC",x"BF",x"99",x"7C",x"56",x"51",x"7C",x"99",
		x"95",x"72",x"80",x"9E",x"BF",x"A7",x"87",x"A3",x"BA",x"99",x"87",x"AC",x"B6",x"90",x"6E",x"6E",
		x"8B",x"B6",x"D2",x"F3",x"E0",x"B6",x"99",x"7C",x"95",x"B6",x"DB",x"E9",x"C4",x"9E",x"95",x"BA",
		x"B6",x"B1",x"C8",x"C4",x"A7",x"8B",x"95",x"C4",x"D7",x"BF",x"99",x"87",x"90",x"8B",x"90",x"87",
		x"87",x"8B",x"8B",x"82",x"87",x"8B",x"95",x"A7",x"99",x"87",x"60",x"4D",x"6E",x"87",x"B6",x"B6",
		x"95",x"77",x"4D",x"56",x"77",x"95",x"BA",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",
		x"72",x"4D",x"4D",x"72",x"99",x"B6",x"A7",x"82",x"60",x"3F",x"22",x"43",x"69",x"87",x"99",x"77",
		x"51",x"4D",x"72",x"95",x"B6",x"AC",x"87",x"64",x"48",x"5B",x"80",x"A3",x"B6",x"9E",x"77",x"51",
		x"48",x"69",x"90",x"90",x"69",x"72",x"95",x"87",x"69",x"7C",x"9E",x"BA",x"C8",x"A7",x"82",x"77",
		x"90",x"BA",x"C8",x"B6",x"99",x"72",x"51",x"56",x"80",x"9E",x"8B",x"6E",x"48",x"1E",x"10",x"2C",
		x"56",x"64",x"3F",x"3F",x"48",x"31",x"35",x"48",x"6E",x"60",x"3F",x"4D",x"48",x"31",x"19",x"35",
		x"60",x"6E",x"56",x"27",x"27",x"48",x"6E",x"90",x"B1",x"A7",x"82",x"5B",x"43",x"56",x"80",x"95",
		x"7C",x"5B",x"35",x"14",x"0B",x"31",x"56",x"7C",x"77",x"56",x"31",x"43",x"64",x"8B",x"A3",x"8B",
		x"6E",x"5B",x"69",x"56",x"4D",x"64",x"69",x"56",x"56",x"6E",x"87",x"AC",x"99",x"77",x"5B",x"72",
		x"87",x"7C",x"8B",x"95",x"82",x"6E",x"48",x"43",x"69",x"8B",x"82",x"80",x"82",x"77",x"69",x"3F",
		x"27",x"43",x"69",x"7C",x"60",x"3A",x"31",x"5B",x"7C",x"95",x"BA",x"B1",x"95",x"6E",x"51",x"69",
		x"87",x"9E",x"82",x"72",x"8B",x"B6",x"BF",x"95",x"95",x"BA",x"B6",x"8B",x"99",x"BA",x"A7",x"87",
		x"6E",x"80",x"A3",x"BF",x"E9",x"F3",x"D2",x"B1",x"82",x"87",x"A3",x"C4",x"EE",x"DB",x"BA",x"99",
		x"AC",x"C4",x"B1",x"C4",x"C8",x"BA",x"9E",x"90",x"AC",x"D2",x"D2",x"AC",x"87",x"90",x"90",x"90",
		x"90",x"87",x"8B",x"90",x"8B",x"82",x"8B",x"90",x"A3",x"A7",x"90",x"7C",x"51",x"5B",x"80",x"99",
		x"BF",x"A7",x"82",x"64",x"48",x"69",x"87",x"AC",x"BA",x"95",x"77",x"51",x"51",x"7C",x"95",x"B6",
		x"AC",x"82",x"69",x"48",x"64",x"82",x"A3",x"B6",x"95",x"77",x"56",x"35",x"31",x"51",x"72",x"95",
		x"8B",x"6E",x"4D",x"60",x"82",x"9E",x"BA",x"99",x"7C",x"5B",x"48",x"72",x"8B",x"B1",x"B1",x"87",
		x"6E",x"48",x"56",x"80",x"95",x"82",x"69",x"82",x"95",x"7C",x"6E",x"87",x"A7",x"C4",x"BA",x"9E",
		x"7C",x"80",x"A7",x"BF",x"C4",x"A7",x"87",x"64",x"4D",x"69",x"90",x"99",x"80",x"56",x"3A",x"14",
		x"19",x"43",x"64",x"5B",x"3A",x"48",x"3F",x"31",x"3F",x"5B",x"72",x"48",x"48",x"51",x"3F",x"1E",
		x"22",x"48",x"69",x"64",x"3F",x"22",x"35",x"60",x"7C",x"9E",x"B1",x"95",x"77",x"51",x"4D",x"6E",
		x"90",x"8B",x"69",x"4D",x"2C",x"0B",x"1E",x"43",x"64",x"80",x"69",x"43",x"31",x"5B",x"77",x"99",
		x"9E",x"7C",x"5B",x"60",x"64",x"4D",x"56",x"69",x"60",x"4D",x"60",x"72",x"9E",x"A7",x"8B",x"6E",
		x"60",x"87",x"82",x"80",x"99",x"8B",x"80",x"5B",x"3F",x"51",x"77",x"8B",x"80",x"87",x"80",x"72",
		x"56",x"31",x"31",x"5B",x"7C",x"77",x"51",x"31",x"43",x"64",x"87",x"B1",x"C4",x"A7",x"82",x"60",
		x"56",x"72",x"9E",x"99",x"90",x"A7",x"C8",x"E9",x"DB",x"B1",x"8B",x"72",x"87",x"AC",x"D2",x"E0",
		x"C4",x"95",x"90",x"B1",x"CD",x"D2",x"A7",x"B1",x"B1",x"B1",x"BA",x"B1",x"B6",x"AC",x"A7",x"AC",
		x"B1",x"C4",x"C8",x"B6",x"95",x"72",x"72",x"95",x"BA",x"D7",x"C8",x"A3",x"7C",x"64",x"7C",x"9E",
		x"C4",x"D2",x"B6",x"87",x"82",x"A3",x"C4",x"D2",x"CD",x"BF",x"99",x"77",x"5B",x"69",x"90",x"B6",
		x"C8",x"AC",x"82",x"60",x"56",x"77",x"9E",x"9E",x"7C",x"56",x"35",x"43",x"69",x"90",x"A7",x"90",
		x"69",x"43",x"3A",x"56",x"80",x"99",x"BF",x"BF",x"95",x"7C",x"51",x"64",x"82",x"72",x"7C",x"77",
		x"69",x"5B",x"6E",x"72",x"72",x"77",x"87",x"8B",x"7C",x"5B",x"60",x"64",x"48",x"31",x"3F",x"6E",
		x"80",x"72",x"77",x"72",x"60",x"5B",x"6E",x"87",x"8B",x"6E",x"48",x"27",x"31",x"56",x"80",x"99",
		x"82",x"60",x"3A",x"2C",x"3A",x"35",x"43",x"51",x"5B",x"48",x"27",x"2C",x"51",x"7C",x"95",x"B6",
		x"9E",x"7C",x"60",x"43",x"69",x"82",x"A7",x"B6",x"8B",x"72",x"4D",x"4D",x"77",x"90",x"B6",x"A3",
		x"80",x"64",x"43",x"64",x"82",x"A3",x"B6",x"90",x"77",x"4D",x"4D",x"72",x"95",x"8B",x"87",x"87",
		x"80",x"82",x"90",x"9E",x"95",x"7C",x"69",x"82",x"A7",x"AC",x"A3",x"A7",x"99",x"8B",x"69",x"77",
		x"95",x"B1",x"9E",x"80",x"60",x"48",x"64",x"80",x"A3",x"B1",x"90",x"72",x"51",x"27",x"31",x"51",
		x"77",x"99",x"87",x"69",x"4D",x"64",x"82",x"9E",x"CD",x"D7",x"B6",x"95",x"6E",x"4D",x"4D",x"72",
		x"95",x"B1",x"A7",x"82",x"60",x"43",x"60",x"82",x"A3",x"B6",x"8B",x"72",x"4D",x"4D",x"72",x"90",
		x"B1",x"D2",x"D7",x"BF",x"9E",x"82",x"95",x"BA",x"D2",x"C8",x"A7",x"8B",x"69",x"60",x"82",x"9E",
		x"C4",x"BA",x"95",x"77",x"87",x"AC",x"C4",x"A7",x"95",x"9E",x"95",x"A3",x"9E",x"9E",x"9E",x"95",
		x"95",x"99",x"A3",x"B6",x"AC",x"95",x"77",x"5B",x"72",x"95",x"AC",x"AC",x"8B",x"72",x"4D",x"48",
		x"6E",x"87",x"AC",x"A3",x"80",x"60",x"72",x"99",x"AC",x"B1",x"A7",x"8B",x"6E",x"4D",x"3F",x"64",
		x"80",x"A3",x"9E",x"80",x"60",x"3F",x"4D",x"72",x"8B",x"77",x"51",x"31",x"1E",x"43",x"60",x"87",
		x"8B",x"69",x"4D",x"27",x"31",x"56",x"77",x"95",x"B1",x"9E",x"7C",x"60",x"43",x"69",x"72",x"69",
		x"6E",x"64",x"51",x"51",x"69",x"64",x"64",x"77",x"82",x"7C",x"64",x"51",x"5B",x"51",x"35",x"2C",
		x"48",x"6E",x"72",x"6E",x"6E",x"64",x"56",x"56",x"6E",x"8B",x"77",x"51",x"35",x"19",x"3F",x"60",
		x"82",x"90",x"6E",x"4D",x"2C",x"2C",x"35",x"35",x"43",x"51",x"51",x"3A",x"1E",x"3A",x"64",x"80",
		x"A3",x"AC",x"90",x"72",x"48",x"4D",x"6E",x"90",x"B6",x"9E",x"82",x"5B",x"43",x"60",x"7C",x"A7",
		x"B1",x"90",x"77",x"48",x"4D",x"6E",x"8B",x"B6",x"A3",x"87",x"60",x"43",x"5B",x"80",x"90",x"87",
		x"8B",x"82",x"80",x"87",x"99",x"9E",x"87",x"6E",x"6E",x"95",x"B6",x"A3",x"A7",x"A3",x"95",x"80",
		x"69",x"87",x"A7",x"B6",x"95",x"72",x"4D",x"4D",x"72",x"95",x"B6",x"A7",x"82",x"60",x"43",x"27",
		x"48",x"69",x"87",x"99",x"77",x"56",x"51",x"72",x"99",x"B6",x"D7",x"CD",x"A3",x"87",x"64",x"4D",
		x"60",x"82",x"A3",x"B6",x"95",x"77",x"56",x"51",x"72",x"8B",x"B1",x"A7",x"87",x"69",x"4D",x"60",
		x"80",x"99",x"C4",x"DB",x"D2",x"BA",x"8B",x"87",x"A7",x"C8",x"D7",x"BF",x"A3",x"80",x"5B",x"72",
		x"8B",x"B6",x"CD",x"B1",x"8B",x"7C",x"95",x"BA",x"C4",x"95",x"9E",x"9E",x"99",x"A7",x"9E",x"A3",
		x"9E",x"95",x"99",x"9E",x"B1",x"BA",x"A7",x"90",x"64",x"64",x"80",x"A3",x"B6",x"A3",x"87",x"64",
		x"43",x"5B",x"77",x"9E",x"B1",x"99",x"77",x"69",x"82",x"A3",x"B6",x"B1",x"A3",x"82",x"64",x"3F",
		x"4D",x"72",x"99",x"AC",x"95",x"72",x"4D",x"3F",x"5B",x"87",x"87",x"69",x"48",x"1E",x"31",x"4D",
		x"77",x"95",x"80",x"64",x"3A",x"27",x"43",x"64",x"87",x"AC",x"B6",x"90",x"6E",x"48",x"51",x"72",
		x"69",x"6E",x"6E",x"60",x"4D",x"60",x"6E",x"64",x"6E",x"7C",x"82",x"72",x"51",x"56",x"60",x"43",
		x"2C",x"31",x"60",x"7C",x"6E",x"72",x"6E",x"5B",x"51",x"60",x"82",x"87",x"69",x"4D",x"22",x"2C",
		x"4D",x"72",x"95",x"80",x"69",x"3A",x"27",x"3A",x"31",x"3F",x"4D",x"56",x"4D",x"27",x"27",x"4D",
		x"6E",x"95",x"B1",x"A7",x"82",x"60",x"43",x"5B",x"80",x"A3",x"B6",x"99",x"72",x"4D",x"48",x"6E",
		x"90",x"B1",x"AC",x"87",x"64",x"48",x"56",x"80",x"A3",x"B6",x"9E",x"7C",x"51",x"4D",x"69",x"95",
		x"8B",x"8B",x"8B",x"80",x"82",x"8B",x"9E",x"99",x"80",x"69",x"80",x"A7",x"B1",x"A3",x"AC",x"9E",
		x"90",x"72",x"72",x"90",x"B6",x"AC",x"82",x"69",x"43",x"60",x"82",x"A3",x"BA",x"95",x"77",x"5B",
		x"35",x"31",x"56",x"72",x"95",x"90",x"6E",x"4D",x"60",x"87",x"A3",x"C4",x"D7",x"BF",x"99",x"77",
		x"51",x"4D",x"72",x"95",x"B6",x"AC",x"87",x"64",x"48",x"5B",x"82",x"A7",x"BA",x"9E",x"7C",x"56",
		x"4D",x"6E",x"90",x"B1",x"D2",x"DB",x"C8",x"A7",x"82",x"95",x"BF",x"D7",x"D2",x"B1",x"90",x"6E",
		x"60",x"82",x"9E",x"C4",x"C4",x"99",x"80",x"82",x"A7",x"C8",x"B1",x"95",x"A3",x"99",x"A3",x"A7",
		x"A3",x"A3",x"99",x"99",x"9E",x"A3",x"B6",x"B6",x"99",x"80",x"60",x"72",x"95",x"B1",x"B6",x"95",
		x"77",x"51",x"43",x"6E",x"87",x"AC",x"AC",x"82",x"64",x"6E",x"90",x"B1",x"B1",x"B1",x"95",x"72",
		x"51",x"3A",x"64",x"80",x"A3",x"A7",x"82",x"64",x"3F",x"48",x"72",x"8B",x"80",x"5B",x"35",x"22",
		x"3A",x"60",x"87",x"90",x"77",x"51",x"2C",x"2C",x"51",x"77",x"95",x"B6",x"A7",x"80",x"64",x"43",
		x"69",x"77",x"69",x"72",x"69",x"56",x"51",x"64",x"69",x"69",x"72",x"82",x"80",x"69",x"51",x"5B",
		x"56",x"3A",x"27",x"43",x"72",x"77",x"6E",x"72",x"69",x"56",x"56",x"6E",x"8B",x"82",x"60",x"3A",
		x"1E",x"35",x"60",x"82",x"95",x"77",x"56",x"2C",x"31",x"3A",x"35",x"43",x"56",x"51",x"3F",x"22",
		x"3A",x"60",x"7C",x"A3",x"B1",x"95",x"77",x"51",x"4D",x"72",x"8B",x"B1",x"A7",x"87",x"69",x"48",
		x"5B",x"80",x"9E",x"B6",x"99",x"7C",x"56",x"4D",x"6E",x"87",x"AC",x"AC",x"8B",x"6E",x"4D",x"5B",
		x"80",x"95",x"8B",x"90",x"87",x"80",x"87",x"99",x"9E",x"90",x"6E",x"6E",x"90",x"AC",x"A7",x"A7",
		x"A7",x"99",x"82",x"69",x"80",x"A7",x"BA",x"99",x"80",x"51",x"4D",x"6E",x"8B",x"B6",x"AC",x"8B",
		x"69",x"43",x"2C",x"3F",x"64",x"8B",x"99",x"82",x"5B",x"51",x"72",x"90",x"B6",x"D7",x"D7",x"AC",
		x"87",x"69",x"48",x"60",x"82",x"9E",x"BA",x"99",x"7C",x"5B",x"48",x"48",x"43",x"43",x"4D",x"56",
		x"56",x"4D",x"51",x"60",x"56",x"4D",x"5B",x"60",x"5B",x"4D",x"43",x"56",x"6E",x"90",x"BA",x"B1",
		x"90",x"72",x"4D",x"60",x"7C",x"A3",x"BF",x"A3",x"82",x"6E",x"8B",x"95",x"87",x"A3",x"9E",x"90",
		x"72",x"77",x"95",x"B6",x"AC",x"80",x"6E",x"77",x"77",x"77",x"72",x"6E",x"77",x"77",x"72",x"72",
		x"7C",x"80",x"90",x"90",x"7C",x"60",x"3A",x"51",x"77",x"95",x"AC",x"8B",x"72",x"4D",x"48",x"69",
		x"87",x"A7",x"A3",x"82",x"64",x"43",x"56",x"77",x"95",x"B1",x"95",x"77",x"56",x"48",x"69",x"87",
		x"A7",x"AC",x"87",x"6E",x"48",x"22",x"3A",x"56",x"82",x"99",x"82",x"60",x"4D",x"6E",x"87",x"AC",
		x"B6",x"90",x"77",x"51",x"5B",x"7C",x"99",x"BA",x"A7",x"87",x"64",x"4D",x"69",x"8B",x"9E",x"77",
		x"72",x"95",x"95",x"6E",x"7C",x"95",x"BA",x"DB",x"C8",x"A3",x"87",x"9E",x"BF",x"E0",x"F3",x"CD",
		x"B1",x"87",x"82",x"A3",x"C8",x"C4",x"99",x"7C",x"5B",x"3F",x"51",x"72",x"8B",x"72",x"60",x"72",
		x"5B",x"5B",x"69",x"87",x"8B",x"64",x"6E",x"72",x"56",x"3A",x"4D",x"72",x"87",x"77",x"51",x"3F",
		x"60",x"82",x"9E",x"C4",x"C4",x"A3",x"82",x"64",x"69",x"8B",x"AC",x"99",x"72",x"56",x"35",x"22",
		x"3F",x"60",x"82",x"8B",x"72",x"4D",x"48",x"72",x"90",x"B6",x"A7",x"80",x"64",x"77",x"69",x"5B",
		x"6E",x"7C",x"64",x"60",x"72",x"87",x"B6",x"AC",x"90",x"6E",x"77",x"95",x"87",x"90",x"A3",x"90",
		x"82",x"56",x"48",x"64",x"87",x"90",x"87",x"90",x"80",x"72",x"51",x"35",x"43",x"69",x"82",x"6E",
		x"48",x"3A",x"51",x"7C",x"99",x"BA",x"C4",x"99",x"80",x"5B",x"64",x"87",x"A3",x"95",x"7C",x"8B",
		x"AC",x"C8",x"A3",x"90",x"B6",x"BF",x"95",x"90",x"B6",x"B6",x"8B",x"72",x"77",x"99",x"BF",x"E0",
		x"FC",x"DB",x"B6",x"95",x"80",x"A3",x"BF",x"E5",x"E9",x"BF",x"9E",x"9E",x"C4",x"B6",x"BA",x"CD",
		x"C4",x"A3",x"90",x"A3",x"CD",x"D7",x"BA",x"95",x"90",x"95",x"8B",x"90",x"87",x"8B",x"90",x"8B",
		x"82",x"8B",x"8B",x"9E",x"A7",x"99",x"82",x"56",x"51",x"72",x"90",x"BA",x"B1",x"90",x"72",x"48",
		x"60",x"7C",x"A3",x"BF",x"9E",x"82",x"56",x"4D",x"6E",x"87",x"B6",x"B1",x"90",x"72",x"48",x"56",
		x"77",x"99",x"BA",x"9E",x"82",x"5B",x"35",x"27",x"43",x"6E",x"90",x"95",x"77",x"4D",x"56",x"77",
		x"95",x"BA",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",x"77",x"4D",x"4D",x"6E",x"90",
		x"87",x"69",x"77",x"90",x"80",x"64",x"7C",x"9E",x"C4",x"C8",x"AC",x"80",x"7C",x"99",x"B6",x"C8",
		x"B1",x"95",x"6E",x"51",x"60",x"87",x"9E",x"82",x"69",x"3F",x"1E",x"14",x"35",x"60",x"60",x"3A",
		x"43",x"43",x"31",x"3A",x"51",x"72",x"56",x"43",x"51",x"48",x"27",x"1E",x"43",x"69",x"6E",x"4D",
		x"22",x"2C",x"51",x"72",x"99",x"B1",x"A3",x"7C",x"56",x"43",x"5B",x"87",x"90",x"77",x"56",x"2C",
		x"0B",x"10",x"35",x"60",x"80",x"72",x"4D",x"31",x"4D",x"69",x"95",x"A3",x"82",x"64",x"5B",x"69",
		x"4D",x"51",x"69",x"64",x"51",x"56",x"6E",x"8B",x"AC",x"90",x"6E",x"5B",x"77",x"82",x"7C",x"90",
		x"90",x"80",x"64",x"3F",x"48",x"72",x"8B",x"80",x"82",x"82",x"72",x"64",x"35",x"2C",x"48",x"6E",
		x"77",x"5B",x"35",x"35",x"60",x"80",x"9E",x"BA",x"AC",x"8B",x"69",x"51",x"6E",x"8B",x"A3",x"7C",
		x"77",x"90",x"B1",x"B6",x"90",x"95",x"B6",x"AC",x"87",x"99",x"B6",x"A3",x"80",x"69",x"87",x"A7",
		x"C4",x"E9",x"EE",x"C8",x"AC",x"87",x"87",x"AC",x"C8",x"E9",x"D7",x"B1",x"90",x"B1",x"C4",x"AC",
		x"C4",x"C4",x"B6",x"95",x"90",x"B6",x"D2",x"D2",x"A7",x"82",x"90",x"8B",x"90",x"8B",x"82",x"8B",
		x"8B",x"87",x"82",x"8B",x"90",x"A3",x"A3",x"8B",x"72",x"4D",x"60",x"82",x"A3",x"BF",x"9E",x"80",
		x"5B",x"48",x"72",x"8B",x"B1",x"B6",x"8B",x"6E",x"48",x"56",x"7C",x"99",x"BA",x"9E",x"7C",x"5B",
		x"43",x"69",x"82",x"A7",x"B1",x"8B",x"6E",x"4D",x"2C",x"35",x"56",x"77",x"95",x"82",x"64",x"48",
		x"64",x"87",x"A7",x"BA",x"90",x"77",x"51",x"4D",x"77",x"90",x"B6",x"A7",x"82",x"64",x"43",x"60",
		x"82",x"95",x"7C",x"69",x"87",x"95",x"72",x"6E",x"8B",x"AC",x"C4",x"B6",x"95",x"72",x"82",x"AC",
		x"BF",x"BF",x"9E",x"80",x"5B",x"4D",x"72",x"95",x"99",x"77",x"51",x"31",x"10",x"1E",x"48",x"64",
		x"51",x"3A",x"48",x"3A",x"31",x"3F",x"60",x"6E",x"48",x"48",x"4D",x"3A",x"22",x"27",x"4D",x"6E",
		x"60",x"35",x"22",x"35",x"64",x"80",x"A3",x"B1",x"8B",x"6E",x"48",x"4D",x"72",x"90",x"8B",x"64",
		x"43",x"22",x"06",x"22",x"48",x"6E",x"80",x"60",x"3A",x"35",x"56",x"7C",x"9E",x"99",x"77",x"56",
		x"64",x"60",x"4D",x"5B",x"69",x"60",x"51",x"60",x"77",x"9E",x"A3",x"82",x"64",x"69",x"8B",x"80",
		x"82",x"95",x"87",x"7C",x"4D",x"3F",x"56",x"80",x"87",x"80",x"87",x"7C",x"6E",x"4D",x"2C",x"35",
		x"60",x"7C",x"72",x"43",x"2C",x"48",x"69",x"8B",x"B6",x"BF",x"9E",x"7C",x"56",x"56",x"7C",x"9E",
		x"95",x"72",x"82",x"A7",x"BF",x"A7",x"90",x"AC",x"BA",x"9E",x"8B",x"B1",x"B6",x"95",x"6E",x"72",
		x"90",x"B1",x"DB",x"F3",x"E5",x"BA",x"90",x"80",x"95",x"BA",x"E0",x"E9",x"C8",x"9E",x"99",x"BF",
		x"B6",x"B6",x"C8",x"C4",x"A7",x"8B",x"9E",x"BF",x"D7",x"BA",x"95",x"87",x"90",x"8B",x"90",x"87",
		x"87",x"8B",x"8B",x"87",x"87",x"8B",x"95",x"A7",x"99",x"82",x"64",x"51",x"6E",x"8B",x"B1",x"B6",
		x"90",x"77",x"51",x"5B",x"7C",x"99",x"B6",x"A3",x"82",x"64",x"4D",x"69",x"82",x"A7",x"B6",x"90",
		x"77",x"51",x"51",x"77",x"90",x"B1",x"A3",x"82",x"69",x"3F",x"27",x"43",x"60",x"8B",x"95",x"7C",
		x"56",x"51",x"77",x"90",x"B6",x"AC",x"87",x"69",x"4D",x"60",x"80",x"9E",x"B6",x"99",x"7C",x"56",
		x"4D",x"6E",x"90",x"90",x"69",x"72",x"95",x"87",x"64",x"7C",x"99",x"BF",x"C4",x"AC",x"80",x"77",
		x"95",x"B6",x"C8",x"B1",x"99",x"72",x"4D",x"60",x"80",x"99",x"87",x"64",x"4D",x"1E",x"14",x"31",
		x"56",x"64",x"3F",x"43",x"48",x"31",x"3A",x"4D",x"6E",x"5B",x"3F",x"51",x"48",x"2C",x"1E",x"35",
		x"64",x"6E",x"51",x"2C",x"2C",x"51",x"6E",x"90",x"B6",x"A3",x"87",x"60",x"43",x"5B",x"80",x"90",
		x"77",x"56",x"3A",x"10",x"10",x"35",x"56",x"80",x"72",x"56",x"35",x"48",x"69",x"8B",x"A3",x"8B",
		x"69",x"56",x"69",x"51",x"4D",x"64",x"69",x"51",x"56",x"69",x"8B",x"AC",x"9E",x"77",x"5B",x"77",
		x"8B",x"7C",x"8B",x"95",x"82",x"69",x"43",x"43",x"69",x"8B",x"82",x"82",x"82",x"77",x"64",x"3F",
		x"2C",x"43",x"6E",x"7C",x"5B",x"3A",x"35",x"56",x"80",x"99",x"BF",x"B6",x"8B",x"72",x"51",x"69",
		x"8B",x"9E",x"90",x"9E",x"B6",x"DB",x"E5",x"BA",x"9E",x"7C",x"7C",x"A3",x"BF",x"E0",x"CD",x"A3",
		x"8B",x"9E",x"C8",x"DB",x"B6",x"A7",x"B1",x"AC",x"B6",x"B6",x"B1",x"B1",x"A7",x"A7",x"B1",x"BA",
		x"C8",x"BA",x"A3",x"80",x"69",x"8B",x"A7",x"CD",x"D2",x"AC",x"90",x"6E",x"72",x"90",x"B1",x"CD",
		x"BA",x"95",x"80",x"95",x"BA",x"D2",x"CD",x"C4",x"A3",x"82",x"64",x"64",x"82",x"A3",x"C4",x"B1",
		x"90",x"72",x"56",x"6E",x"90",x"A3",x"82",x"64",x"3F",x"35",x"60",x"7C",x"A3",x"99",x"77",x"56",
		x"35",x"48",x"72",x"8B",x"AC",x"C4",x"A7",x"87",x"64",x"56",x"80",x"7C",x"77",x"7C",x"6E",x"5B",
		x"64",x"77",x"6E",x"72",x"82",x"8B",x"82",x"69",x"5B",x"64",x"56",x"3A",x"35",x"5B",x"7C",x"77",
		x"77",x"77",x"69",x"5B",x"60",x"7C",x"90",x"77",x"56",x"35",x"22",x"4D",x"69",x"90",x"90",x"69",
		x"4D",x"2C",x"35",x"35",x"3A",x"4D",x"56",x"51",x"35",x"22",x"48",x"69",x"87",x"AC",x"AC",x"8B",
		x"6E",x"4D",x"56",x"77",x"95",x"B1",x"9E",x"80",x"5B",x"48",x"64",x"82",x"A7",x"AC",x"8B",x"72",
		x"4D",x"51",x"77",x"90",x"B1",x"9E",x"82",x"60",x"48",x"60",x"82",x"90",x"87",x"8B",x"80",x"80",
		x"8B",x"99",x"99",x"82",x"64",x"72",x"95",x"AC",x"A3",x"A7",x"9E",x"90",x"77",x"69",x"82",x"AC",
		x"AC",x"8B",x"6E",x"43",x"51",x"77",x"9E",x"B1",x"A3",x"7C",x"56",x"35",x"22",x"4D",x"69",x"90",
		x"95",x"6E",x"4D",x"51",x"7C",x"99",x"BA",x"D7",x"BF",x"99",x"80",x"5B",x"48",x"69",x"82",x"A7",
		x"AC",x"8B",x"72",x"4D",x"51",x"77",x"95",x"B1",x"9E",x"80",x"60",x"48",x"60",x"82",x"9E",x"C8",
		x"DB",x"CD",x"B1",x"82",x"8B",x"A7",x"C8",x"D2",x"B6",x"99",x"72",x"56",x"77",x"90",x"BA",x"C4",
		x"A7",x"82",x"7C",x"99",x"BF",x"BA",x"90",x"9E",x"95",x"9E",x"A3",x"9E",x"9E",x"99",x"95",x"99",
		x"9E",x"B1",x"B6",x"A3",x"87",x"5B",x"69",x"82",x"A3",x"B6",x"9E",x"80",x"56",x"3F",x"60",x"77",
		x"A3",x"AC",x"90",x"6E",x"69",x"87",x"A7",x"B1",x"AC",x"99",x"7C",x"56",x"3A",x"56",x"72",x"99",
		x"AC",x"8B",x"72",x"43",x"3F",x"60",x"82",x"82",x"60",x"43",x"22",x"31",x"56",x"77",x"90",x"77",
		x"5B",x"35",x"27",x"48",x"69",x"87",x"B1",x"AC",x"8B",x"69",x"43",x"56",x"72",x"69",x"6E",x"69",
		x"5B",x"4D",x"60",x"69",x"60",x"6E",x"7C",x"82",x"6E",x"4D",x"56",x"5B",x"3F",x"22",x"35",x"60",
		x"72",x"69",x"6E",x"69",x"56",x"51",x"64",x"87",x"82",x"64",x"43",x"19",x"31",x"51",x"77",x"95",
		x"77",x"60",x"31",x"27",x"35",x"31",x"3F",x"51",x"56",x"43",x"22",x"2C",x"51",x"72",x"99",x"B1",
		x"9E",x"7C",x"56",x"43",x"60",x"82",x"A7",x"B1",x"90",x"69",x"48",x"4D",x"72",x"95",x"B1",x"A3",
		x"80",x"5B",x"43",x"60",x"82",x"A7",x"B1",x"95",x"6E",x"4D",x"4D",x"6E",x"95",x"87",x"8B",x"87",
		x"80",x"82",x"90",x"9E",x"90",x"77",x"69",x"87",x"AC",x"AC",x"A3",x"A7",x"99",x"8B",x"6E",x"77",
		x"99",x"B6",x"9E",x"7C",x"60",x"43",x"69",x"82",x"A7",x"B1",x"8B",x"6E",x"51",x"2C",x"35",x"5B",
		x"7C",x"95",x"87",x"64",x"4D",x"69",x"8B",x"A7",x"CD",x"D7",x"B6",x"95",x"77",x"48",x"56",x"72",
		x"95",x"BA",x"A3",x"87",x"60",x"48",x"64",x"80",x"AC",x"B6",x"95",x"7C",x"4D",x"51",x"72",x"90",
		x"B6",x"D7",x"DB",x"C4",x"99",x"82",x"95",x"BF",x"D7",x"CD",x"B1",x"87",x"64",x"60",x"82",x"A7",
		x"C8",x"BF",x"99",x"77",x"87",x"A7",x"C4",x"A7",x"95",x"A3",x"99",x"A7",x"A3",x"A3",x"9E",x"99",
		x"99",x"9E",x"A7",x"BA",x"AC",x"95",x"77",x"5B",x"7C",x"99",x"B1",x"B1",x"8B",x"72",x"48",x"48",
		x"72",x"8B",x"B1",x"A3",x"7C",x"64",x"72",x"99",x"B6",x"B1",x"AC",x"8B",x"6E",x"48",x"3F",x"69",
		x"82",x"AC",x"A3",x"7C",x"60",x"3F",x"51",x"7C",x"8B",x"7C",x"51",x"2C",x"22",x"43",x"69",x"8B",
		x"8B",x"6E",x"48",x"27",x"31",x"5B",x"80",x"99",x"BA",x"9E",x"7C",x"5B",x"43",x"6E",x"72",x"69",
		x"72",x"64",x"51",x"51",x"69",x"64",x"69",x"77",x"82",x"80",x"60",x"51",x"5B",x"51",x"35",x"27",
		x"4D",x"77",x"72",x"6E",x"72",x"64",x"56",x"5B",x"77",x"8B",x"7C",x"56",x"31",x"1E",x"3F",x"64",
		x"87",x"90",x"72",x"4D",x"27",x"31",x"35",x"35",x"48",x"56",x"51",x"35",x"22",x"3A",x"64",x"82",
		x"A7",x"B1",x"8B",x"72",x"4D",x"4D",x"77",x"90",x"B6",x"A3",x"80",x"60",x"43",x"64",x"82",x"A3",
		x"B6",x"90",x"77",x"51",x"4D",x"77",x"90",x"B6",x"A7",x"82",x"64",x"48",x"5B",x"87",x"95",x"87",
		x"90",x"82",x"82",x"87",x"9E",x"9E",x"8B",x"72",x"72",x"95",x"B1",x"A7",x"A7",x"A3",x"95",x"7C",
		x"69",x"82",x"AC",x"B6",x"90",x"77",x"48",x"56",x"72",x"95",x"BA",x"A3",x"87",x"64",x"3A",x"27",
		x"43",x"6E",x"90",x"99",x"7C",x"51",x"56",x"77",x"95",x"BF",x"DB",x"CD",x"A3",x"82",x"64",x"48",
		x"64",x"87",x"A7",x"BA",x"90",x"77",x"51",x"4D",x"77",x"90",x"B6",x"A7",x"82",x"64",x"48",x"60",
		x"82",x"A3",x"C4",x"DB",x"D2",x"B6",x"90",x"8B",x"AC",x"CD",x"D7",x"BF",x"9E",x"80",x"60",x"72",
		x"90",x"B6",x"C8",x"AC",x"87",x"7C",x"99",x"BF",x"C4",x"99",x"9E",x"9E",x"99",x"A7",x"9E",x"A3",
		x"9E",x"99",x"99",x"9E",x"AC",x"BA",x"A7",x"8B",x"69",x"64",x"82",x"A3",x"B6",x"A3",x"82",x"64",
		x"48",x"5B",x"7C",x"9E",x"B1",x"95",x"72",x"64",x"87",x"A7",x"B6",x"B1",x"9E",x"80",x"60",x"43",
		x"51",x"72",x"90",x"AC",x"90",x"77",x"51",x"43",x"60",x"82",x"8B",x"64",x"48",x"22",x"2C",x"56",
		x"72",x"95",x"80",x"5B",x"3A",x"22",x"43",x"69",x"82",x"A7",x"B1",x"90",x"72",x"4D",x"51",x"77",
		x"6E",x"6E",x"6E",x"60",x"4D",x"60",x"6E",x"64",x"6E",x"80",x"87",x"72",x"51",x"56",x"60",x"43",
		x"27",x"35",x"60",x"77",x"6E",x"72",x"6E",x"5B",x"56",x"64",x"80",x"87",x"69",x"48",x"27",x"2C",
		x"51",x"72",x"90",x"80",x"64",x"3F",x"2C",x"3A",x"35",x"3F",x"51",x"56",x"48",x"2C",x"2C",x"51",
		x"6E",x"90",x"B6",x"A3",x"82",x"60",x"43",x"60",x"7C",x"A7",x"B6",x"95",x"77",x"4D",x"4D",x"6E",
		x"90",x"B6",x"A7",x"87",x"64",x"43",x"60",x"7C",x"A3",x"B6",x"95",x"7C",x"4D",x"4D",x"6E",x"90",
		x"8B",x"8B",x"8B",x"80",x"82",x"90",x"9E",x"95",x"7C",x"69",x"7C",x"A7",x"B1",x"A3",x"AC",x"99",
		x"90",x"6E",x"72",x"99",x"B6",x"AC",x"82",x"60",x"48",x"60",x"82",x"A7",x"B6",x"99",x"72",x"56",
		x"31",x"31",x"5B",x"77",x"99",x"90",x"69",x"4D",x"60",x"87",x"A7",x"C8",x"DB",x"BA",x"95",x"7C",
		x"56",x"51",x"72",x"90",x"B1",x"AC",x"87",x"69",x"48",x"48",x"48",x"48",x"95",x"A7",x"9E",x"A3",
		x"9E",x"9E",x"9E",x"9E",x"9E",x"9E",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"8B",x"8B",
		x"8B",x"8B",x"8B",x"8B",x"8B",x"8B",x"8B",x"8B",x"8B",x"87",x"87",x"87",x"87",x"87",x"87",x"87",
		x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",
		x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",x"7C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
	);

begin
	process (ROM_A)
	begin
		if (ROM_nCS='1') or (ROM_nOE='1') then
			ROM_D <= (others => 'Z');
		else
			ROM_D <= my_rom(conv_integer(ROM_A)) after 10 ns;
		end if;
	end process;
end architecture behavioral;
