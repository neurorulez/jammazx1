library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic23 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic23 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"58",X"14",X"6D",X"FA",X"F0",X"E0",X"90",
		X"0B",X"31",X"99",X"09",X"EB",X"FA",X"58",X"3F",X"10",X"10",X"90",X"70",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"08",X"08",X"04",X"FF",X"FF",X"FF",X"7E",X"3F",X"1C",X"88",X"E4",
		X"E0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4A",X"0F",X"1F",X"3E",X"F4",X"D2",X"80",X"00",X"83",X"2B",X"3F",X"7E",X"F4",X"90",X"02",
		X"06",X"07",X"37",X"53",X"B8",X"D8",X"24",X"D0",X"21",X"5C",X"39",X"2A",X"7C",X"EC",X"E2",X"40",
		X"00",X"8A",X"AD",X"FF",X"FF",X"66",X"29",X"04",X"90",X"40",X"91",X"7F",X"FF",X"EA",X"10",X"40",
		X"9A",X"7C",X"3D",X"98",X"32",X"38",X"1C",X"18",X"24",X"1C",X"38",X"10",X"39",X"5C",X"BA",X"10",
		X"3E",X"99",X"FE",X"E0",X"16",X"C0",X"20",X"00",X"06",X"0F",X"1F",X"3E",X"7D",X"FB",X"F0",X"47",
		X"02",X"30",X"0C",X"8E",X"1F",X"E1",X"BC",X"78",X"76",X"ED",X"BD",X"7F",X"D7",X"C9",X"E4",X"71",
		X"09",X"03",X"66",X"1F",X"BA",X"64",X"58",X"30",X"E3",X"F1",X"F8",X"7C",X"7E",X"3F",X"1F",X"07",
		X"17",X"1F",X"FF",X"7F",X"3F",X"9F",X"8F",X"C7",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",
		X"80",X"E2",X"F4",X"5D",X"1E",X"0A",X"2A",X"10",X"08",X"62",X"78",X"BE",X"5F",X"0B",X"41",X"00",
		X"24",X"4E",X"BC",X"72",X"3E",X"77",X"65",X"20",X"40",X"12",X"38",X"3C",X"9C",X"18",X"21",X"00",
		X"02",X"10",X"44",X"18",X"31",X"80",X"08",X"40",X"20",X"04",X"50",X"12",X"08",X"24",X"01",X"10",
		X"00",X"09",X"00",X"40",X"00",X"02",X"20",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"FC",X"FF",X"F8",X"E0",X"C0",X"80",X"C0",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"C0",
		X"C0",X"C0",X"E0",X"F0",X"F0",X"E0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"00",X"00",
		X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",X"08",X"08",X"1C",X"7F",X"1C",X"08",X"08",X"00",
		X"44",X"AA",X"AA",X"01",X"01",X"AA",X"AA",X"44",X"44",X"AA",X"82",X"01",X"01",X"82",X"AA",X"44",
		X"44",X"82",X"82",X"01",X"01",X"82",X"82",X"44",X"40",X"80",X"80",X"00",X"00",X"80",X"80",X"00",
		X"3C",X"6E",X"EF",X"EF",X"EF",X"EF",X"6E",X"3C",X"3C",X"66",X"E7",X"E7",X"E7",X"E7",X"66",X"3C",
		X"3C",X"66",X"C3",X"C3",X"C3",X"C3",X"66",X"3C",X"E8",X"D0",X"F0",X"5E",X"70",X"30",X"30",X"10",
		X"E8",X"C8",X"E4",X"C3",X"E3",X"C4",X"E8",X"C8",X"10",X"30",X"30",X"70",X"7E",X"D0",X"F0",X"C8",
		X"73",X"06",X"04",X"0C",X"1E",X"30",X"7C",X"C0",X"18",X"18",X"70",X"00",X"00",X"70",X"18",X"18",
		X"C0",X"7C",X"30",X"1E",X"0C",X"04",X"06",X"73",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"C5",X"AB",X"AD",X"9D",X"9C",X"B4",X"B4",X"F0",X"F0",X"B4",X"B4",X"9C",X"9D",X"AD",X"AB",X"C5",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"E0",X"E0",X"80",X"84",X"48",X"30",X"1F",X"30",X"48",X"84",
		X"18",X"24",X"24",X"24",X"24",X"24",X"24",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"F0",X"F8",X"3F",X"00",X"00",X"00",X"00",X"00",X"02",X"3C",X"CC",X"14",X"24",X"48",X"88",
		X"FF",X"FF",X"C1",X"80",X"80",X"00",X"00",X"00",X"08",X"08",X"08",X"0C",X"8F",X"8E",X"C6",X"FF",
		X"08",X"08",X"D0",X"E0",X"78",X"1E",X"00",X"00",X"C0",X"80",X"80",X"E0",X"1B",X"0C",X"34",X"C4",
		X"FF",X"FF",X"C3",X"81",X"80",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"83",X"83",X"C7",X"FF",
		X"FF",X"08",X"10",X"20",X"C0",X"C0",X"60",X"30",X"00",X"30",X"60",X"C0",X"C0",X"A0",X"10",X"08",
		X"FF",X"FF",X"C7",X"83",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"83",X"C7",X"FF",
		X"C0",X"00",X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"00",X"C0",X"FF",
		X"1F",X"7E",X"3C",X"78",X"F0",X"FC",X"00",X"00",X"00",X"FC",X"F0",X"78",X"3C",X"FE",X"1F",X"FF",
		X"1C",X"3E",X"7F",X"1F",X"7F",X"3E",X"1C",X"00",X"00",X"60",X"70",X"FF",X"70",X"60",X"00",X"00",
		X"00",X"00",X"7E",X"07",X"7E",X"00",X"00",X"00",X"00",X"E0",X"F0",X"A0",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"F8",X"F4",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"80",X"10",X"00",X"00",X"00",X"0C",X"0E",X"5F",X"FB",X"B9",X"C8",X"E4",X"60",
		X"00",X"0C",X"0E",X"2F",X"7F",X"7E",X"F2",X"FF",X"D0",X"A0",X"08",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F0",X"D0",X"40",X"20",X"00",X"00",X"00",X"30",X"78",X"68",X"C0",X"40",X"00",X"00",X"00",
		X"1E",X"3E",X"7F",X"FF",X"F5",X"F2",X"6A",X"B0",X"00",X"1C",X"3E",X"7F",X"7F",X"7A",X"FA",X"F0",
		X"00",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"2A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"DC",X"08",X"00",X"00",
		X"00",X"00",X"00",X"1C",X"DC",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"57",X"07",X"57",X"07",X"57",X"07",X"56",X"FC",X"55",X"00",X"55",X"00",X"55",X"00",X"55",X"FF",
		X"01",X"03",X"FF",X"FF",X"57",X"07",X"57",X"07",X"00",X"00",X"FF",X"FF",X"55",X"00",X"55",X"00",
		X"00",X"00",X"FC",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"AA",X"00",X"00",X"00",X"00",X"FF",X"00",X"2A",X"00",X"54",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"04",X"04",X"06",X"06",X"07",X"07",X"00",X"00",
		X"FF",X"FC",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FC",
		X"FF",X"6F",X"C7",X"07",X"0F",X"1F",X"3E",X"00",X"00",X"00",X"3E",X"1F",X"0F",X"07",X"C7",X"6F",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"79",X"00",X"F0",X"00",X"00",X"00",X"00",X"F8",X"00",X"F8",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"80",X"80",X"C0",X"E0",X"C0",X"80",X"80",X"00",X"80",X"80",X"C4",X"EE",X"C4",X"80",X"80",
		X"00",X"80",X"80",X"CE",X"EE",X"CE",X"80",X"80",X"00",X"80",X"8E",X"DF",X"FF",X"DF",X"8E",X"80",
		X"FE",X"88",X"88",X"90",X"E0",X"80",X"80",X"00",X"00",X"00",X"80",X"80",X"E0",X"90",X"88",X"88",
		X"3F",X"08",X"08",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"08",X"08",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",
		X"03",X"0C",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"30",X"C0",
		X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",
		X"00",X"00",X"00",X"00",X"C0",X"30",X"0C",X"03",X"C0",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",
		X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"C0",X"80",X"80",X"80",X"00",X"E0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",X"C0",
		X"80",X"80",X"80",X"C0",X"E0",X"C0",X"80",X"80",X"A0",X"F0",X"60",X"C0",X"80",X"80",X"80",X"00",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"60",X"F0",X"60",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"60",X"F0",X"A0",X"F0",X"80",X"C0",X"60",X"F0",X"A0",X"F0",X"60",X"C0",
		X"60",X"F0",X"A0",X"F0",X"60",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",
		X"E0",X"70",X"78",X"EE",X"B8",X"EE",X"78",X"70",X"78",X"EE",X"B8",X"EE",X"78",X"70",X"E0",X"C0",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"70",X"B8",X"EE",X"78",X"70",X"E0",X"C0",X"C0",X"80",
		X"80",X"80",X"C0",X"C0",X"E0",X"70",X"78",X"EE",X"78",X"70",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"C0",X"C0",X"E0",X"70",X"78",X"EE",X"B8",X"EE",X"70",X"5E",X"E0",X"E0",X"C0",X"C0",X"80",X"80",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"5E",X"03",X"07",X"03",X"01",X"03",X"01",X"03",X"03",
		X"03",X"03",X"03",X"01",X"03",X"01",X"03",X"07",X"7F",X"70",X"7F",X"D0",X"F8",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"D0",X"1E",X"0F",X"1E",X"0C",X"07",X"03",X"0F",X"07",
		X"0E",X"07",X"0F",X"07",X"0F",X"03",X"07",X"0C",X"18",X"0C",X"18",X"0C",X"07",X"03",X"0F",X"07",
		X"F0",X"FF",X"D0",X"F8",X"E0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"F0",X"A0",X"FE",
		X"3C",X"1E",X"3C",X"1D",X"0F",X"07",X"0F",X"03",X"18",X"3C",X"1C",X"3E",X"1F",X"3F",X"0F",X"19",
		X"F0",X"FE",X"A0",X"F0",X"80",X"00",X"00",X"00",X"80",X"80",X"80",X"C0",X"E0",X"F8",X"D0",X"FF",
		X"3C",X"19",X"0F",X"3F",X"1F",X"3E",X"1C",X"3C",X"07",X"03",X"0F",X"07",X"0F",X"1D",X"3C",X"1E",
		X"D0",X"F8",X"E0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"80",X"F0",X"A0",X"FE",X"F0",X"FF",
		X"3C",X"1D",X"0F",X"07",X"0F",X"03",X"07",X"03",X"1C",X"3E",X"1F",X"3F",X"0F",X"19",X"3C",X"1E",
		X"A0",X"F0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F8",X"D0",X"FF",X"F0",X"FE",
		X"0F",X"3F",X"1F",X"3E",X"1C",X"3C",X"18",X"38",X"0F",X"07",X"0F",X"1D",X"3C",X"1E",X"3C",X"19",
		X"80",X"F0",X"A0",X"FE",X"F0",X"FF",X"D0",X"F8",X"0F",X"07",X"0F",X"03",X"07",X"03",X"07",X"03",
		X"1F",X"3F",X"0F",X"19",X"3C",X"1E",X"3C",X"1D",X"E0",X"F8",X"D0",X"FF",X"F0",X"FE",X"A0",X"F0",
		X"1F",X"3E",X"1C",X"3C",X"18",X"38",X"30",X"70",X"0F",X"1D",X"3C",X"1E",X"3C",X"19",X"0F",X"3F",
		X"A0",X"FE",X"F0",X"FF",X"D0",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",
		X"0F",X"19",X"3C",X"1E",X"3C",X"1D",X"0F",X"07",X"30",X"38",X"18",X"3C",X"1C",X"3E",X"1F",X"3F",
		X"D0",X"FF",X"F0",X"FE",X"A0",X"F0",X"80",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"E0",X"F8",
		X"3C",X"1E",X"3C",X"19",X"0F",X"3F",X"1F",X"3E",X"07",X"03",X"07",X"03",X"0F",X"07",X"0F",X"1D",
		X"30",X"B0",X"E0",X"E0",X"C0",X"E0",X"F8",X"D0",X"90",X"A0",X"F0",X"E0",X"E0",X"E0",X"F8",X"D0",
		X"A4",X"EC",X"C8",X"90",X"AC",X"08",X"98",X"50",X"C4",X"8C",X"A8",X"14",X"3C",X"64",X"5C",X"98",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"06",X"06",X"0A",X"0A",X"12",X"34",X"08",X"0A",X"0F",X"0F",X"0E",X"0E",X"0E",X"06",
		X"03",X"07",X"0D",X"2A",X"3A",X"3A",X"76",X"D6",X"08",X"09",X"0E",X"0F",X"0F",X"0E",X"0C",X"06",
		X"48",X"6C",X"3C",X"1C",X"1E",X"0E",X"06",X"02",X"00",X"80",X"80",X"60",X"30",X"98",X"90",X"D8",
		X"8E",X"C6",X"44",X"56",X"72",X"2B",X"0B",X"06",X"00",X"80",X"E0",X"A0",X"B8",X"1C",X"1C",X"08",
		X"0A",X"01",X"0C",X"04",X"0E",X"0E",X"0D",X"0C",X"0E",X"07",X"09",X"00",X"08",X"0C",X"0D",X"0F",
		X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"03",
		X"0C",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",X"07",X"0E",X"06",X"0E",X"0C",X"0C",X"0C",
		X"08",X"08",X"0C",X"0C",X"0C",X"0C",X"0E",X"06",X"80",X"C0",X"C0",X"C0",X"60",X"60",X"60",X"70",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"07",X"03",X"07",X"03",X"03",X"03",X"03",X"03",
		X"C0",X"C0",X"60",X"60",X"60",X"70",X"30",X"38",X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",
		X"18",X"38",X"30",X"70",X"60",X"60",X"60",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"03",
		X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"60",X"60",X"60",X"70",X"30",X"38",X"18",X"3C",X"30",X"70",X"60",X"60",X"60",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"07",X"03",X"07",X"03",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"60",X"70",X"30",X"38",X"18",X"3C",X"1C",X"3E",
		X"80",X"80",X"80",X"C0",X"C0",X"C0",X"60",X"60",X"60",X"60",X"60",X"C0",X"C0",X"C0",X"80",X"80",
		X"03",X"03",X"07",X"03",X"07",X"03",X"0F",X"07",X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"0F",X"03",X"07",X"03",X"07",X"03",X"03",X"03",
		X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"1C",X"3C",X"18",X"38",X"30",X"70",X"60",X"60",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"C0",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
