library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity mayday_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of mayday_prog is
	type rom is array(0 to  28671) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"02",X"FF",X"DE",X"40",X"A7",X"44",X"AF",X"42",X"7E",X"E8",X"7D",X"9E",X"40",X"8D",X"07",X"33",
		X"84",X"7E",X"E8",X"7D",X"AE",X"06",X"34",X"46",X"CE",X"A0",X"3C",X"AC",X"C4",X"26",X"18",X"EC",
		X"84",X"ED",X"C4",X"A6",X"06",X"27",X"06",X"DC",X"46",X"9F",X"46",X"20",X"04",X"DC",X"3E",X"9F",
		X"3E",X"ED",X"84",X"30",X"C4",X"35",X"C6",X"EE",X"C4",X"26",X"E0",X"7E",X"D8",X"16",X"FE",X"34",
		X"62",X"DE",X"46",X"26",X"01",X"BD",X"D0",X"3B",X"10",X"AE",X"C4",X"10",X"9F",X"46",X"86",X"01",
		X"A7",X"46",X"A6",X"E4",X"20",X"11",X"34",X"62",X"DE",X"3E",X"26",X"03",X"BD",X"D0",X"3B",X"10",
		X"AE",X"C4",X"10",X"9F",X"3E",X"6F",X"46",X"AF",X"42",X"A7",X"45",X"86",X"01",X"A7",X"44",X"AE",
		X"9F",X"A0",X"40",X"EF",X"9F",X"A0",X"40",X"AF",X"C4",X"30",X"C4",X"35",X"E2",X"34",X"12",X"8E",
		X"A0",X"3C",X"AE",X"84",X"27",X"0E",X"9C",X"40",X"27",X"F8",X"A6",X"05",X"81",X"02",X"27",X"F2",
		X"8D",X"84",X"20",X"EE",X"35",X"92",X"8D",X"16",X"34",X"66",X"EF",X"06",X"EE",X"66",X"37",X"26",
		X"ED",X"02",X"10",X"AF",X"08",X"37",X"06",X"ED",X"88",X"12",X"EF",X"66",X"35",X"E6",X"34",X"46",
		X"9E",X"44",X"26",X"03",X"BD",X"D0",X"3B",X"EC",X"84",X"DD",X"44",X"DC",X"42",X"ED",X"84",X"4F",
		X"5F",X"ED",X"04",X"A7",X"88",X"14",X"35",X"C6",X"34",X"70",X"CE",X"A0",X"42",X"AC",X"C4",X"26",
		X"10",X"10",X"AE",X"D4",X"10",X"AF",X"C4",X"10",X"9E",X"44",X"9F",X"44",X"10",X"AF",X"84",X"35",
		X"F0",X"EE",X"C4",X"26",X"E8",X"CE",X"A0",X"48",X"AC",X"C4",X"27",X"E5",X"EE",X"C4",X"26",X"F8",
		X"BD",X"D0",X"3B",X"34",X"70",X"CE",X"A0",X"4A",X"20",X"EE",X"34",X"76",X"1F",X"01",X"96",X"36",
		X"34",X"02",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"EC",X"A4",X"10",X"AE",X"22",X"34",X"06",
		X"C5",X"01",X"26",X"17",X"C0",X"02",X"EE",X"A5",X"EF",X"85",X"C0",X"02",X"2A",X"F8",X"E6",X"61",
		X"30",X"89",X"01",X"00",X"31",X"A5",X"4A",X"26",X"EB",X"20",X"1D",X"5A",X"A6",X"A5",X"A7",X"85",
		X"C0",X"02",X"2B",X"08",X"EE",X"A5",X"EF",X"85",X"C0",X"02",X"2A",X"F8",X"E6",X"61",X"30",X"89",
		X"01",X"00",X"31",X"A5",X"6A",X"E4",X"26",X"E3",X"32",X"62",X"35",X"02",X"97",X"36",X"B7",X"D0",
		X"00",X"35",X"F6",X"34",X"56",X"1F",X"01",X"96",X"36",X"34",X"02",X"86",X"02",X"97",X"36",X"B7",
		X"D0",X"00",X"EC",X"A4",X"CE",X"00",X"00",X"34",X"04",X"C5",X"01",X"26",X"13",X"C0",X"02",X"EF",
		X"85",X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",X"89",X"01",X"00",X"4A",X"26",X"EF",X"20",X"16",
		X"5A",X"6F",X"85",X"C0",X"02",X"2B",X"06",X"EF",X"85",X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",
		X"89",X"01",X"00",X"4A",X"26",X"EA",X"35",X"06",X"D7",X"36",X"F7",X"D0",X"00",X"35",X"D6",X"34",
		X"56",X"96",X"36",X"34",X"02",X"A6",X"61",X"20",X"BB",X"34",X"18",X"10",X"DF",X"54",X"24",X"02",
		X"31",X"22",X"10",X"EE",X"22",X"CB",X"08",X"1F",X"03",X"20",X"4E",X"34",X"18",X"CB",X"08",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"20",X"6A",X"34",
		X"18",X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",
		X"00",X"36",X"3F",X"33",X"C9",X"01",X"08",X"20",X"44",X"34",X"18",X"10",X"DF",X"54",X"24",X"02",
		X"31",X"22",X"10",X"EE",X"22",X"CB",X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",
		X"08",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",
		X"08",X"35",X"3F",X"36",X"3F",X"10",X"FE",X"A0",X"54",X"35",X"98",X"34",X"18",X"CB",X"08",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"36",X"3F",X"33",
		X"C9",X"01",X"08",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",
		X"3F",X"35",X"98",X"34",X"18",X"7E",X"EE",X"15",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",
		X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"20",X"9C",X"24",X"02",X"31",
		X"22",X"10",X"AE",X"22",X"1F",X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",X"ED",X"42",X"EC",X"24",
		X"ED",X"C9",X"01",X"00",X"EC",X"26",X"ED",X"C9",X"01",X"02",X"EC",X"28",X"ED",X"C9",X"02",X"00",
		X"EC",X"2A",X"ED",X"C9",X"02",X"02",X"39",X"1F",X"03",X"CC",X"00",X"00",X"ED",X"C4",X"ED",X"42",
		X"ED",X"C9",X"01",X"00",X"ED",X"C9",X"01",X"02",X"ED",X"C9",X"02",X"00",X"ED",X"C9",X"02",X"02",
		X"39",X"24",X"02",X"31",X"22",X"10",X"AE",X"22",X"1F",X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",
		X"A7",X"42",X"E7",X"C9",X"01",X"00",X"EC",X"24",X"ED",X"C9",X"01",X"01",X"39",X"1F",X"03",X"CC",
		X"00",X"00",X"ED",X"C4",X"A7",X"42",X"ED",X"C9",X"01",X"00",X"A7",X"C9",X"01",X"02",X"39",X"34",
		X"56",X"10",X"DF",X"54",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"04",X"1F",X"03",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"10",X"DE",X"54",X"35",X"D6",
		X"34",X"56",X"CB",X"04",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"36",X"16",X"33",X"C9",
		X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",
		X"33",X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"35",X"D6",X"34",X"10",
		X"10",X"DF",X"54",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"10",X"DE",X"54",X"35",X"90",X"34",
		X"10",X"CB",X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"36",X"36",X"33",
		X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",
		X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"35",X"90",X"34",X"10",X"10",X"DF",X"54",
		X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"20",X"89",X"34",X"10",X"CB",
		X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"C2",X"34",X"10",X"10",
		X"DF",X"54",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"7E",X"D3",X"5E",
		X"34",X"10",X"CB",X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"99",
		X"34",X"76",X"1A",X"01",X"09",X"67",X"44",X"34",X"02",X"86",X"00",X"24",X"08",X"58",X"49",X"58",
		X"49",X"58",X"49",X"58",X"49",X"BD",X"D7",X"DC",X"DD",X"50",X"C6",X"03",X"E0",X"E0",X"A6",X"85",
		X"9B",X"51",X"19",X"A7",X"85",X"5A",X"2B",X"0E",X"A6",X"85",X"99",X"50",X"19",X"A7",X"85",X"86",
		X"00",X"97",X"50",X"5A",X"2A",X"F2",X"DC",X"86",X"27",X"2B",X"30",X"01",X"31",X"03",X"8D",X"2A",
		X"25",X"23",X"A6",X"21",X"9B",X"87",X"19",X"A7",X"21",X"A6",X"A4",X"99",X"86",X"19",X"A7",X"A4",
		X"6C",X"06",X"6C",X"08",X"BD",X"D6",X"B9",X"BD",X"D7",X"10",X"CC",X"D5",X"52",X"BD",X"D5",X"ED",
		X"C6",X"05",X"BD",X"F5",X"E0",X"8D",X"12",X"35",X"76",X"39",X"34",X"06",X"EC",X"84",X"10",X"A3",
		X"A4",X"26",X"04",X"A6",X"02",X"A1",X"22",X"35",X"86",X"96",X"68",X"34",X"02",X"4A",X"26",X"08",
		X"8E",X"0F",X"1C",X"CE",X"A1",X"9B",X"20",X"06",X"8E",X"71",X"1C",X"CE",X"A1",X"D8",X"0F",X"50",
		X"C6",X"06",X"96",X"36",X"34",X"02",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"A6",X"C0",X"10",
		X"BE",X"C0",X"00",X"C5",X"01",X"26",X"06",X"33",X"5F",X"44",X"44",X"44",X"44",X"84",X"0F",X"26",
		X"0F",X"C1",X"02",X"23",X"0B",X"0D",X"50",X"26",X"07",X"1E",X"10",X"BD",X"D1",X"53",X"20",X"0B",
		X"0C",X"50",X"48",X"48",X"31",X"A6",X"1E",X"10",X"BD",X"D0",X"FA",X"1E",X"10",X"30",X"89",X"04",
		X"00",X"5A",X"26",X"C9",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"82",X"96",X"92",X"2A",
		X"27",X"BD",X"F5",X"CB",X"BD",X"C0",X"1B",X"20",X"1F",X"96",X"92",X"2A",X"1B",X"1A",X"90",X"7F",
		X"D0",X"00",X"86",X"04",X"B7",X"CC",X"03",X"B6",X"CC",X"02",X"BD",X"F5",X"CB",X"96",X"56",X"44",
		X"25",X"03",X"7E",X"C0",X"27",X"7E",X"C0",X"21",X"7E",X"D0",X"0B",X"8E",X"A0",X"5C",X"C6",X"12",
		X"20",X"0C",X"8E",X"A0",X"5D",X"C6",X"15",X"20",X"05",X"8E",X"A0",X"5E",X"C6",X"18",X"96",X"5B",
		X"26",X"E6",X"A6",X"84",X"26",X"E2",X"86",X"1E",X"A7",X"84",X"86",X"C0",X"ED",X"49",X"86",X"0A",
		X"8E",X"D5",X"46",X"7E",X"D0",X"02",X"96",X"5B",X"26",X"CE",X"BD",X"F5",X"CB",X"AD",X"D8",X"09",
		X"20",X"C6",X"FF",X"03",X"20",X"18",X"00",X"F0",X"02",X"08",X"17",X"01",X"20",X"17",X"00",X"F0",
		X"01",X"40",X"08",X"00",X"F0",X"01",X"10",X"08",X"00",X"E8",X"01",X"04",X"14",X"02",X"06",X"11",
		X"02",X"0A",X"17",X"00",X"E8",X"06",X"04",X"11",X"01",X"10",X"17",X"00",X"F0",X"08",X"05",X"02",
		X"00",X"E0",X"01",X"18",X"1A",X"00",X"20",X"01",X"10",X"01",X"00",X"D8",X"01",X"10",X"1A",X"00",
		X"D0",X"01",X"30",X"11",X"00",X"D0",X"01",X"10",X"05",X"00",X"D0",X"01",X"08",X"11",X"00",X"D0",
		X"01",X"08",X"1A",X"00",X"D0",X"01",X"0A",X"08",X"00",X"D0",X"03",X"03",X"17",X"00",X"D0",X"03",
		X"10",X"08",X"00",X"C8",X"0A",X"01",X"0E",X"00",X"C0",X"01",X"08",X"05",X"00",X"C0",X"01",X"30",
		X"07",X"00",X"C0",X"01",X"20",X"1E",X"00",X"C0",X"01",X"08",X"0C",X"00",X"C0",X"01",X"30",X"1B",
		X"00",X"C0",X"01",X"04",X"03",X"00",X"C0",X"01",X"18",X"0D",X"00",X"34",X"07",X"1A",X"FF",X"7F",
		X"D0",X"00",X"86",X"FF",X"B7",X"CC",X"02",X"53",X"F7",X"CC",X"02",X"35",X"87",X"34",X"17",X"0F",
		X"88",X"1F",X"01",X"A6",X"84",X"91",X"8D",X"25",X"0D",X"97",X"8D",X"30",X"1E",X"1A",X"10",X"9F",
		X"8B",X"CC",X"01",X"01",X"DD",X"8E",X"35",X"97",X"96",X"8E",X"27",X"14",X"0A",X"8E",X"26",X"38",
		X"9E",X"8B",X"0A",X"8F",X"26",X"2C",X"30",X"03",X"9F",X"8B",X"A6",X"84",X"26",X"22",X"97",X"8D",
		X"96",X"58",X"85",X"02",X"26",X"0A",X"96",X"88",X"27",X"1E",X"0F",X"88",X"C6",X"0F",X"20",X"16",
		X"96",X"88",X"26",X"14",X"96",X"92",X"85",X"98",X"26",X"0E",X"C6",X"16",X"D7",X"88",X"20",X"06",
		X"97",X"8F",X"EC",X"01",X"97",X"8E",X"8D",X"93",X"B6",X"CC",X"01",X"85",X"40",X"27",X"04",X"86",
		X"3C",X"97",X"5B",X"96",X"5B",X"27",X"02",X"0A",X"5B",X"96",X"5C",X"27",X"02",X"0A",X"5C",X"96",
		X"5E",X"27",X"02",X"0A",X"5E",X"96",X"5D",X"27",X"02",X"0A",X"5D",X"96",X"57",X"43",X"94",X"56",
		X"D6",X"56",X"D7",X"57",X"F6",X"CC",X"00",X"C4",X"3F",X"D7",X"56",X"94",X"56",X"27",X"05",X"CE",
		X"F8",X"95",X"8D",X"1D",X"96",X"58",X"9A",X"59",X"43",X"D6",X"58",X"D7",X"59",X"7F",X"D0",X"00",
		X"F6",X"CC",X"04",X"D7",X"58",X"F6",X"CC",X"06",X"D7",X"5A",X"94",X"58",X"27",X"1A",X"CE",X"F8",
		X"75",X"5F",X"CB",X"04",X"44",X"24",X"FB",X"33",X"C5",X"37",X"16",X"DE",X"5F",X"26",X"05",X"DD",
		X"5F",X"9F",X"61",X"39",X"DD",X"63",X"9F",X"65",X"39",X"34",X"76",X"8E",X"0F",X"14",X"B6",X"A1",
		X"A1",X"8D",X"0F",X"96",X"69",X"4A",X"27",X"08",X"8E",X"71",X"14",X"B6",X"A1",X"DE",X"8D",X"02",
		X"35",X"F6",X"81",X"05",X"23",X"02",X"86",X"05",X"34",X"02",X"CC",X"20",X"06",X"BD",X"D1",X"9F",
		X"A6",X"E4",X"27",X"0F",X"10",X"8E",X"F9",X"C8",X"1F",X"10",X"BD",X"D0",X"FA",X"8B",X"06",X"6A",
		X"E4",X"26",X"F7",X"35",X"82",X"34",X"76",X"CC",X"22",X"20",X"8E",X"3F",X"08",X"BD",X"D1",X"9F",
		X"8D",X"4A",X"8D",X"B5",X"8D",X"0A",X"96",X"69",X"BD",X"D4",X"8B",X"4A",X"26",X"FA",X"35",X"F6",
		X"34",X"76",X"8E",X"29",X"1B",X"B6",X"A1",X"A3",X"8D",X"0F",X"96",X"69",X"4A",X"27",X"08",X"8E",
		X"8B",X"1B",X"B6",X"A1",X"E0",X"8D",X"02",X"35",X"F6",X"81",X"03",X"23",X"02",X"86",X"03",X"34",
		X"02",X"CC",X"03",X"0B",X"BD",X"D1",X"9F",X"A6",X"E4",X"27",X"0F",X"10",X"8E",X"F9",X"CC",X"1F",
		X"10",X"BD",X"D0",X"FA",X"CB",X"04",X"6A",X"E4",X"26",X"F7",X"35",X"82",X"CC",X"55",X"55",X"8E",
		X"3F",X"28",X"ED",X"84",X"30",X"89",X"01",X"00",X"8C",X"61",X"28",X"25",X"F5",X"8E",X"3F",X"07",
		X"A7",X"84",X"30",X"89",X"01",X"00",X"8C",X"61",X"07",X"26",X"F5",X"8E",X"4C",X"07",X"CC",X"99",
		X"99",X"ED",X"84",X"ED",X"88",X"21",X"30",X"89",X"01",X"00",X"8C",X"54",X"07",X"26",X"F2",X"34",
		X"20",X"8E",X"55",X"55",X"10",X"8E",X"FB",X"FE",X"86",X"2E",X"7E",X"FB",X"D0",X"FF",X"34",X"76",
		X"CE",X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"36",X"36",X"36",X"36",X"36",X"36",
		X"36",X"36",X"36",X"36",X"36",X"10",X"11",X"83",X"00",X"00",X"26",X"EE",X"35",X"F6",X"34",X"7E",
		X"CE",X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"1F",X"8B",X"C6",X"08",X"36",X"3A",
		X"36",X"3A",X"36",X"3A",X"36",X"3A",X"5A",X"26",X"F5",X"36",X"3A",X"36",X"3A",X"36",X"3A",X"36",
		X"30",X"33",X"C8",X"D6",X"11",X"83",X"00",X"00",X"26",X"E2",X"35",X"FE",X"34",X"02",X"96",X"68",
		X"8E",X"A1",X"9A",X"4A",X"27",X"03",X"8E",X"A1",X"D7",X"35",X"82",X"34",X"02",X"20",X"F1",X"34",
		X"04",X"D6",X"B7",X"86",X"03",X"3D",X"CB",X"11",X"96",X"B9",X"44",X"44",X"44",X"98",X"B9",X"44",
		X"06",X"B8",X"06",X"B9",X"DB",X"B9",X"D9",X"B8",X"D7",X"B7",X"96",X"B7",X"35",X"84",X"C0",X"FF",
		X"00",X"80",X"14",X"05",X"34",X"34",X"1A",X"FF",X"10",X"CE",X"BF",X"FF",X"86",X"A0",X"1F",X"8B",
		X"7F",X"D0",X"00",X"C6",X"04",X"CE",X"CC",X"00",X"8E",X"D8",X"0E",X"6F",X"41",X"A6",X"80",X"A7",
		X"C1",X"A6",X"03",X"A7",X"5F",X"5A",X"26",X"F3",X"BD",X"D7",X"8E",X"8E",X"9C",X"00",X"6F",X"80",
		X"C6",X"38",X"F7",X"C3",X"FC",X"8C",X"C0",X"00",X"26",X"F4",X"CC",X"A5",X"5A",X"DD",X"B8",X"CC",
		X"FF",X"70",X"DD",X"7C",X"0F",X"7E",X"C6",X"FF",X"DD",X"56",X"BD",X"F5",X"CB",X"BD",X"C0",X"33",
		X"8D",X"24",X"8D",X"12",X"BD",X"F7",X"EF",X"8E",X"D8",X"E5",X"86",X"01",X"BD",X"D0",X"56",X"03",
		X"92",X"1C",X"00",X"7E",X"E7",X"E5",X"8D",X"3D",X"BD",X"E6",X"C6",X"BD",X"E0",X"9D",X"8D",X"45",
		X"12",X"12",X"12",X"7E",X"E1",X"72",X"34",X"16",X"4F",X"5F",X"8E",X"AA",X"9D",X"9F",X"3E",X"30",
		X"0F",X"AF",X"11",X"8C",X"AE",X"F3",X"26",X"F7",X"ED",X"84",X"DD",X"3C",X"8E",X"AF",X"02",X"9F",
		X"46",X"30",X"88",X"17",X"AF",X"88",X"E9",X"8C",X"AF",X"5E",X"26",X"F5",X"ED",X"84",X"8E",X"A0",
		X"3C",X"9F",X"40",X"35",X"96",X"8E",X"F8",X"B1",X"CE",X"A0",X"26",X"C6",X"10",X"A6",X"80",X"A7",
		X"C0",X"5A",X"26",X"F9",X"39",X"34",X"17",X"1A",X"FF",X"8E",X"A2",X"14",X"9F",X"44",X"30",X"88",
		X"17",X"AF",X"88",X"E9",X"8C",X"AA",X"86",X"26",X"F5",X"4F",X"5F",X"ED",X"84",X"DD",X"48",X"DD",
		X"42",X"DD",X"4A",X"35",X"97",X"BD",X"F5",X"CF",X"7E",X"C0",X"00",X"0C",X"26",X"86",X"28",X"8E",
		X"D8",X"E5",X"7E",X"D0",X"02",X"8E",X"C4",X"95",X"BD",X"F8",X"15",X"4A",X"26",X"04",X"86",X"02",
		X"97",X"37",X"39",X"96",X"92",X"2A",X"0E",X"8D",X"EC",X"96",X"37",X"27",X"08",X"CC",X"D5",X"5F",
		X"BD",X"D5",X"ED",X"8D",X"19",X"7E",X"D0",X"0B",X"96",X"92",X"2A",X"F9",X"8D",X"D7",X"96",X"37",
		X"81",X"02",X"25",X"F1",X"CC",X"D5",X"64",X"BD",X"D5",X"ED",X"8D",X"02",X"20",X"E5",X"96",X"92",
		X"2A",X"58",X"BD",X"D0",X"7D",X"BD",X"D7",X"8E",X"86",X"7F",X"97",X"92",X"86",X"01",X"97",X"68",
		X"97",X"25",X"0F",X"69",X"8E",X"A1",X"9A",X"6F",X"80",X"8C",X"A2",X"14",X"26",X"F9",X"86",X"0A",
		X"B7",X"A1",X"A4",X"8E",X"C4",X"85",X"BD",X"F8",X"15",X"84",X"0F",X"B7",X"A1",X"A1",X"B7",X"A1",
		X"A3",X"8E",X"A1",X"9A",X"BD",X"DE",X"A3",X"8E",X"C4",X"81",X"BD",X"F8",X"2B",X"DD",X"86",X"FD",
		X"A1",X"9E",X"7F",X"A1",X"A0",X"8E",X"A1",X"9A",X"A6",X"80",X"A7",X"88",X"3C",X"8C",X"A1",X"D7",
		X"26",X"F6",X"8E",X"D9",X"97",X"86",X"00",X"BD",X"D0",X"56",X"0C",X"69",X"96",X"37",X"8B",X"99",
		X"19",X"97",X"37",X"BD",X"D6",X"F5",X"39",X"C6",X"07",X"BD",X"F5",X"E0",X"BD",X"DE",X"90",X"4F",
		X"5F",X"DD",X"20",X"DD",X"22",X"BD",X"F5",X"C3",X"BD",X"C0",X"06",X"12",X"12",X"12",X"BD",X"D7",
		X"AE",X"CC",X"03",X"00",X"DD",X"95",X"DD",X"93",X"0F",X"88",X"0F",X"90",X"0F",X"67",X"0F",X"8A",
		X"0F",X"75",X"0F",X"74",X"8E",X"A0",X"F2",X"9F",X"76",X"BD",X"D7",X"DC",X"9F",X"6A",X"A6",X"08",
		X"84",X"07",X"CE",X"DB",X"8F",X"A6",X"C6",X"97",X"2B",X"6A",X"07",X"BD",X"DE",X"50",X"CC",X"20",
		X"80",X"DD",X"99",X"DD",X"97",X"CC",X"20",X"00",X"DD",X"9B",X"CC",X"08",X"00",X"D3",X"20",X"DD",
		X"A4",X"CC",X"80",X"00",X"DD",X"9D",X"4F",X"5F",X"DD",X"9F",X"97",X"A1",X"DD",X"A2",X"8E",X"EA",
		X"0A",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"E7",X"A9",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"F5",
		X"57",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"E9",X"E6",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"F5",
		X"28",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"F5",X"01",X"86",X"00",X"BD",X"D0",X"56",X"96",X"25",
		X"27",X"1E",X"D6",X"69",X"5A",X"27",X"19",X"CE",X"C0",X"EF",X"96",X"68",X"4A",X"27",X"03",X"CE",
		X"C0",X"F1",X"8E",X"3C",X"80",X"BD",X"F5",X"D7",X"86",X"80",X"8E",X"DA",X"50",X"7E",X"D0",X"02",
		X"BD",X"D7",X"AE",X"C6",X"05",X"9E",X"6A",X"A6",X"0A",X"8D",X"15",X"86",X"01",X"8E",X"DA",X"63",
		X"7E",X"D0",X"02",X"BD",X"DC",X"5B",X"8D",X"05",X"0F",X"25",X"7E",X"EF",X"21",X"5F",X"96",X"BA",
		X"26",X"02",X"CA",X"02",X"D7",X"92",X"39",X"C6",X"58",X"8D",X"F3",X"DC",X"20",X"DD",X"22",X"9E",
		X"97",X"CC",X"08",X"06",X"BD",X"D1",X"9F",X"BD",X"DB",X"F2",X"CC",X"D5",X"57",X"BD",X"D5",X"ED",
		X"10",X"8E",X"F9",X"B4",X"96",X"93",X"2A",X"04",X"10",X"8E",X"F9",X"BE",X"8E",X"DB",X"87",X"AF",
		X"47",X"CE",X"AF",X"B5",X"BD",X"DB",X"98",X"1F",X"31",X"DE",X"40",X"AF",X"4B",X"DC",X"99",X"10",
		X"AE",X"4B",X"BD",X"D1",X"53",X"86",X"02",X"8E",X"DA",X"BD",X"7E",X"D0",X"02",X"DC",X"99",X"10",
		X"AE",X"4B",X"BD",X"D0",X"FA",X"AE",X"47",X"A6",X"80",X"27",X"0E",X"97",X"31",X"0F",X"26",X"AF",
		X"47",X"86",X"02",X"8E",X"DA",X"AD",X"7E",X"D0",X"02",X"86",X"7F",X"97",X"92",X"BD",X"D8",X"86",
		X"8E",X"DA",X"EB",X"86",X"00",X"BD",X"D0",X"56",X"7E",X"E7",X"E5",X"86",X"FF",X"97",X"26",X"86",
		X"02",X"8E",X"DA",X"F7",X"7E",X"D0",X"02",X"0F",X"26",X"9E",X"99",X"30",X"89",X"04",X"03",X"BD",
		X"F5",X"C3",X"BD",X"C0",X"0E",X"BD",X"D4",X"89",X"0F",X"8E",X"C6",X"13",X"BD",X"D5",X"DB",X"BD",
		X"DD",X"D8",X"26",X"06",X"BD",X"DE",X"11",X"BD",X"D7",X"AE",X"96",X"68",X"9E",X"6A",X"E6",X"07",
		X"26",X"2F",X"D6",X"69",X"5A",X"27",X"41",X"88",X"03",X"BD",X"D7",X"EB",X"E6",X"07",X"27",X"38",
		X"CE",X"C0",X"EF",X"81",X"02",X"27",X"03",X"CE",X"C0",X"F1",X"8E",X"3C",X"78",X"BD",X"F5",X"D7",
		X"CE",X"C0",X"75",X"8E",X"3E",X"88",X"BD",X"F5",X"D7",X"86",X"60",X"8E",X"DB",X"51",X"7E",X"D0",
		X"02",X"96",X"68",X"4C",X"91",X"69",X"23",X"02",X"86",X"01",X"BD",X"D7",X"EB",X"E6",X"07",X"27",
		X"F2",X"97",X"68",X"0C",X"25",X"7E",X"D9",X"97",X"CE",X"C0",X"75",X"8E",X"3E",X"80",X"86",X"FF",
		X"97",X"92",X"BD",X"F5",X"D7",X"0F",X"8E",X"C6",X"13",X"BD",X"D5",X"DB",X"86",X"28",X"8E",X"DB",
		X"84",X"7E",X"D0",X"02",X"7E",X"D8",X"E5",X"07",X"07",X"07",X"0F",X"3F",X"7F",X"FF",X"FF",X"7E",
		X"81",X"28",X"07",X"16",X"2F",X"84",X"15",X"00",X"34",X"56",X"BD",X"F5",X"C7",X"EC",X"A4",X"ED",
		X"C4",X"3D",X"30",X"4A",X"AF",X"42",X"30",X"8B",X"AF",X"44",X"34",X"10",X"30",X"8B",X"34",X"10",
		X"EC",X"26",X"ED",X"46",X"EC",X"28",X"ED",X"48",X"AE",X"22",X"33",X"4A",X"8D",X"0E",X"AE",X"24",
		X"EE",X"62",X"EC",X"E4",X"ED",X"62",X"8D",X"04",X"32",X"64",X"35",X"D6",X"EC",X"81",X"85",X"F0",
		X"27",X"02",X"8A",X"F0",X"85",X"0F",X"27",X"02",X"8A",X"0F",X"C5",X"F0",X"27",X"02",X"CA",X"F0",
		X"C5",X"0F",X"27",X"02",X"CA",X"0F",X"84",X"BB",X"C4",X"BB",X"ED",X"C1",X"11",X"A3",X"64",X"25",
		X"DB",X"39",X"34",X"56",X"DE",X"6A",X"33",X"4A",X"86",X"33",X"6F",X"C0",X"4A",X"26",X"FB",X"DE",
		X"6A",X"96",X"BA",X"A7",X"4A",X"33",X"4B",X"8E",X"A0",X"BB",X"A6",X"80",X"8C",X"A0",X"C0",X"22",
		X"03",X"AB",X"88",X"16",X"A7",X"C0",X"8C",X"A0",X"D2",X"26",X"EF",X"35",X"D6",X"7E",X"ED",X"CE",
		X"12",X"BD",X"D0",X"96",X"F8",X"F4",X"EE",X"4D",X"66",X"66",X"BD",X"D7",X"EF",X"DC",X"B8",X"84",
		X"1F",X"AB",X"61",X"ED",X"0A",X"54",X"24",X"05",X"CC",X"F8",X"F4",X"ED",X"02",X"86",X"F0",X"A7",
		X"0C",X"86",X"10",X"A7",X"88",X"14",X"4F",X"5F",X"ED",X"06",X"EC",X"0A",X"BD",X"EE",X"77",X"9F",
		X"42",X"AF",X"A1",X"0A",X"51",X"26",X"CA",X"35",X"86",X"FF",X"FF",X"8E",X"ED",X"A6",X"86",X"00",
		X"BD",X"D0",X"56",X"CE",X"A0",X"F2",X"31",X"C4",X"EF",X"07",X"6F",X"C0",X"11",X"83",X"A1",X"1A",
		X"26",X"F8",X"DE",X"6A",X"A6",X"4A",X"97",X"BA",X"27",X"20",X"81",X"07",X"23",X"10",X"44",X"44",
		X"5F",X"8D",X"9A",X"CB",X"40",X"26",X"FA",X"48",X"48",X"40",X"AB",X"4A",X"27",X"0C",X"97",X"50",
		X"D6",X"B8",X"86",X"01",X"8D",X"87",X"0A",X"50",X"26",X"F6",X"DE",X"6A",X"33",X"4B",X"8E",X"A0",
		X"BB",X"A6",X"C0",X"A7",X"80",X"8C",X"A0",X"D2",X"26",X"F7",X"8E",X"A0",X"D2",X"6F",X"80",X"8C",
		X"A0",X"DA",X"26",X"F9",X"BD",X"D0",X"AE",X"96",X"B7",X"44",X"8B",X"2A",X"A7",X"0C",X"BD",X"D7",
		X"EF",X"84",X"3F",X"8B",X"80",X"D3",X"20",X"ED",X"0A",X"96",X"BF",X"27",X"19",X"81",X"06",X"23",
		X"02",X"86",X"06",X"31",X"84",X"BD",X"EC",X"82",X"9E",X"44",X"AF",X"A4",X"10",X"9F",X"44",X"40",
		X"9B",X"BF",X"97",X"BF",X"26",X"CE",X"96",X"BE",X"27",X"05",X"BD",X"EF",X"F1",X"0F",X"BE",X"96",
		X"BD",X"97",X"D4",X"27",X"05",X"0F",X"BD",X"BD",X"EC",X"1B",X"96",X"BC",X"97",X"D3",X"27",X"13",
		X"81",X"03",X"23",X"02",X"86",X"03",X"34",X"02",X"BD",X"F3",X"63",X"96",X"BC",X"A0",X"E0",X"97",
		X"BC",X"26",X"ED",X"39",X"DE",X"40",X"86",X"28",X"A7",X"47",X"96",X"CF",X"97",X"D8",X"86",X"01",
		X"97",X"D7",X"96",X"92",X"85",X"08",X"26",X"6E",X"BD",X"E8",X"D0",X"26",X"14",X"86",X"77",X"97",
		X"92",X"BD",X"D0",X"7D",X"BD",X"DB",X"F2",X"BD",X"DE",X"11",X"9E",X"6A",X"6C",X"07",X"7E",X"D9",
		X"9C",X"81",X"08",X"22",X"0F",X"D6",X"CF",X"54",X"81",X"03",X"22",X"01",X"54",X"5C",X"D1",X"D8",
		X"24",X"02",X"D7",X"D8",X"0A",X"D8",X"26",X"18",X"81",X"04",X"96",X"CF",X"24",X"05",X"44",X"44",
		X"BD",X"DD",X"C8",X"97",X"D8",X"96",X"D9",X"81",X"0C",X"24",X"05",X"BD",X"EB",X"68",X"0C",X"D9",
		X"0A",X"D7",X"27",X"04",X"96",X"D2",X"26",X"1E",X"96",X"C0",X"97",X"D7",X"96",X"BB",X"27",X"16",
		X"96",X"D2",X"81",X"08",X"24",X"10",X"96",X"C1",X"91",X"BB",X"23",X"02",X"96",X"BB",X"BD",X"F6",
		X"62",X"40",X"9B",X"BB",X"97",X"BB",X"96",X"89",X"81",X"10",X"24",X"02",X"0C",X"89",X"96",X"24",
		X"4C",X"81",X"F0",X"23",X"06",X"C6",X"06",X"BD",X"F5",X"E0",X"4F",X"97",X"24",X"DE",X"40",X"6A",
		X"47",X"26",X"0D",X"C6",X"02",X"10",X"8E",X"A0",X"BB",X"BD",X"DF",X"0D",X"86",X"28",X"A7",X"47",
		X"86",X"0F",X"8E",X"DD",X"22",X"7E",X"D0",X"02",X"34",X"02",X"BD",X"D7",X"EF",X"A1",X"E4",X"23",
		X"03",X"44",X"20",X"F9",X"4C",X"32",X"61",X"39",X"96",X"D2",X"9B",X"BB",X"9B",X"D3",X"9B",X"D4",
		X"9B",X"D6",X"9B",X"D5",X"9B",X"BE",X"39",X"34",X"04",X"5F",X"81",X"10",X"25",X"06",X"CB",X"0A",
		X"80",X"10",X"20",X"F6",X"34",X"04",X"AB",X"E0",X"35",X"84",X"34",X"04",X"1F",X"89",X"4F",X"C1",
		X"0A",X"25",X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",
		X"84",X"0F",X"26",X"DE",X"40",X"35",X"10",X"AF",X"4D",X"12",X"12",X"12",X"CE",X"C0",X"F9",X"8E",
		X"38",X"50",X"BD",X"F5",X"D7",X"9E",X"6A",X"A6",X"08",X"8D",X"CF",X"1F",X"89",X"4F",X"BE",X"B2",
		X"16",X"BD",X"C0",X"0E",X"8E",X"3D",X"60",X"CE",X"C0",X"FB",X"BD",X"F5",X"D7",X"9E",X"6A",X"BD",
		X"DE",X"A3",X"CC",X"D5",X"C2",X"BD",X"D5",X"ED",X"86",X"80",X"8E",X"DE",X"A0",X"7E",X"D0",X"02",
		X"BD",X"D6",X"F5",X"BD",X"F6",X"F5",X"34",X"20",X"10",X"8E",X"FB",X"3E",X"12",X"12",X"12",X"48",
		X"48",X"E6",X"A6",X"D7",X"1A",X"4C",X"E6",X"A6",X"E7",X"0A",X"4C",X"E6",X"A6",X"D7",X"1E",X"4C",
		X"E6",X"A6",X"D7",X"1F",X"C6",X"02",X"DA",X"92",X"D7",X"92",X"96",X"36",X"34",X"02",X"86",X"07",
		X"97",X"36",X"B7",X"D0",X"00",X"BD",X"C0",X"00",X"35",X"22",X"97",X"36",X"B7",X"D0",X"00",X"39",
		X"BD",X"F5",X"C3",X"BD",X"CB",X"A0",X"BD",X"D8",X"76",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6E",X"D8",X"0D",X"34",X"56",X"6C",X"08",X"8E",X"C4",X"9D",X"BD",X"F8",X"15",X"97",X"50",X"AE",
		X"62",X"A6",X"08",X"90",X"50",X"25",X"06",X"26",X"FA",X"86",X"0A",X"A7",X"0A",X"A6",X"08",X"34",
		X"02",X"84",X"03",X"BD",X"F7",X"99",X"12",X"CE",X"DF",X"35",X"8B",X"04",X"30",X"0B",X"E6",X"C6",
		X"E7",X"80",X"33",X"48",X"11",X"83",X"DF",X"ED",X"26",X"F4",X"35",X"02",X"80",X"04",X"24",X"01",
		X"4F",X"97",X"50",X"8E",X"C4",X"97",X"BD",X"F8",X"2B",X"BD",X"DD",X"E7",X"9B",X"50",X"97",X"50",
		X"27",X"19",X"1F",X"98",X"BD",X"DD",X"E7",X"91",X"50",X"24",X"02",X"97",X"50",X"96",X"50",X"C6",
		X"03",X"BD",X"D7",X"DC",X"31",X"0B",X"8D",X"05",X"4A",X"26",X"F4",X"35",X"D6",X"34",X"32",X"8E",
		X"DF",X"35",X"A6",X"85",X"2B",X"0A",X"AB",X"A4",X"25",X"10",X"A1",X"84",X"22",X"0C",X"20",X"08",
		X"AB",X"A4",X"24",X"06",X"A1",X"01",X"25",X"02",X"A7",X"A4",X"31",X"21",X"30",X"08",X"8C",X"DF",
		X"ED",X"26",X"DF",X"35",X"B2",X"14",X"00",X"00",X"00",X"0A",X"02",X"00",X"00",X"03",X"00",X"00",
		X"00",X"06",X"06",X"00",X"06",X"06",X"00",X"00",X"00",X"04",X"00",X"00",X"02",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"02",X"0A",X"00",X"1E",X"00",X"00",
		X"00",X"1E",X"19",X"14",X"10",X"05",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"60",X"00",X"03",
		X"02",X"20",X"28",X"30",X"38",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"FF",X"00",X"10",
		X"04",X"70",X"B0",X"00",X"00",X"80",X"10",X"FC",X"FE",X"40",X"30",X"20",X"20",X"30",X"00",X"00",
		X"00",X"20",X"28",X"2C",X"30",X"02",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"01",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"FF",X"00",X"08",X"06",X"80",X"00",X"20",X"30",X"60",X"00",X"08",
		X"04",X"20",X"30",X"38",X"3C",X"FF",X"08",X"FE",X"FE",X"20",X"18",X"14",X"12",X"60",X"00",X"08",
		X"02",X"20",X"28",X"2A",X"2C",X"28",X"0A",X"FE",X"FF",X"14",X"14",X"14",X"14",X"3F",X"00",X"00",
		X"00",X"1F",X"1F",X"1F",X"3F",X"C0",X"18",X"F4",X"FC",X"C0",X"B0",X"90",X"80",X"0A",X"03",X"FF",
		X"FF",X"0A",X"08",X"07",X"05",X"C8",X"28",X"F4",X"F8",X"C8",X"B4",X"A0",X"A0",X"7F",X"D0",X"00",
		X"86",X"A0",X"1F",X"8B",X"86",X"04",X"B7",X"CC",X"03",X"B6",X"CC",X"02",X"B6",X"C8",X"00",X"81",
		X"80",X"25",X"32",X"96",X"6C",X"26",X"7F",X"0C",X"6C",X"0F",X"6D",X"BD",X"D6",X"08",X"BD",X"E2",
		X"8C",X"BD",X"E0",X"C9",X"B6",X"C8",X"00",X"80",X"08",X"81",X"A8",X"23",X"02",X"86",X"A8",X"97",
		X"7D",X"86",X"02",X"B7",X"D0",X"00",X"DC",X"7D",X"BD",X"E3",X"C8",X"DC",X"7D",X"BD",X"E2",X"3C",
		X"BD",X"E4",X"7C",X"20",X"51",X"D6",X"6D",X"26",X"4D",X"0C",X"6D",X"0F",X"6C",X"F6",X"CC",X"00",
		X"0C",X"3A",X"C6",X"38",X"F7",X"C3",X"FC",X"81",X"08",X"22",X"1B",X"CE",X"C0",X"10",X"DC",X"30",
		X"9E",X"32",X"10",X"9E",X"34",X"36",X"36",X"DC",X"2A",X"9E",X"2C",X"10",X"9E",X"2E",X"36",X"36",
		X"DC",X"26",X"9E",X"28",X"36",X"16",X"86",X"07",X"B7",X"D0",X"00",X"96",X"92",X"85",X"02",X"26",
		X"03",X"BD",X"C0",X"03",X"86",X"02",X"B7",X"D0",X"00",X"DC",X"7C",X"BD",X"E2",X"3C",X"DC",X"7C",
		X"BD",X"E3",X"C8",X"BD",X"E3",X"9F",X"1A",X"FF",X"7F",X"D0",X"00",X"86",X"05",X"B7",X"CC",X"03",
		X"96",X"36",X"B7",X"D0",X"00",X"A6",X"E4",X"84",X"6F",X"A7",X"E4",X"35",X"FF",X"8E",X"AF",X"75",
		X"C6",X"10",X"D7",X"89",X"5F",X"BD",X"D7",X"EF",X"81",X"9C",X"24",X"F9",X"A7",X"84",X"BD",X"D7",
		X"EF",X"81",X"A8",X"22",X"F9",X"81",X"2A",X"23",X"F5",X"A7",X"01",X"E7",X"02",X"CB",X"11",X"C4",
		X"77",X"30",X"04",X"8C",X"AF",X"B5",X"26",X"DD",X"39",X"96",X"92",X"85",X"20",X"26",X"F9",X"7E",
		X"E8",X"C3",X"DC",X"20",X"C4",X"80",X"DD",X"4C",X"DC",X"22",X"C4",X"80",X"93",X"4C",X"58",X"49",
		X"97",X"4C",X"C6",X"F0",X"96",X"21",X"85",X"40",X"26",X"01",X"53",X"D7",X"4E",X"4F",X"A7",X"94",
		X"A7",X"98",X"04",X"A7",X"98",X"08",X"A7",X"98",X"0C",X"A7",X"98",X"10",X"A7",X"98",X"14",X"A7",
		X"98",X"18",X"A7",X"98",X"1C",X"A7",X"98",X"20",X"A7",X"98",X"24",X"A7",X"98",X"28",X"A7",X"98",
		X"2C",X"A7",X"98",X"30",X"A7",X"98",X"34",X"A7",X"98",X"38",X"A7",X"98",X"3C",X"D6",X"89",X"A6",
		X"84",X"9B",X"4C",X"81",X"9C",X"25",X"0A",X"81",X"C0",X"23",X"04",X"86",X"9B",X"20",X"02",X"86",
		X"00",X"A7",X"84",X"A6",X"02",X"94",X"4E",X"A7",X"98",X"00",X"30",X"04",X"5A",X"26",X"E0",X"D6",
		X"B7",X"C4",X"3C",X"8E",X"AF",X"75",X"3A",X"A6",X"02",X"8B",X"11",X"84",X"77",X"A7",X"02",X"96",
		X"B7",X"85",X"01",X"27",X"1C",X"81",X"98",X"25",X"02",X"80",X"84",X"6F",X"98",X"00",X"A7",X"84",
		X"96",X"92",X"85",X"02",X"27",X"0B",X"96",X"B9",X"84",X"3F",X"C6",X"03",X"3D",X"CB",X"2A",X"E7",
		X"01",X"39",X"8E",X"A1",X"3A",X"9F",X"7A",X"BD",X"D7",X"EF",X"A7",X"88",X"20",X"A7",X"80",X"8C",
		X"A1",X"5B",X"26",X"F3",X"39",X"9E",X"7A",X"DE",X"97",X"33",X"C9",X"FF",X"01",X"EC",X"84",X"ED",
		X"C4",X"A6",X"05",X"E6",X"09",X"ED",X"42",X"A6",X"0C",X"A7",X"44",X"96",X"58",X"85",X"02",X"27",
		X"36",X"A6",X"03",X"E6",X"06",X"ED",X"C9",X"FF",X"01",X"ED",X"C9",X"FE",X"01",X"A6",X"0A",X"A7",
		X"C9",X"FE",X"03",X"A7",X"C9",X"FF",X"03",X"A6",X"04",X"E6",X"07",X"ED",X"C9",X"FD",X"01",X"ED",
		X"C9",X"FC",X"01",X"A6",X"0B",X"A7",X"C9",X"FD",X"03",X"A7",X"C9",X"FC",X"03",X"A6",X"08",X"A7",
		X"C9",X"FA",X"02",X"A7",X"C9",X"FB",X"02",X"39",X"41",X"08",X"02",X"4B",X"08",X"41",X"02",X"08",
		X"01",X"10",X"AF",X"89",X"01",X"02",X"37",X"26",X"10",X"AF",X"89",X"02",X"01",X"A7",X"89",X"02",
		X"03",X"E7",X"89",X"03",X"02",X"39",X"DE",X"97",X"5F",X"8E",X"00",X"00",X"31",X"84",X"33",X"C9",
		X"FF",X"06",X"36",X"34",X"AF",X"C9",X"FF",X"01",X"E7",X"C9",X"FF",X"03",X"AF",X"C9",X"FE",X"01",
		X"E7",X"C9",X"FE",X"03",X"AF",X"C9",X"FD",X"01",X"E7",X"C9",X"FD",X"03",X"AF",X"C9",X"FC",X"01",
		X"E7",X"C9",X"FC",X"03",X"AF",X"C9",X"FB",X"02",X"E7",X"C9",X"FA",X"02",X"39",X"FF",X"03",X"AF",
		X"C9",X"FE",X"01",X"E7",X"C9",X"FE",X"03",X"E7",X"C9",X"FD",X"02",X"39",X"97",X"54",X"96",X"92",
		X"85",X"10",X"26",X"28",X"96",X"54",X"91",X"98",X"23",X"22",X"D1",X"98",X"22",X"1E",X"BD",X"E2",
		X"87",X"BD",X"E1",X"F6",X"20",X"0A",X"E2",X"19",X"20",X"06",X"BD",X"E2",X"87",X"BD",X"E1",X"F6",
		X"DC",X"93",X"BD",X"E2",X"73",X"BD",X"E1",X"85",X"39",X"BD",X"E1",X"85",X"39",X"BD",X"E2",X"81",
		X"7E",X"E1",X"C4",X"10",X"8E",X"F9",X"B4",X"96",X"9C",X"48",X"DC",X"99",X"DD",X"97",X"7E",X"D3",
		X"3E",X"10",X"8E",X"F9",X"BE",X"20",X"F0",X"DC",X"97",X"7E",X"D3",X"8F",X"96",X"92",X"85",X"40",
		X"10",X"26",X"01",X"0A",X"0F",X"4C",X"DC",X"9F",X"43",X"53",X"C3",X"00",X"01",X"2A",X"02",X"03",
		X"4C",X"58",X"49",X"58",X"49",X"D3",X"A0",X"DD",X"A0",X"96",X"4C",X"99",X"9F",X"97",X"9F",X"DC",
		X"9F",X"96",X"58",X"85",X"02",X"27",X"12",X"0F",X"4C",X"DC",X"95",X"2A",X"02",X"03",X"4C",X"D3",
		X"A0",X"DD",X"A0",X"96",X"4C",X"99",X"9F",X"97",X"9F",X"DC",X"9F",X"47",X"56",X"47",X"56",X"4F",
		X"57",X"46",X"97",X"6F",X"D7",X"6E",X"96",X"95",X"2B",X"07",X"86",X"20",X"5D",X"2B",X"07",X"20",
		X"09",X"86",X"70",X"5D",X"2B",X"04",X"0F",X"6F",X"0F",X"6E",X"D6",X"6F",X"9B",X"6E",X"97",X"6E",
		X"93",X"9B",X"27",X"26",X"25",X"12",X"10",X"83",X"01",X"00",X"23",X"1E",X"CC",X"00",X"40",X"DD",
		X"70",X"CC",X"01",X"00",X"D3",X"9B",X"20",X"18",X"10",X"83",X"FF",X"00",X"2E",X"0C",X"CC",X"FF",
		X"C0",X"DD",X"70",X"CC",X"FF",X"00",X"D3",X"9B",X"20",X"06",X"4F",X"5F",X"DD",X"70",X"DC",X"6E",
		X"DD",X"9B",X"97",X"99",X"DC",X"20",X"DD",X"22",X"DC",X"9F",X"10",X"83",X"01",X"00",X"2D",X"03",
		X"CC",X"01",X"00",X"10",X"83",X"FF",X"00",X"2E",X"03",X"CC",X"00",X"04",X"DD",X"9F",X"D3",X"20",
		X"93",X"70",X"DD",X"20",X"DC",X"9B",X"44",X"56",X"44",X"56",X"C4",X"E0",X"D3",X"20",X"DD",X"A4",
		X"D6",X"9D",X"96",X"5A",X"44",X"25",X"09",X"96",X"58",X"2B",X"20",X"CC",X"00",X"00",X"20",X"36",
		X"C1",X"2B",X"23",X"3A",X"DC",X"A2",X"2A",X"0E",X"C3",X"FF",X"F8",X"10",X"83",X"FE",X"00",X"2C",
		X"25",X"CC",X"FE",X"00",X"20",X"20",X"CC",X"FF",X"00",X"20",X"1B",X"C1",X"EE",X"24",X"1F",X"DC",
		X"A2",X"2F",X"0E",X"C3",X"00",X"08",X"10",X"83",X"02",X"00",X"23",X"0A",X"CC",X"02",X"00",X"20",
		X"05",X"CC",X"01",X"00",X"20",X"00",X"DD",X"A2",X"D3",X"9D",X"DD",X"9D",X"97",X"9A",X"39",X"BD",
		X"E9",X"D9",X"12",X"26",X"22",X"8E",X"A0",X"42",X"20",X"19",X"EC",X"0A",X"E3",X"0E",X"ED",X"0A",
		X"EC",X"88",X"10",X"BD",X"E9",X"53",X"EC",X"0C",X"E3",X"88",X"10",X"12",X"12",X"12",X"12",X"12",
		X"12",X"ED",X"0C",X"AE",X"84",X"26",X"E3",X"39",X"34",X"06",X"96",X"92",X"85",X"20",X"26",X"4A",
		X"8E",X"A0",X"42",X"20",X"41",X"EC",X"04",X"27",X"12",X"E1",X"E4",X"22",X"39",X"E1",X"61",X"23",
		X"35",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"4F",X"5F",X"ED",X"04",X"E6",X"0C",X"E1",X"E4",X"22",
		X"25",X"E1",X"61",X"23",X"21",X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",X"80",X"24",X"17",X"10",
		X"AE",X"02",X"58",X"49",X"58",X"49",X"AB",X"A4",X"81",X"9C",X"22",X"0A",X"A0",X"A4",X"58",X"E6",
		X"0C",X"ED",X"04",X"AD",X"B8",X"06",X"AE",X"84",X"26",X"BB",X"35",X"86",X"34",X"66",X"96",X"74",
		X"81",X"14",X"24",X"4F",X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",X"80",X"24",X"45",X"58",X"49",
		X"58",X"49",X"E6",X"0C",X"C1",X"2A",X"23",X"3B",X"9E",X"44",X"27",X"37",X"ED",X"04",X"ED",X"0A",
		X"1E",X"89",X"ED",X"0C",X"EF",X"06",X"4F",X"5F",X"ED",X"0E",X"ED",X"88",X"10",X"EE",X"66",X"37",
		X"26",X"ED",X"88",X"12",X"10",X"AF",X"02",X"37",X"06",X"EF",X"66",X"ED",X"08",X"86",X"14",X"A7",
		X"88",X"15",X"A7",X"88",X"16",X"EC",X"84",X"DD",X"44",X"DC",X"4A",X"ED",X"84",X"0C",X"74",X"9F",
		X"4A",X"35",X"E6",X"EE",X"66",X"33",X"46",X"EF",X"66",X"4F",X"35",X"E6",X"96",X"92",X"85",X"20",
		X"26",X"3E",X"DC",X"20",X"C4",X"E0",X"DD",X"78",X"DC",X"22",X"C4",X"E0",X"93",X"78",X"58",X"49",
		X"58",X"49",X"DD",X"78",X"8E",X"A0",X"4A",X"20",X"23",X"10",X"AE",X"04",X"EC",X"88",X"10",X"E3",
		X"0C",X"81",X"2A",X"23",X"4A",X"ED",X"0C",X"EC",X"0E",X"D3",X"78",X"E3",X"0A",X"81",X"98",X"24",
		X"3E",X"ED",X"0A",X"E6",X"0C",X"ED",X"04",X"EE",X"04",X"6E",X"98",X"12",X"AE",X"84",X"26",X"D9",
		X"39",X"DE",X"81",X"E6",X"0B",X"2A",X"02",X"33",X"46",X"CC",X"00",X"00",X"ED",X"A4",X"A7",X"22",
		X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"10",X"AE",X"04",X"EC",X"C4",X"ED",X"A4",X"EC",
		X"42",X"A7",X"22",X"E7",X"A9",X"01",X"00",X"EC",X"44",X"ED",X"A9",X"01",X"01",X"20",X"CD",X"4F",
		X"5F",X"A7",X"88",X"16",X"BD",X"E5",X"17",X"20",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"BA",X"8D",X"13",X"EC",X"04",X"10",X"AE",X"02",X"8D",X"1F",X"27",X"04",X"10",X"8E",X"F9",
		X"DA",X"BD",X"D0",X"FA",X"7E",X"E4",X"BC",X"34",X"10",X"EC",X"98",X"02",X"8D",X"0C",X"27",X"03",
		X"FC",X"F9",X"DA",X"1F",X"21",X"BD",X"D1",X"9F",X"35",X"90",X"34",X"02",X"B6",X"A1",X"8A",X"84",
		X"01",X"35",X"82",X"FF",X"BD",X"D4",X"10",X"CC",X"D5",X"74",X"BD",X"D5",X"ED",X"39",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",X"25",X"BD",X"D4",X"10",X"0A",X"74",X"BD",
		X"D0",X"F3",X"BD",X"F4",X"C2",X"EC",X"0A",X"44",X"56",X"44",X"56",X"D3",X"20",X"ED",X"0A",X"A6",
		X"0C",X"80",X"02",X"A7",X"0C",X"CC",X"F9",X"44",X"ED",X"02",X"BD",X"FC",X"83",X"CC",X"D5",X"86",
		X"7E",X"D5",X"ED",X"FF",X"FF",X"34",X"02",X"A6",X"0C",X"91",X"1B",X"24",X"06",X"96",X"1B",X"A7",
		X"0C",X"20",X"08",X"91",X"1C",X"23",X"04",X"96",X"1C",X"A7",X"0C",X"35",X"02",X"E3",X"0C",X"39",
		X"FF",X"FF",X"FF",X"FF",X"8E",X"A0",X"4A",X"20",X"1B",X"A6",X"88",X"16",X"27",X"05",X"6A",X"88",
		X"15",X"26",X"11",X"EE",X"84",X"EF",X"A4",X"DE",X"44",X"EF",X"84",X"9F",X"44",X"BD",X"F4",X"C2",
		X"0A",X"74",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"DF",X"39",X"4F",X"20",X"02",X"86",X"01",
		X"7E",X"F2",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"34",X"46",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"06",
		X"CE",X"F9",X"62",X"BD",X"E6",X"E1",X"35",X"C0",X"BD",X"EF",X"52",X"12",X"AF",X"47",X"AF",X"49",
		X"AF",X"4B",X"96",X"92",X"85",X"40",X"26",X"50",X"86",X"04",X"AE",X"47",X"C6",X"11",X"8C",X"98",
		X"00",X"24",X"45",X"E7",X"84",X"BD",X"ED",X"BC",X"12",X"4A",X"26",X"F7",X"C6",X"99",X"E7",X"84",
		X"AF",X"47",X"10",X"9E",X"7F",X"10",X"8C",X"A1",X"37",X"25",X"04",X"10",X"8E",X"A1",X"1A",X"AE",
		X"49",X"86",X"03",X"E6",X"A0",X"E7",X"84",X"BD",X"ED",X"BC",X"12",X"4A",X"26",X"F5",X"10",X"9F",
		X"7F",X"AF",X"49",X"BD",X"FA",X"7E",X"12",X"12",X"EC",X"47",X"80",X"06",X"8D",X"97",X"26",X"08",
		X"7E",X"EF",X"5A",X"12",X"12",X"12",X"12",X"12",X"AE",X"4B",X"4F",X"A7",X"84",X"BD",X"ED",X"BC",
		X"12",X"AC",X"47",X"23",X"F6",X"20",X"6A",X"30",X"04",X"AF",X"47",X"AF",X"49",X"AF",X"4B",X"96",
		X"92",X"85",X"40",X"26",X"4F",X"86",X"04",X"AE",X"47",X"C6",X"11",X"8C",X"05",X"00",X"23",X"44",
		X"E7",X"84",X"30",X"89",X"FF",X"00",X"4A",X"26",X"F7",X"C6",X"99",X"E7",X"84",X"AF",X"47",X"10",
		X"9E",X"7F",X"10",X"8C",X"A1",X"37",X"25",X"04",X"10",X"8E",X"A1",X"1A",X"AE",X"49",X"86",X"03",
		X"E6",X"A0",X"E7",X"84",X"30",X"89",X"FF",X"00",X"4A",X"26",X"F5",X"10",X"9F",X"7F",X"AF",X"49",
		X"6F",X"D8",X"0B",X"6A",X"4B",X"EC",X"47",X"BD",X"E5",X"D5",X"26",X"08",X"86",X"01",X"8E",X"E6",
		X"5F",X"7E",X"D0",X"02",X"AE",X"4B",X"4F",X"A7",X"84",X"30",X"89",X"FF",X"00",X"AC",X"47",X"24",
		X"F6",X"0A",X"90",X"7E",X"D0",X"0B",X"8E",X"A1",X"1A",X"9F",X"7F",X"BD",X"D7",X"EF",X"5F",X"44",
		X"24",X"02",X"CB",X"01",X"44",X"24",X"02",X"CB",X"10",X"E7",X"80",X"8C",X"A1",X"3A",X"26",X"EB",
		X"39",X"8E",X"A0",X"42",X"DD",X"AE",X"E3",X"C4",X"DD",X"B0",X"20",X"17",X"EC",X"04",X"27",X"13",
		X"91",X"B0",X"24",X"0F",X"D1",X"B1",X"24",X"0B",X"E3",X"98",X"02",X"91",X"AE",X"23",X"04",X"D1",
		X"AF",X"22",X"05",X"AE",X"84",X"26",X"E5",X"39",X"DF",X"B4",X"10",X"AE",X"02",X"A3",X"A4",X"DD",
		X"50",X"4F",X"5F",X"DD",X"A8",X"DD",X"AA",X"DC",X"50",X"D0",X"AF",X"22",X"05",X"50",X"D7",X"A9",
		X"20",X"02",X"D7",X"AB",X"90",X"AE",X"22",X"05",X"40",X"97",X"A8",X"20",X"02",X"97",X"AA",X"DC",
		X"50",X"E3",X"A4",X"D0",X"B1",X"22",X"01",X"5F",X"90",X"B0",X"22",X"01",X"4F",X"DD",X"B2",X"EC",
		X"A4",X"93",X"A8",X"93",X"B2",X"DD",X"A6",X"A6",X"41",X"97",X"AD",X"D6",X"AA",X"3D",X"EE",X"42",
		X"33",X"CB",X"A6",X"21",X"97",X"AC",X"10",X"AE",X"22",X"D6",X"A8",X"3D",X"31",X"AB",X"96",X"A9",
		X"31",X"A6",X"96",X"AB",X"33",X"C6",X"D6",X"A7",X"5A",X"A6",X"C5",X"27",X"2A",X"A6",X"A5",X"27",
		X"26",X"31",X"A5",X"1F",X"20",X"EE",X"02",X"A3",X"42",X"10",X"AE",X"04",X"E0",X"41",X"82",X"00",
		X"25",X"06",X"31",X"A9",X"01",X"00",X"20",X"F4",X"EB",X"41",X"89",X"00",X"31",X"A5",X"10",X"9F",
		X"F0",X"AD",X"98",X"08",X"86",X"01",X"39",X"5A",X"2A",X"CF",X"DC",X"AC",X"31",X"A6",X"33",X"C5",
		X"0A",X"A6",X"26",X"C2",X"DE",X"B4",X"7E",X"E7",X"03",X"0F",X"91",X"8E",X"E7",X"C0",X"96",X"91",
		X"E6",X"86",X"27",X"F5",X"0C",X"91",X"D7",X"27",X"86",X"02",X"8E",X"E7",X"AB",X"7E",X"D0",X"02",
		X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",
		X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",X"CA",X"DA",X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",
		X"BF",X"3F",X"3E",X"3C",X"00",X"8E",X"A0",X"3C",X"9F",X"40",X"96",X"3A",X"27",X"FC",X"0F",X"3A",
		X"D6",X"92",X"C5",X"7D",X"27",X"04",X"0F",X"3B",X"20",X"47",X"48",X"9B",X"3B",X"80",X"04",X"2A",
		X"01",X"4F",X"97",X"3B",X"81",X"02",X"25",X"39",X"C6",X"03",X"D7",X"89",X"81",X"02",X"23",X"31",
		X"86",X"02",X"97",X"3B",X"10",X"8E",X"A0",X"42",X"AE",X"A4",X"27",X"25",X"A6",X"88",X"14",X"12",
		X"12",X"31",X"84",X"20",X"F3",X"EE",X"84",X"EF",X"A4",X"DC",X"B7",X"84",X"3F",X"8B",X"60",X"E3",
		X"0A",X"ED",X"0A",X"BD",X"F4",X"C2",X"CC",X"00",X"00",X"ED",X"04",X"DE",X"48",X"9F",X"48",X"EF",
		X"84",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"8D",X"3E",X"BD",X"FC",X"86",X"BD",X"D7",X"EF",
		X"9E",X"5F",X"26",X"0C",X"9E",X"63",X"27",X"17",X"DC",X"65",X"0F",X"63",X"0F",X"64",X"20",X"06",
		X"DC",X"61",X"0F",X"5F",X"0F",X"60",X"D4",X"92",X"26",X"E6",X"BD",X"D0",X"56",X"20",X"E1",X"CE",
		X"A0",X"3C",X"20",X"09",X"6A",X"44",X"26",X"05",X"DF",X"40",X"6E",X"D8",X"02",X"EE",X"C4",X"26",
		X"F3",X"10",X"CE",X"BF",X"FF",X"7E",X"E7",X"E5",X"96",X"92",X"85",X"10",X"26",X"2D",X"DC",X"97",
		X"CE",X"F9",X"B4",X"0D",X"95",X"2A",X"03",X"CE",X"F9",X"BE",X"34",X"46",X"0C",X"B6",X"BD",X"E6",
		X"E1",X"35",X"46",X"26",X"08",X"8E",X"A0",X"4A",X"BD",X"F6",X"B5",X"27",X"0E",X"8E",X"DA",X"77",
		X"86",X"00",X"BD",X"D0",X"56",X"96",X"92",X"8A",X"08",X"97",X"92",X"0F",X"B6",X"39",X"0F",X"8A",
		X"7E",X"D0",X"0B",X"96",X"1A",X"81",X"7F",X"26",X"01",X"39",X"8E",X"AF",X"75",X"7E",X"E0",X"D2",
		X"BD",X"DD",X"D8",X"9B",X"BA",X"39",X"C3",X"30",X"07",X"81",X"40",X"25",X"05",X"81",X"60",X"24",
		X"01",X"39",X"32",X"62",X"7E",X"EB",X"61",X"FF",X"96",X"75",X"26",X"1C",X"9E",X"6A",X"A6",X"09",
		X"27",X"16",X"0C",X"75",X"6A",X"09",X"BD",X"D7",X"10",X"8E",X"48",X"18",X"CE",X"C0",X"AD",X"BD",
		X"F6",X"A7",X"86",X"01",X"97",X"19",X"12",X"12",X"7E",X"D0",X"0B",X"0D",X"19",X"27",X"0B",X"CC",
		X"04",X"7F",X"FD",X"BC",X"10",X"F7",X"BC",X"12",X"0F",X"19",X"7D",X"BC",X"12",X"27",X"06",X"7A",
		X"BC",X"12",X"7E",X"E0",X"95",X"FC",X"BC",X"10",X"27",X"16",X"7F",X"D0",X"00",X"BD",X"EF",X"42",
		X"BD",X"FC",X"20",X"26",X"0B",X"8E",X"48",X"18",X"CE",X"C0",X"AD",X"BD",X"F6",X"AE",X"0F",X"75",
		X"7E",X"DF",X"ED",X"FF",X"FF",X"FF",X"7E",X"E5",X"BE",X"EC",X"88",X"10",X"58",X"49",X"58",X"49",
		X"58",X"49",X"39",X"8D",X"1F",X"BD",X"E5",X"75",X"91",X"1B",X"24",X"09",X"63",X"88",X"10",X"63",
		X"88",X"11",X"12",X"20",X"0E",X"91",X"1C",X"23",X"0A",X"63",X"88",X"10",X"63",X"88",X"11",X"12",
		X"12",X"12",X"12",X"39",X"34",X"06",X"96",X"1A",X"27",X"0B",X"81",X"FF",X"26",X"14",X"CC",X"2A",
		X"F0",X"DD",X"1B",X"20",X"1C",X"7E",X"F3",X"31",X"12",X"BD",X"EE",X"36",X"80",X"08",X"97",X"1C",
		X"20",X"0F",X"BD",X"EE",X"36",X"34",X"02",X"80",X"08",X"97",X"1C",X"35",X"02",X"90",X"1A",X"97",
		X"1B",X"35",X"86",X"34",X"18",X"10",X"DF",X"54",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",
		X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"7E",X"D1",X"F9",X"34",X"18",
		X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",
		X"36",X"3F",X"33",X"C9",X"01",X"08",X"7E",X"D2",X"2D",X"0D",X"1D",X"27",X"01",X"39",X"96",X"92",
		X"85",X"20",X"39",X"FF",X"FF",X"FF",X"9E",X"7A",X"30",X"01",X"8C",X"A1",X"5A",X"23",X"03",X"8E",
		X"A1",X"3A",X"9F",X"7A",X"9E",X"83",X"30",X"01",X"8C",X"A1",X"92",X"23",X"03",X"8E",X"A1",X"7A",
		X"9F",X"83",X"86",X"04",X"8E",X"E9",X"E6",X"7E",X"D0",X"02",X"BD",X"EA",X"57",X"86",X"02",X"8E",
		X"EA",X"15",X"7E",X"D0",X"02",X"BD",X"EA",X"2E",X"BD",X"E5",X"94",X"86",X"02",X"8E",X"EA",X"23",
		X"7E",X"D0",X"02",X"BD",X"EA",X"A3",X"86",X"04",X"8E",X"EA",X"0A",X"7E",X"D0",X"02",X"DC",X"20",
		X"83",X"0C",X"80",X"DD",X"50",X"8E",X"A0",X"42",X"20",X"16",X"EC",X"0A",X"93",X"50",X"10",X"83",
		X"3E",X"80",X"25",X"0C",X"EE",X"84",X"EF",X"A4",X"DE",X"48",X"EF",X"84",X"9F",X"48",X"30",X"A4",
		X"31",X"84",X"AE",X"84",X"26",X"E4",X"39",X"DC",X"20",X"83",X"0C",X"80",X"DD",X"50",X"8E",X"A0",
		X"48",X"20",X"39",X"EC",X"88",X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"EC",X"88",X"10",X"BD",
		X"E9",X"53",X"BD",X"E9",X"49",X"E3",X"0C",X"12",X"12",X"12",X"ED",X"0C",X"EC",X"0E",X"58",X"49",
		X"58",X"49",X"58",X"49",X"E3",X"0A",X"ED",X"0A",X"93",X"50",X"10",X"83",X"3E",X"80",X"24",X"0C",
		X"EE",X"84",X"EF",X"A4",X"DE",X"42",X"EF",X"84",X"9F",X"42",X"30",X"A4",X"31",X"84",X"AE",X"84",
		X"26",X"C1",X"39",X"CE",X"00",X"00",X"C6",X"08",X"8E",X"B0",X"35",X"EF",X"94",X"EF",X"98",X"02",
		X"EF",X"98",X"04",X"EF",X"98",X"06",X"3A",X"9C",X"72",X"25",X"F0",X"AE",X"9F",X"A0",X"72",X"27",
		X"08",X"EF",X"84",X"6F",X"02",X"EF",X"89",X"FF",X"00",X"86",X"07",X"97",X"36",X"B7",X"D0",X"00",
		X"DC",X"20",X"83",X"6D",X"40",X"DD",X"50",X"20",X"1F",X"7F",X"D0",X"00",X"C6",X"04",X"CE",X"CC",
		X"00",X"8E",X"D8",X"0E",X"6F",X"41",X"A6",X"80",X"A7",X"C1",X"A6",X"03",X"A7",X"5F",X"5A",X"26",
		X"F3",X"86",X"02",X"97",X"36",X"7E",X"E8",X"45",X"34",X"16",X"8E",X"C1",X"24",X"BD",X"F7",X"00",
		X"BE",X"A1",X"95",X"E7",X"82",X"35",X"16",X"12",X"12",X"8E",X"4C",X"09",X"CC",X"90",X"90",X"ED",
		X"84",X"ED",X"88",X"1D",X"8E",X"53",X"09",X"CC",X"09",X"09",X"ED",X"84",X"ED",X"88",X"1D",X"8E",
		X"A0",X"42",X"CE",X"B0",X"35",X"8D",X"3A",X"8E",X"A0",X"48",X"8D",X"35",X"DF",X"72",X"DC",X"97",
		X"44",X"44",X"44",X"44",X"54",X"54",X"54",X"C3",X"4B",X"07",X"ED",X"C4",X"AE",X"C4",X"CC",X"90",
		X"99",X"ED",X"84",X"A7",X"02",X"86",X"09",X"A7",X"89",X"FF",X"01",X"39",X"EC",X"0A",X"93",X"50",
		X"44",X"44",X"E6",X"0C",X"54",X"54",X"54",X"BD",X"E8",X"D6",X"ED",X"C4",X"EC",X"88",X"12",X"ED",
		X"D1",X"AE",X"84",X"26",X"E7",X"39",X"FF",X"FF",X"8E",X"EB",X"9C",X"86",X"00",X"BD",X"D0",X"56",
		X"33",X"84",X"BD",X"D0",X"96",X"F9",X"96",X"EC",X"11",X"22",X"22",X"AF",X"47",X"EF",X"06",X"DC",
		X"B7",X"84",X"1F",X"D3",X"20",X"ED",X"0A",X"54",X"CB",X"2A",X"E7",X"0C",X"4F",X"5F",X"ED",X"88",
		X"10",X"ED",X"0E",X"86",X"08",X"A7",X"49",X"8D",X"42",X"7E",X"FC",X"80",X"AE",X"47",X"EC",X"02",
		X"10",X"83",X"F8",X"DF",X"27",X"27",X"6A",X"49",X"26",X"12",X"96",X"D0",X"BD",X"DD",X"C8",X"A7",
		X"49",X"BD",X"EF",X"97",X"27",X"06",X"CC",X"D5",X"D1",X"BD",X"D5",X"ED",X"EE",X"02",X"33",X"4A",
		X"11",X"83",X"F9",X"AA",X"23",X"05",X"CE",X"F9",X"96",X"8D",X"0A",X"EF",X"02",X"86",X"06",X"8E",
		X"EB",X"9C",X"7E",X"D0",X"02",X"96",X"B7",X"91",X"D1",X"23",X"35",X"CC",X"40",X"01",X"DD",X"50",
		X"EC",X"0A",X"93",X"A4",X"2B",X"02",X"00",X"50",X"C3",X"02",X"80",X"10",X"83",X"05",X"00",X"23",
		X"07",X"D6",X"50",X"1D",X"D3",X"9F",X"ED",X"0E",X"A6",X"0C",X"90",X"98",X"2B",X"02",X"00",X"51",
		X"8B",X"0A",X"81",X"14",X"23",X"0A",X"5F",X"96",X"51",X"D3",X"A2",X"47",X"56",X"ED",X"88",X"10",
		X"39",X"0A",X"D9",X"BD",X"F4",X"DA",X"01",X"20",X"D5",X"9F",X"39",X"97",X"50",X"BD",X"D0",X"96",
		X"F8",X"EA",X"EC",X"59",X"CC",X"CC",X"BD",X"D7",X"EF",X"DC",X"B8",X"84",X"3F",X"8B",X"10",X"ED",
		X"0A",X"54",X"CB",X"2A",X"E7",X"0C",X"D6",X"B7",X"C4",X"3F",X"CB",X"E0",X"1D",X"ED",X"0E",X"D6",
		X"B9",X"C4",X"7F",X"C0",X"40",X"1D",X"2B",X"04",X"CA",X"20",X"20",X"02",X"C4",X"DF",X"ED",X"88",
		X"10",X"BD",X"FC",X"80",X"0A",X"50",X"26",X"C5",X"39",X"BD",X"F4",X"E1",X"02",X"10",X"D5",X"95",
		X"86",X"06",X"BD",X"DD",X"C8",X"31",X"84",X"BD",X"EC",X"82",X"0A",X"D4",X"39",X"BD",X"D7",X"EF",
		X"D6",X"B7",X"1D",X"58",X"49",X"ED",X"88",X"10",X"D6",X"B9",X"C4",X"3F",X"CB",X"E0",X"1D",X"ED",
		X"0E",X"39",X"34",X"76",X"97",X"50",X"96",X"D6",X"4C",X"81",X"14",X"22",X"3A",X"97",X"D6",X"8E",
		X"EC",X"F6",X"86",X"00",X"BD",X"D0",X"56",X"33",X"84",X"BD",X"F8",X"FE",X"12",X"12",X"12",X"12",
		X"12",X"12",X"EC",X"2A",X"ED",X"0A",X"EC",X"2C",X"ED",X"0C",X"AF",X"47",X"EF",X"06",X"8D",X"BD",
		X"DC",X"B8",X"D4",X"CE",X"E7",X"49",X"84",X"1F",X"A7",X"44",X"96",X"CD",X"BD",X"DD",X"C8",X"A7",
		X"4B",X"9F",X"42",X"0A",X"50",X"26",X"BF",X"35",X"F6",X"0A",X"D6",X"BD",X"F4",X"BF",X"34",X"10",
		X"BD",X"D0",X"14",X"35",X"10",X"EC",X"0A",X"83",X"00",X"40",X"ED",X"0A",X"EC",X"0C",X"80",X"02",
		X"A7",X"0C",X"CE",X"F8",X"D5",X"EF",X"02",X"BD",X"FC",X"83",X"CC",X"01",X"15",X"BD",X"D4",X"10",
		X"CC",X"D5",X"B8",X"7E",X"D5",X"ED",X"AE",X"47",X"D6",X"CC",X"10",X"9E",X"A4",X"10",X"AC",X"0A",
		X"24",X"01",X"50",X"BD",X"F2",X"62",X"20",X"54",X"E6",X"49",X"AE",X"47",X"96",X"98",X"A1",X"0C",
		X"22",X"01",X"50",X"1D",X"E3",X"88",X"10",X"10",X"83",X"02",X"00",X"2D",X"03",X"CC",X"02",X"00",
		X"10",X"83",X"FE",X"00",X"2E",X"03",X"CC",X"FE",X"00",X"ED",X"88",X"10",X"43",X"53",X"58",X"49",
		X"58",X"49",X"1F",X"89",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"D6",X"B7",X"C4",X"1F",X"CB",
		X"F0",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"DC",X"A4",X"A3",X"0A",X"C3",X"15",X"00",X"10",
		X"83",X"25",X"80",X"22",X"A1",X"6A",X"4B",X"26",X"03",X"BD",X"ED",X"64",X"86",X"03",X"7E",X"F3",
		X"12",X"12",X"12",X"12",X"34",X"10",X"DC",X"A4",X"A3",X"0A",X"A8",X"0E",X"12",X"12",X"31",X"84",
		X"BD",X"E4",X"1C",X"E5",X"02",X"F9",X"4E",X"E5",X"47",X"27",X"22",X"EC",X"2E",X"BD",X"F3",X"4D",
		X"12",X"58",X"49",X"ED",X"0E",X"CC",X"D5",X"D6",X"BD",X"D5",X"ED",X"5F",X"96",X"98",X"A0",X"0C",
		X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",X"88",X"10",X"96",X"CD",X"BD",
		X"DD",X"C8",X"A7",X"4B",X"35",X"90",X"AE",X"47",X"30",X"02",X"8C",X"A1",X"12",X"25",X"03",X"8E",
		X"A0",X"F2",X"AF",X"47",X"86",X"02",X"8E",X"ED",X"A6",X"7E",X"D0",X"02",X"34",X"02",X"30",X"89",
		X"01",X"00",X"B6",X"A1",X"8A",X"84",X"01",X"27",X"02",X"30",X"01",X"35",X"82",X"FF",X"8D",X"12",
		X"26",X"1D",X"34",X"06",X"97",X"51",X"7E",X"DC",X"21",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"34",X"02",X"B6",X"A1",X"8A",X"84",X"02",X"35",X"82",X"FF",X"FF",X"FF",X"FF",X"34",
		X"04",X"D6",X"36",X"34",X"04",X"C6",X"07",X"D7",X"36",X"F7",X"D0",X"00",X"BD",X"C9",X"A0",X"35",
		X"04",X"D7",X"36",X"F7",X"D0",X"00",X"35",X"84",X"FF",X"FF",X"FF",X"05",X"08",X"CD",X"30",X"CD",
		X"58",X"D2",X"43",X"D1",X"CF",X"34",X"02",X"BD",X"ED",X"E2",X"27",X"0A",X"A6",X"0D",X"1C",X"FE",
		X"85",X"01",X"26",X"02",X"1A",X"01",X"35",X"02",X"10",X"DF",X"54",X"7E",X"D2",X"48",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"34",X"14",X"EC",X"0A",X"44",X"56",X"44",X"56",X"44",X"56",
		X"44",X"56",X"44",X"56",X"44",X"56",X"8E",X"B3",X"00",X"A6",X"8B",X"35",X"94",X"CC",X"01",X"30",
		X"BD",X"E5",X"34",X"12",X"8D",X"4B",X"BD",X"F4",X"BF",X"CC",X"F8",X"CB",X"ED",X"02",X"EC",X"0A",
		X"83",X"00",X"40",X"ED",X"0A",X"BD",X"FC",X"83",X"CC",X"D5",X"86",X"7E",X"D5",X"ED",X"EE",X"06",
		X"27",X"DB",X"8D",X"D9",X"7E",X"D0",X"14",X"10",X"83",X"20",X"00",X"23",X"06",X"10",X"83",X"E0",
		X"00",X"23",X"05",X"C3",X"40",X"00",X"ED",X"0A",X"7E",X"FA",X"EE",X"03",X"00",X"00",X"60",X"01",
		X"00",X"00",X"20",X"03",X"00",X"00",X"60",X"02",X"00",X"00",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"31",X"84",X"34",X"52",X"CE",X"A0",X"F2",X"86",X"40",X"10",X"AC",X"C1",X"27",X"06",X"4A",
		X"26",X"F8",X"BD",X"D0",X"3B",X"4F",X"5F",X"ED",X"5E",X"0A",X"BA",X"BE",X"A1",X"95",X"A6",X"82",
		X"B1",X"A1",X"93",X"27",X"02",X"35",X"02",X"35",X"D2",X"8A",X"02",X"97",X"92",X"6F",X"47",X"BD",
		X"F5",X"C3",X"BD",X"C0",X"09",X"8E",X"B0",X"FD",X"CE",X"00",X"00",X"86",X"40",X"EF",X"91",X"4A",
		X"26",X"FB",X"9E",X"44",X"CC",X"F9",X"E4",X"ED",X"02",X"C6",X"02",X"D7",X"50",X"BD",X"D7",X"EF",
		X"84",X"3F",X"D3",X"20",X"ED",X"0A",X"96",X"B7",X"12",X"8A",X"40",X"A7",X"0C",X"BD",X"FC",X"83",
		X"0A",X"50",X"26",X"E9",X"96",X"B7",X"84",X"1F",X"8E",X"E7",X"C0",X"A6",X"86",X"97",X"26",X"CC",
		X"D5",X"86",X"BD",X"D5",X"ED",X"8E",X"EF",X"28",X"86",X"02",X"C6",X"08",X"D7",X"3B",X"7E",X"D0",
		X"02",X"86",X"17",X"97",X"1D",X"7E",X"EE",X"E2",X"0A",X"1D",X"26",X"B6",X"BD",X"EF",X"7C",X"12",
		X"8E",X"E1",X"D8",X"84",X"07",X"A6",X"86",X"97",X"26",X"86",X"01",X"8E",X"DD",X"14",X"7E",X"D0",
		X"02",X"0B",X"34",X"04",X"10",X"83",X"00",X"3F",X"24",X"02",X"C6",X"C6",X"F7",X"C0",X"00",X"35",
		X"04",X"39",X"BD",X"EF",X"6F",X"30",X"89",X"07",X"04",X"39",X"7A",X"A1",X"7B",X"27",X"03",X"7E",
		X"E5",X"F2",X"86",X"01",X"8E",X"EF",X"6A",X"7E",X"D0",X"02",X"8D",X"03",X"7E",X"E5",X"F2",X"86",
		X"01",X"7D",X"BC",X"12",X"27",X"02",X"86",X"07",X"B7",X"A1",X"7B",X"39",X"96",X"36",X"34",X"02",
		X"86",X"01",X"97",X"36",X"B7",X"D0",X"00",X"BD",X"C9",X"27",X"35",X"02",X"97",X"36",X"9E",X"6A",
		X"A6",X"08",X"39",X"FF",X"FF",X"FF",X"FF",X"34",X"10",X"BD",X"E4",X"1C",X"E5",X"02",X"F9",X"4E",
		X"E5",X"47",X"27",X"35",X"D6",X"B7",X"C4",X"1F",X"CB",X"F0",X"DB",X"97",X"E0",X"04",X"1D",X"58",
		X"49",X"58",X"49",X"ED",X"0E",X"D6",X"B7",X"C1",X"78",X"23",X"0A",X"DC",X"9F",X"58",X"49",X"58",
		X"49",X"E3",X"0E",X"ED",X"0E",X"D6",X"B9",X"C4",X"1F",X"CB",X"F0",X"DB",X"98",X"E0",X"05",X"1D",
		X"58",X"49",X"58",X"49",X"ED",X"88",X"10",X"86",X"01",X"35",X"90",X"6A",X"4D",X"26",X"11",X"96",
		X"C5",X"BD",X"DD",X"C8",X"A7",X"4D",X"8D",X"AF",X"27",X"06",X"CC",X"D5",X"C7",X"BD",X"D5",X"ED",
		X"39",X"34",X"02",X"97",X"50",X"8E",X"F2",X"2B",X"86",X"00",X"BD",X"D0",X"56",X"33",X"84",X"BD",
		X"D0",X"96",X"F8",X"C1",X"F0",X"47",X"CC",X"55",X"BD",X"D7",X"EF",X"DC",X"20",X"83",X"25",X"80",
		X"DD",X"52",X"DC",X"B8",X"93",X"52",X"10",X"83",X"4B",X"00",X"24",X"03",X"C3",X"80",X"00",X"D3",
		X"52",X"ED",X"0A",X"96",X"B7",X"44",X"8B",X"2A",X"A7",X"0C",X"4F",X"5F",X"ED",X"88",X"10",X"ED",
		X"0E",X"96",X"CB",X"BD",X"DD",X"C8",X"A7",X"47",X"BD",X"FC",X"80",X"EF",X"06",X"AF",X"47",X"0C",
		X"D5",X"0A",X"50",X"26",X"B0",X"35",X"82",X"0A",X"D5",X"BD",X"F4",X"DA",X"01",X"15",X"D5",X"9A",
		X"39",X"34",X"10",X"96",X"BA",X"27",X"1C",X"9E",X"76",X"30",X"02",X"8C",X"A1",X"32",X"25",X"03",
		X"8E",X"A0",X"F2",X"EC",X"84",X"26",X"06",X"9C",X"76",X"26",X"EE",X"35",X"90",X"9F",X"76",X"ED",
		X"49",X"AF",X"4B",X"35",X"90",X"34",X"02",X"97",X"50",X"0D",X"BA",X"26",X"03",X"7E",X"EF",X"F5",
		X"8E",X"F0",X"CB",X"86",X"00",X"BD",X"D0",X"56",X"33",X"84",X"BD",X"D0",X"96",X"F9",X"78",X"F2",
		X"D2",X"33",X"22",X"BD",X"D7",X"EF",X"7E",X"F6",X"86",X"12",X"86",X"2C",X"A7",X"0C",X"DC",X"C3",
		X"ED",X"88",X"10",X"96",X"C5",X"BD",X"DD",X"C8",X"A7",X"4D",X"96",X"C2",X"BD",X"DD",X"C8",X"1F",
		X"89",X"4F",X"C5",X"01",X"27",X"02",X"53",X"43",X"ED",X"0E",X"EF",X"06",X"BD",X"F6",X"9C",X"AF",
		X"47",X"8D",X"8E",X"0C",X"D2",X"0A",X"50",X"26",X"B0",X"35",X"82",X"AE",X"47",X"10",X"AE",X"49",
		X"EC",X"D8",X"0B",X"27",X"16",X"A6",X"29",X"81",X"4D",X"26",X"10",X"A6",X"0A",X"84",X"FC",X"97",
		X"50",X"A6",X"2A",X"84",X"FC",X"91",X"50",X"27",X"4F",X"20",X"0F",X"A6",X"88",X"14",X"84",X"FE",
		X"A7",X"88",X"14",X"BD",X"F0",X"51",X"10",X"27",X"01",X"14",X"BD",X"EE",X"36",X"80",X"32",X"A0",
		X"0C",X"22",X"0E",X"81",X"EC",X"2D",X"04",X"4F",X"5F",X"20",X"08",X"DC",X"C3",X"43",X"53",X"20",
		X"02",X"DC",X"C3",X"ED",X"88",X"10",X"EC",X"02",X"10",X"83",X"F8",X"DF",X"27",X"12",X"BD",X"EF",
		X"DB",X"EE",X"02",X"33",X"4A",X"11",X"83",X"F9",X"8C",X"23",X"03",X"CE",X"F9",X"78",X"EF",X"02",
		X"86",X"06",X"8E",X"F0",X"CB",X"7E",X"D0",X"02",X"4F",X"5F",X"6C",X"88",X"14",X"ED",X"0E",X"ED",
		X"88",X"10",X"CC",X"F9",X"78",X"ED",X"02",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"27",
		X"9A",X"A6",X"29",X"81",X"4D",X"26",X"94",X"EC",X"2A",X"C4",X"E0",X"DD",X"52",X"EC",X"0A",X"C4",
		X"E0",X"10",X"93",X"52",X"27",X"0D",X"2D",X"04",X"C6",X"E0",X"20",X"02",X"C6",X"20",X"1D",X"E3",
		X"0A",X"ED",X"0A",X"A6",X"2C",X"80",X"0C",X"A1",X"0C",X"27",X"15",X"DC",X"C3",X"24",X"02",X"43",
		X"53",X"12",X"12",X"12",X"12",X"BD",X"EF",X"DB",X"86",X"01",X"8E",X"F1",X"47",X"7E",X"D0",X"02",
		X"EC",X"0A",X"C3",X"00",X"40",X"A3",X"2A",X"10",X"83",X"00",X"80",X"22",X"E8",X"CC",X"F2",X"A7",
		X"ED",X"08",X"DC",X"C3",X"53",X"43",X"ED",X"88",X"10",X"ED",X"A8",X"10",X"CC",X"D5",X"AE",X"BD",
		X"D5",X"ED",X"CC",X"EE",X"6E",X"ED",X"28",X"DE",X"40",X"AE",X"47",X"BD",X"F6",X"3A",X"12",X"25",
		X"0B",X"BD",X"EF",X"DB",X"86",X"04",X"8E",X"F1",X"B7",X"7E",X"D0",X"02",X"CC",X"D5",X"B3",X"BD",
		X"D5",X"ED",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"26",X"0A",X"BD",X"F4",X"BF",X"0A",
		X"D2",X"0C",X"BB",X"7E",X"D0",X"0B",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"A8",X"10",X"A6",X"2C",
		X"A1",X"0C",X"23",X"0F",X"6A",X"2C",X"86",X"12",X"BD",X"D5",X"DB",X"86",X"01",X"8E",X"F1",X"D2",
		X"7E",X"D0",X"02",X"30",X"A4",X"EC",X"24",X"8B",X"01",X"DD",X"F0",X"BD",X"F6",X"6C",X"0A",X"D2",
		X"0C",X"D5",X"AE",X"47",X"6F",X"88",X"14",X"CC",X"F8",X"C1",X"ED",X"02",X"CC",X"55",X"33",X"ED",
		X"88",X"12",X"CC",X"F0",X"47",X"ED",X"08",X"96",X"CB",X"A7",X"49",X"96",X"36",X"34",X"02",X"86",
		X"07",X"97",X"36",X"B7",X"D0",X"00",X"BD",X"C8",X"00",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",
		X"7E",X"F2",X"78",X"34",X"02",X"96",X"90",X"81",X"04",X"24",X"14",X"0C",X"90",X"CC",X"D5",X"BD",
		X"BD",X"D5",X"ED",X"9E",X"99",X"A6",X"E0",X"26",X"03",X"7E",X"E5",X"E8",X"7E",X"E6",X"57",X"7E",
		X"D0",X"0B",X"1D",X"10",X"9E",X"A4",X"0D",X"1A",X"26",X"04",X"58",X"49",X"58",X"49",X"ED",X"0E",
		X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D6",X"C7",X"96",X"B7",X"2B",X"01",X"50",X"EB",
		X"0C",X"C1",X"2A",X"24",X"02",X"C6",X"2F",X"E7",X"0C",X"6A",X"49",X"26",X"12",X"96",X"CB",X"BD",
		X"DD",X"C8",X"A7",X"49",X"BD",X"EF",X"97",X"27",X"06",X"CC",X"D5",X"CC",X"BD",X"D5",X"ED",X"86",
		X"0F",X"8E",X"F2",X"2B",X"7E",X"D0",X"02",X"EE",X"06",X"EC",X"D8",X"0B",X"27",X"24",X"CC",X"00",
		X"00",X"CC",X"00",X"00",X"34",X"10",X"8E",X"F2",X"DC",X"86",X"00",X"BD",X"D0",X"56",X"EE",X"49",
		X"EF",X"07",X"CC",X"D5",X"8B",X"BD",X"D5",X"ED",X"CC",X"00",X"00",X"ED",X"C8",X"10",X"AF",X"46",
		X"35",X"10",X"0A",X"D2",X"BD",X"F4",X"DA",X"01",X"15",X"D5",X"A9",X"39",X"AE",X"47",X"CC",X"00",
		X"08",X"E3",X"88",X"10",X"10",X"83",X"03",X"00",X"24",X"03",X"ED",X"88",X"10",X"BD",X"F6",X"34",
		X"A1",X"0C",X"22",X"16",X"EC",X"88",X"10",X"10",X"83",X"00",X"E0",X"12",X"12",X"EC",X"04",X"C3",
		X"01",X"07",X"DD",X"F0",X"BD",X"EE",X"54",X"7E",X"D0",X"0B",X"86",X"04",X"8E",X"F2",X"DC",X"7E",
		X"D0",X"02",X"F6",X"A1",X"8A",X"C4",X"01",X"27",X"12",X"34",X"40",X"CE",X"F9",X"BE",X"6D",X"0E",
		X"2B",X"03",X"CE",X"F9",X"D0",X"EF",X"02",X"35",X"40",X"86",X"03",X"8E",X"ED",X"08",X"7E",X"D0",
		X"02",X"B6",X"A1",X"8A",X"84",X"01",X"26",X"07",X"86",X"2A",X"97",X"1B",X"7E",X"E9",X"89",X"BD",
		X"EE",X"36",X"80",X"08",X"97",X"1B",X"86",X"E0",X"97",X"1C",X"7E",X"E9",X"A1",X"34",X"02",X"B6",
		X"A1",X"8A",X"84",X"01",X"27",X"02",X"35",X"82",X"35",X"02",X"58",X"49",X"58",X"49",X"39",X"FF",
		X"FF",X"FF",X"FF",X"97",X"50",X"D6",X"C6",X"03",X"85",X"2B",X"01",X"50",X"D7",X"51",X"8E",X"F3",
		X"BC",X"86",X"00",X"BD",X"D0",X"3F",X"33",X"84",X"96",X"50",X"A7",X"4F",X"4F",X"5F",X"ED",X"47",
		X"ED",X"49",X"ED",X"4B",X"ED",X"4D",X"BD",X"D0",X"96",X"F9",X"1C",X"F4",X"81",X"55",X"55",X"D6",
		X"51",X"1D",X"ED",X"0E",X"4F",X"5F",X"ED",X"88",X"10",X"96",X"50",X"44",X"56",X"9B",X"50",X"D3",
		X"A4",X"8B",X"80",X"ED",X"0A",X"86",X"50",X"A7",X"0C",X"A7",X"C8",X"10",X"EF",X"06",X"9F",X"42",
		X"96",X"50",X"48",X"8B",X"05",X"AF",X"C6",X"0A",X"50",X"26",X"CB",X"39",X"96",X"B7",X"84",X"06",
		X"8B",X"07",X"AE",X"C6",X"10",X"27",X"00",X"B1",X"D6",X"B7",X"86",X"0A",X"C4",X"3F",X"CB",X"E0",
		X"2B",X"01",X"40",X"10",X"AE",X"02",X"31",X"A6",X"10",X"8C",X"F9",X"1C",X"24",X"04",X"10",X"8E",
		X"F9",X"1C",X"10",X"8C",X"F9",X"3A",X"23",X"04",X"10",X"8E",X"F9",X"3A",X"10",X"AF",X"02",X"1D",
		X"E3",X"88",X"10",X"ED",X"88",X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"1F",X"89",X"50",X"1D",
		X"E3",X"88",X"10",X"ED",X"88",X"10",X"A6",X"05",X"26",X"3B",X"96",X"B7",X"81",X"40",X"22",X"16",
		X"84",X"03",X"8B",X"FE",X"AB",X"C8",X"10",X"81",X"40",X"24",X"02",X"86",X"40",X"81",X"68",X"25",
		X"02",X"86",X"68",X"A7",X"C8",X"10",X"A6",X"C8",X"10",X"A0",X"0C",X"8B",X"10",X"81",X"20",X"23",
		X"48",X"80",X"10",X"2B",X"05",X"CC",X"FF",X"F0",X"20",X"03",X"CC",X"00",X"10",X"E3",X"88",X"10",
		X"ED",X"88",X"10",X"20",X"34",X"90",X"98",X"2B",X"12",X"81",X"20",X"25",X"05",X"CC",X"FF",X"F0",
		X"20",X"19",X"81",X"10",X"22",X"1B",X"CC",X"00",X"10",X"20",X"10",X"81",X"E0",X"2E",X"05",X"CC",
		X"00",X"10",X"20",X"07",X"81",X"F0",X"2D",X"09",X"CC",X"FF",X"F0",X"E3",X"88",X"10",X"ED",X"88",
		X"10",X"96",X"B9",X"84",X"07",X"26",X"02",X"8D",X"27",X"86",X"01",X"8E",X"F3",X"BC",X"7E",X"D0",
		X"02",X"BD",X"F4",X"E1",X"01",X"25",X"D5",X"A4",X"0A",X"D3",X"EE",X"06",X"31",X"47",X"AC",X"A1",
		X"26",X"FC",X"4F",X"5F",X"ED",X"3E",X"6A",X"4F",X"26",X"05",X"30",X"C4",X"BD",X"D0",X"16",X"39",
		X"96",X"74",X"81",X"0A",X"24",X"18",X"BD",X"E4",X"1C",X"E4",X"C1",X"F9",X"4E",X"E5",X"47",X"27",
		X"0D",X"D6",X"B8",X"1D",X"58",X"49",X"96",X"B7",X"84",X"1F",X"4C",X"A7",X"88",X"15",X"39",X"BD",
		X"D0",X"C8",X"34",X"76",X"BD",X"F5",X"C7",X"EC",X"04",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"35",
		X"F6",X"34",X"10",X"BD",X"D0",X"14",X"35",X"10",X"20",X"0A",X"34",X"10",X"BD",X"D0",X"14",X"35",
		X"10",X"BD",X"D0",X"C8",X"34",X"46",X"EE",X"64",X"37",X"06",X"BD",X"D4",X"10",X"8D",X"09",X"37",
		X"06",X"EF",X"64",X"BD",X"D5",X"ED",X"35",X"C6",X"34",X"76",X"8D",X"C6",X"BD",X"FC",X"83",X"35",
		X"F6",X"8E",X"F5",X"1F",X"AF",X"47",X"86",X"06",X"8E",X"F5",X"0E",X"7E",X"D0",X"02",X"AE",X"47",
		X"EC",X"81",X"DD",X"33",X"A6",X"80",X"97",X"35",X"8C",X"F5",X"28",X"25",X"E7",X"20",X"E2",X"81",
		X"81",X"2F",X"81",X"2F",X"07",X"2F",X"81",X"07",X"86",X"FF",X"97",X"30",X"0F",X"32",X"86",X"03",
		X"8E",X"F5",X"36",X"7E",X"D0",X"02",X"96",X"B7",X"84",X"1F",X"8E",X"E7",X"C0",X"A6",X"86",X"97",
		X"30",X"97",X"32",X"8E",X"CC",X"B0",X"9C",X"81",X"26",X"03",X"8E",X"CC",X"BC",X"9F",X"81",X"86",
		X"06",X"8E",X"F5",X"28",X"7E",X"D0",X"02",X"96",X"67",X"26",X"24",X"8E",X"0F",X"1C",X"96",X"68",
		X"4A",X"27",X"03",X"8E",X"71",X"1C",X"CC",X"18",X"08",X"BD",X"D1",X"9F",X"86",X"08",X"8E",X"F5",
		X"74",X"7E",X"D0",X"02",X"BD",X"D4",X"89",X"86",X"0C",X"8E",X"F5",X"57",X"7E",X"D0",X"02",X"7E",
		X"D0",X"0B",X"DE",X"40",X"AF",X"4D",X"D6",X"36",X"E7",X"4C",X"8E",X"F5",X"90",X"7E",X"D0",X"02",
		X"A6",X"4C",X"8D",X"3D",X"6E",X"D8",X"0D",X"32",X"7D",X"34",X"42",X"96",X"36",X"A7",X"65",X"EE",
		X"66",X"A6",X"42",X"EE",X"C4",X"EF",X"63",X"8D",X"28",X"35",X"42",X"AD",X"F4",X"34",X"42",X"A6",
		X"65",X"8D",X"1E",X"EE",X"66",X"33",X"43",X"EF",X"66",X"35",X"42",X"32",X"63",X"39",X"8D",X"03",
		X"7E",X"C0",X"00",X"86",X"07",X"20",X"0A",X"86",X"02",X"20",X"06",X"86",X"03",X"20",X"02",X"86",
		X"01",X"97",X"36",X"B7",X"D0",X"00",X"39",X"34",X"7F",X"8D",X"EC",X"BD",X"C0",X"02",X"35",X"FF",
		X"8D",X"E9",X"7E",X"C0",X"0F",X"FF",X"FF",X"7F",X"D0",X"00",X"8E",X"CC",X"00",X"6F",X"01",X"6F",
		X"03",X"6F",X"05",X"6F",X"07",X"86",X"C0",X"A7",X"84",X"86",X"00",X"A7",X"02",X"6F",X"04",X"6F",
		X"06",X"86",X"04",X"A7",X"03",X"A7",X"05",X"A7",X"07",X"8A",X"10",X"A7",X"01",X"8E",X"C0",X"00",
		X"86",X"C0",X"A7",X"80",X"C6",X"B5",X"3D",X"8C",X"C0",X"10",X"26",X"F6",X"1A",X"80",X"1C",X"EF",
		X"10",X"8E",X"00",X"01",X"4F",X"1F",X"8B",X"1C",X"BF",X"86",X"9E",X"1F",X"8B",X"10",X"CE",X"C0",
		X"00",X"7E",X"FB",X"20",X"BD",X"EE",X"36",X"80",X"10",X"39",X"EC",X"10",X"BD",X"E9",X"53",X"A6",
		X"0C",X"90",X"1B",X"8B",X"10",X"81",X"20",X"39",X"4F",X"97",X"1A",X"BD",X"F5",X"C3",X"BD",X"C0",
		X"06",X"BD",X"C0",X"00",X"BD",X"F5",X"CF",X"BD",X"F7",X"99",X"7E",X"F7",X"87",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"32",X"7F",X"6F",X"E4",X"BD",X"F0",X"75",X"32",X"61",X"39",X"BD",X"EE",X"54",X"34",
		X"40",X"AE",X"47",X"A6",X"0C",X"34",X"02",X"EC",X"0A",X"34",X"06",X"86",X"01",X"34",X"02",X"BD",
		X"F0",X"75",X"32",X"64",X"35",X"C0",X"6D",X"63",X"26",X"07",X"DC",X"B8",X"ED",X"0A",X"7E",X"F0",
		X"9A",X"EC",X"64",X"ED",X"0A",X"A6",X"66",X"A7",X"0C",X"7E",X"F0",X"9E",X"6D",X"65",X"26",X"04",
		X"BD",X"FC",X"80",X"39",X"9F",X"42",X"39",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"39",X"BD",X"FF",
		X"CE",X"C0",X"05",X"02",X"39",X"BD",X"E6",X"E4",X"26",X"0C",X"BD",X"F7",X"36",X"26",X"07",X"0D",
		X"1A",X"27",X"03",X"BD",X"F7",X"68",X"39",X"40",X"33",X"30",X"30",X"2F",X"40",X"32",X"35",X"30",
		X"2F",X"40",X"32",X"30",X"30",X"2F",X"40",X"31",X"35",X"30",X"2F",X"40",X"31",X"30",X"30",X"2F",
		X"BD",X"E6",X"E4",X"27",X"01",X"39",X"B6",X"A1",X"8A",X"84",X"01",X"26",X"03",X"7E",X"F6",X"BA",
		X"BD",X"F7",X"68",X"4A",X"39",X"34",X"10",X"9E",X"6A",X"A6",X"08",X"4A",X"84",X"07",X"35",X"90",
		X"34",X"20",X"96",X"36",X"34",X"02",X"10",X"BE",X"A1",X"98",X"B6",X"A1",X"97",X"97",X"36",X"B7",
		X"D4",X"9E",X"E6",X"A9",X"00",X"D9",X"A6",X"A9",X"00",X"95",X"E6",X"A9",X"07",X"50",X"A6",X"84",
		X"E6",X"A9",X"03",X"56",X"35",X"02",X"97",X"36",X"B7",X"DE",X"98",X"35",X"A0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8D",X"23",X"34",X"06",X"8E",X"BC",X"F1",X"E6",X"8B",X"27",
		X"17",X"5C",X"D0",X"B1",X"35",X"06",X"23",X"0D",X"C3",X"00",X"10",X"E6",X"8B",X"C0",X"05",X"D0",
		X"AF",X"23",X"02",X"4F",X"39",X"86",X"01",X"39",X"4F",X"35",X"86",X"4F",X"C6",X"98",X"D0",X"B0",
		X"58",X"49",X"58",X"49",X"C3",X"00",X"08",X"39",X"8D",X"F1",X"34",X"06",X"8E",X"BC",X"F3",X"E6",
		X"8B",X"27",X"E5",X"5C",X"D0",X"B1",X"35",X"06",X"24",X"DB",X"C3",X"00",X"10",X"E6",X"8B",X"C0",
		X"05",X"D0",X"AF",X"24",X"D0",X"4F",X"39",X"34",X"16",X"8E",X"C3",X"A6",X"BD",X"F7",X"00",X"BE",
		X"A1",X"95",X"E7",X"84",X"35",X"16",X"7E",X"D0",X"7D",X"34",X"32",X"8E",X"A1",X"92",X"10",X"8E",
		X"F7",X"AD",X"A6",X"A0",X"A7",X"80",X"8C",X"A1",X"9A",X"26",X"F7",X"35",X"B2",X"31",X"62",X"E2",
		X"A1",X"91",X"09",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"86",X"03",X"97",X"36",X"B7",X"D0",
		X"00",X"BD",X"C0",X"00",X"BD",X"C0",X"09",X"7E",X"D8",X"16",X"34",X"03",X"96",X"36",X"34",X"02",
		X"0F",X"36",X"7F",X"D0",X"00",X"E7",X"84",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"83",
		X"34",X"03",X"96",X"36",X"34",X"02",X"0F",X"36",X"7F",X"D0",X"00",X"E6",X"84",X"20",X"E8",X"34",
		X"06",X"7F",X"B2",X"18",X"7F",X"B2",X"0F",X"86",X"03",X"97",X"36",X"B7",X"B2",X"0E",X"CC",X"FF",
		X"FF",X"FD",X"B2",X"1F",X"35",X"86",X"A6",X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",
		X"48",X"48",X"AB",X"E0",X"39",X"34",X"04",X"D6",X"36",X"34",X"04",X"0F",X"36",X"7F",X"D0",X"00",
		X"8D",X"E4",X"35",X"04",X"D7",X"36",X"F7",X"D0",X"00",X"35",X"84",X"8D",X"E8",X"34",X"02",X"8D",
		X"E4",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",X"A7",X"81",X"35",
		X"82",X"34",X"04",X"D6",X"36",X"34",X"04",X"0F",X"36",X"7F",X"D0",X"00",X"8D",X"E7",X"35",X"04",
		X"D7",X"36",X"F7",X"D0",X"00",X"35",X"84",X"8D",X"E8",X"34",X"02",X"1F",X"98",X"8D",X"E2",X"35",
		X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E5",X"BB",X"00",X"E8",X"00",X"00",X"00",
		X"00",X"E8",X"E8",X"00",X"F8",X"E9",X"46",X"00",X"F8",X"D9",X"18",X"00",X"00",X"D9",X"03",X"00",
		X"00",X"E8",X"BE",X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"F9",X"00",
		X"00",X"D5",X"22",X"02",X"00",X"D4",X"ED",X"00",X"00",X"D5",X"1B",X"02",X"00",X"D5",X"29",X"02",
		X"00",X"00",X"00",X"07",X"28",X"2F",X"81",X"A4",X"15",X"C7",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"08",X"F9",X"EE",X"FA",X"16",X"D2",X"43",X"D1",X"CF",X"04",X"08",X"FA",X"3E",X"FA",
		X"3E",X"D1",X"E9",X"D2",X"1B",X"04",X"08",X"FA",X"5E",X"FA",X"5E",X"D1",X"E9",X"D2",X"1B",X"01",
		X"01",X"F8",X"E9",X"F8",X"E9",X"D9",X"96",X"D9",X"96",X"00",X"05",X"08",X"FA",X"A6",X"FA",X"A6",
		X"E9",X"A3",X"E9",X"BE",X"02",X"08",X"FA",X"CE",X"FA",X"DE",X"D1",X"A9",X"D1",X"BB",X"B6",X"A1",
		X"8A",X"84",X"01",X"26",X"0A",X"BD",X"D0",X"96",X"F9",X"6E",X"EC",X"C9",X"88",X"88",X"39",X"BD",
		X"D0",X"96",X"F9",X"BE",X"EC",X"C9",X"33",X"33",X"39",X"FF",X"FF",X"FF",X"04",X"08",X"FB",X"5E",
		X"FB",X"5E",X"D1",X"E9",X"D2",X"1B",X"04",X"08",X"FB",X"5E",X"FB",X"5E",X"D1",X"E9",X"D2",X"1B",
		X"04",X"08",X"FB",X"5E",X"FB",X"5E",X"D1",X"E9",X"D2",X"1B",X"04",X"08",X"FB",X"5E",X"FB",X"5E",
		X"D1",X"E9",X"D2",X"1B",X"04",X"08",X"CC",X"90",X"CC",X"90",X"D1",X"E9",X"D2",X"1B",X"02",X"03",
		X"CC",X"B0",X"CC",X"B6",X"D2",X"A1",X"D2",X"BD",X"02",X"03",X"CC",X"BC",X"CC",X"C2",X"D2",X"A1",
		X"D2",X"BD",X"08",X"01",X"F9",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"04",
		X"CC",X"C8",X"CC",X"C8",X"D2",X"5D",X"D2",X"87",X"04",X"08",X"CC",X"E0",X"CD",X"08",X"D2",X"43",
		X"D1",X"CF",X"04",X"08",X"CC",X"E0",X"CD",X"08",X"D2",X"43",X"D1",X"CF",X"04",X"08",X"CC",X"E0",
		X"CD",X"08",X"D2",X"43",X"D1",X"CF",X"06",X"04",X"CD",X"D0",X"CD",X"D0",X"D2",X"CF",X"D3",X"10",
		X"06",X"04",X"CD",X"D0",X"CD",X"D0",X"D2",X"CF",X"D3",X"10",X"06",X"04",X"CD",X"D0",X"CD",X"D0",
		X"D2",X"CF",X"D3",X"10",X"08",X"06",X"CE",X"60",X"CE",X"60",X"D3",X"3E",X"D3",X"8F",X"08",X"06",
		X"CE",X"C0",X"CE",X"C0",X"D3",X"3E",X"D3",X"8F",X"05",X"04",X"CF",X"20",X"03",X"03",X"CF",X"34",
		X"08",X"06",X"CE",X"F0",X"CE",X"F0",X"D3",X"3E",X"D3",X"8F",X"02",X"08",X"CF",X"3D",X"CF",X"3D",
		X"D1",X"A9",X"D1",X"BB",X"08",X"06",X"CF",X"CD",X"CF",X"CD",X"D0",X"FA",X"D1",X"53",X"C0",X"C0",
		X"0C",X"00",X"08",X"88",X"00",X"00",X"00",X"00",X"08",X"82",X"23",X"88",X"83",X"08",X"00",X"88",
		X"22",X"33",X"33",X"22",X"33",X"33",X"00",X"00",X"50",X"15",X"31",X"55",X"35",X"50",X"0C",X"0C",
		X"C0",X"00",X"50",X"55",X"00",X"00",X"C0",X"C0",X"0C",X"00",X"05",X"55",X"00",X"00",X"00",X"00",
		X"05",X"52",X"23",X"55",X"53",X"05",X"00",X"55",X"22",X"33",X"33",X"22",X"33",X"33",X"00",X"00",
		X"80",X"18",X"31",X"88",X"38",X"80",X"0C",X"0C",X"C0",X"00",X"80",X"88",X"00",X"00",X"00",X"00",
		X"0D",X"6C",X"6C",X"0D",X"00",X"00",X"06",X"E6",X"C8",X"83",X"82",X"C8",X"EC",X"06",X"60",X"6D",
		X"8C",X"28",X"28",X"8C",X"6D",X"60",X"00",X"00",X"E0",X"C6",X"C6",X"E0",X"00",X"00",X"00",X"00",
		X"02",X"22",X"24",X"02",X"00",X"00",X"02",X"22",X"44",X"44",X"24",X"42",X"22",X"00",X"20",X"22",
		X"44",X"44",X"24",X"42",X"22",X"00",X"00",X"00",X"20",X"22",X"22",X"20",X"00",X"00",X"34",X"02",
		X"6F",X"D8",X"0B",X"B6",X"A1",X"8A",X"84",X"01",X"26",X"04",X"6C",X"4B",X"35",X"82",X"CC",X"01",
		X"01",X"E3",X"4B",X"ED",X"4B",X"35",X"82",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"5C",X"5C",X"5C",X"5C",X"50",X"50",X"00",X"00",
		X"06",X"CC",X"CC",X"06",X"00",X"00",X"00",X"66",X"00",X"FF",X"FF",X"00",X"66",X"00",X"00",X"00",
		X"60",X"CC",X"CC",X"60",X"00",X"00",X"05",X"05",X"C5",X"C5",X"C5",X"C5",X"05",X"05",X"05",X"15",
		X"55",X"06",X"66",X"06",X"06",X"06",X"50",X"51",X"55",X"60",X"66",X"60",X"60",X"60",X"05",X"15",
		X"55",X"06",X"66",X"06",X"60",X"60",X"50",X"51",X"55",X"60",X"66",X"60",X"06",X"06",X"34",X"40",
		X"DE",X"6A",X"A6",X"48",X"84",X"03",X"48",X"48",X"34",X"02",X"CE",X"EE",X"8B",X"EC",X"C6",X"ED",
		X"88",X"10",X"35",X"02",X"33",X"42",X"EC",X"C6",X"7C",X"A1",X"7C",X"34",X"02",X"B6",X"A1",X"7C",
		X"85",X"01",X"35",X"02",X"26",X"05",X"43",X"53",X"C3",X"00",X"01",X"ED",X"0E",X"35",X"C0",X"12",
		X"86",X"09",X"B7",X"D7",X"49",X"8E",X"C0",X"00",X"86",X"AA",X"A7",X"84",X"A7",X"84",X"A7",X"84",
		X"8E",X"C0",X"04",X"86",X"55",X"A7",X"84",X"A7",X"84",X"A7",X"84",X"7E",X"F7",X"BA",X"7F",X"10",
		X"DD",X"CC",X"00",X"02",X"EE",X"88",X"6F",X"08",X"BB",X"44",X"FF",X"00",X"77",X"77",X"6F",X"10",
		X"AA",X"66",X"00",X"02",X"CC",X"88",X"5F",X"0A",X"99",X"44",X"FF",X"00",X"77",X"77",X"00",X"00",
		X"55",X"00",X"00",X"55",X"00",X"00",X"05",X"50",X"0D",X"DE",X"DE",X"0D",X"50",X"05",X"50",X"05",
		X"D0",X"ED",X"ED",X"D0",X"05",X"50",X"00",X"00",X"55",X"00",X"00",X"55",X"00",X"00",X"F8",X"EA",
		X"F8",X"F4",X"F9",X"1C",X"F9",X"96",X"F9",X"6E",X"F8",X"C1",X"F9",X"78",X"FB",X"AA",X"FB",X"AC",
		X"FB",X"AE",X"FB",X"B0",X"FB",X"B2",X"FB",X"B4",X"FB",X"B6",X"FB",X"B8",X"FB",X"BA",X"FB",X"BC",
		X"FB",X"BE",X"FB",X"C0",X"FB",X"C2",X"FB",X"C4",X"FB",X"C6",X"C5",X"01",X"FB",X"C6",X"C3",X"6E",
		X"C3",X"5A",X"C5",X"76",X"C4",X"B2",X"C4",X"84",X"C4",X"C9",X"F6",X"C7",X"F6",X"CC",X"F6",X"D1",
		X"F6",X"D6",X"F6",X"D6",X"F6",X"DB",X"44",X"52",X"4F",X"4E",X"45",X"2F",X"33",X"30",X"30",X"2F",
		X"E6",X"A0",X"8D",X"18",X"E6",X"A0",X"8D",X"1B",X"81",X"3F",X"26",X"F4",X"86",X"61",X"E6",X"A2",
		X"8D",X"0A",X"E6",X"A2",X"8D",X"0D",X"81",X"72",X"26",X"F4",X"35",X"A0",X"1E",X"10",X"ED",X"84",
		X"1E",X"01",X"39",X"1E",X"10",X"ED",X"84",X"1E",X"01",X"4C",X"39",X"FF",X"FF",X"FF",X"18",X"18",
		X"17",X"19",X"16",X"1A",X"15",X"1B",X"14",X"1C",X"13",X"1D",X"12",X"1E",X"11",X"1F",X"10",X"20",
		X"0F",X"21",X"0E",X"22",X"0D",X"23",X"0C",X"24",X"0B",X"25",X"0A",X"26",X"09",X"27",X"08",X"28",
		X"CC",X"D5",X"B3",X"BD",X"D5",X"ED",X"86",X"7F",X"B7",X"BC",X"12",X"FC",X"BC",X"10",X"83",X"00",
		X"01",X"FD",X"BC",X"10",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"FC",X"89",X"7E",X"FC",X"EC",X"7E",X"FD",X"4D",X"34",X"66",X"EC",X"02",X"34",X"06",X"FC",
		X"FF",X"A0",X"ED",X"02",X"9F",X"42",X"EC",X"0A",X"93",X"20",X"10",X"83",X"26",X"00",X"22",X"17",
		X"10",X"9E",X"DA",X"27",X"09",X"31",X"A8",X"40",X"10",X"8C",X"A0",X"00",X"26",X"04",X"10",X"8E",
		X"9C",X"00",X"10",X"9C",X"DA",X"26",X"06",X"35",X"06",X"ED",X"02",X"20",X"2D",X"A6",X"A4",X"2B",
		X"E4",X"27",X"03",X"BD",X"FD",X"F5",X"96",X"92",X"85",X"80",X"26",X"06",X"FC",X"FF",X"DD",X"BD",
		X"FF",X"DA",X"A6",X"88",X"14",X"8A",X"02",X"A7",X"88",X"14",X"CC",X"AF",X"00",X"ED",X"A4",X"35",
		X"06",X"ED",X"22",X"33",X"A8",X"40",X"EF",X"24",X"AF",X"2A",X"35",X"E6",X"34",X"66",X"EC",X"0A",
		X"93",X"20",X"81",X"26",X"22",X"55",X"DD",X"E1",X"10",X"9E",X"DA",X"27",X"09",X"31",X"A8",X"40",
		X"10",X"8C",X"A0",X"00",X"26",X"04",X"10",X"8E",X"9C",X"00",X"10",X"9C",X"DA",X"27",X"3C",X"A6",
		X"A4",X"2B",X"EA",X"27",X"03",X"BD",X"FD",X"F5",X"10",X"9F",X"DA",X"CC",X"01",X"00",X"ED",X"A4",
		X"EC",X"02",X"ED",X"22",X"33",X"A8",X"40",X"EF",X"24",X"DC",X"E1",X"58",X"49",X"58",X"49",X"E6",
		X"0C",X"ED",X"28",X"93",X"F0",X"EE",X"22",X"AB",X"C4",X"24",X"08",X"EB",X"41",X"24",X"04",X"DC",
		X"F0",X"20",X"06",X"EC",X"C4",X"44",X"54",X"E3",X"28",X"ED",X"26",X"35",X"E6",X"10",X"8E",X"9C",
		X"00",X"96",X"92",X"85",X"04",X"27",X"0C",X"A6",X"A4",X"2B",X"56",X"CC",X"00",X"00",X"ED",X"A4",
		X"7E",X"FD",X"E9",X"EC",X"A4",X"10",X"27",X"00",X"80",X"2B",X"33",X"C3",X"00",X"AA",X"ED",X"A4",
		X"81",X"30",X"23",X"0A",X"BD",X"FD",X"F5",X"CC",X"00",X"00",X"ED",X"A4",X"20",X"6B",X"DC",X"20",
		X"C4",X"C0",X"34",X"06",X"DC",X"22",X"C4",X"C0",X"A3",X"E1",X"58",X"49",X"58",X"49",X"34",X"02",
		X"A6",X"26",X"AB",X"E4",X"A7",X"26",X"A6",X"28",X"AB",X"E0",X"A7",X"28",X"20",X"45",X"83",X"01",
		X"00",X"ED",X"A4",X"2A",X"0C",X"AE",X"2A",X"EC",X"0A",X"93",X"20",X"8B",X"0C",X"85",X"C0",X"27",
		X"18",X"CC",X"00",X"00",X"ED",X"A4",X"EC",X"22",X"AE",X"2A",X"ED",X"02",X"A6",X"88",X"14",X"84",
		X"FD",X"A7",X"88",X"14",X"BD",X"FD",X"F5",X"20",X"20",X"80",X"0C",X"58",X"49",X"58",X"49",X"E6",
		X"0C",X"ED",X"28",X"C6",X"DA",X"3D",X"48",X"EE",X"22",X"E6",X"C4",X"3D",X"E6",X"41",X"54",X"E3",
		X"28",X"ED",X"26",X"BD",X"FD",X"F5",X"BD",X"FE",X"0F",X"31",X"A8",X"40",X"10",X"8C",X"A0",X"00",
		X"10",X"26",X"FF",X"5D",X"39",X"34",X"16",X"CC",X"00",X"00",X"30",X"A8",X"40",X"9F",X"EB",X"AE",
		X"24",X"9C",X"EB",X"27",X"08",X"ED",X"91",X"9C",X"EB",X"26",X"FA",X"AF",X"24",X"35",X"96",X"34",
		X"76",X"10",X"9F",X"EE",X"A6",X"A4",X"84",X"7F",X"97",X"DF",X"33",X"A8",X"40",X"0F",X"DE",X"AE",
		X"22",X"EC",X"02",X"DD",X"EB",X"EC",X"84",X"97",X"E9",X"D7",X"EA",X"C5",X"01",X"26",X"05",X"8E",
		X"FF",X"47",X"20",X"03",X"8E",X"FF",X"13",X"9F",X"E5",X"EC",X"26",X"A3",X"28",X"97",X"DC",X"54",
		X"D7",X"DD",X"09",X"DE",X"96",X"DF",X"D6",X"DC",X"3D",X"DD",X"E1",X"E6",X"26",X"4F",X"93",X"E1",
		X"DD",X"E1",X"4D",X"27",X"18",X"DC",X"EB",X"DB",X"EA",X"89",X"00",X"DD",X"EB",X"0A",X"E9",X"10",
		X"27",X"00",X"F2",X"DC",X"E1",X"DB",X"DF",X"89",X"00",X"DD",X"E1",X"20",X"E5",X"C1",X"98",X"10",
		X"22",X"00",X"E2",X"96",X"DF",X"48",X"97",X"E0",X"D6",X"DD",X"3D",X"DD",X"E3",X"E6",X"27",X"4F",
		X"93",X"E3",X"D0",X"DE",X"89",X"00",X"0F",X"ED",X"4D",X"26",X"04",X"C1",X"2A",X"24",X"10",X"0C",
		X"ED",X"0A",X"EA",X"0A",X"EA",X"10",X"2F",X"00",X"BC",X"DB",X"E0",X"89",X"00",X"20",X"E9",X"DD",
		X"E3",X"96",X"EA",X"84",X"FE",X"8E",X"FF",X"68",X"AE",X"86",X"9F",X"E7",X"9E",X"EB",X"08",X"ED",
		X"96",X"E2",X"D6",X"ED",X"3A",X"D6",X"E4",X"6E",X"9F",X"A0",X"E7",X"ED",X"C3",X"10",X"AE",X"81",
		X"10",X"AF",X"D4",X"DB",X"E0",X"25",X"56",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",
		X"E0",X"25",X"50",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E0",X"25",X"4A",X"ED",
		X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E0",X"25",X"44",X"ED",X"C3",X"10",X"AE",X"81",
		X"10",X"AF",X"D4",X"DB",X"E0",X"25",X"3E",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",
		X"E0",X"25",X"38",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E0",X"25",X"32",X"6E",
		X"9F",X"A0",X"E5",X"25",X"30",X"ED",X"C3",X"E6",X"80",X"E7",X"D4",X"20",X"2A",X"30",X"0C",X"6E",
		X"9F",X"A0",X"E5",X"30",X"0A",X"6E",X"9F",X"A0",X"E5",X"30",X"08",X"6E",X"9F",X"A0",X"E5",X"30",
		X"06",X"6E",X"9F",X"A0",X"E5",X"30",X"04",X"6E",X"9F",X"A0",X"E5",X"30",X"02",X"6E",X"9F",X"A0",
		X"E5",X"6E",X"9F",X"A0",X"E5",X"30",X"01",X"0A",X"E9",X"27",X"0A",X"9B",X"DF",X"25",X"06",X"81",
		X"98",X"10",X"23",X"FF",X"5D",X"9E",X"EE",X"EF",X"04",X"EC",X"06",X"81",X"98",X"22",X"07",X"D0",
		X"DE",X"8E",X"00",X"00",X"AF",X"8B",X"35",X"F6",X"FF",X"0F",X"FF",X"03",X"FE",X"F7",X"FE",X"EB",
		X"FE",X"DF",X"FE",X"D3",X"FE",X"C7",X"FE",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"DF",X"F8",X"61",X"7E",X"F8",X"15",X"7E",X"F8",X"2D",X"7E",X"F8",X"2B",X"7E",X"F8",X"41",
		X"7E",X"F8",X"59",X"7E",X"F8",X"57",X"7E",X"D0",X"FA",X"7E",X"D1",X"53",X"7E",X"D7",X"8E",X"7E",
		X"F7",X"22",X"7E",X"F7",X"78",X"7E",X"F6",X"2A",X"7E",X"F7",X"C4",X"7E",X"F5",X"BE",X"7E",X"F5",
		X"97",X"7E",X"F5",X"82",X"7E",X"F7",X"CA",X"7E",X"F7",X"E0",X"7E",X"D5",X"ED",X"D5",X"90",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F5",X"E7",X"F5",X"E7",X"F5",X"E7",X"F5",X"E7",X"E9",X"0B",X"F5",X"E7",X"F5",X"E7",X"F5",X"E7",
		X"BD",X"D0",X"7D",X"86",X"FF",X"B7",X"A0",X"92",X"BD",X"E0",X"9D",X"B6",X"A0",X"37",X"B7",X"A1",
		X"59",X"4F",X"B7",X"A1",X"5A",X"B7",X"A1",X"4E",X"8E",X"C8",X"D8",X"86",X"00",X"BD",X"D0",X"56",
		X"10",X"8E",X"A1",X"9A",X"86",X"01",X"B7",X"A0",X"06",X"10",X"BF",X"A1",X"51",X"8E",X"B2",X"90",
		X"BD",X"C1",X"38",X"10",X"24",X"00",X"E3",X"7C",X"A1",X"4E",X"BD",X"D7",X"AE",X"C6",X"85",X"F7",
		X"A0",X"27",X"86",X"FE",X"8E",X"B2",X"60",X"BD",X"C1",X"38",X"24",X"02",X"86",X"FD",X"8E",X"CC",
		X"02",X"C6",X"FF",X"BD",X"FF",X"D4",X"C6",X"E4",X"BD",X"FF",X"D4",X"5A",X"26",X"FD",X"C6",X"FF",
		X"BD",X"FF",X"D4",X"1F",X"89",X"BD",X"C6",X"AA",X"CE",X"C0",X"ED",X"B6",X"A0",X"06",X"48",X"33",
		X"C6",X"8E",X"3E",X"38",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"CE",X"C0",X"FD",X"8E",X"14",X"58",
		X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"CC",X"41",X"2F",X"FD",X"A0",X"00",X"86",X"40",X"FD",X"A0",
		X"02",X"FD",X"A0",X"04",X"BD",X"C1",X"49",X"86",X"28",X"B7",X"A1",X"53",X"8E",X"C1",X"CD",X"86",
		X"00",X"BD",X"D0",X"56",X"8E",X"C1",X"D8",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"C1",X"EE",X"86",
		X"00",X"BD",X"D0",X"56",X"7F",X"A1",X"50",X"BD",X"C1",X"5C",X"4F",X"B7",X"A1",X"5C",X"B7",X"A1",
		X"5B",X"86",X"01",X"8E",X"C0",X"C9",X"7E",X"F5",X"82",X"B6",X"A0",X"58",X"85",X"01",X"26",X"14",
		X"7D",X"A1",X"53",X"27",X"29",X"7C",X"A1",X"5C",X"B6",X"A1",X"5C",X"81",X"05",X"26",X"E2",X"B7",
		X"A1",X"5B",X"20",X"DD",X"7F",X"A1",X"5C",X"7D",X"A1",X"5B",X"27",X"D5",X"86",X"14",X"B7",X"A1",
		X"53",X"7C",X"A1",X"50",X"BD",X"C1",X"5C",X"B6",X"A1",X"50",X"81",X"03",X"26",X"BC",X"BD",X"D0",
		X"7D",X"8E",X"B2",X"84",X"CE",X"B2",X"54",X"BD",X"C1",X"85",X"8E",X"C4",X"71",X"8D",X"29",X"24",
		X"09",X"8E",X"C4",X"65",X"CE",X"C4",X"11",X"BD",X"C1",X"85",X"10",X"8E",X"A1",X"D7",X"B6",X"A0",
		X"06",X"4C",X"81",X"03",X"10",X"26",X"FE",X"FE",X"7D",X"A1",X"4E",X"26",X"08",X"86",X"FF",X"8E",
		X"C1",X"35",X"7E",X"F5",X"82",X"7E",X"C2",X"59",X"34",X"16",X"BD",X"F8",X"2B",X"10",X"A3",X"21",
		X"26",X"05",X"BD",X"F8",X"15",X"A1",X"23",X"35",X"96",X"8E",X"46",X"AC",X"CC",X"14",X"08",X"BD",
		X"D1",X"9F",X"CE",X"C0",X"FF",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"39",X"7F",X"A1",X"3A",X"8E",
		X"45",X"B7",X"CE",X"11",X"11",X"B6",X"A1",X"3A",X"B1",X"A1",X"50",X"26",X"03",X"CE",X"DD",X"DD",
		X"CC",X"04",X"00",X"EF",X"8B",X"4A",X"26",X"FB",X"7C",X"A1",X"3A",X"30",X"89",X"08",X"00",X"8C",
		X"5D",X"B7",X"26",X"DE",X"39",X"FF",X"A1",X"3C",X"10",X"BE",X"A1",X"51",X"8D",X"AA",X"24",X"09",
		X"8D",X"24",X"30",X"14",X"BC",X"A1",X"3C",X"22",X"F3",X"30",X"0C",X"EC",X"21",X"BD",X"F8",X"57",
		X"A6",X"23",X"BD",X"F8",X"41",X"CE",X"A0",X"00",X"A6",X"C4",X"BD",X"F8",X"41",X"33",X"42",X"11",
		X"83",X"A0",X"06",X"26",X"F3",X"39",X"34",X"10",X"BD",X"F8",X"2B",X"30",X"08",X"BD",X"F8",X"57",
		X"30",X"88",X"E8",X"AC",X"E4",X"27",X"04",X"30",X"0C",X"20",X"ED",X"35",X"90",X"7A",X"A1",X"53",
		X"86",X"3C",X"8E",X"C1",X"CD",X"7E",X"F5",X"82",X"B6",X"A0",X"33",X"26",X"05",X"B6",X"A0",X"27",
		X"20",X"01",X"4F",X"B7",X"A0",X"33",X"86",X"0F",X"8E",X"C1",X"D8",X"7E",X"F5",X"82",X"7F",X"A1",
		X"4F",X"B6",X"A0",X"58",X"85",X"80",X"27",X"04",X"86",X"FF",X"20",X"10",X"B6",X"A0",X"5A",X"85",
		X"01",X"27",X"04",X"86",X"01",X"20",X"05",X"7F",X"A1",X"4F",X"20",X"34",X"B1",X"A1",X"4F",X"26",
		X"37",X"7A",X"A1",X"55",X"26",X"2A",X"8E",X"A0",X"00",X"F6",X"A1",X"50",X"58",X"3A",X"A6",X"84",
		X"BB",X"A1",X"4F",X"81",X"3F",X"26",X"02",X"86",X"5A",X"81",X"5B",X"26",X"02",X"86",X"40",X"A7",
		X"84",X"BD",X"C1",X"49",X"B6",X"A1",X"54",X"44",X"8B",X"05",X"B7",X"A1",X"54",X"B7",X"A1",X"55",
		X"86",X"01",X"8E",X"C1",X"F1",X"7E",X"F5",X"82",X"B7",X"A1",X"4F",X"86",X"37",X"B7",X"A1",X"54",
		X"86",X"03",X"B7",X"A1",X"55",X"20",X"E9",X"FF",X"FF",X"BD",X"D0",X"7D",X"BD",X"C8",X"53",X"BD",
		X"D7",X"8E",X"7F",X"A0",X"27",X"8E",X"C8",X"D8",X"86",X"00",X"BD",X"D0",X"56",X"12",X"12",X"12",
		X"7E",X"C2",X"90",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"CE",X"11",X"11",X"8E",
		X"1E",X"7B",X"CC",X"5F",X"00",X"EF",X"8B",X"81",X"41",X"26",X"02",X"86",X"1F",X"4A",X"2A",X"F5",
		X"86",X"2F",X"B7",X"A0",X"07",X"B7",X"A0",X"0B",X"B7",X"A0",X"12",X"CE",X"C1",X"03",X"8E",X"38",
		X"86",X"BF",X"A1",X"57",X"8E",X"B2",X"60",X"BF",X"A1",X"3C",X"8D",X"48",X"7E",X"C2",X"BA",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"86",X"3F",X"BD",X"C9",X"A9",X"10",
		X"8E",X"B3",X"00",X"CC",X"3C",X"18",X"ED",X"A4",X"CC",X"B4",X"12",X"ED",X"22",X"CC",X"30",X"38",
		X"BD",X"C9",X"B7",X"8E",X"E7",X"A9",X"86",X"00",X"BD",X"D0",X"56",X"86",X"3C",X"B7",X"A1",X"53",
		X"7D",X"A1",X"5A",X"26",X"0D",X"7A",X"A1",X"53",X"27",X"08",X"86",X"0A",X"8E",X"C2",X"E0",X"7E",
		X"F5",X"82",X"20",X"50",X"86",X"31",X"B7",X"A0",X"06",X"4F",X"10",X"8E",X"A0",X"0C",X"BE",X"A1",
		X"3C",X"BD",X"FF",X"D7",X"30",X"01",X"C4",X"0F",X"26",X"07",X"4D",X"26",X"04",X"C6",X"40",X"20",
		X"03",X"4C",X"CB",X"30",X"E7",X"A0",X"10",X"8C",X"A0",X"12",X"26",X"E5",X"BD",X"F8",X"2B",X"FD",
		X"A0",X"08",X"BD",X"F8",X"15",X"B7",X"A0",X"0A",X"BF",X"A1",X"3C",X"BE",X"A1",X"57",X"BD",X"FF",
		X"CE",X"C0",X"02",X"02",X"30",X"0A",X"BF",X"A1",X"57",X"7C",X"A0",X"06",X"B6",X"A0",X"06",X"81",
		X"36",X"26",X"B6",X"39",X"BD",X"F6",X"48",X"BD",X"C4",X"32",X"86",X"D9",X"B7",X"A0",X"92",X"BD",
		X"C9",X"1B",X"8E",X"C8",X"D8",X"86",X"00",X"BD",X"D0",X"56",X"BD",X"D7",X"4C",X"8E",X"CC",X"49",
		X"BF",X"A1",X"6C",X"8E",X"E7",X"A9",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"F5",X"28",X"86",X"00",
		X"BD",X"D0",X"56",X"8E",X"F5",X"01",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"EA",X"0A",X"86",X"00",
		X"BD",X"D0",X"56",X"8E",X"C6",X"4D",X"86",X"00",X"BD",X"D0",X"56",X"BD",X"D0",X"AE",X"7E",X"C5",
		X"48",X"ED",X"0E",X"ED",X"88",X"10",X"CC",X"1E",X"00",X"ED",X"0A",X"CC",X"DB",X"00",X"ED",X"0C",
		X"CC",X"F8",X"F4",X"ED",X"02",X"BF",X"A0",X"42",X"CC",X"66",X"66",X"ED",X"88",X"12",X"BF",X"A1",
		X"5F",X"CC",X"00",X"00",X"ED",X"0E",X"CC",X"00",X"00",X"ED",X"88",X"10",X"CC",X"04",X"00",X"ED",
		X"0A",X"CC",X"40",X"00",X"ED",X"0C",X"CC",X"F9",X"B4",X"ED",X"02",X"BF",X"A0",X"42",X"CC",X"00",
		X"00",X"ED",X"88",X"12",X"BF",X"A1",X"61",X"BD",X"D0",X"AE",X"7E",X"C5",X"48",X"ED",X"02",X"CC",
		X"1D",X"A0",X"ED",X"0A",X"CC",X"40",X"00",X"ED",X"0C",X"CC",X"00",X"A0",X"ED",X"88",X"10",X"CC",
		X"00",X"00",X"ED",X"0E",X"CC",X"44",X"33",X"ED",X"88",X"12",X"BD",X"FC",X"80",X"BF",X"A1",X"63",
		X"86",X"E6",X"8E",X"C4",X"08",X"7E",X"F5",X"82",X"CC",X"FF",X"50",X"BE",X"A1",X"63",X"ED",X"88",
		X"10",X"BE",X"A1",X"5F",X"ED",X"88",X"10",X"86",X"A0",X"8E",X"C4",X"1F",X"7E",X"F5",X"82",X"8E",
		X"C5",X"F1",X"86",X"00",X"BD",X"D0",X"56",X"BF",X"A1",X"5D",X"86",X"15",X"8E",X"C4",X"70",X"7E",
		X"F5",X"82",X"86",X"FF",X"B7",X"A0",X"92",X"BD",X"D8",X"C5",X"BD",X"D7",X"8E",X"CC",X"00",X"00",
		X"FD",X"A0",X"20",X"FD",X"A0",X"22",X"BD",X"FF",X"CE",X"F5",X"BE",X"00",X"BD",X"D8",X"B5",X"86",
		X"DB",X"B7",X"A0",X"92",X"8E",X"10",X"30",X"BF",X"A0",X"97",X"39",X"BE",X"A1",X"5D",X"FE",X"A1",
		X"6A",X"4F",X"A7",X"C4",X"33",X"C9",X"01",X"00",X"11",X"A3",X"07",X"23",X"F5",X"7E",X"D0",X"16",
		X"8D",X"E9",X"BE",X"A1",X"63",X"BD",X"D0",X"C8",X"BD",X"FC",X"83",X"BE",X"A1",X"61",X"CC",X"00",
		X"40",X"ED",X"0E",X"CC",X"00",X"D4",X"ED",X"88",X"10",X"86",X"2D",X"B7",X"A1",X"65",X"BE",X"A1",
		X"5F",X"CC",X"00",X"00",X"ED",X"88",X"10",X"BE",X"A1",X"5F",X"EC",X"88",X"10",X"C3",X"00",X"08",
		X"ED",X"88",X"10",X"7A",X"A1",X"65",X"27",X"08",X"86",X"02",X"8E",X"C4",X"97",X"7E",X"F5",X"82",
		X"BD",X"D0",X"AE",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",X"10",X"CC",X"1D",X"FF",X"ED",X"0A",
		X"CC",X"90",X"00",X"ED",X"0C",X"CC",X"F9",X"DA",X"ED",X"02",X"BF",X"A0",X"42",X"CC",X"00",X"00",
		X"ED",X"88",X"12",X"BF",X"A1",X"66",X"CC",X"00",X"00",X"CE",X"00",X"C0",X"BE",X"A1",X"61",X"ED",
		X"0E",X"EF",X"88",X"10",X"BE",X"A1",X"5F",X"CC",X"1E",X"80",X"ED",X"0A",X"CC",X"A2",X"E0",X"ED",
		X"0C",X"EF",X"88",X"10",X"86",X"50",X"8E",X"C4",X"FC",X"7E",X"F5",X"82",X"BE",X"A1",X"66",X"CC",
		X"E0",X"00",X"ED",X"0C",X"CC",X"1C",X"00",X"ED",X"0A",X"BE",X"A1",X"5F",X"CC",X"00",X"00",X"ED",
		X"88",X"10",X"BE",X"A1",X"61",X"CC",X"F9",X"BE",X"ED",X"02",X"CC",X"FF",X"C0",X"ED",X"0E",X"CC",
		X"FE",X"80",X"ED",X"88",X"10",X"86",X"60",X"8E",X"C5",X"2D",X"7E",X"F5",X"82",X"BE",X"A1",X"61",
		X"CC",X"F9",X"B4",X"ED",X"02",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",X"10",X"BE",X"A1",X"66",
		X"EC",X"04",X"BD",X"D0",X"C8",X"BD",X"D4",X"00",X"CE",X"FB",X"7E",X"8E",X"28",X"60",X"FF",X"A1",
		X"63",X"BF",X"A1",X"68",X"86",X"20",X"8E",X"C5",X"5C",X"7E",X"F5",X"82",X"FE",X"A1",X"63",X"BE",
		X"A1",X"68",X"1F",X"10",X"10",X"AE",X"C4",X"BD",X"D0",X"FA",X"86",X"20",X"8E",X"C5",X"72",X"7E",
		X"F5",X"82",X"FE",X"A1",X"63",X"BE",X"A1",X"68",X"30",X"89",X"18",X"00",X"33",X"4E",X"BD",X"F6",
		X"A7",X"86",X"20",X"8E",X"C5",X"89",X"7E",X"F5",X"82",X"FE",X"A1",X"63",X"BE",X"A1",X"68",X"30",
		X"89",X"3C",X"00",X"33",X"C8",X"1C",X"BD",X"F6",X"A7",X"FE",X"A1",X"63",X"BE",X"A1",X"68",X"30",
		X"88",X"10",X"33",X"42",X"11",X"83",X"FB",X"8C",X"26",X"A4",X"20",X"35",X"EC",X"C1",X"ED",X"0C",
		X"CC",X"00",X"00",X"ED",X"88",X"10",X"ED",X"0E",X"BD",X"FC",X"80",X"FF",X"A1",X"68",X"86",X"20",
		X"8E",X"C5",X"C6",X"7E",X"F5",X"82",X"BE",X"A1",X"6C",X"30",X"02",X"BF",X"A1",X"6C",X"86",X"20",
		X"8E",X"C5",X"D6",X"7E",X"F5",X"82",X"FE",X"A1",X"68",X"11",X"83",X"CC",X"6F",X"10",X"26",X"FF",
		X"6A",X"86",X"FF",X"8E",X"C5",X"E9",X"7E",X"F5",X"82",X"86",X"FF",X"8E",X"C6",X"75",X"7E",X"F5",
		X"82",X"BE",X"A1",X"61",X"AE",X"04",X"30",X"89",X"07",X"04",X"AF",X"47",X"AF",X"49",X"BF",X"A1",
		X"6A",X"86",X"04",X"AE",X"47",X"C6",X"11",X"E7",X"84",X"30",X"89",X"01",X"00",X"4A",X"26",X"F7",
		X"C6",X"99",X"E7",X"84",X"AF",X"47",X"10",X"BE",X"A0",X"7F",X"10",X"8C",X"A1",X"37",X"25",X"04",
		X"10",X"8E",X"A1",X"1A",X"AE",X"49",X"86",X"03",X"E6",X"A0",X"E7",X"84",X"30",X"89",X"01",X"00",
		X"4A",X"26",X"F5",X"10",X"BF",X"A0",X"7F",X"AF",X"49",X"BE",X"A1",X"6A",X"6F",X"84",X"30",X"89",
		X"01",X"00",X"BF",X"A1",X"6A",X"86",X"01",X"8E",X"C6",X"01",X"7E",X"F5",X"82",X"10",X"8E",X"CC",
		X"47",X"EE",X"A9",X"00",X"0E",X"AE",X"A1",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"10",X"BF",X"A1",
		X"6E",X"86",X"06",X"8E",X"C6",X"69",X"7E",X"F5",X"82",X"10",X"BE",X"A1",X"6E",X"10",X"BC",X"A1",
		X"6C",X"26",X"DE",X"20",X"D8",X"BD",X"D0",X"7D",X"7F",X"A1",X"5A",X"86",X"FB",X"B7",X"A0",X"92",
		X"BD",X"D7",X"8E",X"7F",X"B2",X"18",X"CC",X"FF",X"FF",X"FD",X"B2",X"1F",X"8E",X"E7",X"A9",X"86",
		X"00",X"BD",X"D0",X"56",X"8E",X"F5",X"01",X"86",X"00",X"BD",X"D0",X"56",X"86",X"3F",X"B7",X"A0",
		X"32",X"7E",X"C6",X"A4",X"BD",X"C8",X"53",X"7E",X"C7",X"2F",X"CC",X"D5",X"7C",X"BD",X"D5",X"ED",
		X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8E",
		X"C7",X"4B",X"86",X"00",X"BD",X"D0",X"56",X"8E",X"32",X"58",X"CE",X"C0",X"ED",X"BD",X"FF",X"CE",
		X"C0",X"02",X"02",X"86",X"05",X"8E",X"C7",X"37",X"BD",X"F5",X"82",X"BE",X"A1",X"95",X"A6",X"84",
		X"B1",X"A1",X"94",X"26",X"03",X"8E",X"C7",X"B7",X"86",X"30",X"7E",X"F5",X"82",X"A1",X"45",X"CC",
		X"00",X"00",X"FD",X"A0",X"20",X"CC",X"0C",X"00",X"FD",X"A1",X"47",X"CC",X"B3",X"04",X"FD",X"A1",
		X"49",X"BE",X"A1",X"49",X"10",X"BE",X"A1",X"43",X"CC",X"04",X"0C",X"ED",X"A4",X"FC",X"A1",X"45",
		X"ED",X"22",X"C3",X"00",X"60",X"FD",X"A1",X"45",X"10",X"AF",X"02",X"FC",X"A1",X"47",X"ED",X"0A",
		X"C3",X"01",X"00",X"FD",X"A1",X"47",X"CC",X"98",X"00",X"ED",X"0C",X"BD",X"FC",X"80",X"30",X"0E",
		X"BF",X"A1",X"49",X"31",X"24",X"10",X"BF",X"A1",X"43",X"10",X"8C",X"B4",X"12",X"26",X"C2",X"86",
		X"2E",X"8E",X"C7",X"B7",X"7E",X"F5",X"82",X"8E",X"B3",X"00",X"CC",X"3C",X"18",X"ED",X"84",X"CC",
		X"B4",X"12",X"ED",X"02",X"8E",X"C8",X"2C",X"86",X"00",X"BD",X"D0",X"56",X"86",X"28",X"8E",X"C7",
		X"D4",X"7E",X"F5",X"82",X"8E",X"F5",X"28",X"86",X"00",X"BD",X"D0",X"56",X"12",X"12",X"12",X"7E",
		X"C8",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8E",X"C8",X"D8",X"86",X"00",X"BD",X"D0",X"56",
		X"86",X"3C",X"B7",X"A1",X"53",X"7D",X"A1",X"5A",X"10",X"26",X"FB",X"28",X"7A",X"A1",X"53",X"27",
		X"08",X"86",X"0A",X"8E",X"C8",X"15",X"7E",X"F5",X"82",X"7E",X"C2",X"59",X"10",X"8E",X"B3",X"00",
		X"CC",X"30",X"90",X"BD",X"D0",X"FA",X"7D",X"9C",X"00",X"26",X"10",X"7D",X"9C",X"40",X"26",X"0B",
		X"8E",X"C9",X"06",X"86",X"00",X"BD",X"C9",X"BD",X"7E",X"D0",X"0B",X"86",X"01",X"8E",X"C8",X"2C",
		X"7E",X"F5",X"82",X"8E",X"B4",X"12",X"10",X"8E",X"CA",X"86",X"4F",X"B7",X"A1",X"4D",X"B7",X"A1",
		X"4C",X"A6",X"A4",X"44",X"44",X"44",X"44",X"8D",X"0C",X"A6",X"A0",X"84",X"0F",X"8D",X"06",X"10",
		X"8C",X"CB",X"A8",X"26",X"EC",X"85",X"0C",X"26",X"09",X"BB",X"A1",X"4C",X"48",X"48",X"B7",X"A1",
		X"4C",X"39",X"34",X"02",X"84",X"03",X"BB",X"A1",X"4C",X"B7",X"A1",X"4C",X"35",X"02",X"84",X"0C",
		X"44",X"44",X"CE",X"CB",X"A7",X"E6",X"C6",X"F7",X"A1",X"4B",X"8C",X"B9",X"B2",X"25",X"04",X"30",
		X"89",X"FA",X"61",X"B6",X"A1",X"4D",X"27",X"14",X"A6",X"84",X"84",X"F0",X"A7",X"84",X"B6",X"A1",
		X"4B",X"84",X"0F",X"AA",X"84",X"A7",X"84",X"B6",X"A1",X"4B",X"20",X"0D",X"73",X"A1",X"4D",X"B6",
		X"A1",X"4B",X"A7",X"84",X"7A",X"A1",X"4C",X"2B",X"0B",X"30",X"88",X"18",X"7A",X"A1",X"4C",X"2A",
		X"F1",X"7F",X"A1",X"4D",X"7F",X"A1",X"4C",X"39",X"F6",X"A0",X"37",X"27",X"21",X"F1",X"A1",X"59",
		X"23",X"06",X"F7",X"A1",X"59",X"7C",X"A1",X"5A",X"CE",X"C0",X"E9",X"8E",X"28",X"E5",X"BD",X"FF",
		X"CE",X"C0",X"02",X"02",X"4F",X"8E",X"48",X"E5",X"BD",X"FF",X"CE",X"C0",X"0E",X"02",X"86",X"10",
		X"8E",X"C8",X"D8",X"7E",X"F5",X"82",X"86",X"FF",X"B7",X"A1",X"40",X"86",X"02",X"8E",X"C9",X"13",
		X"7E",X"F5",X"82",X"86",X"0A",X"B7",X"A1",X"40",X"7E",X"D0",X"0B",X"B6",X"A0",X"69",X"27",X"06",
		X"BD",X"D4",X"8B",X"4A",X"20",X"F8",X"39",X"BD",X"C9",X"8F",X"CC",X"08",X"06",X"34",X"02",X"86",
		X"66",X"A7",X"1E",X"A7",X"1F",X"A7",X"84",X"30",X"89",X"01",X"00",X"6F",X"1E",X"6F",X"1F",X"5A",
		X"26",X"F3",X"C6",X"06",X"6A",X"E4",X"26",X"E9",X"A7",X"1E",X"A7",X"1F",X"A7",X"84",X"35",X"02",
		X"9E",X"6A",X"A6",X"08",X"1F",X"89",X"81",X"50",X"23",X"04",X"80",X"50",X"20",X"F8",X"4A",X"44",
		X"44",X"44",X"8E",X"C9",X"9F",X"A6",X"86",X"5A",X"C4",X"07",X"5C",X"34",X"04",X"BD",X"C9",X"8F",
		X"30",X"89",X"01",X"00",X"C6",X"05",X"6D",X"E4",X"27",X"13",X"A7",X"1E",X"A7",X"1F",X"30",X"89",
		X"01",X"00",X"5A",X"26",X"F5",X"30",X"89",X"01",X"00",X"6A",X"E4",X"20",X"E7",X"35",X"82",X"34",
		X"02",X"8E",X"08",X"29",X"96",X"68",X"81",X"01",X"27",X"03",X"8E",X"66",X"29",X"35",X"82",X"22",
		X"44",X"88",X"55",X"33",X"FF",X"EE",X"AA",X"DD",X"CC",X"B7",X"A0",X"32",X"86",X"81",X"97",X"33",
		X"97",X"34",X"86",X"2F",X"97",X"35",X"39",X"BD",X"D0",X"FA",X"8D",X"07",X"39",X"8D",X"04",X"BD",
		X"D0",X"56",X"39",X"34",X"36",X"10",X"8E",X"FB",X"7E",X"8E",X"10",X"20",X"34",X"30",X"10",X"AE",
		X"A4",X"1F",X"10",X"BD",X"D0",X"FA",X"35",X"30",X"34",X"30",X"10",X"AE",X"A4",X"30",X"89",X"00",
		X"B0",X"1F",X"10",X"BD",X"D0",X"FA",X"35",X"30",X"31",X"22",X"10",X"8C",X"FB",X"8C",X"25",X"04",
		X"10",X"8E",X"FB",X"7E",X"30",X"89",X"08",X"00",X"8C",X"90",X"20",X"23",X"CF",X"10",X"8E",X"FB",
		X"80",X"8E",X"10",X"30",X"34",X"30",X"10",X"AE",X"A4",X"1F",X"10",X"BD",X"D0",X"FA",X"35",X"30",
		X"34",X"30",X"10",X"AE",X"A4",X"30",X"89",X"80",X"00",X"1F",X"10",X"BD",X"D0",X"FA",X"35",X"30",
		X"31",X"22",X"10",X"8C",X"FB",X"8C",X"25",X"04",X"10",X"8E",X"FB",X"7E",X"30",X"88",X"10",X"8C",
		X"10",X"C0",X"23",X"D0",X"35",X"B6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"8E",X"CB",X"AB",X"8E",X"3B",X"38",X"86",X"02",X"34",X"02",X"EC",X"A1",X"FD",X"A1",X"3C",
		X"86",X"01",X"5F",X"B5",X"A1",X"3C",X"27",X"02",X"C6",X"10",X"B5",X"A1",X"3D",X"27",X"02",X"CA",
		X"01",X"E7",X"80",X"48",X"26",X"EC",X"6A",X"E4",X"26",X"E1",X"35",X"02",X"30",X"89",X"00",X"F0",
		X"10",X"8C",X"CC",X"43",X"26",X"D1",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"13",X"1F",X"20",X"E1",X"6D",X"16",X"D2",X"4F",X"24",X"D1",
		X"72",X"0E",X"13",X"C3",X"4C",X"24",X"C2",X"5E",X"12",X"61",X"2E",X"11",X"E2",X"24",X"D2",X"04",
		X"11",X"C1",X"0D",X"11",X"14",X"10",X"C3",X"C1",X"13",X"53",X"C2",X"E1",X"A7",X"1A",X"15",X"18",
		X"5B",X"14",X"B5",X"29",X"17",X"18",X"51",X"87",X"18",X"41",X"85",X"18",X"2E",X"2E",X"1A",X"71",
		X"A1",X"51",X"94",X"18",X"61",X"85",X"2A",X"15",X"19",X"6B",X"7B",X"51",X"85",X"18",X"2E",X"2E",
		X"1A",X"71",X"A1",X"41",X"A5",X"18",X"41",X"86",X"2B",X"14",X"1A",X"6B",X"5B",X"61",X"85",X"18",
		X"2E",X"2E",X"1A",X"71",X"A1",X"41",X"B4",X"18",X"41",X"85",X"CB",X"14",X"B6",X"1B",X"7A",X"5A",
		X"71",X"85",X"18",X"2E",X"2E",X"1B",X"51",X"B7",X"B4",X"B5",X"28",X"5D",X"B1",X"4B",X"62",X"86",
		X"1B",X"71",X"85",X"18",X"2E",X"2E",X"B4",X"A5",X"A4",X"B7",X"A6",X"B5",X"1B",X"4E",X"B1",X"4B",
		X"51",X"84",X"B7",X"19",X"14",X"18",X"51",X"82",X"E2",X"EB",X"4A",X"5A",X"4B",X"6B",X"6B",X"61",
		X"94",X"FB",X"14",X"B5",X"B6",X"B6",X"19",X"14",X"18",X"51",X"82",X"E2",X"EB",X"4A",X"5A",X"4B",
		X"62",X"B6",X"B5",X"FB",X"14",X"B4",X"18",X"6B",X"7B",X"16",X"A7",X"A2",X"F2",X"EB",X"41",X"B4",
		X"B5",X"38",X"6B",X"41",X"C2",X"BD",X"38",X"6B",X"16",X"A7",X"A2",X"F2",X"EB",X"51",X"95",X"B5",
		X"39",X"5B",X"41",X"C2",X"AD",X"39",X"6B",X"16",X"A7",X"A2",X"F2",X"EB",X"51",X"95",X"B4",X"18",
		X"5E",X"18",X"5B",X"1D",X"29",X"E1",X"81",X"C1",X"85",X"B1",X"6A",X"7A",X"2F",X"2E",X"B5",X"19",
		X"5B",X"41",X"84",X"FA",X"13",X"CA",X"1C",X"18",X"5B",X"C3",X"63",X"C2",X"EB",X"6B",X"6B",X"49",
		X"30",X"E9",X"5B",X"D7",X"18",X"51",X"82",X"E2",X"EB",X"6B",X"69",X"33",X"D9",X"E6",X"18",X"51",
		X"82",X"E2",X"EB",X"6B",X"10",X"2E",X"18",X"D1",X"82",X"E2",X"EB",X"51",X"10",X"DA",X"D1",X"82",
		X"E2",X"EA",X"11",X"2F",X"A2",X"E1",X"31",X"F0",X"22",X"EE",X"00",X"FC",X"FE",X"01",X"03",X"FF",
		X"01",X"07",X"04",X"42",X"CF",X"02",X"07",X"40",X"00",X"00",X"00",X"FF",X"FF",X"07",X"07",X"FF",
		X"21",X"07",X"00",X"21",X"21",X"00",X"00",X"FF",X"00",X"07",X"00",X"FF",X"FF",X"07",X"07",X"FF",
		X"06",X"07",X"00",X"38",X"06",X"00",X"00",X"FF",X"00",X"07",X"00",X"FF",X"FF",X"07",X"07",X"FF",
		X"21",X"07",X"04",X"F9",X"03",X"04",X"06",X"8F",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"07",X"07",X"FF",X"21",X"07",X"00",X"21",X"21",X"00",X"00",X"1E",X"00",X"00",X"00",X"FF",
		X"FF",X"07",X"07",X"FF",X"00",X"07",X"04",X"00",X"00",X"04",X"06",X"80",X"00",X"07",X"00",X"FF",
		X"FF",X"07",X"07",X"FF",X"21",X"07",X"00",X"21",X"21",X"00",X"00",X"FF",X"00",X"07",X"00",X"FF",
		X"FF",X"07",X"07",X"FF",X"06",X"07",X"00",X"38",X"C0",X"00",X"01",X"FF",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"04",X"01",X"02",X"F2",X"FA",X"04",X"05",X"0A",X"92",X"05",X"04",X"04",
		X"F8",X"02",X"01",X"FF",X"FF",X"FF",X"FF",X"43",X"30",X"1C",X"70",X"3C",X"70",X"5F",X"70",X"1C",
		X"A8",X"40",X"A8",X"5C",X"A8",X"C0",X"EB",X"C0",X"DD",X"C0",X"DF",X"C0",X"E7",X"C0",X"E3",X"C0",
		X"E1",X"C0",X"E5",X"60",X"00",X"60",X"00",X"62",X"00",X"98",X"00",X"98",X"00",X"9A",X"00",X"F9",
		X"78",X"F8",X"C1",X"F9",X"96",X"F9",X"1C",X"F8",X"EA",X"F9",X"6E",X"09",X"00",X"11",X"00",X"19",
		X"80",X"09",X"60",X"11",X"60",X"19",X"E0",X"33",X"22",X"CC",X"55",X"22",X"22",X"55",X"55",X"CC",
		X"CC",X"88",X"88",X"FF",X"FF",X"CC",X"0C",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"00",
		X"A0",X"0A",X"A0",X"A0",X"00",X"A0",X"0A",X"00",X"0A",X"0A",X"A0",X"0A",X"0A",X"AA",X"0A",X"00",
		X"A0",X"00",X"00",X"0A",X"00",X"A0",X"AA",X"A0",X"00",X"02",X"23",X"02",X"20",X"22",X"23",X"22",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"02",X"22",X"32",X"22",X"00",X"20",X"32",X"20",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"04",X"34",X"30",X"30",X"34",X"30",X"00",X"00",
		X"44",X"44",X"33",X"33",X"34",X"30",X"30",X"30",X"00",X"30",X"03",X"03",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"33",X"33",X"03",X"03",X"30",X"00",X"44",X"44",X"03",X"03",X"43",X"03",X"03",X"03",
		X"40",X"43",X"30",X"30",X"43",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"04",X"34",X"03",X"03",X"34",X"30",X"00",X"00",
		X"44",X"44",X"30",X"30",X"34",X"30",X"30",X"30",X"00",X"30",X"33",X"33",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"30",X"30",X"03",X"03",X"30",X"00",X"44",X"44",X"33",X"33",X"43",X"03",X"03",X"03",
		X"40",X"43",X"03",X"03",X"43",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"00",X"33",X"33",X"33",X"33",X"30",X"00",X"00",
		X"00",X"33",X"03",X"03",X"33",X"30",X"30",X"30",X"00",X"30",X"33",X"33",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"33",X"33",X"03",X"03",X"30",X"00",X"00",X"33",X"30",X"30",X"03",X"03",X"03",X"03",
		X"00",X"33",X"33",X"33",X"33",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"03",X"34",X"03",X"33",X"70",X"40",X"33",X"33",X"07",X"44",X"33",X"33",X"00",X"04",X"33",
		X"30",X"73",X"40",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"37",X"44",X"33",
		X"33",X"00",X"04",X"33",X"33",X"70",X"40",X"33",X"33",X"07",X"44",X"33",X"00",X"30",X"03",X"30",
		X"00",X"03",X"30",X"03",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"33",X"07",X"40",X"33",
		X"30",X"03",X"44",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"04",X"33",
		X"33",X"07",X"40",X"33",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"00",X"30",X"43",X"30",
		X"00",X"03",X"34",X"03",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"33",X"70",X"44",X"33",
		X"30",X"03",X"04",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"40",X"33",
		X"33",X"70",X"44",X"33",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"00",X"30",X"43",X"30",
		X"00",X"06",X"26",X"06",X"26",X"00",X"66",X"66",X"66",X"88",X"88",X"88",X"00",X"60",X"66",X"66",
		X"88",X"86",X"00",X"00",X"00",X"66",X"66",X"93",X"00",X"00",X"00",X"6D",X"66",X"00",X"00",X"00",
		X"00",X"EF",X"66",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"06",X"66",X"66",X"28",X"68",X"08",X"60",X"66",X"66",X"86",
		X"88",X"88",X"00",X"00",X"60",X"66",X"86",X"69",X"00",X"00",X"00",X"66",X"66",X"30",X"00",X"00",
		X"00",X"DE",X"66",X"00",X"00",X"00",X"00",X"F0",X"66",X"00",X"00",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"0F",X"66",X"00",X"00",X"00",X"00",X"ED",
		X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"03",X"00",X"00",X"06",X"66",X"68",X"96",X"06",X"66",
		X"66",X"68",X"88",X"88",X"60",X"66",X"66",X"83",X"86",X"80",X"00",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"00",X"FE",
		X"66",X"00",X"00",X"00",X"00",X"D6",X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"39",X"00",X"06",
		X"66",X"66",X"88",X"68",X"66",X"66",X"66",X"88",X"88",X"88",X"00",X"60",X"63",X"30",X"63",X"00",
		X"06",X"26",X"68",X"28",X"60",X"66",X"66",X"86",X"00",X"00",X"66",X"66",X"00",X"00",X"ED",X"66",
		X"00",X"00",X"00",X"63",X"90",X"09",X"90",X"99",X"99",X"99",X"90",X"CC",X"90",X"11",X"00",X"11",
		X"10",X"11",X"00",X"10",X"10",X"10",X"00",X"10",X"00",X"11",X"10",X"11",X"00",X"11",X"00",X"10",
		X"00",X"10",X"10",X"10",X"00",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"10",
		X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"11",X"01",X"11",X"00",X"11",X"00",X"01",X"01",X"01",
		X"00",X"01",X"00",X"11",X"00",X"11",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"01",X"01",X"01",X"11",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"F0",
		X"00",X"EE",X"E0",X"E0",X"E0",X"EE",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"DD",X"D0",X"D0",
		X"D0",X"DD",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"00",X"FF",
		X"00",X"FF",X"0F",X"FF",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"0E",X"EE",
		X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"DD",X"0D",X"0D",X"0D",X"DD",X"00",X"1C",X"0D",X"7F",
		X"E7",X"70",X"00",X"0F",X"71",X"71",X"07",X"DC",X"77",X"7C",X"0D",X"71",X"C7",X"77",X"DE",X"07",
		X"71",X"17",X"17",X"DE",X"F7",X"71",X"17",X"71",X"7C",X"DE",X"F0",X"07",X"77",X"C7",X"71",X"17",
		X"70",X"70",X"7C",X"D7",X"77",X"77",X"70",X"01",X"CD",X"FF",X"D7",X"70",X"F0",X"00",X"00",X"00",
		X"C6",X"27",X"7E",X"CA",X"D4",X"7E",X"CA",X"DF",X"7E",X"CA",X"EA",X"7E",X"CA",X"F5",X"7E",X"CB",
		X"FC",X"7E",X"CC",X"07",X"7E",X"CC",X"12",X"7E",X"CC",X"1D",X"7E",X"CA",X"9D",X"7E",X"CA",X"A5",
		X"7E",X"CA",X"75",X"7E",X"CA",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"C0",X"BD",X"C0",X"BF",X"C0",X"C1",X"00",X"00",X"C0",X"C1",X"00",X"00",X"C0",X"C3",X"00",
		X"00",X"C0",X"C5",X"00",X"00",X"C0",X"C5",X"00",X"00",X"C0",X"C7",X"00",X"00",X"C0",X"C3",X"00",
		X"00",X"C0",X"C9",X"00",X"00",X"C0",X"CB",X"C0",X"CD",X"C0",X"CF",X"00",X"00",X"C0",X"BD",X"C0",
		X"D1",X"C0",X"D3",X"C0",X"D5",X"C0",X"DB",X"00",X"00",X"C1",X"07",X"C1",X"0D",X"C1",X"11",X"C1",
		X"13",X"C1",X"15",X"C1",X"19",X"C1",X"1D",X"C1",X"21",X"C1",X"27",X"C1",X"2B",X"C1",X"33",X"C1",
		X"4D",X"C1",X"53",X"C1",X"6D",X"C1",X"88",X"C1",X"92",X"C1",X"96",X"C1",X"9C",X"C1",X"A0",X"C1",
		X"A2",X"C1",X"A6",X"C1",X"A8",X"C1",X"AC",X"C1",X"B0",X"C1",X"B2",X"C1",X"B4",X"C1",X"B6",X"C1",
		X"B8",X"C1",X"BC",X"C1",X"BE",X"C1",X"C2",X"C1",X"C6",X"C1",X"C8",X"C1",X"CA",X"C1",X"CC",X"C1",
		X"CE",X"C1",X"D0",X"C1",X"D2",X"C1",X"D4",X"C1",X"D6",X"C1",X"D8",X"C1",X"DA",X"C1",X"EA",X"C1",
		X"F8",X"C2",X"00",X"C2",X"08",X"C2",X"10",X"C2",X"1A",X"C2",X"24",X"C2",X"2C",X"C2",X"34",X"C2",
		X"3E",X"C2",X"48",X"C2",X"52",X"C2",X"5A",X"C2",X"64",X"C2",X"68",X"C2",X"74",X"C2",X"7E",X"C2",
		X"85",X"C2",X"8C",X"C2",X"93",X"C2",X"9A",X"C2",X"A1",X"C2",X"A8",X"C2",X"AA",X"C2",X"AC",X"C2",
		X"B4",X"C2",X"B8",X"C2",X"BC",X"C2",X"BE",X"C2",X"C6",X"C2",X"D2",X"C2",X"D6",X"C2",X"D8",X"C3",
		X"01",X"C3",X"0B",X"C3",X"21",X"C3",X"2B",X"C4",X"64",X"C5",X"91",X"C4",X"50",X"C5",X"BF",X"C4",
		X"D5",X"C5",X"31",X"C5",X"1F",X"C5",X"31",X"C4",X"04",X"C5",X"1F",X"C4",X"04",X"C4",X"15",X"C4",
		X"E4",X"C3",X"3E",X"C5",X"35",X"C4",X"D5",X"C5",X"1F",X"C5",X"85",X"C4",X"CE",X"C5",X"1F",X"C3",
		X"F8",X"C3",X"C6",X"C3",X"93",X"C5",X"1F",X"C4",X"04",X"06",X"28",X"A0",X"C5",X"85",X"C4",X"AD",
		X"C3",X"66",X"C3",X"F0",X"07",X"C5",X"DE",X"C3",X"98",X"C3",X"CF",X"C4",X"DC",X"C3",X"93",X"C5",
		X"1F",X"C4",X"D5",X"C4",X"A4",X"C5",X"1F",X"C4",X"04",X"03",X"FE",X"C3",X"81",X"04",X"10",X"02",
		X"F8",X"C3",X"93",X"C5",X"1F",X"C3",X"7D",X"C4",X"D1",X"C3",X"66",X"C5",X"8A",X"C3",X"9D",X"C5",
		X"1F",X"C5",X"85",X"04",X"30",X"02",X"E8",X"C5",X"C7",X"C3",X"9D",X"C3",X"61",X"C4",X"50",X"07",
		X"03",X"FC",X"C3",X"9D",X"C5",X"1F",X"C4",X"04",X"C3",X"49",X"C5",X"85",X"07",X"07",X"03",X"04",
		X"C5",X"58",X"C5",X"7E",X"C5",X"85",X"C4",X"9C",X"C5",X"85",X"C4",X"E9",X"C3",X"55",X"C5",X"C4",
		X"C3",X"36",X"C5",X"2B",X"C3",X"98",X"C4",X"35",X"C4",X"8B",X"C3",X"98",X"C3",X"85",X"C3",X"98",
		X"C4",X"75",X"C4",X"75",X"C4",X"0C",X"C5",X"A0",X"C5",X"52",X"C3",X"69",X"C4",X"45",X"C5",X"BB",
		X"C4",X"F9",X"C4",X"D8",X"C4",X"F2",X"C5",X"23",X"C3",X"D4",X"C5",X"C4",X"C5",X"D5",X"C4",X"75",
		X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C5",X"0F",X"C3",X"36",X"C5",X"DE",
		X"C5",X"7E",X"C5",X"49",X"C4",X"11",X"03",X"FE",X"C3",X"83",X"C3",X"55",X"C4",X"11",X"C3",X"4F",
		X"03",X"FE",X"C3",X"81",X"C4",X"15",X"C3",X"2B",X"C4",X"95",X"C4",X"11",X"C5",X"31",X"C5",X"85",
		X"C3",X"55",X"C4",X"11",X"C5",X"1F",X"C5",X"85",X"C3",X"55",X"C5",X"B1",X"C3",X"FF",X"C5",X"85",
		X"C3",X"55",X"C4",X"11",X"C3",X"93",X"C5",X"1F",X"C5",X"85",X"C3",X"55",X"C4",X"11",X"C3",X"9D",
		X"C5",X"1F",X"C5",X"85",X"C3",X"55",X"C4",X"11",X"C3",X"49",X"C5",X"85",X"C3",X"55",X"C4",X"11",
		X"C5",X"7E",X"C5",X"85",X"C4",X"95",X"C5",X"B1",X"C5",X"85",X"C4",X"59",X"C5",X"5E",X"C3",X"55",
		X"C4",X"11",X"C4",X"9C",X"C5",X"85",X"C4",X"E9",X"C4",X"95",X"C5",X"B1",X"C5",X"6B",X"C5",X"9B",
		X"C4",X"E9",X"C3",X"55",X"C4",X"11",X"C4",X"15",X"C4",X"E4",X"C4",X"95",X"C5",X"B1",X"C5",X"6B",
		X"C5",X"9B",X"C3",X"2B",X"C5",X"D5",X"C3",X"BD",X"C5",X"0F",X"C3",X"36",X"C5",X"B1",X"C5",X"6B",
		X"C5",X"9B",X"C5",X"85",X"C5",X"0F",X"C4",X"35",X"C5",X"B1",X"C4",X"90",X"C3",X"8C",X"C4",X"84",
		X"07",X"03",X"06",X"C4",X"B9",X"C4",X"B2",X"07",X"03",X"06",X"C4",X"BD",X"C5",X"01",X"07",X"03",
		X"00",X"C4",X"C9",X"C3",X"6E",X"07",X"03",X"06",X"C4",X"C5",X"C5",X"76",X"07",X"03",X"08",X"C4",
		X"BD",X"C3",X"5A",X"07",X"03",X"06",X"C4",X"C1",X"C3",X"B4",X"C5",X"3A",X"C3",X"D9",X"07",X"07",
		X"03",X"0C",X"C5",X"06",X"C4",X"F2",X"C4",X"D8",X"C4",X"F2",X"C5",X"BB",X"C3",X"75",X"C5",X"0F",
		X"C4",X"D8",X"C4",X"F2",X"C5",X"65",X"C5",X"0F",X"C4",X"D8",X"C4",X"E1",X"C5",X"BB",X"C4",X"F2",
		X"C5",X"65",X"C3",X"A3",X"C3",X"42",X"C3",X"42",X"C5",X"E3",X"C4",X"30",X"C5",X"15",X"C4",X"11",
		X"07",X"C5",X"97",X"C3",X"BD",X"C4",X"23",X"07",X"07",X"C5",X"42",X"C4",X"6C",X"C5",X"DE",X"C5",
		X"C4",X"C3",X"D4",X"C5",X"70",X"07",X"07",X"C5",X"0F",X"C4",X"0C",X"C5",X"B1",X"C3",X"EA",X"C4",
		X"64",X"A0",X"00",X"02",X"08",X"A0",X"02",X"02",X"10",X"A0",X"04",X"C4",X"1A",X"06",X"22",X"70",
		X"C5",X"B4",X"02",X"3E",X"C3",X"3E",X"C5",X"AC",X"07",X"03",X"FC",X"C4",X"1A",X"02",X"3D",X"C4",
		X"1A",X"A0",X"06",X"02",X"05",X"A0",X"08",X"02",X"13",X"A0",X"0C",X"41",X"44",X"4A",X"55",X"53",
		X"54",X"4D",X"45",X"4E",X"54",X"2F",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"2F",X"41",X"4C",
		X"4C",X"2F",X"20",X"20",X"20",X"20",X"20",X"20",X"2F",X"41",X"55",X"44",X"49",X"4F",X"2F",X"41",
		X"55",X"44",X"49",X"54",X"2F",X"41",X"55",X"54",X"4F",X"2F",X"50",X"52",X"4F",X"42",X"45",X"52",
		X"2F",X"42",X"41",X"52",X"53",X"2F",X"42",X"45",X"2F",X"42",X"4F",X"4D",X"42",X"2F",X"43",X"41",
		X"4E",X"4E",X"4F",X"4E",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"20",X"58",X"2F",X"43",X"41",X"4E",
		X"2F",X"2C",X"2F",X"3A",X"2F",X"43",X"45",X"4E",X"54",X"45",X"52",X"2F",X"43",X"48",X"41",X"4E",
		X"47",X"45",X"2F",X"43",X"4D",X"4F",X"53",X"2F",X"43",X"4F",X"49",X"4E",X"2F",X"43",X"4F",X"4C",
		X"4F",X"52",X"2F",X"20",X"20",X"4D",X"49",X"53",X"53",X"49",X"4F",X"4E",X"2F",X"43",X"52",X"45",
		X"44",X"49",X"54",X"2F",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"3A",X"2F",X"20",X"4D",X"41",
		X"59",X"44",X"41",X"59",X"20",X"2F",X"44",X"45",X"54",X"45",X"43",X"54",X"45",X"44",X"2F",X"44",
		X"4F",X"4F",X"52",X"2F",X"44",X"4F",X"57",X"4E",X"2F",X"4D",X"41",X"59",X"44",X"41",X"59",X"20",
		X"4D",X"2C",X"41",X"49",X"44",X"45",X"5A",X"2F",X"2F",X"2F",X"45",X"4E",X"54",X"45",X"52",X"2F",
		X"45",X"4E",X"54",X"45",X"52",X"45",X"44",X"2F",X"45",X"52",X"52",X"4F",X"52",X"53",X"2F",X"45",
		X"58",X"49",X"54",X"2F",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",X"2F",X"46",X"49",X"52",X"45",
		X"2F",X"46",X"4F",X"52",X"2F",X"47",X"41",X"4D",X"45",X"2F",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"2F",X"48",X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",X"41",X"4D",X"45",X"2F",
		X"48",X"41",X"56",X"45",X"2F",X"48",X"49",X"47",X"48",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",
		X"45",X"53",X"45",X"54",X"2F",X"48",X"59",X"50",X"45",X"52",X"53",X"50",X"41",X"43",X"45",X"2F",
		X"49",X"4E",X"44",X"49",X"43",X"41",X"54",X"45",X"2F",X"49",X"4E",X"44",X"49",X"56",X"49",X"44",
		X"55",X"41",X"4C",X"2F",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"2F",X"49",X"4E",X"49",X"54",
		X"49",X"41",X"4C",X"53",X"2F",X"49",X"4E",X"56",X"41",X"4C",X"49",X"44",X"20",X"53",X"57",X"49",
		X"54",X"43",X"48",X"2F",X"52",X"4F",X"43",X"4B",X"45",X"54",X"2F",X"4C",X"45",X"46",X"54",X"2F",
		X"4D",X"41",X"4B",X"45",X"2F",X"4D",X"41",X"4E",X"55",X"41",X"4C",X"2F",X"4D",X"4F",X"4E",X"49",
		X"54",X"4F",X"52",X"2F",X"4D",X"55",X"4C",X"54",X"49",X"50",X"4C",X"45",X"2F",X"4D",X"55",X"53",
		X"54",X"2F",X"4C",X"41",X"53",X"45",X"52",X"20",X"2F",X"31",X"30",X"30",X"2F",X"31",X"35",X"30",
		X"2F",X"32",X"30",X"30",X"2F",X"32",X"35",X"30",X"2F",X"31",X"30",X"30",X"30",X"2F",X"4E",X"4F",
		X"2F",X"4E",X"4F",X"54",X"2F",X"4F",X"4B",X"2F",X"4F",X"4E",X"45",X"2F",X"4F",X"50",X"45",X"4E",
		X"2F",X"4F",X"52",X"2F",X"4F",X"56",X"45",X"52",X"2F",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",
		X"53",X"2F",X"50",X"4C",X"41",X"59",X"45",X"52",X"2F",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",
		X"2F",X"4D",X"49",X"4E",X"45",X"2F",X"2F",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"2F",X"50",
		X"52",X"45",X"53",X"53",X"2F",X"51",X"55",X"41",X"4C",X"49",X"46",X"49",X"45",X"44",X"2F",X"52",
		X"41",X"4D",X"2F",X"52",X"45",X"56",X"45",X"52",X"53",X"45",X"2F",X"52",X"49",X"47",X"48",X"54",
		X"2F",X"52",X"4F",X"4D",X"2F",X"52",X"4F",X"4D",X"53",X"2F",X"20",X"52",X"41",X"44",X"41",X"52",
		X"20",X"2F",X"53",X"45",X"4C",X"45",X"43",X"54",X"2F",X"53",X"45",X"54",X"2F",X"53",X"4C",X"41",
		X"4D",X"2F",X"53",X"4D",X"41",X"52",X"54",X"2F",X"53",X"4F",X"55",X"4E",X"44",X"2F",X"53",X"4F",
		X"55",X"4E",X"44",X"53",X"2F",X"53",X"54",X"41",X"52",X"54",X"2F",X"53",X"54",X"45",X"50",X"2F",
		X"53",X"54",X"49",X"43",X"4B",X"2F",X"52",X"41",X"4D",X"4D",X"45",X"52",X"20",X"2F",X"53",X"57",
		X"49",X"54",X"43",X"48",X"2F",X"54",X"45",X"53",X"54",X"2F",X"54",X"45",X"53",X"54",X"45",X"44",
		X"2F",X"54",X"45",X"53",X"54",X"53",X"2F",X"54",X"48",X"45",X"2F",X"54",X"48",X"52",X"55",X"2F",
		X"54",X"48",X"52",X"55",X"53",X"54",X"2F",X"54",X"49",X"4C",X"54",X"2F",X"54",X"49",X"4D",X"45",
		X"2F",X"54",X"4F",X"2F",X"54",X"4F",X"44",X"41",X"59",X"53",X"2F",X"54",X"57",X"4F",X"2F",X"55",
		X"4E",X"49",X"54",X"2F",X"55",X"50",X"2F",X"56",X"45",X"52",X"54",X"49",X"43",X"41",X"4C",X"2F",
		X"20",X"20",X"20",X"20",X"2F",X"4D",X"41",X"59",X"44",X"41",X"59",X"2F",X"40",X"40",X"57",X"49",
		X"54",X"48",X"2F",X"59",X"4F",X"55",X"2F",X"01",X"08",X"C5",X"EF",X"01",X"08",X"C6",X"D3",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",X"C6",X"DB",X"00",X"00",X"00",X"00",X"01",
		X"08",X"C6",X"E3",X"00",X"00",X"00",X"00",X"03",X"08",X"C6",X"EB",X"03",X"08",X"C7",X"03",X"03",
		X"08",X"C7",X"1B",X"03",X"08",X"C7",X"33",X"03",X"08",X"C7",X"4B",X"03",X"08",X"C7",X"63",X"03",
		X"08",X"C7",X"7B",X"03",X"08",X"C7",X"93",X"03",X"08",X"C7",X"AB",X"03",X"08",X"C7",X"C3",X"01",
		X"08",X"C7",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"08",X"C7",X"E3",X"03",X"08",X"C5",X"EF",X"03",X"08",X"C7",X"FB",X"03",
		X"08",X"C8",X"13",X"03",X"08",X"C8",X"2B",X"03",X"08",X"C8",X"43",X"03",X"08",X"C8",X"5B",X"03",
		X"08",X"C8",X"73",X"03",X"08",X"C8",X"8B",X"03",X"08",X"C8",X"A3",X"02",X"08",X"C8",X"BB",X"03",
		X"08",X"C8",X"CB",X"03",X"08",X"C8",X"E3",X"03",X"08",X"C8",X"FB",X"04",X"08",X"C9",X"13",X"03",
		X"08",X"C9",X"33",X"03",X"08",X"C9",X"4B",X"03",X"08",X"C9",X"63",X"03",X"08",X"C9",X"7B",X"03",
		X"08",X"C9",X"93",X"03",X"08",X"C9",X"AB",X"03",X"08",X"C9",X"C3",X"03",X"08",X"C9",X"DB",X"03",
		X"08",X"C9",X"F3",X"04",X"08",X"CA",X"0B",X"03",X"08",X"CA",X"2B",X"03",X"08",X"CA",X"43",X"03",
		X"08",X"CA",X"5B",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"01",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"01",X"01",X"01",X"01",
		X"01",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"10",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"01",X"01",X"00",X"00",X"00",
		X"01",X"01",X"00",X"11",X"00",X"00",X"01",X"10",X"00",X"11",X"00",X"11",X"01",X"01",X"10",X"00",
		X"00",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"11",X"01",X"01",X"11",X"01",X"01",X"11",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"01",X"10",X"00",X"11",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"11",X"10",
		X"10",X"10",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"01",
		X"01",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",
		X"10",X"10",X"00",X"11",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",X"01",X"01",X"10",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"11",X"01",X"01",X"11",X"01",X"01",X"11",X"00",X"00",X"00",X"01",X"00",X"00",
		X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"01",
		X"00",X"01",X"00",X"11",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"11",X"01",
		X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"11",X"01",X"01",X"11",X"01",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"10",X"01",X"01",X"01",X"01",X"01",X"10",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"10",X"00",
		X"00",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"11",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"11",X"01",
		X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"10",X"01",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"01",X"01",X"01",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"01",X"01",X"01",X"01",
		X"11",X"11",X"10",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"11",X"01",X"01",X"11",X"10",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"00",
		X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"01",
		X"01",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"10",X"10",X"10",X"10",X"10",
		X"10",X"01",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"10",X"01",X"10",X"00",X"00",X"00",X"01",X"01",X"10",X"00",X"10",
		X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"01",
		X"01",X"01",X"00",X"01",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"01",X"01",X"00",X"11",X"00",X"01",X"10",X"00",X"00",X"11",X"00",X"11",X"10",X"00",X"00",X"00",
		X"00",X"11",X"00",X"FF",X"FF",X"34",X"70",X"CE",X"C0",X"D9",X"20",X"05",X"34",X"70",X"CE",X"C0",
		X"BB",X"8E",X"18",X"CE",X"BD",X"CA",X"D4",X"EE",X"A1",X"27",X"06",X"8E",X"10",X"DA",X"BD",X"CA",
		X"D4",X"EE",X"A1",X"27",X"06",X"8E",X"10",X"E4",X"BD",X"CA",X"D4",X"35",X"F0",X"34",X"77",X"10",
		X"8E",X"FF",X"B9",X"20",X"06",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CC",X"CB",X"22",X"10",X"BF",
		X"B2",X"03",X"FD",X"B2",X"05",X"BF",X"B2",X"16",X"BF",X"B2",X"14",X"8E",X"01",X"0A",X"BF",X"B2",
		X"12",X"7F",X"B2",X"1E",X"EE",X"65",X"FF",X"B2",X"1A",X"33",X"C8",X"20",X"FF",X"B2",X"1C",X"FF",
		X"B2",X"18",X"20",X"4E",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CC",X"CB",X"22",X"20",X"1F",X"34",
		X"77",X"10",X"8E",X"FF",X"B9",X"CC",X"CB",X"22",X"20",X"14",X"34",X"77",X"10",X"8E",X"FF",X"B6",
		X"CC",X"CB",X"85",X"20",X"09",X"34",X"77",X"10",X"8E",X"FF",X"B9",X"CC",X"CB",X"85",X"10",X"BF",
		X"B2",X"03",X"FD",X"B2",X"05",X"7D",X"B2",X"18",X"26",X"18",X"BF",X"B2",X"16",X"BF",X"B2",X"14",
		X"8E",X"01",X"0A",X"BF",X"B2",X"12",X"7F",X"B2",X"1E",X"AE",X"42",X"BF",X"B2",X"1C",X"AE",X"C4",
		X"20",X"28",X"7D",X"B2",X"1E",X"26",X"10",X"BE",X"B2",X"1A",X"E6",X"80",X"C1",X"2F",X"26",X"33",
		X"C6",X"20",X"F7",X"B2",X"1E",X"20",X"2C",X"7F",X"B2",X"1E",X"BE",X"B2",X"18",X"BC",X"B2",X"1C",
		X"26",X"08",X"7F",X"B2",X"18",X"35",X"77",X"1A",X"01",X"39",X"EE",X"81",X"2B",X"0D",X"30",X"1F",
		X"1F",X"30",X"48",X"10",X"8E",X"CB",X"8A",X"AD",X"B6",X"20",X"E2",X"BF",X"B2",X"18",X"FF",X"B2",
		X"1A",X"20",X"BF",X"BF",X"B2",X"1A",X"C0",X"20",X"58",X"58",X"8E",X"C5",X"E7",X"3A",X"1F",X"12",
		X"FC",X"B2",X"16",X"BE",X"B2",X"03",X"AD",X"84",X"AB",X"A4",X"BB",X"B2",X"12",X"B7",X"B2",X"16",
		X"BE",X"B2",X"05",X"6E",X"84",X"35",X"77",X"1C",X"FE",X"39",X"CB",X"9C",X"CB",X"A2",X"CB",X"A8",
		X"CB",X"B1",X"CB",X"BA",X"CB",X"C3",X"CB",X"CC",X"CB",X"D5",X"CB",X"E2",X"A6",X"80",X"B7",X"B2",
		X"12",X"39",X"E6",X"80",X"F7",X"B2",X"13",X"39",X"B6",X"B2",X"14",X"AB",X"80",X"B7",X"B2",X"16",
		X"39",X"B6",X"B2",X"16",X"AB",X"80",X"B7",X"B2",X"16",X"39",X"F6",X"B2",X"15",X"EB",X"80",X"F7",
		X"B2",X"17",X"39",X"F6",X"B2",X"17",X"EB",X"80",X"F7",X"B2",X"17",X"39",X"EC",X"81",X"FD",X"B2",
		X"14",X"FD",X"B2",X"16",X"39",X"B6",X"B2",X"14",X"F6",X"B2",X"17",X"FB",X"B2",X"13",X"FD",X"B2",
		X"16",X"39",X"10",X"AE",X"81",X"BF",X"B2",X"18",X"BE",X"B2",X"03",X"AD",X"84",X"AB",X"A4",X"BB",
		X"B2",X"12",X"B7",X"B2",X"16",X"32",X"62",X"BE",X"B2",X"05",X"6E",X"84",X"34",X"77",X"10",X"8E",
		X"FF",X"B6",X"CE",X"CC",X"51",X"20",X"1F",X"34",X"77",X"10",X"8E",X"FF",X"B9",X"CE",X"CC",X"51",
		X"20",X"14",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CE",X"CC",X"83",X"20",X"09",X"34",X"77",X"10",
		X"8E",X"FF",X"B9",X"CE",X"CC",X"83",X"10",X"BF",X"B2",X"03",X"FF",X"B2",X"05",X"FE",X"B2",X"1F",
		X"11",X"83",X"FF",X"FF",X"26",X"18",X"BF",X"B2",X"16",X"FD",X"B2",X"1F",X"26",X"05",X"CC",X"0F",
		X"FF",X"20",X"08",X"85",X"F0",X"26",X"04",X"8D",X"3F",X"20",X"F8",X"FD",X"B2",X"1F",X"FC",X"B2",
		X"1F",X"84",X"F0",X"81",X"F0",X"26",X"08",X"35",X"77",X"BE",X"B2",X"16",X"1A",X"01",X"39",X"44",
		X"44",X"8E",X"C6",X"27",X"31",X"86",X"FC",X"B2",X"16",X"BE",X"B2",X"03",X"AD",X"84",X"AB",X"A4",
		X"BB",X"B2",X"12",X"B7",X"B2",X"16",X"FC",X"B2",X"1F",X"8D",X"0D",X"FD",X"B2",X"1F",X"BE",X"B2",
		X"05",X"6E",X"84",X"35",X"77",X"1C",X"FE",X"39",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",
		X"CA",X"0F",X"39",X"CC",X"CC",X"CC",X"0C",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"08",X"82",X"82",X"08",X"00",X"33",X"33",X"00",
		X"80",X"28",X"28",X"80",X"02",X"28",X"28",X"02",X"00",X"33",X"33",X"00",X"20",X"82",X"82",X"20",
		X"00",X"00",X"02",X"22",X"22",X"28",X"20",X"02",X"03",X"35",X"35",X"33",X"88",X"00",X"00",X"00",
		X"30",X"53",X"53",X"33",X"88",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"22",X"82",X"02",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"82",X"80",X"08",
		X"03",X"35",X"35",X"33",X"22",X"00",X"00",X"00",X"30",X"53",X"53",X"33",X"22",X"00",X"00",X"00",
		X"00",X"00",X"80",X"88",X"88",X"28",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"82",X"82",X"82",X"08",X"00",X"00",X"80",X"22",X"22",X"20",X"20",X"22",X"80",X"00",
		X"80",X"22",X"26",X"02",X"26",X"22",X"80",X"00",X"00",X"00",X"60",X"66",X"60",X"03",X"00",X"00",
		X"00",X"22",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"08",X"82",X"82",X"82",X"08",X"00",X"00",
		X"80",X"22",X"00",X"06",X"22",X"22",X"80",X"00",X"80",X"22",X"22",X"66",X"68",X"68",X"66",X"00",
		X"00",X"00",X"20",X"00",X"80",X"02",X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"20",X"00",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"00",X"33",X"33",X"33",X"33",X"30",X"00",X"00",
		X"00",X"33",X"03",X"03",X"33",X"30",X"30",X"30",X"00",X"30",X"33",X"33",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"33",X"33",X"03",X"03",X"30",X"00",X"00",X"33",X"30",X"30",X"03",X"03",X"03",X"03",
		X"00",X"33",X"33",X"33",X"33",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"02",X"22",X"02",X"22",X"20",X"66",X"22",X"06",X"05",X"05",X"06",X"60",X"50",X"50",X"60",
		X"22",X"02",X"66",X"22",X"00",X"20",X"22",X"20",X"00",X"03",X"33",X"03",X"33",X"30",X"66",X"33",
		X"06",X"02",X"02",X"06",X"60",X"20",X"20",X"60",X"33",X"03",X"66",X"33",X"00",X"30",X"33",X"30",
		X"00",X"03",X"30",X"03",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"33",X"07",X"40",X"33",
		X"30",X"03",X"44",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"04",X"33",
		X"33",X"07",X"40",X"33",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"00",X"30",X"43",X"30",
		X"00",X"03",X"34",X"03",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"33",X"70",X"44",X"33",
		X"30",X"03",X"04",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"40",X"33",
		X"33",X"70",X"44",X"33",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"00",X"30",X"43",X"30",
		X"60",X"66",X"66",X"66",X"55",X"05",X"00",X"00",X"60",X"66",X"56",X"50",X"00",X"00",X"00",X"66",
		X"65",X"00",X"00",X"00",X"06",X"66",X"55",X"55",X"00",X"06",X"66",X"66",X"55",X"50",X"00",X"66",
		X"6C",X"6C",X"55",X"55",X"00",X"00",X"C0",X"CC",X"66",X"60",X"00",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"06",X"66",X"66",X"28",X"68",X"08",X"60",X"66",X"66",X"86",
		X"88",X"88",X"00",X"00",X"60",X"66",X"86",X"69",X"00",X"00",X"00",X"66",X"66",X"30",X"00",X"00",
		X"00",X"DE",X"66",X"00",X"00",X"00",X"00",X"F0",X"66",X"00",X"00",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"00",X"03",X"33",X"03",X"00",X"00",X"00",X"33",X"E3",X"33",X"02",X"02",X"6E",X"33",
		X"E3",X"33",X"00",X"60",X"E6",X"33",X"E3",X"33",X"00",X"00",X"60",X"33",X"E3",X"33",X"00",X"00",
		X"00",X"33",X"E3",X"33",X"00",X"00",X"00",X"33",X"E3",X"33",X"00",X"00",X"00",X"0C",X"30",X"0C",
		X"00",X"00",X"00",X"C0",X"03",X"C0",X"00",X"00",X"00",X"33",X"3E",X"33",X"00",X"00",X"00",X"33",
		X"3E",X"33",X"00",X"00",X"06",X"33",X"3E",X"33",X"00",X"06",X"6E",X"33",X"3E",X"33",X"20",X"20",
		X"E6",X"33",X"3E",X"33",X"00",X"00",X"00",X"33",X"3E",X"33",X"00",X"00",X"00",X"30",X"33",X"30",
		X"60",X"56",X"33",X"05",X"00",X"00",X"55",X"50",X"00",X"06",X"55",X"33",X"66",X"6C",X"55",X"35",
		X"00",X"C0",X"52",X"00",X"06",X"06",X"06",X"FF",X"FF",X"FF",X"60",X"60",X"60",X"00",X"00",X"00",
		X"00",X"03",X"03",X"03",X"03",X"C0",X"80",X"80",X"80",X"83",X"03",X"03",X"03",X"11",X"00",X"10",
		X"00",X"10",X"10",X"10",X"00",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"10",
		X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"11",X"01",X"11",X"00",X"11",X"00",X"01",X"01",X"01",
		X"00",X"01",X"00",X"11",X"00",X"11",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"01",X"01",X"01",X"11",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"F0",
		X"00",X"EE",X"E0",X"E0",X"E0",X"EE",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"DD",X"D0",X"D0",
		X"D0",X"DD",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"00",X"FF",
		X"00",X"FF",X"0F",X"FF",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"0E",X"EE",
		X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"DD",X"0D",X"0D",X"0D",X"DD",X"00",X"00",X"0E",X"CF",
		X"CE",X"0C",X"00",X"CC",X"AB",X"CD",X"EF",X"DC",X"CE",X"00",X"B0",X"EC",X"CF",X"C0",X"00",X"0D",
		X"CF",X"CE",X"AC",X"CE",X"0B",X"E0",X"DC",X"CE",X"DE",X"EC",X"F0",X"00",X"0A",X"CD",X"EC",X"0F",
		X"FC",X"AF",X"BC",X"CE",X"DC",X"CF",X"B0",X"EC",X"FE",X"D0",X"00",X"70",X"F0",X"00",X"00",X"00",
		X"7E",X"C0",X"76",X"7E",X"C0",X"9F",X"7E",X"C0",X"BE",X"7E",X"C0",X"F1",X"7E",X"CB",X"DC",X"7E",
		X"CB",X"D6",X"7E",X"CC",X"1E",X"7E",X"CC",X"12",X"7E",X"CC",X"18",X"7E",X"CC",X"A9",X"7E",X"CB",
		X"A5",X"7E",X"C7",X"9A",X"7E",X"C1",X"12",X"7E",X"C1",X"43",X"7E",X"C2",X"5C",X"7E",X"C2",X"EF",
		X"7E",X"C4",X"3C",X"7E",X"CC",X"BB",X"7E",X"FF",X"D4",X"7E",X"FF",X"D7",X"BD",X"FF",X"CE",X"C0",
		X"02",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"05",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"0E",X"02",
		X"39",X"BD",X"FF",X"CE",X"C0",X"11",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"1A",X"02",X"39",X"BD",
		X"FF",X"CE",X"C0",X"1D",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"20",X"02",X"39",X"BD",X"FF",X"CE",
		X"C0",X"23",X"02",X"39",X"FF",X"FF",X"BD",X"CA",X"E9",X"BD",X"CA",X"0A",X"C6",X"7A",X"BD",X"C7",
		X"94",X"CE",X"C0",X"69",X"8E",X"28",X"70",X"BD",X"C0",X"3C",X"CE",X"C0",X"6B",X"8E",X"40",X"90",
		X"BD",X"C0",X"3C",X"C6",X"0F",X"BD",X"CA",X"B3",X"10",X"8E",X"0B",X"B8",X"7E",X"CA",X"24",X"BD",
		X"CA",X"E9",X"BD",X"CA",X"0A",X"C6",X"57",X"BD",X"C7",X"94",X"CE",X"C0",X"69",X"8E",X"28",X"70",
		X"BD",X"C0",X"3C",X"CE",X"C0",X"73",X"8E",X"38",X"90",X"BD",X"C0",X"3C",X"20",X"2C",X"BD",X"CA",
		X"E9",X"BD",X"CA",X"0A",X"C6",X"57",X"BD",X"C7",X"94",X"CE",X"C0",X"69",X"8E",X"28",X"60",X"BD",
		X"C0",X"3C",X"CE",X"C0",X"71",X"8E",X"38",X"80",X"BD",X"C0",X"3C",X"1F",X"B8",X"81",X"9E",X"27",
		X"09",X"CE",X"C0",X"73",X"8E",X"38",X"A0",X"BD",X"C0",X"3C",X"10",X"8E",X"75",X"30",X"7E",X"CA",
		X"24",X"1C",X"EF",X"8E",X"C4",X"7F",X"BD",X"FF",X"A7",X"7E",X"C1",X"23",X"12",X"8E",X"C4",X"7D",
		X"BD",X"FF",X"A7",X"34",X"04",X"5F",X"8E",X"C4",X"7D",X"BD",X"FF",X"B0",X"35",X"04",X"C1",X"15",
		X"26",X"04",X"1C",X"7F",X"20",X"2D",X"C1",X"35",X"26",X"05",X"BD",X"CB",X"B5",X"20",X"0C",X"C1",
		X"45",X"26",X"08",X"32",X"62",X"BD",X"CB",X"C5",X"7E",X"C7",X"9A",X"39",X"CA",X"0A",X"C6",X"A5",
		X"BD",X"C7",X"94",X"CE",X"C0",X"75",X"8E",X"38",X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"31",
		X"7E",X"C0",X"6D",X"1A",X"10",X"BD",X"CA",X"0A",X"BD",X"FF",X"BF",X"34",X"40",X"FE",X"FF",X"A2",
		X"33",X"C8",X"18",X"FF",X"B2",X"09",X"35",X"40",X"11",X"B3",X"B2",X"09",X"10",X"27",X"00",X"8A",
		X"FF",X"B2",X"21",X"C6",X"08",X"BD",X"CA",X"95",X"C6",X"57",X"BD",X"C7",X"94",X"CE",X"C0",X"71",
		X"8E",X"38",X"60",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"35",X"BD",X"C0",X"6D",X"CC",X"42",X"66",
		X"FD",X"B2",X"10",X"BE",X"B2",X"10",X"30",X"0A",X"BF",X"B2",X"10",X"CE",X"C0",X"6D",X"BD",X"C0",
		X"3C",X"FE",X"FF",X"A2",X"FF",X"B2",X"09",X"FE",X"B2",X"21",X"FC",X"B2",X"21",X"B3",X"B2",X"09",
		X"54",X"25",X"02",X"33",X"41",X"5C",X"BD",X"CB",X"13",X"BE",X"B2",X"16",X"BD",X"CB",X"FC",X"BD",
		X"CA",X"4E",X"BD",X"FF",X"C2",X"FF",X"B2",X"21",X"FE",X"FF",X"A2",X"33",X"C8",X"18",X"11",X"B3",
		X"B2",X"21",X"26",X"BF",X"BD",X"C9",X"EE",X"7D",X"B2",X"0F",X"26",X"40",X"34",X"40",X"FE",X"FF",
		X"A2",X"FF",X"B2",X"09",X"35",X"40",X"FC",X"B2",X"21",X"B3",X"B2",X"09",X"54",X"5C",X"BD",X"CA",
		X"95",X"10",X"8E",X"C0",X"39",X"BD",X"C0",X"6D",X"20",X"1F",X"1F",X"A9",X"5D",X"2A",X"40",X"C6",
		X"7A",X"BD",X"C7",X"94",X"CE",X"C0",X"77",X"8E",X"38",X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",
		X"39",X"BD",X"C0",X"6D",X"C6",X"08",X"BD",X"CA",X"B3",X"BD",X"CA",X"18",X"BD",X"CA",X"0A",X"5F",
		X"BD",X"CA",X"95",X"C6",X"A5",X"BD",X"C7",X"94",X"CE",X"C0",X"79",X"8E",X"40",X"80",X"BD",X"C0",
		X"3C",X"10",X"8E",X"C0",X"3D",X"BD",X"C0",X"6D",X"10",X"8E",X"13",X"88",X"BD",X"CA",X"24",X"BD",
		X"CA",X"38",X"7D",X"B2",X"0F",X"10",X"26",X"00",X"E5",X"7D",X"B2",X"0D",X"26",X"F1",X"8E",X"C0",
		X"00",X"C6",X"C0",X"BD",X"C0",X"36",X"86",X"B5",X"3D",X"1E",X"89",X"30",X"01",X"8C",X"C0",X"10",
		X"26",X"F1",X"CC",X"00",X"00",X"10",X"8E",X"00",X"0A",X"7E",X"FF",X"C5",X"1F",X"20",X"E8",X"82",
		X"A8",X"82",X"FD",X"B2",X"07",X"BF",X"B2",X"09",X"BD",X"CA",X"E9",X"BD",X"FF",X"BC",X"BD",X"CA",
		X"CF",X"BD",X"CA",X"4E",X"C6",X"04",X"BD",X"CA",X"95",X"C6",X"57",X"BD",X"C7",X"94",X"CE",X"C0",
		X"73",X"8E",X"38",X"70",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"41",X"BD",X"C0",X"6D",X"FC",X"B2",
		X"07",X"4D",X"26",X"02",X"1F",X"98",X"5F",X"5C",X"44",X"24",X"FC",X"F7",X"B2",X"00",X"FC",X"B2",
		X"09",X"80",X"03",X"24",X"FC",X"8B",X"04",X"B7",X"B2",X"01",X"CE",X"C0",X"6F",X"8E",X"42",X"90",
		X"BD",X"C0",X"3C",X"F6",X"B2",X"01",X"58",X"58",X"58",X"58",X"FB",X"B2",X"00",X"4F",X"BE",X"B2",
		X"16",X"BD",X"C0",X"4A",X"BD",X"C9",X"EE",X"7D",X"B2",X"0F",X"26",X"52",X"B6",X"B2",X"01",X"C6",
		X"10",X"54",X"4A",X"26",X"FC",X"BD",X"CA",X"95",X"BD",X"C9",X"EE",X"7D",X"B2",X"0F",X"26",X"3E",
		X"F6",X"B2",X"00",X"BD",X"CA",X"95",X"10",X"8E",X"C0",X"45",X"BD",X"C0",X"6D",X"20",X"2C",X"BD",
		X"CA",X"E9",X"BD",X"FF",X"BC",X"BD",X"CA",X"CF",X"BD",X"CA",X"4E",X"10",X"8C",X"00",X"0A",X"27",
		X"1D",X"C6",X"7A",X"BD",X"C7",X"94",X"CE",X"C0",X"7B",X"8E",X"28",X"80",X"BD",X"C0",X"3C",X"10",
		X"8E",X"C0",X"45",X"BD",X"C0",X"6D",X"C6",X"04",X"BD",X"CA",X"B3",X"BD",X"CA",X"18",X"BD",X"CA",
		X"0A",X"1F",X"B8",X"81",X"A2",X"26",X"1D",X"C6",X"02",X"BD",X"CA",X"95",X"C6",X"57",X"BD",X"C7",
		X"94",X"CE",X"C0",X"81",X"8E",X"28",X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"49",X"BD",X"C0",
		X"6D",X"7E",X"C3",X"EE",X"8B",X"03",X"5F",X"FD",X"B2",X"07",X"FE",X"B2",X"07",X"8E",X"C4",X"00",
		X"BD",X"C0",X"39",X"E7",X"C0",X"30",X"01",X"8C",X"C5",X"00",X"26",X"F4",X"CC",X"00",X"10",X"F7",
		X"B2",X"00",X"8E",X"C4",X"00",X"F6",X"B2",X"00",X"BD",X"C0",X"36",X"30",X"01",X"5C",X"F1",X"B2",
		X"00",X"26",X"F5",X"BD",X"C0",X"39",X"F7",X"B2",X"01",X"30",X"01",X"BD",X"C0",X"39",X"F0",X"B2",
		X"01",X"5A",X"C4",X"0F",X"26",X"10",X"4C",X"26",X"EA",X"BD",X"CA",X"4E",X"7D",X"B2",X"0F",X"26",
		X"05",X"7A",X"B2",X"00",X"26",X"CC",X"FE",X"B2",X"07",X"8E",X"C4",X"00",X"E6",X"C0",X"BD",X"C0",
		X"36",X"30",X"01",X"8C",X"C5",X"00",X"26",X"F4",X"7D",X"B2",X"0F",X"26",X"44",X"B6",X"B2",X"00",
		X"27",X"22",X"C6",X"02",X"BD",X"CA",X"95",X"C6",X"57",X"BD",X"C7",X"94",X"BD",X"CA",X"4E",X"CE",
		X"C0",X"7D",X"8E",X"30",X"80",X"BD",X"C0",X"3C",X"BD",X"CA",X"4E",X"10",X"8E",X"C0",X"49",X"BD",
		X"C0",X"6D",X"20",X"1A",X"C6",X"7A",X"BD",X"C7",X"94",X"CE",X"C0",X"7F",X"8E",X"38",X"80",X"BD",
		X"C0",X"3C",X"10",X"8E",X"C0",X"49",X"BD",X"C0",X"6D",X"C6",X"02",X"BD",X"CA",X"B3",X"BD",X"CA",
		X"18",X"BD",X"CA",X"0A",X"C6",X"01",X"BD",X"CA",X"95",X"C6",X"A5",X"BD",X"C7",X"94",X"CE",X"C0",
		X"83",X"8E",X"38",X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"4D",X"BD",X"C0",X"6D",X"10",X"8E",
		X"13",X"88",X"BD",X"CA",X"24",X"BD",X"CB",X"5A",X"10",X"8E",X"07",X"D0",X"CE",X"C9",X"BA",X"E6",
		X"C0",X"8E",X"C0",X"00",X"BD",X"C0",X"36",X"30",X"01",X"8C",X"C0",X"10",X"26",X"F6",X"BD",X"CA",
		X"24",X"11",X"83",X"C9",X"C2",X"26",X"E8",X"7D",X"B2",X"0F",X"27",X"E0",X"BD",X"CA",X"E9",X"BD",
		X"CA",X"0A",X"5F",X"F7",X"B2",X"07",X"F7",X"B2",X"08",X"BD",X"CA",X"95",X"C6",X"A5",X"BD",X"C7",
		X"94",X"CE",X"C0",X"85",X"8E",X"40",X"78",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"55",X"BD",X"C0",
		X"6D",X"10",X"8E",X"00",X"01",X"CE",X"C9",X"D2",X"4F",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",
		X"01",X"26",X"09",X"C5",X"02",X"26",X"16",X"BD",X"CA",X"38",X"20",X"ED",X"BD",X"CA",X"24",X"4C",
		X"A1",X"C4",X"26",X"04",X"33",X"41",X"20",X"F7",X"B7",X"B2",X"00",X"88",X"3F",X"C6",X"13",X"BD",
		X"CA",X"FB",X"7D",X"B2",X"0F",X"26",X"33",X"F6",X"B2",X"00",X"BD",X"CA",X"FB",X"10",X"8E",X"03",
		X"E8",X"FC",X"B2",X"07",X"8E",X"5A",X"8C",X"BD",X"C0",X"51",X"F6",X"B2",X"00",X"BD",X"CB",X"13",
		X"4F",X"FD",X"B2",X"07",X"8E",X"5A",X"8C",X"BD",X"C0",X"4A",X"B6",X"B2",X"00",X"81",X"1F",X"26",
		X"A8",X"1F",X"A9",X"5D",X"10",X"2A",X"00",X"B4",X"20",X"9B",X"BD",X"CA",X"0A",X"CE",X"C0",X"87",
		X"8E",X"38",X"20",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"59",X"BD",X"C0",X"6D",X"CC",X"B2",X"26",
		X"FD",X"B2",X"07",X"CC",X"B2",X"36",X"1F",X"01",X"86",X"FF",X"A7",X"82",X"BC",X"B2",X"07",X"26",
		X"F9",X"7F",X"B2",X"36",X"7F",X"B2",X"37",X"7F",X"B2",X"38",X"8E",X"CC",X"00",X"FE",X"B2",X"07",
		X"33",X"C8",X"10",X"4F",X"BD",X"C0",X"39",X"F7",X"B2",X"00",X"E8",X"C0",X"26",X"1E",X"8B",X"08",
		X"30",X"02",X"8C",X"CC",X"02",X"27",X"F9",X"8C",X"CC",X"08",X"26",X"E8",X"7C",X"B2",X"02",X"26",
		X"00",X"BD",X"CA",X"4E",X"7D",X"B2",X"0F",X"27",X"D1",X"7E",X"C5",X"7C",X"F7",X"B2",X"01",X"C6",
		X"01",X"F5",X"B2",X"01",X"26",X"04",X"4C",X"58",X"20",X"F7",X"BE",X"B2",X"07",X"F5",X"B2",X"00",
		X"26",X"10",X"E8",X"C2",X"E7",X"C4",X"A1",X"80",X"26",X"FC",X"63",X"82",X"10",X"8E",X"C0",X"43",
		X"20",X"13",X"E8",X"C2",X"E7",X"C4",X"C6",X"08",X"BD",X"CA",X"FB",X"6D",X"80",X"2A",X"FC",X"A7",
		X"82",X"10",X"8E",X"C0",X"3C",X"CE",X"C0",X"8B",X"48",X"33",X"C6",X"1F",X"10",X"B3",X"B2",X"07",
		X"86",X"0A",X"3D",X"C3",X"38",X"30",X"1F",X"01",X"AD",X"A4",X"20",X"A0",X"BD",X"CA",X"0A",X"CE",
		X"C0",X"89",X"8E",X"28",X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"5D",X"BD",X"C0",X"6D",X"8E",
		X"CC",X"00",X"CE",X"C9",X"D4",X"BD",X"C0",X"39",X"C5",X"01",X"27",X"15",X"10",X"8E",X"13",X"88",
		X"BD",X"CA",X"24",X"7D",X"B2",X"0F",X"10",X"26",X"01",X"F0",X"BD",X"C0",X"39",X"C5",X"01",X"26",
		X"0A",X"BD",X"C9",X"EE",X"7D",X"B2",X"0F",X"10",X"26",X"01",X"DF",X"34",X"70",X"AD",X"D4",X"35",
		X"70",X"33",X"42",X"11",X"83",X"C9",X"DE",X"26",X"CC",X"10",X"8E",X"13",X"88",X"BD",X"CA",X"24",
		X"1F",X"A9",X"5D",X"10",X"2A",X"FB",X"6C",X"20",X"B9",X"BD",X"CA",X"4E",X"BD",X"FF",X"BC",X"BD",
		X"CA",X"E9",X"8E",X"C0",X"01",X"C6",X"FF",X"BD",X"C0",X"36",X"8E",X"C0",X"02",X"C6",X"C0",X"BD",
		X"C0",X"36",X"8E",X"C0",X"03",X"C6",X"38",X"BD",X"C0",X"36",X"8E",X"C0",X"04",X"C6",X"07",X"BD",
		X"C0",X"36",X"BD",X"CA",X"4E",X"10",X"8E",X"C6",X"FA",X"CC",X"01",X"01",X"AE",X"A4",X"ED",X"81",
		X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"C7",X"22",X"26",X"F0",X"BD",X"CA",X"4E",X"86",
		X"11",X"10",X"8E",X"C6",X"DA",X"AE",X"A4",X"BF",X"B2",X"0B",X"A7",X"84",X"7C",X"B2",X"0B",X"BE",
		X"B2",X"0B",X"AC",X"22",X"26",X"F4",X"31",X"24",X"10",X"8C",X"C6",X"FA",X"26",X"E7",X"BD",X"CA",
		X"4E",X"10",X"8E",X"C7",X"22",X"AE",X"A4",X"BF",X"B2",X"0B",X"A6",X"24",X"A7",X"84",X"7C",X"B2",
		X"0B",X"BE",X"B2",X"0B",X"AC",X"22",X"26",X"F4",X"31",X"25",X"10",X"8C",X"C7",X"5E",X"26",X"E5",
		X"BD",X"CA",X"4E",X"10",X"8E",X"C7",X"5E",X"AE",X"A4",X"A6",X"24",X"A7",X"80",X"AC",X"22",X"26",
		X"FA",X"31",X"25",X"10",X"8C",X"C7",X"72",X"26",X"EE",X"BD",X"CA",X"4E",X"86",X"21",X"B7",X"46",
		X"7E",X"86",X"20",X"B7",X"96",X"7E",X"8E",X"4E",X"0A",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"A7",
		X"80",X"8C",X"4E",X"6D",X"26",X"F3",X"8E",X"4E",X"90",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"A7",
		X"80",X"8C",X"4E",X"F3",X"26",X"F3",X"BD",X"CA",X"4E",X"8E",X"0E",X"18",X"BF",X"B2",X"0B",X"BE",
		X"B2",X"0B",X"A6",X"84",X"84",X"F0",X"8A",X"01",X"A7",X"84",X"F6",X"B2",X"0C",X"CB",X"22",X"25",
		X"05",X"F7",X"B2",X"0C",X"20",X"E9",X"C6",X"18",X"F7",X"B2",X"0C",X"F6",X"B2",X"0B",X"CB",X"10",
		X"F7",X"B2",X"0B",X"C1",X"9E",X"26",X"D8",X"7E",X"CA",X"4E",X"07",X"07",X"97",X"07",X"07",X"29",
		X"97",X"29",X"07",X"4B",X"97",X"4B",X"07",X"6D",X"97",X"6D",X"07",X"8F",X"97",X"8F",X"07",X"B1",
		X"97",X"B1",X"07",X"D3",X"97",X"D3",X"07",X"F5",X"97",X"F5",X"06",X"07",X"06",X"F5",X"16",X"07",
		X"16",X"F5",X"26",X"07",X"26",X"F5",X"36",X"07",X"36",X"F5",X"46",X"07",X"46",X"F5",X"56",X"07",
		X"56",X"F5",X"66",X"07",X"66",X"F5",X"76",X"07",X"76",X"F5",X"86",X"07",X"86",X"F5",X"96",X"07",
		X"96",X"F5",X"48",X"05",X"55",X"05",X"44",X"48",X"06",X"55",X"06",X"44",X"48",X"07",X"55",X"07",
		X"00",X"48",X"08",X"55",X"08",X"33",X"48",X"09",X"55",X"09",X"33",X"48",X"F3",X"55",X"F3",X"33",
		X"48",X"F4",X"55",X"F4",X"33",X"48",X"F5",X"55",X"F5",X"00",X"48",X"F6",X"55",X"F6",X"44",X"48",
		X"F7",X"55",X"F7",X"44",X"07",X"7E",X"46",X"7E",X"22",X"57",X"7E",X"96",X"7E",X"22",X"05",X"6F",
		X"05",X"8E",X"04",X"06",X"6F",X"06",X"8E",X"30",X"96",X"6F",X"96",X"8E",X"00",X"97",X"6F",X"97",
		X"8E",X"34",X"BD",X"FF",X"BC",X"C6",X"05",X"8E",X"C0",X"00",X"8D",X"03",X"8E",X"C0",X"0C",X"7E",
		X"C0",X"36",X"C6",X"28",X"20",X"F1",X"C6",X"80",X"20",X"ED",X"10",X"8E",X"C9",X"DE",X"BD",X"CA",
		X"82",X"7E",X"CB",X"2B",X"8E",X"C0",X"01",X"7E",X"C0",X"36",X"8E",X"CC",X"06",X"BD",X"FF",X"D7",
		X"54",X"C4",X"1F",X"86",X"03",X"C5",X"10",X"27",X"02",X"86",X"05",X"1E",X"89",X"8E",X"C4",X"85",
		X"BD",X"F8",X"59",X"84",X"0F",X"34",X"02",X"AB",X"E4",X"AB",X"E4",X"10",X"8E",X"C7",X"D8",X"E6",
		X"A6",X"4C",X"8E",X"C4",X"89",X"BD",X"F8",X"59",X"E6",X"A6",X"4C",X"BD",X"F8",X"59",X"E6",X"A6",
		X"30",X"02",X"BD",X"F8",X"59",X"7E",X"D8",X"16",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"03",
		X"01",X"01",X"06",X"01",X"01",X"02",X"02",X"01",X"04",X"02",X"01",X"06",X"02",X"01",X"12",X"02",
		X"01",X"03",X"03",X"01",X"06",X"03",X"01",X"09",X"03",X"01",X"18",X"03",X"01",X"04",X"04",X"01",
		X"08",X"04",X"01",X"12",X"04",X"01",X"24",X"04",X"34",X"02",X"AB",X"E4",X"34",X"02",X"AB",X"E4",
		X"AB",X"E4",X"35",X"24",X"7E",X"C7",X"BB",X"26",X"27",X"32",X"E8",X"20",X"BD",X"CA",X"4E",X"BD",
		X"C1",X"2B",X"7E",X"FF",X"C8",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",X"01",X"26",X"11",X"C5",
		X"02",X"27",X"0D",X"7C",X"B2",X"01",X"7A",X"B2",X"02",X"2A",X"05",X"C6",X"1B",X"F7",X"B2",X"02",
		X"BD",X"C9",X"69",X"7D",X"B2",X"01",X"27",X"B5",X"F6",X"B2",X"02",X"C1",X"09",X"26",X"25",X"8E",
		X"C4",X"87",X"BD",X"FF",X"A7",X"5D",X"27",X"1C",X"C1",X"08",X"22",X"05",X"BD",X"CB",X"8F",X"20",
		X"13",X"8E",X"C4",X"87",X"34",X"10",X"C6",X"01",X"BD",X"FF",X"B0",X"BD",X"CB",X"8F",X"5F",X"35",
		X"10",X"BD",X"FF",X"B0",X"8D",X"05",X"7F",X"B2",X"01",X"20",X"82",X"31",X"62",X"8E",X"10",X"80",
		X"BD",X"C0",X"58",X"BD",X"C9",X"0C",X"B6",X"B2",X"02",X"4C",X"BD",X"C8",X"EF",X"BD",X"C8",X"FD",
		X"ED",X"84",X"F6",X"B2",X"02",X"58",X"58",X"8E",X"CC",X"D0",X"3A",X"10",X"AE",X"84",X"EE",X"02",
		X"30",X"6E",X"A6",X"A0",X"81",X"2F",X"27",X"04",X"A7",X"80",X"20",X"F6",X"1F",X"30",X"33",X"62",
		X"8E",X"C4",X"00",X"3A",X"BD",X"FF",X"A7",X"34",X"06",X"F6",X"B2",X"02",X"5C",X"C1",X"07",X"22",
		X"13",X"35",X"06",X"1F",X"98",X"BD",X"C8",X"FD",X"ED",X"47",X"BD",X"FF",X"A4",X"BD",X"C8",X"FD",
		X"ED",X"49",X"20",X"13",X"C1",X"08",X"26",X"09",X"CC",X"30",X"30",X"ED",X"49",X"33",X"5E",X"20",
		X"E0",X"35",X"06",X"1F",X"98",X"20",X"E6",X"8E",X"10",X"80",X"31",X"62",X"7E",X"C0",X"5F",X"34",
		X"04",X"1F",X"89",X"86",X"99",X"8B",X"01",X"19",X"5A",X"2A",X"FA",X"35",X"84",X"1F",X"89",X"84",
		X"F0",X"44",X"44",X"44",X"44",X"8B",X"30",X"C4",X"0F",X"CB",X"30",X"39",X"86",X"20",X"1F",X"89",
		X"5A",X"30",X"64",X"A7",X"80",X"5A",X"26",X"FB",X"86",X"2F",X"A7",X"80",X"30",X"64",X"39",X"02",
		X"00",X"00",X"4D",X"49",X"54",X"01",X"50",X"00",X"4E",X"4F",X"42",X"01",X"00",X"00",X"4E",X"55",
		X"4E",X"00",X"70",X"00",X"48",X"4F",X"4E",X"00",X"50",X"00",X"49",X"4B",X"55",X"FF",X"B3",X"BD",
		X"FF",X"A4",X"8B",X"01",X"19",X"30",X"1E",X"7C",X"B2",X"01",X"7E",X"FF",X"AD",X"8C",X"C4",X"81",
		X"26",X"10",X"BD",X"FF",X"AA",X"30",X"1C",X"1E",X"89",X"8B",X"90",X"19",X"1E",X"89",X"89",X"99",
		X"20",X"D2",X"BD",X"FF",X"A4",X"8B",X"99",X"20",X"DB",X"F6",X"B2",X"02",X"5C",X"C1",X"07",X"22",
		X"01",X"39",X"C1",X"09",X"23",X"11",X"C1",X"10",X"22",X"0D",X"C1",X"0A",X"27",X"09",X"8E",X"C4",
		X"87",X"BD",X"FF",X"A4",X"4D",X"26",X"EA",X"5A",X"58",X"58",X"8E",X"CC",X"D0",X"3A",X"E6",X"03",
		X"8E",X"C4",X"00",X"3A",X"34",X"10",X"BD",X"CA",X"38",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",
		X"02",X"27",X"02",X"35",X"90",X"C5",X"08",X"27",X"ED",X"10",X"8E",X"00",X"20",X"BD",X"CA",X"24",
		X"35",X"10",X"54",X"10",X"25",X"FF",X"68",X"7E",X"C9",X"4D",X"02",X"03",X"04",X"10",X"18",X"20",
		X"40",X"80",X"00",X"FF",X"11",X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",
		X"77",X"88",X"13",X"00",X"C5",X"D9",X"C7",X"72",X"C7",X"82",X"C7",X"86",X"C7",X"8A",X"05",X"05",
		X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",X"8E",X"CC",
		X"00",X"10",X"8E",X"00",X"64",X"BD",X"CA",X"24",X"BD",X"C0",X"39",X"C5",X"02",X"26",X"F6",X"BD",
		X"CA",X"24",X"BD",X"C0",X"39",X"C5",X"02",X"27",X"F6",X"39",X"BD",X"FF",X"BC",X"8D",X"3F",X"7A",
		X"B2",X"0F",X"2A",X"03",X"7F",X"B2",X"0F",X"39",X"10",X"8E",X"00",X"01",X"8D",X"06",X"7D",X"B2",
		X"0F",X"27",X"F9",X"39",X"34",X"23",X"8D",X"26",X"7D",X"B2",X"0F",X"26",X"09",X"86",X"B2",X"4A",
		X"26",X"FD",X"31",X"3F",X"26",X"F0",X"35",X"A3",X"34",X"24",X"F6",X"B2",X"0F",X"7F",X"B2",X"0F",
		X"10",X"8E",X"00",X"0A",X"8D",X"DE",X"FB",X"B2",X"0F",X"F7",X"B2",X"0F",X"35",X"A4",X"34",X"15",
		X"C6",X"38",X"8E",X"C3",X"FC",X"BD",X"C0",X"36",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"53",X"C4",
		X"03",X"27",X"02",X"1C",X"FE",X"F6",X"B2",X"0D",X"56",X"F7",X"B2",X"0D",X"26",X"03",X"F7",X"B2",
		X"0E",X"53",X"26",X"0C",X"F6",X"B2",X"0E",X"26",X"07",X"53",X"F7",X"B2",X"0E",X"7C",X"B2",X"0F",
		X"35",X"95",X"34",X"34",X"8E",X"C0",X"00",X"E6",X"A0",X"BD",X"C0",X"36",X"30",X"01",X"8C",X"C0",
		X"10",X"26",X"F4",X"35",X"B4",X"34",X"14",X"54",X"56",X"56",X"56",X"2A",X"01",X"5C",X"56",X"56",
		X"8E",X"CC",X"00",X"BD",X"C0",X"36",X"58",X"58",X"58",X"CA",X"3F",X"8E",X"CC",X"02",X"BD",X"C0",
		X"36",X"35",X"94",X"34",X"26",X"86",X"02",X"10",X"8E",X"01",X"F4",X"BD",X"CA",X"95",X"BD",X"CA",
		X"24",X"5F",X"BD",X"CA",X"95",X"BD",X"CA",X"24",X"E6",X"61",X"4A",X"26",X"EE",X"35",X"26",X"34",
		X"06",X"7F",X"B2",X"18",X"7F",X"B2",X"0F",X"86",X"01",X"B7",X"B2",X"0E",X"86",X"03",X"B7",X"A0",
		X"36",X"CC",X"FF",X"FF",X"FD",X"B2",X"1F",X"35",X"86",X"34",X"14",X"5F",X"8E",X"C0",X"00",X"BD",
		X"C0",X"36",X"30",X"01",X"8C",X"C0",X"10",X"26",X"F6",X"35",X"94",X"34",X"14",X"53",X"C4",X"3F",
		X"8E",X"CC",X"02",X"BD",X"C0",X"36",X"BD",X"CA",X"38",X"C6",X"3F",X"BD",X"C0",X"36",X"BD",X"CA",
		X"38",X"35",X"94",X"34",X"02",X"1F",X"98",X"84",X"0F",X"8B",X"00",X"19",X"C4",X"F0",X"27",X"07",
		X"8B",X"16",X"19",X"C0",X"10",X"20",X"F7",X"1F",X"89",X"35",X"82",X"34",X"16",X"CC",X"00",X"00",
		X"8E",X"00",X"00",X"BF",X"B2",X"03",X"30",X"89",X"0F",X"00",X"ED",X"83",X"BC",X"B2",X"03",X"26",
		X"F9",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0F",X"00",X"BD",X"CA",X"4E",X"7D",X"B2",
		X"0F",X"26",X"05",X"C3",X"11",X"11",X"24",X"DB",X"35",X"96",X"BD",X"CA",X"E9",X"8E",X"00",X"00",
		X"10",X"8E",X"C9",X"C2",X"BF",X"B2",X"03",X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",
		X"83",X"BC",X"B2",X"03",X"26",X"F9",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0F",X"00",
		X"BD",X"CA",X"4E",X"7D",X"B2",X"0F",X"26",X"06",X"10",X"8C",X"C9",X"D2",X"26",X"D6",X"39",X"8E",
		X"C4",X"87",X"BD",X"FF",X"B0",X"58",X"34",X"04",X"58",X"EB",X"E0",X"8E",X"CF",X"0A",X"3A",X"10",
		X"8E",X"C4",X"89",X"C6",X"06",X"34",X"02",X"A6",X"80",X"1E",X"12",X"BD",X"FF",X"AD",X"1E",X"12",
		X"5A",X"26",X"F4",X"35",X"82",X"C6",X"0E",X"20",X"01",X"5F",X"8E",X"C4",X"01",X"4F",X"BD",X"FF",
		X"AD",X"5A",X"26",X"FA",X"39",X"34",X"36",X"8D",X"F0",X"8E",X"CE",X"C9",X"10",X"8E",X"C4",X"1D",
		X"C6",X"47",X"8D",X"D1",X"35",X"B6",X"34",X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"07",
		X"27",X"1F",X"58",X"58",X"8E",X"C3",X"FD",X"3A",X"BD",X"FF",X"A7",X"34",X"04",X"BD",X"FF",X"A7",
		X"34",X"04",X"AB",X"E0",X"19",X"1E",X"89",X"35",X"02",X"89",X"00",X"19",X"30",X"1C",X"BD",X"FF",
		X"B3",X"35",X"96",X"34",X"02",X"BB",X"A0",X"37",X"19",X"24",X"02",X"86",X"99",X"B7",X"A0",X"37",
		X"35",X"82",X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",
		X"C6",X"01",X"BD",X"CB",X"D6",X"58",X"8E",X"C4",X"87",X"3A",X"BD",X"FF",X"A7",X"8D",X"6A",X"B6",
		X"A0",X"39",X"34",X"04",X"AB",X"E4",X"B7",X"A0",X"39",X"B6",X"A0",X"38",X"AB",X"E0",X"B7",X"A0",
		X"38",X"8E",X"C4",X"93",X"BD",X"FF",X"A7",X"8D",X"50",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",
		X"96",X"8E",X"C4",X"8F",X"BD",X"FF",X"A7",X"8D",X"40",X"8D",X"28",X"34",X"02",X"F7",X"A0",X"38",
		X"8E",X"C4",X"91",X"BD",X"FF",X"A7",X"B6",X"A0",X"39",X"8D",X"2E",X"8D",X"16",X"4D",X"27",X"06",
		X"7F",X"A0",X"38",X"7F",X"A0",X"39",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"CB",X"DC",X"BD",X"CC",
		X"03",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",
		X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",X"1E",X"89",X"5F",X"4D",X"26",
		X"02",X"35",X"82",X"8B",X"99",X"19",X"5C",X"20",X"F5",X"34",X"36",X"8E",X"CE",X"C9",X"10",X"8E",
		X"C4",X"1D",X"C6",X"30",X"BD",X"CB",X"A5",X"8D",X"02",X"35",X"B6",X"34",X"36",X"10",X"8E",X"C9",
		X"1F",X"8E",X"B2",X"60",X"C6",X"1E",X"A6",X"A0",X"BD",X"F8",X"35",X"5A",X"26",X"F8",X"35",X"B6",
		X"CD",X"40",X"00",X"01",X"CD",X"4B",X"00",X"05",X"CD",X"58",X"00",X"09",X"CD",X"64",X"00",X"0D",
		X"CD",X"6F",X"00",X"11",X"CD",X"79",X"00",X"15",X"CD",X"84",X"00",X"19",X"CD",X"90",X"00",X"81",
		X"CD",X"A1",X"00",X"85",X"CD",X"B1",X"00",X"87",X"CD",X"C0",X"00",X"89",X"CD",X"CF",X"00",X"8B",
		X"CD",X"E0",X"00",X"8D",X"CD",X"F0",X"00",X"8F",X"CE",X"01",X"00",X"91",X"CE",X"11",X"00",X"93",
		X"CE",X"1F",X"00",X"95",X"CE",X"29",X"00",X"97",X"CE",X"37",X"00",X"99",X"CE",X"45",X"00",X"9B",
		X"CE",X"53",X"00",X"9D",X"CE",X"61",X"00",X"9F",X"CE",X"6F",X"00",X"A1",X"CE",X"7D",X"00",X"A3",
		X"CE",X"8B",X"00",X"A5",X"CE",X"99",X"00",X"A7",X"CE",X"A7",X"00",X"A9",X"CE",X"B6",X"00",X"7D",
		X"43",X"4F",X"49",X"4E",X"53",X"20",X"4C",X"45",X"46",X"54",X"2F",X"43",X"4F",X"49",X"4E",X"53",
		X"20",X"43",X"45",X"4E",X"54",X"45",X"52",X"2F",X"43",X"4F",X"49",X"4E",X"53",X"20",X"52",X"49",
		X"47",X"48",X"54",X"2F",X"54",X"4F",X"54",X"41",X"4C",X"20",X"50",X"41",X"49",X"44",X"2F",X"53",
		X"48",X"49",X"50",X"53",X"20",X"57",X"4F",X"4E",X"2F",X"54",X"4F",X"54",X"41",X"4C",X"20",X"54",
		X"49",X"4D",X"45",X"2F",X"54",X"4F",X"54",X"41",X"4C",X"20",X"53",X"48",X"49",X"50",X"53",X"2F",
		X"42",X"4F",X"4E",X"55",X"53",X"20",X"53",X"48",X"49",X"50",X"20",X"4C",X"45",X"56",X"45",X"4C",
		X"2F",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",X"20",X"53",X"48",X"49",X"50",X"53",
		X"2F",X"43",X"4F",X"49",X"4E",X"41",X"47",X"45",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"2F",
		X"4C",X"45",X"46",X"54",X"20",X"43",X"4F",X"49",X"4E",X"20",X"4D",X"55",X"4C",X"54",X"2F",X"43",
		X"45",X"4E",X"54",X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",X"20",X"4D",X"55",X"4C",X"54",X"2F",
		X"52",X"49",X"47",X"48",X"54",X"20",X"43",X"4F",X"49",X"4E",X"20",X"4D",X"55",X"4C",X"54",X"2F",
		X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",X"4F",X"52",X"20",X"43",X"52",X"45",X"44",X"49",X"54",
		X"2F",X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",X"4F",X"52",X"20",X"42",X"4F",X"4E",X"55",X"53",
		X"2F",X"4D",X"49",X"4E",X"49",X"4D",X"55",X"4D",X"20",X"43",X"4F",X"49",X"4E",X"53",X"2F",X"46",
		X"52",X"45",X"45",X"20",X"50",X"4C",X"41",X"59",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",
		X"4A",X"55",X"53",X"54",X"20",X"31",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",
		X"53",X"54",X"20",X"32",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",
		X"20",X"33",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"34",
		X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"35",X"2F",X"47",
		X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"36",X"2F",X"47",X"41",X"4D",
		X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"37",X"2F",X"47",X"41",X"4D",X"45",X"20",
		X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"38",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",
		X"4A",X"55",X"53",X"54",X"20",X"39",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",
		X"53",X"54",X"20",X"31",X"30",X"2F",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"46",X"55",
		X"4E",X"43",X"54",X"49",X"4F",X"4E",X"2F",X"FF",X"FF",X"02",X"00",X"00",X"44",X"52",X"4A",X"01",
		X"80",X"00",X"53",X"43",X"44",X"01",X"60",X"00",X"4C",X"45",X"44",X"01",X"40",X"00",X"50",X"47",
		X"44",X"01",X"20",X"00",X"43",X"52",X"42",X"01",X"00",X"00",X"4D",X"52",X"53",X"00",X"80",X"00",
		X"4B",X"4A",X"46",X"00",X"60",X"00",X"54",X"4D",X"48",X"00",X"5A",X"01",X"00",X"03",X"03",X"01",
		X"04",X"01",X"01",X"00",X"00",X"00",X"00",X"10",X"01",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"01",
		X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",X"01",X"02",X"00",X"00",X"01",X"00",
		X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"01",X"00",X"02",X"02",X"00",X"00",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"30",X"20",X"2D",
		X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",
		X"4F",X"4E",X"49",X"43",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C0",X"11",X"7E",X"C1",X"70",X"7E",X"C2",X"5E",X"7E",X"C1",X"7E",X"C4",X"4C",X"7E",X"C5",
		X"CC",X"DC",X"20",X"C4",X"E0",X"DD",X"17",X"C3",X"26",X"10",X"DD",X"15",X"0F",X"0F",X"BD",X"CA",
		X"50",X"9F",X"09",X"BD",X"CC",X"00",X"12",X"BD",X"C2",X"A6",X"8E",X"00",X"10",X"9C",X"15",X"27",
		X"12",X"96",X"0D",X"2A",X"04",X"0A",X"11",X"20",X"02",X"0C",X"11",X"BD",X"C2",X"A6",X"30",X"88",
		X"20",X"20",X"EA",X"DC",X"09",X"DD",X"03",X"96",X"0F",X"97",X"00",X"96",X"0D",X"97",X"01",X"96",
		X"11",X"97",X"02",X"8E",X"B7",X"00",X"9F",X"05",X"8E",X"B9",X"60",X"9F",X"07",X"DC",X"15",X"83",
		X"00",X"20",X"DD",X"15",X"10",X"93",X"17",X"2B",X"05",X"BD",X"C1",X"C9",X"20",X"EF",X"DC",X"03",
		X"DD",X"0B",X"96",X"00",X"97",X"10",X"96",X"01",X"97",X"0E",X"96",X"02",X"97",X"12",X"10",X"8E",
		X"BC",X"00",X"8E",X"00",X"00",X"AF",X"A1",X"10",X"8C",X"BF",X"50",X"26",X"F8",X"39",X"DC",X"20",
		X"C4",X"E0",X"93",X"15",X"58",X"49",X"58",X"49",X"58",X"49",X"97",X"00",X"27",X"20",X"2B",X"10",
		X"DC",X"15",X"C3",X"00",X"20",X"DD",X"15",X"BD",X"C1",X"C9",X"0A",X"00",X"26",X"F2",X"20",X"0E",
		X"DC",X"15",X"83",X"00",X"20",X"DD",X"15",X"BD",X"C1",X"C9",X"0C",X"00",X"26",X"F2",X"DC",X"20",
		X"C4",X"E0",X"DD",X"15",X"8E",X"00",X"00",X"10",X"8E",X"BC",X"F0",X"10",X"DF",X"13",X"10",X"DE",
		X"05",X"C5",X"20",X"26",X"03",X"10",X"DE",X"07",X"DE",X"1E",X"12",X"86",X"98",X"AF",X"B4",X"35",
		X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",
		X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",
		X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"4A",
		X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",
		X"4A",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",
		X"B1",X"4A",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",X"A4",
		X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",X"ED",
		X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"04",X"ED",X"A4",X"EF",X"B1",X"AF",X"B4",X"35",X"04",
		X"ED",X"A4",X"EF",X"B1",X"4A",X"10",X"26",X"FF",X"74",X"10",X"DE",X"13",X"39",X"11",X"CC",X"77",
		X"7C",X"BC",X"00",X"B6",X"BC",X"00",X"85",X"01",X"27",X"03",X"7E",X"C0",X"8E",X"39",X"8E",X"00",
		X"00",X"10",X"8E",X"BC",X"F0",X"AF",X"B4",X"AF",X"A1",X"10",X"8C",X"BF",X"50",X"26",X"F6",X"10",
		X"8E",X"B0",X"FD",X"86",X"40",X"AF",X"B4",X"EE",X"A1",X"33",X"C8",X"ED",X"AF",X"C4",X"4A",X"26",
		X"F4",X"86",X"FF",X"97",X"1A",X"39",X"05",X"39",X"96",X"11",X"A7",X"84",X"A7",X"89",X"01",X"C8",
		X"4C",X"97",X"11",X"CC",X"77",X"77",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"30",X"03",X"8C",X"B8",
		X"C8",X"26",X"03",X"8E",X"B7",X"00",X"9F",X"05",X"39",X"96",X"0D",X"2A",X"04",X"0A",X"11",X"20",
		X"02",X"0C",X"11",X"BD",X"C2",X"A6",X"86",X"20",X"95",X"16",X"27",X"41",X"9E",X"07",X"30",X"1E",
		X"8C",X"B9",X"5E",X"26",X"03",X"8E",X"BA",X"8E",X"9F",X"07",X"96",X"0E",X"2A",X"17",X"0A",X"12",
		X"96",X"12",X"A7",X"80",X"A7",X"89",X"01",X"2F",X"90",X"1A",X"A7",X"84",X"A7",X"89",X"01",X"30",
		X"7E",X"C2",X"CC",X"12",X"12",X"96",X"12",X"A7",X"80",X"A7",X"89",X"01",X"2F",X"4C",X"97",X"12",
		X"90",X"1A",X"A7",X"84",X"A7",X"89",X"01",X"30",X"7E",X"C2",X"CC",X"12",X"12",X"9E",X"05",X"30",
		X"1E",X"8C",X"B6",X"FE",X"26",X"03",X"8E",X"B8",X"2E",X"9F",X"05",X"96",X"0E",X"2A",X"17",X"0A",
		X"12",X"96",X"12",X"A7",X"80",X"A7",X"89",X"01",X"2F",X"90",X"1A",X"A7",X"84",X"A7",X"89",X"01",
		X"30",X"7E",X"C2",X"CC",X"12",X"12",X"96",X"12",X"A7",X"80",X"A7",X"89",X"01",X"2F",X"4C",X"97",
		X"12",X"90",X"1A",X"A7",X"84",X"A7",X"89",X"01",X"30",X"20",X"71",X"12",X"12",X"12",X"BD",X"CA",
		X"79",X"9F",X"0B",X"A6",X"84",X"97",X"0E",X"86",X"07",X"97",X"10",X"BD",X"CC",X"05",X"12",X"8E",
		X"B3",X"00",X"96",X"12",X"A7",X"80",X"96",X"0E",X"2A",X"04",X"0A",X"12",X"20",X"02",X"0C",X"12",
		X"BD",X"C2",X"CC",X"96",X"0E",X"2A",X"04",X"0A",X"12",X"20",X"02",X"0C",X"12",X"BD",X"C2",X"CC",
		X"8C",X"B7",X"00",X"26",X"DD",X"39",X"8E",X"00",X"00",X"10",X"8E",X"BC",X"F0",X"AF",X"B1",X"10",
		X"8C",X"BF",X"50",X"26",X"F8",X"39",X"96",X"0F",X"27",X"0A",X"0A",X"0F",X"96",X"0D",X"48",X"89",
		X"00",X"97",X"0D",X"39",X"DE",X"09",X"33",X"41",X"BD",X"CA",X"5E",X"12",X"12",X"12",X"12",X"12",
		X"12",X"DF",X"09",X"86",X"07",X"97",X"0F",X"A6",X"C4",X"97",X"0D",X"39",X"96",X"10",X"27",X"0A",
		X"0A",X"10",X"96",X"0E",X"48",X"89",X"00",X"97",X"0E",X"39",X"DE",X"0B",X"33",X"41",X"BD",X"CA",
		X"5E",X"12",X"12",X"12",X"12",X"12",X"12",X"DF",X"0B",X"86",X"07",X"97",X"10",X"A6",X"C4",X"97",
		X"0E",X"39",X"96",X"0F",X"81",X"07",X"27",X"0C",X"0C",X"0F",X"96",X"0D",X"44",X"24",X"02",X"8B",
		X"80",X"97",X"0D",X"39",X"DE",X"09",X"11",X"83",X"C3",X"4C",X"26",X"03",X"CE",X"C4",X"4C",X"33",
		X"5F",X"DF",X"09",X"0F",X"0F",X"A6",X"C4",X"44",X"24",X"02",X"8B",X"80",X"97",X"0D",X"39",X"96",
		X"10",X"81",X"07",X"27",X"0C",X"0C",X"10",X"96",X"0E",X"44",X"24",X"02",X"8B",X"80",X"97",X"0E",
		X"39",X"DE",X"0B",X"11",X"83",X"C3",X"4C",X"26",X"03",X"CE",X"C4",X"4C",X"33",X"5F",X"DF",X"0B",
		X"0F",X"10",X"A6",X"C4",X"44",X"24",X"02",X"8B",X"80",X"97",X"0E",X"39",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"6B",X"6D",X"DD",X"DD",X"EF",X"7D",X"F7",X"EF",X"77",X"6D",X"55",X"55",X"55",X"2A",X"54",X"A5",
		X"24",X"91",X"22",X"21",X"08",X"20",X"81",X"02",X"4A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"6E",X"EE",X"EE",X"EE",X"ED",X"B6",X"D4",X"92",
		X"49",X"10",X"84",X"44",X"49",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"DB",X"77",X"7F",X"EA",X"AA",X"EA",X"BA",X"FF",X"D5",X"54",
		X"0A",X"00",X"02",X"A0",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"B6",X"AD",X"AB",X"AE",X"EF",
		X"7B",X"DF",X"7E",X"FF",X"FF",X"EE",X"EA",X"A9",X"10",X"80",X"50",X"11",X"88",X"88",X"88",X"89",
		X"54",X"44",X"44",X"91",X"24",X"AA",X"AA",X"AA",X"AF",X"FF",X"F0",X"0F",X"FF",X"FF",X"FF",X"F0",
		X"00",X"1F",X"FF",X"FF",X"F0",X"00",X"00",X"AA",X"80",X"00",X"55",X"55",X"55",X"00",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AD",X"DE",X"FB",X"FB",X"FD",X"FF",X"7F",
		X"D5",X"00",X"02",X"AB",X"FF",X"55",X"00",X"2A",X"AF",X"FF",X"FF",X"F5",X"22",X"10",X"40",X"80",
		X"80",X"40",X"10",X"02",X"24",X"AD",X"B7",X"77",X"BD",X"F7",X"DF",X"BF",X"7F",X"7F",X"7F",X"55",
		X"FF",X"D5",X"22",X"10",X"40",X"80",X"81",X"12",X"DD",X"EF",X"BF",X"02",X"08",X"44",X"44",X"44",
		X"49",X"25",X"6D",X"B7",X"77",X"77",X"7B",X"DF",X"7D",X"EF",X"7B",X"BB",X"55",X"22",X"21",X"08",
		X"20",X"81",X"02",X"08",X"20",X"82",X"10",X"88",X"89",X"2A",X"AA",X"AA",X"25",X"70",X"07",X"26",
		X"77",X"00",X"26",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",X"70",X"07",X"24",X"07",
		X"70",X"25",X"70",X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",
		X"21",X"07",X"70",X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",X"26",X"77",X"00",X"26",
		X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"70",
		X"07",X"25",X"77",X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"07",X"70",
		X"23",X"07",X"70",X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",X"23",X"70",X"07",X"25",
		X"70",X"07",X"25",X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",X"77",X"00",X"22",X"07",
		X"70",X"20",X"07",X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",X"07",X"1F",X"70",X"07",
		X"21",X"70",X"07",X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",X"26",X"77",X"00",X"26",
		X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",
		X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",
		X"23",X"70",X"07",X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",X"25",X"70",X"07",X"26",
		X"77",X"00",X"26",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",X"70",X"07",X"24",X"07",
		X"70",X"25",X"70",X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",
		X"21",X"07",X"70",X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",X"26",X"77",X"00",X"26",
		X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"70",
		X"07",X"25",X"77",X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"07",X"70",
		X"23",X"07",X"70",X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",X"23",X"70",X"07",X"25",
		X"70",X"07",X"25",X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",X"77",X"00",X"22",X"07",
		X"70",X"20",X"07",X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",X"07",X"1F",X"70",X"07",
		X"21",X"70",X"07",X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",X"26",X"77",X"00",X"26",
		X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",
		X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",
		X"23",X"70",X"07",X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",X"34",X"76",X"9F",X"00",
		X"BD",X"C6",X"C0",X"DD",X"04",X"CC",X"17",X"32",X"DD",X"06",X"10",X"8E",X"B3",X"00",X"96",X"00",
		X"5F",X"ED",X"22",X"96",X"01",X"ED",X"24",X"96",X"05",X"44",X"98",X"05",X"44",X"44",X"06",X"04",
		X"06",X"05",X"96",X"04",X"84",X"01",X"80",X"01",X"D6",X"05",X"ED",X"26",X"2A",X"02",X"43",X"53",
		X"34",X"06",X"96",X"07",X"44",X"98",X"07",X"44",X"44",X"06",X"06",X"06",X"07",X"96",X"06",X"84",
		X"03",X"80",X"02",X"D6",X"07",X"ED",X"28",X"2A",X"02",X"43",X"53",X"44",X"56",X"E3",X"E1",X"10",
		X"83",X"01",X"6A",X"24",X"B9",X"8E",X"00",X"00",X"AF",X"A4",X"31",X"2A",X"10",X"8C",X"B8",X"00",
		X"26",X"AC",X"8E",X"C6",X"9C",X"9F",X"02",X"86",X"38",X"97",X"01",X"8E",X"00",X"00",X"10",X"8E",
		X"B3",X"00",X"A6",X"9F",X"A0",X"02",X"97",X"31",X"27",X"50",X"EE",X"A4",X"AF",X"C4",X"AF",X"C9",
		X"01",X"00",X"EC",X"28",X"E3",X"24",X"81",X"2A",X"25",X"28",X"ED",X"24",X"A7",X"21",X"EC",X"26",
		X"E3",X"22",X"81",X"98",X"22",X"1C",X"ED",X"22",X"A7",X"A4",X"5D",X"2B",X"07",X"10",X"AF",X"B4",
		X"12",X"12",X"20",X"0E",X"EE",X"A4",X"CC",X"00",X"7F",X"83",X"00",X"01",X"26",X"FB",X"12",X"12",
		X"12",X"12",X"31",X"2A",X"10",X"8C",X"B8",X"00",X"26",X"C0",X"0A",X"01",X"26",X"B0",X"DE",X"02",
		X"33",X"41",X"DF",X"02",X"86",X"04",X"97",X"01",X"20",X"A4",X"20",X"14",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"86",X"81",X"97",X"33",X"86",X"81",X"97",X"34",X"86",X"2F",X"97",X"35",X"35",X"F6",X"FF",X"FF",
		X"CC",X"00",X"01",X"FD",X"BC",X"10",X"86",X"00",X"B7",X"BC",X"12",X"CC",X"08",X"08",X"39",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B6",X"A1",X"80",X"85",X"01",X"27",X"0A",X"85",X"02",X"26",X"1D",X"85",X"04",X"26",X"30",X"20",
		X"40",X"8A",X"01",X"B7",X"A1",X"80",X"86",X"01",X"B7",X"A1",X"81",X"CC",X"00",X"BF",X"FD",X"A1",
		X"83",X"86",X"00",X"B7",X"A1",X"82",X"20",X"29",X"84",X"FD",X"B7",X"A1",X"80",X"86",X"02",X"B7",
		X"A1",X"81",X"CC",X"00",X"7F",X"FD",X"A1",X"83",X"86",X"00",X"B7",X"A1",X"82",X"20",X"12",X"84",
		X"FB",X"B7",X"A1",X"80",X"86",X"03",X"B7",X"A1",X"81",X"96",X"D5",X"B7",X"A1",X"87",X"7F",X"A1",
		X"7F",X"B6",X"A1",X"81",X"4A",X"48",X"8E",X"C8",X"5B",X"6E",X"96",X"C8",X"61",X"C8",X"B0",X"C8",
		X"F6",X"AE",X"47",X"D6",X"CA",X"10",X"9E",X"B7",X"10",X"AC",X"0A",X"2C",X"01",X"50",X"1D",X"ED",
		X"0E",X"7C",X"A1",X"7E",X"26",X"03",X"7C",X"A1",X"7D",X"B6",X"A1",X"7D",X"81",X"80",X"25",X"17",
		X"F6",X"A1",X"7E",X"C4",X"07",X"96",X"B7",X"5D",X"27",X"04",X"46",X"5A",X"20",X"F9",X"84",X"7F",
		X"6D",X"0E",X"27",X"01",X"43",X"A7",X"0F",X"DC",X"B7",X"84",X"01",X"C5",X"01",X"27",X"01",X"43",
		X"ED",X"88",X"10",X"8D",X"43",X"26",X"08",X"B6",X"A1",X"80",X"8A",X"02",X"B7",X"A1",X"80",X"39",
		X"AE",X"47",X"D6",X"CA",X"10",X"9E",X"A4",X"31",X"A9",X"10",X"00",X"10",X"AC",X"0A",X"2C",X"01",
		X"50",X"1D",X"ED",X"0E",X"96",X"98",X"A1",X"0C",X"DC",X"C8",X"24",X"02",X"43",X"53",X"ED",X"88",
		X"10",X"96",X"D5",X"B1",X"A1",X"87",X"12",X"12",X"B7",X"A1",X"87",X"8D",X"0B",X"26",X"08",X"B6",
		X"A1",X"80",X"8A",X"04",X"B7",X"A1",X"80",X"39",X"7E",X"C9",X"80",X"26",X"08",X"7A",X"A1",X"83",
		X"26",X"03",X"39",X"A1",X"82",X"39",X"7D",X"A1",X"7F",X"26",X"3C",X"AE",X"47",X"10",X"BE",X"A1",
		X"85",X"10",X"8C",X"C9",X"44",X"25",X"06",X"10",X"8C",X"C9",X"6C",X"25",X"04",X"10",X"8E",X"C9",
		X"44",X"7D",X"A1",X"87",X"27",X"0F",X"EC",X"A1",X"ED",X"0E",X"EC",X"A1",X"ED",X"88",X"10",X"BD",
		X"C9",X"70",X"12",X"20",X"1E",X"86",X"01",X"B7",X"A1",X"7F",X"CC",X"00",X"2F",X"FD",X"A1",X"83",
		X"86",X"00",X"B7",X"A1",X"82",X"20",X"0C",X"8D",X"AF",X"26",X"08",X"B6",X"A1",X"80",X"84",X"FE",
		X"B7",X"A1",X"80",X"39",X"00",X"00",X"FE",X"00",X"00",X"40",X"FE",X"00",X"00",X"40",X"00",X"00",
		X"00",X"40",X"02",X"00",X"00",X"00",X"02",X"00",X"FF",X"C0",X"02",X"00",X"FF",X"C0",X"00",X"00",
		X"FF",X"C0",X"FE",X"00",X"FF",X"E0",X"FE",X"00",X"FF",X"E0",X"02",X"00",X"FF",X"FF",X"FF",X"FF",
		X"10",X"BF",X"A1",X"85",X"7A",X"A1",X"87",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7D",X"A1",X"84",X"26",X"10",X"7D",X"A1",X"83",X"26",X"08",X"7D",X"A1",X"82",X"27",X"0C",X"7A",
		X"A1",X"82",X"7A",X"A1",X"83",X"7A",X"A1",X"84",X"86",X"01",X"39",X"4F",X"39",X"FF",X"FF",X"FF",
		X"34",X"06",X"97",X"51",X"FC",X"A1",X"88",X"26",X"03",X"CC",X"C9",X"F1",X"10",X"83",X"CA",X"41",
		X"25",X"03",X"CC",X"C9",X"F1",X"FD",X"A1",X"88",X"BD",X"D0",X"96",X"EE",X"0B",X"EE",X"4D",X"66",
		X"66",X"34",X"20",X"10",X"BE",X"A1",X"88",X"EC",X"A1",X"ED",X"0A",X"EC",X"A1",X"ED",X"0C",X"EC",
		X"A1",X"ED",X"0E",X"EC",X"A1",X"ED",X"88",X"10",X"10",X"BF",X"A1",X"88",X"35",X"20",X"86",X"10",
		X"A7",X"88",X"14",X"4F",X"5F",X"ED",X"06",X"9F",X"42",X"AF",X"A1",X"0A",X"51",X"26",X"B5",X"35",
		X"86",X"54",X"00",X"70",X"00",X"FF",X"40",X"FF",X"F1",X"52",X"00",X"80",X"00",X"FF",X"40",X"FF",
		X"F1",X"50",X"00",X"90",X"00",X"FF",X"40",X"FF",X"F1",X"52",X"00",X"A0",X"00",X"FF",X"40",X"FF",
		X"F1",X"54",X"00",X"B0",X"00",X"FF",X"40",X"FF",X"F1",X"A0",X"00",X"40",X"00",X"FF",X"48",X"FF",
		X"01",X"A0",X"00",X"60",X"00",X"FF",X"20",X"01",X"01",X"A0",X"00",X"80",X"00",X"FF",X"10",X"FF",
		X"21",X"A0",X"00",X"A0",X"00",X"FF",X"50",X"00",X"E1",X"A0",X"00",X"C0",X"00",X"FF",X"54",X"00",
		X"A1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B6",X"A1",X"8A",X"8E",X"C3",X"4B",X"84",X"01",X"27",X"03",X"8E",X"CA",X"9B",X"39",X"B6",X"A1",
		X"8A",X"84",X"01",X"26",X"0A",X"11",X"83",X"C4",X"4C",X"26",X"03",X"CE",X"C3",X"4C",X"39",X"11",
		X"83",X"CB",X"9C",X"26",X"03",X"CE",X"CA",X"9C",X"39",X"B6",X"A1",X"8A",X"8E",X"C3",X"4C",X"84",
		X"01",X"27",X"03",X"8E",X"CA",X"9C",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"B6",X"DD",X"EF",X"F0",
		X"08",X"44",X"92",X"B6",X"DB",X"BB",X"DD",X"A4",X"42",X"22",X"49",X"2A",X"FF",X"FF",X"FF",X"FF",
		X"34",X"06",X"5F",X"BD",X"CB",X"D0",X"81",X"01",X"27",X"0E",X"81",X"05",X"27",X"0A",X"81",X"02",
		X"27",X"0A",X"81",X"06",X"27",X"06",X"20",X"06",X"CA",X"01",X"20",X"02",X"CA",X"02",X"F7",X"A1",
		X"8A",X"35",X"86",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"34",X"10",X"BD",X"D7",X"DC",X"9F",X"6A",X"A6",X"08",X"4A",X"84",X"07",X"35",X"90",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8D",X"08",X"97",X"11",X"39",X"8D",X"03",X"97",X"12",X"39",X"34",X"10",X"8E",X"CC",X"16",X"BD",
		X"F6",X"F5",X"A6",X"86",X"35",X"90",X"F0",X"98",X"E0",X"F0",X"E0",X"98",X"D0",X"F0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
