-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_PGM_1 is

	signal rom_addr : std_logic_vector(13 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(13 downto 0) <= ADDR;
	end process;

	ROM_PGM_1_0 : RAMB16_S1
	generic map (
		INIT_00 => x"747FB557CE90AA7D9D20080F7756C943A329C1212E6D756C94766C3D6F322F1D",
		INIT_01 => x"E6DE95137F7BF7BEE4920E855FF0369DBB76ED818181010808090951A39DD1FF",
		INIT_02 => x"DDF8C5DBD9BF8C7FA53657ED635B97F6BEB10FD0EEBD818BEB7E7CFA947E8007",
		INIT_03 => x"F25AA23BEFA7FA8DBB6DA77F9CE3177FC99818726465F3030E4C0C3EFAF65ECB",
		INIT_04 => x"D885B7225DB8F69877237180261C7B5D998038A0F64366CD9B37A183F26887E7",
		INIT_05 => x"EDDB1D3ED51E27B31D15E8D7A35BA6E5EB96C2E6B2912BD9AEC33310B6216C42",
		INIT_06 => x"6F61016CD9D3A474732FBED8FDB7D63755B3D90CE5308E90928402C6C6EFA2B6",
		INIT_07 => x"76EDDBDBB76F6EDDBDBB76EABAA5114C13A510F64888F65BB76EDDBCDA6B18E3",
		INIT_08 => x"ADCEDEC6BAE5D72F118E71ACCDF9C8A1CE3C99AC796E3CA11E58877287CFEDC6",
		INIT_09 => x"8CC56A3AD9FA43A8F62073A660063FDA8B42B0DD65BC68237DFD9CC3C76777B2",
		INIT_0A => x"3E945A1401D35877601C9D263FDA8B42B8F6D479A1D01A8BA548CD42B8ED9D12",
		INIT_0B => x"0DC436F9F2EF5AD27C387A974C558BEE9757A17E5F8E7BDA6D369D361507BA8B",
		INIT_0C => x"FFFFFFFFFFFFFFFFFFFFFFFFD55E2A2DDBB76EE21B7A0A9EF256F7C45C6C371B",
		INIT_0D => x"2946294629462946294629462946294629462946294629462946294629462946",
		INIT_0E => x"2946294629462946294629462946294629462946294629462946294629462946",
		INIT_0F => x"2946294629462946294629462946294629462946294629462946294629462946",
		INIT_10 => x"15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4",
		INIT_11 => x"15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4",
		INIT_12 => x"15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4",
		INIT_13 => x"15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4",
		INIT_14 => x"2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC",
		INIT_15 => x"2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC",
		INIT_16 => x"2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC",
		INIT_17 => x"2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC",
		INIT_18 => x"7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E",
		INIT_19 => x"7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E",
		INIT_1A => x"7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E",
		INIT_1B => x"7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E",
		INIT_1C => x"074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A",
		INIT_1D => x"074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A",
		INIT_1E => x"074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A",
		INIT_1F => x"074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A",
		INIT_20 => x"00081182008826000000110001080A000104080000800A000000000000000100",
		INIT_21 => x"00C20ACF0000154F40A84A9C0088153301000A4F00980937818018D000802A3C",
		INIT_22 => x"04080947040D0A9D05800D1B00400AB728220C2C001A295838300E70000809A3",
		INIT_23 => x"07E1F84007E1F82000000A0201000C0006000A00040105000100002704010E0F",
		INIT_24 => x"DE06DDBB400F3FFC000060BFFD03FFEE1CC03FFFFFFFFFFFFFFF185E15800000",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE000000000003FFFFC7401F7063803CDF",
		INIT_26 => x"FFFFF1800000FF87FC80003FEFC4FFFC00003FFFFF7FF5FFFFFFFFDFF8000000",
		INIT_27 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAF80000000038001FFCF7FFFFFFF",
		INIT_28 => x"FFB002100100901042108210810865BFFFEE836B772EFDFBFBF7FFF7FAFFFDFF",
		INIT_29 => x"02AFBEFFFFFFFFF7FFFF556AA4914449529A291308445E56F7DEFDBAB52A4927",
		INIT_2A => x"5555FEFFFFFFFFC00020000DFFFFFA6EFE2001C0049800000600001F54FFFF72",
		INIT_2B => x"BDEFDEF78F7BDFBFBFBEFEFBEF7DEFDFEFF7FFBD9D2A949C924889042108410B",
		INIT_2C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9B",
		INIT_2D => x"AAAAAAAA9010040200001008AFFF91BA13BB8ED0ACAB7636D2AD0A8AEEFDF7DF",
		INIT_2E => x"FFFDFFEFFFFDFFF7BDAA0880495B7FBFFFFFFFFFFFFFFDF775EFEFEFBFFFFBFF",
		INIT_2F => x"3AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9FCFE",
		INIT_30 => x"7E154327FFFFFFFFFFFFFFFDAAABFFFDAAAB6A0BFFF81A00FFFA1220FFF09220",
		INIT_31 => x"C443903BFE50104BFFFFFF91111111111111111111111139FFFFFFF940401591",
		INIT_32 => x"FFFFFFFF341041313041043331041031FFFFFFE0001BFF80049BFFFFFE111111",
		INIT_33 => x"EC60606060726243FFFE44444449FFB0808080828080804BFFF8001BFFFFFFFF",
		INIT_34 => x"FFFFFFF9100000E1FFFFFFF8411111E1FFFFFFFFAD5555E14C0000E30C0000E3",
		INIT_35 => x"555005455154555555540155555005E1FFFFFFFFFFFFFFFFFFFFFFF8011111E1",
		INIT_36 => x"5154555555540155555005E30014451555441515450511455541451555E10015",
		INIT_37 => x"FFFFFFFFE0D54063E0D5406383050461FFFFFFFFFB3FEA41FFFF001555500545",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB054220D905040345157D4B1501540563",
		INIT_39 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC1515151551517440404040404040423",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC1504040540407551514040404040421",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFE4441093FFFFFFFFFFFFFFFFFFF9040410104091",
		INIT_3E => x"6666666666CC150015001500150015E3FFFFFFFFFFFFFFFFFFFFFFFFFE400591",
		INIT_3F => x"4400FFFFFFFFFFFF1504104104104161333333333315400550015000540015E1"
	)
	port map (
		DO   => DATA(0 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_1 : RAMB16_S1
	generic map (
		INIT_00 => x"11422FF95EA65D89264A2223590986655C4295757633909864A98950A2E35B71",
		INIT_01 => x"8A0B2228014113C8018417088B45B9200000000C8C8C0C00000000050A004508",
		INIT_02 => x"10F9133AB29FDA000FC598218A62D818C1C452C5898B352D8040BF7A695256B2",
		INIT_03 => x"4503474013C9A336801004AAE739D7C51452D2A14B4A8A5A5429E9D3BC040180",
		INIT_04 => x"011E080000E21A091001C40000710D048800E222B49B88102040893545219289",
		INIT_05 => x"A34273CA6228D417A46623588D6093160C1830972666922BCD1A2823C047808F",
		INIT_06 => x"40183F1512D819D158C4104BA69101A1980D6C72362138465C32E5989989CCD0",
		INIT_07 => x"90A34242CD898A36262CD0AEDCDE03C60772890A13D080E08102040367B052B0",
		INIT_08 => x"F1FF78EFC09800C376508A09DE1E664A11403BC07FBC3FDA1FED0BBF6207E434",
		INIT_09 => x"15CE0442154D8A1110DAA2D8EDD46104D0642D10494157FEA4C2010A207FDE27",
		INIT_0A => x"53668331696C12810DA916CE6144D0642D0808A6D504A4D0891AB6642D00C034",
		INIT_0B => x"8011B800416318C464E9CC3891996CDA6E7A32EDE49CE044A6D12451972E0112",
		INIT_0C => x"FFFFFFFFFFFFFFFFFFFFFFFFB880867102040808DC04BE25BF981410E4000000",
		INIT_0D => x"44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0",
		INIT_0E => x"44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0",
		INIT_0F => x"44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0",
		INIT_10 => x"89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF",
		INIT_11 => x"89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF",
		INIT_12 => x"89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF",
		INIT_13 => x"89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF",
		INIT_14 => x"9425942594259425942594259425942594259425942594259425942594259425",
		INIT_15 => x"9425942594259425942594259425942594259425942594259425942594259425",
		INIT_16 => x"9425942594259425942594259425942594259425942594259425942594259425",
		INIT_17 => x"9425942594259425942594259425942594259425942594259425942594259425",
		INIT_18 => x"8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95",
		INIT_19 => x"8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95",
		INIT_1A => x"8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95",
		INIT_1B => x"8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95",
		INIT_1C => x"8233823382338233823382338233823382338233823382338233823382338233",
		INIT_1D => x"8233823382338233823382338233823382338233823382338233823382338233",
		INIT_1E => x"8233823382338233823382338233823382338233823382338233823382338233",
		INIT_1F => x"8233823382338233823382338233823382338233823382338233823382338233",
		INIT_20 => x"FF80037CFF0812FFFF8814FFFE8809FFFF800BFF7F040BFF0000000000000100",
		INIT_21 => x"3F30134B7F90598F7F104D5D3EB007B47E1852507F1840477F0050C0FE002104",
		INIT_22 => x"070825D907002013078006872342038F2782011C0FE006380FE825303FF83362",
		INIT_23 => x"08E0E43C0071E01C00000BFC010009F002000DE0000006E2060101E4078103C0",
		INIT_24 => x"DEF6C3293CCC87FA00007EB402BFFDE10245BFFFFFFFFFFFFD004541D5A0007F",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA40000000000040000193FE9001B909C1F",
		INIT_26 => x"FFFFF003F8FE807C607BC23BE002100200003FE80079F1FFFFFFFFDFF800FFFF",
		INIT_27 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA8400000401DA005FFF07FFFF7FF",
		INIT_28 => x"001FFDFEFFFFFFFFFFFFFFFFEFFFBFFD30017EFFFFFFFFFFFFFFF7FFFFFFFFFF",
		INIT_29 => x"F9504000002296BE7DEF7FFFFFFFFFFFFFFFFFFFEFFFF8FFFFFF7FFEDFFFFFFF",
		INIT_2A => x"0000007F9B6DB6FFFFDFFFF3093FFBFFEFFFFFFFFFFFFFFFFFFFFFE300FFFFF7",
		INIT_2B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF3FFFF3FFFFFFFFFFFFFFFF",
		INIT_2C => x"000000000000000000000000000000000000000000000000000000000000003F",
		INIT_2D => x"000000000FFFFFFFFFFFFFFFFBE463FFEC44712F5FFFFF3FFFF3FFFFFFFFFFFF",
		INIT_2E => x"FFFFFFFFFFFFFFFFFFFFFE7FB6A48020AAF77FFFFFEFFFFFFFFFFFFFB7EEFF5B",
		INIT_2F => x"550000000000000000000000000000000000000000000000000000000000003E",
		INIT_30 => x"FFBBAC57FFFFFFFFFFFFFFFD2283FFFD0A234AA3FFFA92A0FFF89280FFF81280",
		INIT_31 => x"AA1FC04DFF90109FFFFFFFD414141414141414141414140DFFFFFFFC2EAEAC6F",
		INIT_32 => x"FFFFFFFF641041476041044561041045FFFFFFF4450DFFD1148DFFFFFF050505",
		INIT_33 => x"F117711771155315FFFF0505051FFFC44CC44CC44CC44C1DFFFC088DFFFFFFFF",
		INIT_34 => x"FFFFFFFDEAAAAA1FFFFFFFFCFAEFFB1FFFFFFFFFBBFFFF17BAAAAA15BAAAAA17",
		INIT_35 => x"451145511B16C50F9144516B45114597FFFFFFFFFFFFFFFFFFFFFFFCAAEFFB1F",
		INIT_36 => x"1B16C50F9144516B45114597047F555145505B56D55FD554517F55514595047E",
		INIT_37 => x"FFFFFFFFF0844095F0844095C24A0097FFFFFFFFFE91041FFFFF047E45114551",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAFEDCE77E62EB9AAABD3A1B8AAE2AB9F",
		INIT_39 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFAAFFBDBBFBDAAABFEAAAAAAAAAA95",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFBBEEADAAEADAAABFEAAAAAAAAAA97",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFF9841065FFFFFFFFFFFFFFFFFFFD041410104067",
		INIT_3E => x"6666666666CC405F555F550A000A0097FFFFFFFFFFFFFFFFFFFFFFFFFF800567",
		INIT_3F => x"0100FFFFFFFFFFFF6836F3CF63A69A97333333333340404F4013D040A0102897"
	)
	port map (
		DO   => DATA(1 downto 1),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_2 : RAMB16_S1
	generic map (
		INIT_00 => x"4933BAA95EF44F4DB52AAAAE0CCCEB69662655656C99CCCEB52CCDC89999EF78",
		INIT_01 => x"1CDC733B2E1486E2418613882618BDB3972E5C880008000E060E0624C91924CE",
		INIT_02 => x"C8D891A02A20171D8A66DDC9E9F35DFCEEF65390CFE5E4AE49EFFD78B324A527",
		INIT_03 => x"AF6B6766FE5E1BBFE259228AA5294A2EBD4BCABD2F2AE97957A5E55C50BAD65A",
		INIT_04 => x"C9CF96198C729F902318E50CC6394FC8118C72F7EDDBDE7CF9F2B887AF79171F",
		INIT_05 => x"4C996CB7B33A1097B73779DDE779E7A74E9E50F7BFF0984BC9E91A39F273E4E7",
		INIT_06 => x"6C2F0A6C18EB4DA3795C71C367D582B5FD17E56A5719B562C51626575665EAE7",
		INIT_07 => x"074C991D326474C991D3267E8EEB102200E1019F587C12B9B366CD9EF7E95AF8",
		INIT_08 => x"5C550009606C0763631CE885131F46639D10A262AFBD57DCABEE177F62000D59",
		INIT_09 => x"BD9F0E6BC496C9399413B16EE9D27D96DB6BB5F77FE52A2229870519F32A8004",
		INIT_0A => x"05B6DB5508B7DADD43258B6EFD96DB6BB5AF9CCB64B476DB7CDA5B6BBDBBFB15",
		INIT_0B => x"BC95BE44715EF7BC01D7B02F19DDCE3EFD7FB4DFF17AD93FDB6DB3CD874D939B",
		INIT_0C => x"FFFFFFFFFFFFFFFFFFFFFFFFBCD4ACFACD9B364ADF2F86B2F7DE5695F1E6F379",
		INIT_0D => x"4000400040004000400040004000400040004000400040004000400040004000",
		INIT_0E => x"4000400040004000400040004000400040004000400040004000400040004000",
		INIT_0F => x"4000400040004000400040004000400040004000400040004000400040004000",
		INIT_10 => x"0736073607360736073607360736073607360736073607360736073607360736",
		INIT_11 => x"0736073607360736073607360736073607360736073607360736073607360736",
		INIT_12 => x"0736073607360736073607360736073607360736073607360736073607360736",
		INIT_13 => x"0736073607360736073607360736073607360736073607360736073607360736",
		INIT_14 => x"34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA",
		INIT_15 => x"34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA",
		INIT_16 => x"34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA",
		INIT_17 => x"34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA",
		INIT_18 => x"3080308030803080308030803080308030803080308030803080308030803080",
		INIT_19 => x"3080308030803080308030803080308030803080308030803080308030803080",
		INIT_1A => x"3080308030803080308030803080308030803080308030803080308030803080",
		INIT_1B => x"3080308030803080308030803080308030803080308030803080308030803080",
		INIT_1C => x"0310031003100310031003100310031003100310031003100310031003100310",
		INIT_1D => x"0310031003100310031003100310031003100310031003100310031003100310",
		INIT_1E => x"0310031003100310031003100310031003100310031003100310031003100310",
		INIT_1F => x"0310031003100310031003100310031003100310031003100310031003100310",
		INIT_20 => x"0008330200083600000814000008080081800800008008000000000000000100",
		INIT_21 => x"0042120800005050000040E3410048C801804DA001804187819843FF00081303",
		INIT_22 => x"040121680085206000882040200A2440206A268110280480102A0600000A3201",
		INIT_23 => x"388003C0300007E000000C0501000E0F05000E1F0200073E0400013C04800278",
		INIT_24 => x"0000004000001002000210000001000200008000000000000000000888000040",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000004080820000001000",
		INIT_26 => x"0012000202025000400000000000000000000080000020000000000000004000",
		INIT_27 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0200000000080000010000000008",
		INIT_28 => x"00104211010010104210A210910865FD10117F9488D102040408080805000203",
		INIT_29 => x"FD524000002296BE7FFFD52AA493444952922913184559AD0821824555AA4927",
		INIT_2A => x"000000004000003FFFDFFFE20937FE6EFE2001C00C980000060000030000008D",
		INIT_2B => x"42102108608420404041010410821020100C00426DEA949C924889C42108410B",
		INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000004",
		INIT_2D => x"000000000010040200001008AFE46245EC44412F535489C92D5EF57511020823",
		INIT_2E => x"00020010000200084255F7FFB6A48020AAF77FFFFFEFFDF775EFEDEFF7FEFF5B",
		INIT_2F => x"0500000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => x"7E015077FFFFFFFFFFFFFFFD2003FFFD00234003FFF89A28FFF89A28FFF89A28",
		INIT_31 => x"40159A4FFE54541FFFFFFF8015400015400015400015400DFFFFFFFBD0505645",
		INIT_32 => x"FFFFFFFF1FBEFB4F1EFBEF4D1BEFBE4DFFFFFFE4E70FFF939C8FFFFFFE005500",
		INIT_33 => x"E511177771333317FFFE0550021DFF94444CCCC6444CCC1DFFF8AA8FFFFFFFFF",
		INIT_34 => x"FFFFFFF95400009FFFFFFFF90114559FFFFFFFFF2555559D4555559D0400009F",
		INIT_35 => x"AFAAAAABA0B82EADABEAAAA2AFAAAA1DFFFFFFFFFFFFFFFFFFFFFFF80114559F",
		INIT_36 => x"A0B82EADABEAAAA2AFAAAA1D0277EABAAFEBE1FC6BBDFAAEABF7EABAAF1D0276",
		INIT_37 => x"FFFFFFFFEA7CEA17EA7CEA17A9B7EA17FFFFFFFFF9015015FFFF0276AFAAAAAB",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB1111555555C44541110000024449111D",
		INIT_39 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC404015155151544040551515151515D",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC515115155151544040440404040405F",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFE44EBF45FFFFFFFFFFFFFFFFFFF9EFA7BE9EFA45",
		INIT_3E => x"6666666666CC3FA03FA03FA03FA03F15FFFFFFFFFFFFFFFFFFFFFFFFFE5AEF47",
		INIT_3F => x"1401FFFFFFFFFFFF17CD1C718C18619733333333333FEEA5FBA97EAA5FAA9715"
	)
	port map (
		DO   => DATA(2 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_3 : RAMB16_S1
	generic map (
		INIT_00 => x"C7D19006F57FEA6671DD00039DFD61B299D7EA9A85E76666F2FF66BC61DAA5B0",
		INIT_01 => x"348D888322BF01257AE9A9C0737303AA97363FAAD5D5AAA85657A8A2C7DFE2E2",
		INIT_02 => x"5BADEB80EF0A09ACFFD967AEA4F5E7A6839B28FA5786838AE783575278F6BBA3",
		INIT_03 => x"D2CEB1AB4B757BA83E793C08ED7BC2864BB5400BD4D42A8AABDA2A0E43F52191",
		INIT_04 => x"CEFE87AAAAB4E2EA3AAA71C488946A60EAEE34A23DDF2E2EFADB27E978668BC5",
		INIT_05 => x"BD7AA9A1B55BC44E5C4C910299484180A9530ABCF6BD1DFB86F7228C91950230",
		INIT_06 => x"DC5B80FA07DBC0E1D30661A86DBCD6367B39B9C8FF5BCF839EB7AB271620BAAF",
		INIT_07 => x"3EBD0686F56B99E2ADAF81BF7BB3AA21077F20AA3C9D86047375FA00FB699A97",
		INIT_08 => x"F8EE8129F554DFF7FF0993CE8B07AAB6C8D3E6352DBA43864B6F522ED6D50A79",
		INIT_09 => x"4F75EEF959F7BABBA52902E8F547238B0DD08EC0F8B4AAAA5AEDFAB2F2A23540",
		INIT_0A => x"97576C8EFFDD6A66FAB6F9FF9E29A9B27A7EE679DB131BA9DDEBF9B27A61A98B",
		INIT_0B => x"BC8F013BAEBD3603977F3ABF1F56466257D6D0A65FEF24AEFF75A820199F4BB8",
		INIT_0C => x"0000555500005555000055557FCD3AAF47FD2E4389906936D9FF69C6F7EEBA39",
		INIT_0D => x"54A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA02",
		INIT_0E => x"7C0028007C0028007C0028007C0028007C0028007C0028007C0028007C002800",
		INIT_0F => x"54A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA02",
		INIT_10 => x"4AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B6",
		INIT_11 => x"4AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E58",
		INIT_12 => x"4AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B6",
		INIT_13 => x"4AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E58",
		INIT_14 => x"6BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB9674",
		INIT_15 => x"6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E",
		INIT_16 => x"6BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB9674",
		INIT_17 => x"6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E",
		INIT_18 => x"2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C",
		INIT_19 => x"2AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB5572",
		INIT_1A => x"2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C",
		INIT_1B => x"2AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB5572",
		INIT_1C => x"522B857C522B857C522B857C522B857C522B857C522B857C522B857C522B857C",
		INIT_1D => x"522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82",
		INIT_1E => x"522B857C522B857C522B857C522B857C522B857C522B857C522B857C522B857C",
		INIT_1F => x"522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82",
		INIT_20 => x"FF77A829FF77A8AAFF77A8AAFF77A0AA7FF3A0AAFF7BA0AAFFFFAAAAFFFFABAA",
		INIT_21 => x"551FA9EE157DABFA157DAA49157DAA66555DAA1A554DAA67554DAB7A55DDAAD6",
		INIT_22 => x"FF73AAFBFFFFAAB8FF7FAAAEFFB7AAA2FF97AAF9DFC7ABEEDFC7ABAAFFE7ABF9",
		INIT_23 => x"5DC48EEA5DC58E8A5555A2AC5555A2AA5555A2BA5555AA895555AA8E55D5AAEA",
		INIT_24 => x"210D5FF561117951FFFFD5F7FEC2555FFFAD55550000555501FFFFFF162FAAD5",
		INIT_25 => x"AAAA5555AAAA5555AAAA5555AAAA55145555AAAA55FF5555FBAA55547EFF5475",
		INIT_26 => x"0000579F0785FFD78B4447D70FFAFFFDFFFFD55FFF8757550000557583DFD555",
		INIT_27 => x"AAAA5555AAAA5555AAAA5555AAAA5555AAAA0555FFFB6AA5FFFC55552AAA5155",
		INIT_28 => x"FFFFEAABFFFFAAAAFFFFAAAAFFFFEAEAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAA",
		INIT_29 => x"5157AAAA5555AAA257552AEA5557BAAA555DAAA85555AAAE5555AAAB5555AAAB",
		INIT_2A => x"FFFFABAABFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAABFFFFAAAA",
		INIT_2B => x"5555AAAA7555AAAA5555AAAA5555AAAA5553AAAA5555AAAE5555AAEA5555AAAB",
		INIT_2C => x"FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAEA",
		INIT_2D => x"5555AAAA5555AAAA5555AAAA5555A2AA7555BAAA5555AAEA5555AABA5555AAAB",
		INIT_2E => x"FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFABAAFFFFAAAB",
		INIT_2F => x"0055AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAB",
		INIT_30 => x"55FF00025555AAAA5555AAA84441AAA851010546555005745550443055504574",
		INIT_31 => x"EAFF2FE255FFFFB25555002AFFFFEABFFFEABFFFAAAAFFE255550003FFFFFEE2",
		INIT_32 => x"5555AAAAFFFF5500FFFE5500FFFA55005555AAA2FFFFAA88FEBFAAAA55AA5555",
		INIT_33 => x"5FBBEEEEBBBB8CBA5555AFFFAAFF002BEEEEBBB3EEEE33B25556BEEA55550000",
		INIT_34 => x"5555AAABAAEB51005555AAAAFEEB51005555AAAA1EFB5100FEFB5100FEFB5100",
		INIT_35 => x"AAAFFABBAEABAEAFAAABFEAAAAAFFABA555500005555000055550001AAEBFFBA",
		INIT_36 => x"AEAB5555AAAB0155AAAF0500AFEA5555AAAA5555AAAA5555AAAA5555AAFF5015",
		INIT_37 => x"555500005FFFFFB25FFFFFB26BAAFBB25555000057FFFFB25555FAFEAAAFFABB",
		INIT_38 => x"5555AAAA5555AAAA5555AAAA5555AAAAFFFF0000FFFF0000FFFF1440FFFF0000",
		INIT_39 => x"555500005555000055550000555500007FBFAFFFBFFBFFBFBBBBFBFBBBBBFBFA",
		INIT_3A => x"5555AAAA5555AAAA5555AAAA5555AAAA7BBB4444BFBB4415AAAB4444BBBB4440",
		INIT_3B => x"5555000055550000555500005555000055550000555500005555000055550000",
		INIT_3C => x"5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA",
		INIT_3D => x"5555000055550000555500005FFBFFE255550000555500005557EFEFFFEBFFE2",
		INIT_3E => x"CCCC3333CC661455AAAAD555AAAAD5085555AAAA5555AAAA5555AAAA55FF0508",
		INIT_3F => x"FEAB000055550000EBAAFFFFAAAAFFB29999CCCC99EBEEEFAEEEFEEEAAEEBFB2"
	)
	port map (
		DO   => DATA(3 downto 3),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_4 : RAMB16_S1
	generic map (
		INIT_00 => x"B9B8FA8450310E01064088882CCCCB446608413130D9CCCCB08CC80E1C116C08",
		INIT_01 => x"2D41B77C2B60B8E4575F73BA80649C90102040848484040606060602855AE6E2",
		INIT_02 => x"30D6182522A0121548081D51C5741D5CEAE777A610F1E2E69B6AC08524A135E0",
		INIT_03 => x"1790646C58AC81DB601001FC11846A805E2BAB80AEAE05757015D5C0104DC9B9",
		INIT_04 => x"898F18BB99CF1DB367339E5DCCE78ED9B399CF0006E9C0408102181417BD702C",
		INIT_05 => x"12246A03C3305B547777FB9FEE71FCE7CFDC5301C3A2BD8AABA50C31E263C4C7",
		INIT_06 => x"404A0410810451A082504903500B64A0A624321307013543721B91018191E4E9",
		INIT_07 => x"0912242408101120404089104EECF6FDFD8C6400514514C142850A1427D26124",
		INIT_08 => x"53772B1D4C82641072DEF941128F0C5BDF2922532C459620CB10699884371522",
		INIT_09 => x"58AA066848824919C25380260A934D961B45B5D385C12022861B6CA902BB8ACD",
		INIT_0A => x"6090DA233812DACC250781214D961B45B58D8CC130A4121B0A304905B59ADB00",
		INIT_0B => x"509A9C59155294A48250A64009DC6E5CF51F825EF04AD10B45A2D041242D1198",
		INIT_0C => x"FFFFFFFFFFFFFFFFFFFFFFFF9CCBC4780810204D4E2014A8CFDC557AF68742A1",
		INIT_0D => x"11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE",
		INIT_0E => x"11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE",
		INIT_0F => x"11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE",
		INIT_10 => x"8811881188118811881188118811881188118811881188118811881188118811",
		INIT_11 => x"8811881188118811881188118811881188118811881188118811881188118811",
		INIT_12 => x"8811881188118811881188118811881188118811881188118811881188118811",
		INIT_13 => x"8811881188118811881188118811881188118811881188118811881188118811",
		INIT_14 => x"849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F",
		INIT_15 => x"849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F",
		INIT_16 => x"849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F",
		INIT_17 => x"849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F",
		INIT_18 => x"9011901190119011901190119011901190119011901190119011901190119011",
		INIT_19 => x"9011901190119011901190119011901190119011901190119011901190119011",
		INIT_1A => x"9011901190119011901190119011901190119011901190119011901190119011",
		INIT_1B => x"9011901190119011901190119011901190119011901190119011901190119011",
		INIT_1C => x"8003800380038003800380038003800380038003800380038003800380038003",
		INIT_1D => x"8003800380038003800380038003800380038003800380038003800380038003",
		INIT_1E => x"8003800380038003800380038003800380038003800380038003800380038003",
		INIT_1F => x"8003800380038003800380038003800380038003800380038003800380038003",
		INIT_20 => x"0000600300086500000005000100080000080900010008000000000000000000",
		INIT_21 => x"00422240002044C0002044C3002004880000042000100087001000E001006040",
		INIT_22 => x"0401060104050282048A06A4244206A8286206D318302560182227A0001207C3",
		INIT_23 => x"001104000000000000000A0600000A0006010A00020102000401040404812600",
		INIT_24 => x"DF03FD9BE00F5BF80000705DFEC3FFF61E503FFFFFFFFFFFFF7F585F0BC00000",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE000000000001FFFFC3801F70F100AC7F",
		INIT_26 => x"FFFFF98000047FC5F800083DF7E6F7FC00003FFFFF7EFFFFFFFFFFDF7C200000",
		INIT_27 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFC0000400038003FFCFFFFFFBFF",
		INIT_28 => x"0008000000000000000020000000010020100100001000000000000000000001",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => x"0000000010000000000000000400100020002000080000800008002000000002",
		INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => x"FF400157FFFFFFFFFFFFFFFFAEABFFFFBAABEEFBFFFABAAAFFFAFAAAFFFABAAA",
		INIT_31 => x"5555F455FF400055FFFFFFD5555540000015555540000015FFFFFFFD00000055",
		INIT_32 => x"FFFFFFFF554054555501505554054055FFFFFFF44555FFD55515FFFFFF000000",
		INIT_33 => x"F511111111111555FFFF55555055FFD44444444444444455FFFC4555FFFFFFFF",
		INIT_34 => x"FFFFFFFD54410455FFFFFFFC01145155FFFFFFFF350451555504515555045155",
		INIT_35 => x"55500555515455555554015555500555FFFFFFFFFFFFFFFFFFFFFFFC01145155",
		INIT_36 => x"5154555555540155555005550555505555555555515554155555505555550555",
		INIT_37 => x"FFFFFFFFF5400455F5400455D5555555FFFFFFFFFD400055FFFF055555500555",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF50155555551155555555411455515555",
		INIT_39 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0404040540405444444444444444455",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4040404144041511110000000000015",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFF7651555FFFFFFFFFFFFFFFFFFFF555840355555",
		INIT_3E => x"6666666666CC41554055405540554055FFFFFFFFFFFFFFFFFFFFFFFFFF610555",
		INIT_3F => x"5501FFFFFFFFFFFF410000000000005533333333334111100444011100444055"
	)
	port map (
		DO   => DATA(4 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_5 : RAMB16_S1
	generic map (
		INIT_00 => x"B52ED2AC54C53AF5EE37F7F2131355D7FE39D1216BF975754B3174FF3EE476E5",
		INIT_01 => x"3971F77141DFE31AB1C7645FFC255C776051D455575755545555557D543C3D45",
		INIT_02 => x"9C59C8C058555F2C822B954D164E1557EBF15D77B9F9939B9C6B682CE3B9C593",
		INIT_03 => x"5590151514B984574D345001D4B57FF55601959806077D4D1DB03500548DCEC5",
		INIT_04 => x"9FDCDBDD0067F69591FFFBD55DEDF97537443AFF653B7E5CEC66F447D7B85B37",
		INIT_05 => x"8342155C46680AA16664C47755C61C1D9171C3C46567C2EF996CF1714D5DFDC4",
		INIT_06 => x"FAB4D4452F7E0C78B4EDB2E79658EF5B9CC6E02B94C6BE56214EF2FE3A22273E",
		INIT_07 => x"D0837B7B0D09ED6724209EC0141C85D4F4555847E17754BF0D1847F4678417E9",
		INIT_08 => x"595582346FB1AE2566645497646CDD616546806457F0C01C55FD3CC0541D01A3",
		INIT_09 => x"149E91131C65C54410559F1C1F703C61164D743F1D4F5FD5F51E3DD564FF8BBE",
		INIT_0A => x"59CF4A87D1C74D762759477A51D61DD4C191D54F74E7529DB515DFD4C99E4DD2",
		INIT_0B => x"D1795FDCCD47E4F0E441502D5198B15CEC595BD166505F7186517514656CB443",
		INIT_0C => x"AAAAAAAAAAAAAAAAAAAAAAAA9139A57F9CCA374A2E6FCF3B1F127BEFCDB3F279",
		INIT_0D => x"D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400",
		INIT_0E => x"55FD54A855FD54A855FD54A855FD54A855FD54A855FD54A855FD54A855FD54A8",
		INIT_0F => x"D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400",
		INIT_10 => x"AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555",
		INIT_11 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_12 => x"AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555",
		INIT_13 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_14 => x"AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555",
		INIT_15 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_16 => x"AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555",
		INIT_17 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_18 => x"AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555",
		INIT_19 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_1A => x"AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555",
		INIT_1B => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_1C => x"AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5",
		INIT_1D => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_1E => x"AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5",
		INIT_1F => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_20 => x"54DD555654DD515554DD535554DD5F5554555F5554555F555555555555555455",
		INIT_21 => x"555D547D157D50D5157D51F6147D51DD545D51F554DD55DAD45D54F554DD55FD",
		INIT_22 => x"50D5735454D577D754DD73D1715773DD7D5773C44D5551554D57535555577356",
		INIT_23 => x"5DC471155DC57175555551535455515D51555155545551765055517150D5515D",
		INIT_24 => x"8AAA9FAF2AAABEAFAAAA2BAFAAAAABAE8AABAAAAAAAAAAAAAAAA7A9FA8A5552A",
		INIT_25 => x"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA4B555555555500FFFF38AABEFF8C10BB6A",
		INIT_26 => x"AAAAA6FEAAAABFAFAAEA9FEAAA9AFFFEAAAAEABFAA2BA4AAAAAAAA8AAA9AAAAA",
		INIT_27 => x"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA57FF0000955AB008AAAF2AAAAEAA",
		INIT_28 => x"550557555555D55551557555455555555555575555D5555555555D5551555557",
		INIT_29 => x"555555555555555D5555D5555555555555555555455455555555555555555555",
		INIT_2A => x"555555555555555555555555555555555555555555555555555555555555555D",
		INIT_2B => x"5555555565555555555555555555555555555555551555555555555555555555",
		INIT_2C => x"5555555555555555555555555555555555555555555555555555555555555555",
		INIT_2D => x"5555555555555555555555555555555545555555515555555551555555555555",
		INIT_2E => x"5555555555555555555554D55555557555555555555D555515555555755D5755",
		INIT_2F => x"0155555555555555555555555555555555555555555555555555555555555755",
		INIT_30 => x"55AA54025555AAAA5555AAAAEFA9AAAAFEA9ABFA555EAEBE555AEAAE555EAABE",
		INIT_31 => x"EAFF2FAA55EAFFAA5555003FAAAAFFFFAAAAFFFFAAAAFFEA55550003AAAAFFAA",
		INIT_32 => x"5555AAAAFAAA5500FAAA5500FAAA55005555AAA1EFBFAA84BEBFAAAA55AA5555",
		INIT_33 => x"5FBBEEEEBBBBEEAA5555FFFFAAFF002BEEEEBBBBEEEEBBAA5556BEEA55550000",
		INIT_34 => x"5555AAA9AAEB51005555AAA9AAAA55005555AAAA9EAA5500BEAA5500BEAA5500",
		INIT_35 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFAA555500005555000055550003AAAAFFAA",
		INIT_36 => x"AAAA5555AAAA5555AAAA5500AFEA5555AAAA5555AAAA5555AAAA5555AAFF5015",
		INIT_37 => x"555500005AEAFFAA5AEAFFAA6BAAFFAA5555000057AAFFAA5555FABFAAAAFFFF",
		INIT_38 => x"5555AAAA5555AAAA5555AAAA5555AAAAEAAA5555AFAA5405AAAA5555AAAA5540",
		INIT_39 => x"555500005555000055550000555500007AAAFFFFBEAAFEBFAAAAFFFFAAAAFFEA",
		INIT_3A => x"5555AAAA5555AAAA5555AAAA5555AAAA7AAA5555BEAA5415AAAA5555AAAA5540",
		INIT_3B => x"5555000055550000555500005555000055550000555500005555000055550000",
		INIT_3C => x"5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA",
		INIT_3D => x"5555000055550000555500005FEBFFAA55550000555500005556EFEFEAABFFAA",
		INIT_3E => x"CCCC3333CC661455AAAA5555AAAA55005555AAAA5555AAAA5555AAAA55EB5500",
		INIT_3F => x"AEAB000055550000EBAAFFFFAAAAFFAA9999CCCC99EBEEEFAEEEFEEEAAEEBFAA"
	)
	port map (
		DO   => DATA(5 downto 5),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_6 : RAMB16_S1
	generic map (
		INIT_00 => x"717BBAAA403022FEFBFF77718E46C3A223BEFEDED39C646C384476DC49B16C20",
		INIT_01 => x"8FC631163EB769786AA2A8C55182CDBD5AB4688000000000000000458BC5C5EF",
		INIT_02 => x"9F54EF85098018A41FF247FC4B1907C63E200BCBE425C5C3DB7EE1C7FF77D6E1",
		INIT_03 => x"C6ED7577D94FB8CB32492601BDEF75531B9C5C327170D38B864E2E1BEB2664CC",
		INIT_04 => x"888B1388449DC4C180013BC4224EE260C0009DF59CECFD7AF1E32180C6CD398C",
		INIT_05 => x"F9F3DFFCB1120A10B919488522112DA1428440C990B00D28CDDB37116A22D445",
		INIT_06 => x"BF6300F848EF416A631C79C2F1C4D65FCBB0C79841F2EE03661B30F4F4CF3A3C",
		INIT_07 => x"BCF9F3F3E7CFCF9F3F3E7CEBE323007001F008E60809F631AB568D1DF24B98EB",
		INIT_08 => x"5D77AE057BE0DF053221081E222984442103C4462AC115608AB14DD580680C44",
		INIT_09 => x"9D46A239C5D6CB88E600336F809625C759A0B59161D17F75FA63D45B8B3BAB81",
		INIT_0A => x"15BACD0401B65AE6602C9B68258759A0B5C4C46B65903759E1C2DBA0B5C91B11",
		INIT_0B => x"28EECC7078FBDEF31FBF606E9C4603AC33ACD1B6BFF7B5F6FB7DBD343B1B1889",
		INIT_0C => x"FFFFFFFFFFFFFFFFFFFFFFFFC467745EAD5A347766320312C24468EEB954AA51",
		INIT_0D => x"7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00",
		INIT_0E => x"7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00",
		INIT_0F => x"7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00",
		INIT_10 => x"1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE",
		INIT_11 => x"1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE",
		INIT_12 => x"1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE",
		INIT_13 => x"1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE",
		INIT_14 => x"3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE",
		INIT_15 => x"3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE",
		INIT_16 => x"3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE",
		INIT_17 => x"3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE",
		INIT_18 => x"7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE",
		INIT_19 => x"7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE",
		INIT_1A => x"7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE",
		INIT_1B => x"7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE",
		INIT_1C => x"077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E",
		INIT_1D => x"077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E",
		INIT_1E => x"077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E",
		INIT_1F => x"077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E",
		INIT_20 => x"00887880008078000088180000880000000C0000008400000000000000000000",
		INIT_21 => x"004A396C002859D0002858E0002858C40008589000984848001859F0008878FC",
		INIT_22 => x"008D2858008D2890008A28A0004A28A0006A28C0003A2964003A29A8001A39D0",
		INIT_23 => x"0000000000000000000000000000000801010010040108200001082000812848",
		INIT_24 => x"0000040040200100400000000000000002201000000000000000400010200000",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000008000000001000000000000",
		INIT_26 => x"0000010000100020020004000008000000000000000401000000000042000000",
		INIT_27 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000002000000000002400003000",
		INIT_28 => x"0048000000000000000020000000010020100100001000000000000000000001",
		INIT_29 => x"0400010000000000801000000002000000000002000001000000800000800002",
		INIT_2A => x"0000018040000000002000100008040010000000080000000000000281000000",
		INIT_2B => x"0000000020000000000000000000000000040000008000080000008000000002",
		INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000060",
		INIT_2D => x"0000000030000000000000000400100020002000080000800008002000000002",
		INIT_2E => x"0000000000000000000001000000004000000000001000008000020040100402",
		INIT_2F => x"D100000000000000000000000000000000000000000000000000000000020301",
		INIT_30 => x"FF000157FFFFFFFFFFFFFFFFFFBBFFFFFEFBFBEFFFFABBEFFFFABEABFFFABAAB",
		INIT_31 => x"4055D055FF400055FFFFFFC0000000000000000000000015FFFFFFFC00000055",
		INIT_32 => x"FFFFFFFF500000555000005550000055FFFFFFF44515FFD11415FFFFFF000000",
		INIT_33 => x"F511111111111155FFFF55555555FFD44444444444444455FFFD5115FFFFFFFF",
		INIT_34 => x"FFFFFFFC00410455FFFFFFFC00000055FFFFFFFF340000551400005514000055",
		INIT_35 => x"00000000000000000000000000000055FFFFFFFFFFFFFFFFFFFFFFFC00000055",
		INIT_36 => x"0000000000000000000000550540000000000000000000000000000000550540",
		INIT_37 => x"FFFFFFFFF0400055F0400055C1000055FFFFFFFFFD000055FFFF054000000000",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40000000050001500000144000000015",
		INIT_39 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0000000140001400000000000000015",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0000000140001400000000000000015",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3C => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFF5410055FFFFFFFFFFFFFFFFFFFC101040010055",
		INIT_3E => x"6666666666CC55555555555555555555FFFFFFFFFFFFFFFFFFFFFFFFFF410055",
		INIT_3F => x"4401FFFFFFFFFFFF410000000000005533333333334111100444011100444055"
	)
	port map (
		DO   => DATA(6 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_PGM_1_7 : RAMB16_S1
	generic map (
		INIT_00 => x"E0CFE5F7EA9BDC9A15827770B5FDB0AC898F2AAAFEB78A8B587F9A61E51BDBE7",
		INIT_01 => x"0D9D611AAA02D07177D77DBFAE5C88EC932E19D70000575500005518D3C17489",
		INIT_02 => x"57A31A7FEB2A96537D8CAAA2FDF5EAA9809432275696565D63801E7E3EC74340",
		INIT_03 => x"A748656F5E0C5D9E335DE2009CC6354B9D9FCAAB7E7FABDBD67F6F69437F61DA",
		INIT_04 => x"6235685511532B1DC5DD9A0055778CA41D550655CE6719A333D9C33E0DE5E0F2",
		INIT_05 => x"DFFB0C39B11754407D57DDCF227964BBD7BE540DF0F9DD9C1DA75A157227D455",
		INIT_06 => x"9A8766B2B2CEFC978DE0DF5F7FF62D234CDF58E46BFE30F6C8E9FD194C45CDC1",
		INIT_07 => x"3EDF87873FEF1CA8BFB3A1C4226BFCD500404A09DC528FC432E4BC42B65F5821",
		INIT_08 => x"BDBF79F7F36C28D841745762B9133B9175B219D97AE6FE8F0AB8FBBA68CAE6B7",
		INIT_09 => x"9CDB777A45B2BEDDB517A5391AA651F61954C5C420E628285193C92E1B8AF58D",
		INIT_0A => x"A61E3249263CB318FBE7B6DAEE5CB6AF3B6E3BA48F7CCCB6917E36AF3B67F67F",
		INIT_0B => x"5CD4893C6D9D12070672255C8D767621FF5C96A67D67A483C97CEA6954B34DDA",
		INIT_0C => x"5555000055550000555500007FF48BB36539C198CD193E09EDFC966B51CF8D26",
		INIT_0D => x"444493BB444493BB444493BB444493BB444493BB444493BB444493BB444493BB",
		INIT_0E => x"EEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBB",
		INIT_0F => x"444493BB444493BB444493BB444493BB444493BB444493BB444493BB444493BB",
		INIT_10 => x"D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105",
		INIT_11 => x"D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041",
		INIT_12 => x"D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105",
		INIT_13 => x"D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041",
		INIT_14 => x"C7341041C7341041C7341041C7341041C7341041C7341041C7341041C7341041",
		INIT_15 => x"C734C101C734C101C734C101C734C101C734C101C734C101C734C101C734C101",
		INIT_16 => x"C7341041C7341041C7341041C7341041C7341041C7341041C7341041C7341041",
		INIT_17 => x"C734C101C734C101C734C101C734C101C734C101C734C101C734C101C734C101",
		INIT_18 => x"FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005",
		INIT_19 => x"FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041",
		INIT_1A => x"FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005",
		INIT_1B => x"FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041",
		INIT_1C => x"D1280455D1280455D1280455D1280455D1280455D1280455D1280455D1280455",
		INIT_1D => x"D128F881D128F881D128F881D128F881D128F881D128F881D128F881D128F881",
		INIT_1E => x"D1280455D1280455D1280455D1280455D1280455D1280455D1280455D1280455",
		INIT_1F => x"D128F881D128F881D128F881D128F881D128F881D128F881D128F881D128F881",
		INIT_20 => x"ABAAEE7CABAAEBFFABAAEBFFAAAAFFFF2B2AFFFFAA2AFFFFAAAAFFFFAAAAFFFF",
		INIT_21 => x"00C0555500805345000042570180021D01800275018014D78180074500004685",
		INIT_22 => x"ABABFFA7ABAFFE6DABAAFE5B8E6AFF5782EAFF6D92AAFEDF92BAFE57AAAAFA7D",
		INIT_23 => x"0880751508907175000059530000595503015955030151560101555101015515",
		INIT_24 => x"545C0200544560005555002255150000F4D500005555000055D58000554AFF80",
		INIT_25 => x"FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAE10000555500FD0000FFFFA801F97FC90A",
		INIT_26 => x"5555004055D50002555500424D540801D555400055D500005555000051550000",
		INIT_27 => x"FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFF800FFFB1548EFEFAA00FFFFA2AA",
		INIT_28 => x"AABABDFEAAAA7FFFAEAAFFFFBAAABEBFAAAAFDFFAA2AFFFFAAAAF7FFAEAAFFFD",
		INIT_29 => x"0402555500005555021055150000455500085555100155510000555400005554",
		INIT_2A => x"AAAAFFFFEAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFE2AAAFFF7",
		INIT_2B => x"0000555510005555000055550000555500065555004055510000551500005554",
		INIT_2C => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_2D => x"0000555520005555000055550600515510004555040055150004554500005554",
		INIT_2E => x"AAAAFFFFAAAAFFFFAAAAFE7FAAAAFFDFAAAAFFFFAAA2FFFFEAAAFEFF8AA2FDFE",
		INIT_2F => x"D000555500005555000055550000555500005555000055550000555500025555",
		INIT_30 => x"AA410117AAAAFFFFAAAAFFFD5556FFFD55564003AAAF1000AAAF1000AAAF1000",
		INIT_31 => x"1518F455AA155555AAAAFFD5155555555540000040150015AAAAFFFD55555555",
		INIT_32 => x"AAAAFFFF055500150555001505550015AAAAFFF418C8FFD163C8FFFFAA550055",
		INIT_33 => x"A044111142021155AAAA00005018FFD41111444499994455AAAB4115AAAAFFFF",
		INIT_34 => x"AAAAFFFC55140445AAAAFFFC55550045AAAAFFFF615500454155004541550045",
		INIT_35 => x"05055000041100000141540005055055AAAAFFFFAAAAFFFFAAAAFFFC55550455",
		INIT_36 => x"0411515001410155050505455055050505551401515501410155050505100501",
		INIT_37 => x"AAAAFFFFA5165555A516555594550055AAAAFFFFA8415555AAAA054005055000",
		INIT_38 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFE11150000545500545100411554410445",
		INIT_39 => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFC4041515515551515555111151511115",
		INIT_3A => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFC5154000515500514445040451510405",
		INIT_3B => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_3C => x"AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF",
		INIT_3D => x"AAAAFFFFAAAAFFFFAAAAFFFFA2144055AAAAFFFFAAAAFFFFAAA9555515540055",
		INIT_3E => x"3333666633994100D5550000D5550045AAAAFFFFAAAAFFFFAAAAFFFFAA140015",
		INIT_3F => x"5054FFFFAAAAFFFF145500005555005566663333661411105111011155114055"
	)
	port map (
		DO   => DATA(7 downto 7),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
