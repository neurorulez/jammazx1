-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9BF3D52AAE560788A410940F1E0D405690B300FF7A9E00A0C1FEA7A3D3F3EDB5";
    attribute INIT_01 of inst : label is "09AD1A420D4758A728FEBE80A631D951D3861FCAC640054CA52C09AB149B71B9";
    attribute INIT_02 of inst : label is "A3BB7988EE6CEEBFD3F7FA7EFF49878CF1A52D8168B74A53000947E4DA6DF65A";
    attribute INIT_03 of inst : label is "5BDFC55CDF77CC90D74C0000092480012480480DD2B57F8747EE11FC54D2E9FD";
    attribute INIT_04 of inst : label is "DEF3EF0A090410A1492BFF7E94A5C055FA7F0CB517C5C40C625C4B75535E87D8";
    attribute INIT_05 of inst : label is "0FF00FE30FFFFE030000030301F1C363A84359B3F8D0A9ABBFFAEA944026F5E6";
    attribute INIT_06 of inst : label is "7FAD3ED399BFC4C782A8812EC85FD6B13E8D94A2AAFAA3577FFFFFE30E7999F3";
    attribute INIT_07 of inst : label is "27C0C91B02127861C8CE4C70C39D1C6CF88845BC7ACEB6DB25880411C33EED9B";
    attribute INIT_08 of inst : label is "D1DBA5DAA9235A4D2AFD9A3CA40B9301A480451CFC51A46023A881428C0563C5";
    attribute INIT_09 of inst : label is "C89E644A12A80063546D1A33C255C020049ACA0BF8B5D72546CA344614B7C7C4";
    attribute INIT_0A of inst : label is "5003EA0223E46800A02840CD00548C4410A13C94FED0622C25A1A7A5B26AA448";
    attribute INIT_0B of inst : label is "10C4310CE310C43108621886310C431086218CC6802090C421886310D06A0003";
    attribute INIT_0C of inst : label is "CCA70F283DF3DDBA59098C041533EAC25684561E11A1511E10BBAED4AD22CC43";
    attribute INIT_0D of inst : label is "3AFFCCD06A2A434A211880D5A778749AA99348D2112A147811A39D1427B58881";
    attribute INIT_0E of inst : label is "94502F822A2832AEA997A1F5DBE0E6D4EE15725FC1F1572EFE40616F13A55ADD";
    attribute INIT_0F of inst : label is "A216E3A2007D9E5FE64820760FD503CB8029FEC842AA8DF44893F9C2A0BE2F05";
    attribute INIT_10 of inst : label is "E0422DD569040D57EF79DE175170A11EF605CC95069222EABE3DB0DF6D0EABFC";
    attribute INIT_11 of inst : label is "093CA333CB961E5A4D54E0C4153944A29A7FE94B53FE6CBB418D7136704A365B";
    attribute INIT_12 of inst : label is "2B9334F6C3A81C5F68701134598F08CAA5DD75ECC3496E2B9D9F59A5D33B892D";
    attribute INIT_13 of inst : label is "9F5BD64DD35381EC42E0C7D7409E97FF955575194C9A2C0EEEA20B370789E901";
    attribute INIT_14 of inst : label is "DBD6E70B9621A4DEB3585C21B2E0000557EDDFD8D773EB7AD15F79BBFB1ADD07";
    attribute INIT_15 of inst : label is "BB7E7921A1A1A1F1338AA743F3E253A01FFB2B42DF85EB771868137ADDC61A14";
    attribute INIT_16 of inst : label is "101010101010101010101010101010101144400510501010101AAA800006664B";
    attribute INIT_17 of inst : label is "5043A085410B9454545010101010101010101010101010101010101010101010";
    attribute INIT_18 of inst : label is "D68D77E876CB25965B2C9659116CB25965B2C9659116CB25965B2C9659116821";
    attribute INIT_19 of inst : label is "1C000001C0001C8889C0001C8889C0001C00001410141155555B6FFBFDFD0590";
    attribute INIT_1A of inst : label is "5C000001D1111C8889D1111C8889D1111C000001D1111C8889D1111C8889D111";
    attribute INIT_1B of inst : label is "1C000001C4445C8889D5555C8889D1111C000001D5555C8889C0001C8889C444";
    attribute INIT_1C of inst : label is "1C000001D1111C8889D1111C8889D1111C000001D1111C8889D5555C8889D111";
    attribute INIT_1D of inst : label is "0000000004000100000400010000040000000001C0001D1111C0001D1111C000";
    attribute INIT_1E of inst : label is "0000000004000100000400010000040000000000000001110100000110110000";
    attribute INIT_1F of inst : label is "0000000000000140000000010000040000000000000001110111000110110000";
    attribute INIT_20 of inst : label is "0000000004000100000400010000040000000000000001110100000111010000";
    attribute INIT_21 of inst : label is "71C34E14853153C03AEEEEE15111551014EF8000000000880000000088000000";
    attribute INIT_22 of inst : label is "DB718AB938AE03C968FAD63B7172299D862D4B8B9785BFB6AACB50C61C0ABDCC";
    attribute INIT_23 of inst : label is "810374D0A4318C000F8001F0001E0007C00078001F0001E0007C00078003F5A5";
    attribute INIT_24 of inst : label is "0D0F9D0D0D0D0E1F8FE47583390E5F2DEEF39CB7B5FA6F30055A1B0155A1B01E";
    attribute INIT_25 of inst : label is "822D14D2C07640EFE5ECFB3243434343E74343434387E3F91D60EF97B3ECD50D";
    attribute INIT_26 of inst : label is "C9D0C217B32761A723B32761DBB7349EF3CD5570E8A82AE28B4536442E82A02B";
    attribute INIT_27 of inst : label is "95FEBDA4E27491D3EA91FCB9A4E27491C47B21927617B21849D85ECC9D0C85EC";
    attribute INIT_28 of inst : label is "F853320A7C9143C8A9E50810197793E2821C5DBA040C52C45FEDDD2713A493EA";
    attribute INIT_29 of inst : label is "82512AA23094462233E7CC7AB3E7CC7A33F9734E24246281091FF5450977E7E5";
    attribute INIT_2A of inst : label is "3012324172CF7121349338909B2FEA1289C582513BA2B0944622BB2FE2128944";
    attribute INIT_2B of inst : label is "F3335BAC6AF6F7B79D9A9DB764D6374C048C905CB3DC494D24CE2426D99318DD";
    attribute INIT_2C of inst : label is "00398671C6400F4F4A31C6400F4F4A31C66618DEB320EE37822A3E3D8D5EDEF6";
    attribute INIT_2D of inst : label is "CE7D6E83FBBB7AA00FFF5A9D8B4FBBFC6E66CDDA7B89D36148B4935073800000";
    attribute INIT_2E of inst : label is "CE63550FD2CA4E881E6F9ADD3A21E6F972D3A7440F37CB969F3A21E6F9AD10DA";
    attribute INIT_2F of inst : label is "6953B9530FFFA596E239DC636BAFD2DB4A07939B87346B741C6B7B408F9F381C";
    attribute INIT_30 of inst : label is "05965A49165957C46B740C5A3D029E5DAE2C6CC2A35BA0480977953226143F4B";
    attribute INIT_31 of inst : label is "0C954B6DB7E9A7B6FF776746BB439B5D8EB679728D7E8550544DE8E47C97D600";
    attribute INIT_32 of inst : label is "EDB1AED0E46373635DA1E3759D1AD902F42A399B9B1C75BAEDEBA5364FF90D10";
    attribute INIT_33 of inst : label is "EFB7DF53800013A19B1ADD2D08A31BB7CD36824C49D7DF7FBEDF7DFAFA1042FE";
    attribute INIT_34 of inst : label is "3A1D0E86870A1D7475F6E9E444440C070002301E9A1D347A6874D111FBE9F7DF";
    attribute INIT_35 of inst : label is "0AECFC518ACC21C6A6A3A02B30871A9A8FC58A8FE26FB56528E8686874347434";
    attribute INIT_36 of inst : label is "01E23725BAC9992C6318C28A0470025E16161617340D76EF6FEC42C0AECEC42C";
    attribute INIT_37 of inst : label is "999ADD263DD93264CB9F2F134D8737098F764C9932E7CF339789A680EC981232";
    attribute INIT_38 of inst : label is "8BF648665F37C3BF8148657C6FD740A730CF30CD8D5EDEF6F3335BAC6AF6F7B7";
    attribute INIT_39 of inst : label is "0D0D0D0F9D0D0D0D0E1F8FE579733EED50D0D0F9D0D0D0D0E1F8FE57762FD9DD";
    attribute INIT_3A of inst : label is "222000010106020400040002A802A0062002200000020000000000079733EEC9";
    attribute INIT_3B of inst : label is "324A01649258E14E5F2DECF8282C3034282FC3C000040004000400040002A2A6";
    attribute INIT_3C of inst : label is "0CA134F54D177691CA5E3DE45A0A548A3B77A80029AFDE8F7C58406EC0193733";
    attribute INIT_3D of inst : label is "A05971F4F4C670A1C2853B7FC36DFF8997ED38E38FA3C1F63C9F04E0580A5414";
    attribute INIT_3E of inst : label is "4EC23DA4725F4AE7C702D452A4552AAE84D70FE49AA28035FD6057EB832EA1DB";
    attribute INIT_3F of inst : label is "F778057F5E000E06368919D1D7FEB93A7DDDF4DE0801844D8E75391D9D3B0F67";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "F2F71E3EF96E3F6D0086CCDD7747BDEBC40080FA5D28592DCAFBCD6603E38D93";
    attribute INIT_01 of inst : label is "C8A4E93AC459F28FD7A1CA593F7C21CAC24E277C2824F0B0428CC0C3A061C72C";
    attribute INIT_02 of inst : label is "2E8D4AC6818834FCF53F9EA7F3D461411E8C67B24D9918C765425AA926DB0C3A";
    attribute INIT_03 of inst : label is "6333EF21404601B4405004804000124924800800544753F7E22C7AB348FFA365";
    attribute INIT_04 of inst : label is "30679ED325B24408000600023199D9B12BFF2DEFBFCC76D32B8D793FE7A43412";
    attribute INIT_05 of inst : label is "7F00FFCE6FFFFFFE7FFFF3FEFFF0038EACD0BF1803B5021400038D596DEB1251";
    attribute INIT_06 of inst : label is "80024088CCE00239D8D5EB7B23700127402802EC0AFD75A07FFFFFEE619E1E0E";
    attribute INIT_07 of inst : label is "930626E9F7A93081C04E8A7103891C8CF7D755F596ABE906186473EB041824B1";
    attribute INIT_08 of inst : label is "16E3621932FC04D0B4004B8F03BF347490372A636EC7EA8D991F34EE4070DCB8";
    attribute INIT_09 of inst : label is "4B89B1A77843DB7723E442C7C8F719ED97B7216E0006A5561402869E8668581C";
    attribute INIT_0A of inst : label is "8D9A1E8CF905D5E17F57FF7EF7BAB785C9BFC719C07E06BD19085B0C570561AB";
    attribute INIT_0B of inst : label is "F77BEE777EE77DDEFF9CFF79EE77FCE7BDCEFB7AED35777BFE73DFEF23B19BBC";
    attribute INIT_0C of inst : label is "0D074343C00BFFFDB2541135E89003E6CDDFCDE0AC2CE57D40AAEFAA006C3FBC";
    attribute INIT_0D of inst : label is "A446AA559D0F36D4FAC8A630065E800A64BD7389262E53A95AAC1562B406AD95";
    attribute INIT_0E of inst : label is "B489DB3CDA4BB495742CAC08040D43B9F16FFF1C74027C224D348BA67BC2A582";
    attribute INIT_0F of inst : label is "95A9D2156DFDB6F00549AC1C5266346E582D0112BAEF16D1FDBC01194C6CD469";
    attribute INIT_10 of inst : label is "8F29F10F8CA0A9A000A0EF7FDD3A637D45DF85B0D241955ACE62374EDB45AC01";
    attribute INIT_11 of inst : label is "B68294A4D0A28EC005323C933CA0602C02DB725396DB97E47295BE0005AF90CD";
    attribute INIT_12 of inst : label is "2BE5470E3C528E0526E33E32622B2B2ED6134B03B9814476D364929219001292";
    attribute INIT_13 of inst : label is "2ED6BD8041E7ECE7741069219A4C7D291685AC4A5006F59D8A91CDD99E2E0001";
    attribute INIT_14 of inst : label is "B68020D0AB5A5BB40146815A6E39BF5321E032B30085DAD7A6213C06566014D4";
    attribute INIT_15 of inst : label is "AE5ECC3232323205FFE3FFB4002EB48CD257783590EB52411C2682D4904709B0";
    attribute INIT_16 of inst : label is "001011001011001011001011001011001151511115401011001AAAAAAAA44402";
    attribute INIT_17 of inst : label is "D24BA405480BC011001011001011001011001011001011001011001011001011";
    attribute INIT_18 of inst : label is "F932402682DB6DB6DB6D96DB1424B6C96D92D925B142492C9259249249142925";
    attribute INIT_19 of inst : label is "9C000001C0001C4445C0001C4445C0001C0000BFEEBFEEAAAAC000FF7FA52049";
    attribute INIT_1A of inst : label is "9C000001C8889C4445C8889C4445C0001C000001C8889C4445C8889C4445C888";
    attribute INIT_1B of inst : label is "DC000001C8889C4445C8889C0001C4445C000001C8889C4445C8889C4445D999";
    attribute INIT_1C of inst : label is "9C000001C8889C4445C8889D5555C0001C000001CCCCDC0001C8889C0001CCCC";
    attribute INIT_1D of inst : label is "0400000000000080000000008000000000000001D9999C4445D9999C4445D999";
    attribute INIT_1E of inst : label is "0400000010000080001000008000100000000000151004880095011000000400";
    attribute INIT_1F of inst : label is "0000000004000080001400008000100000000000151004880084040000000400";
    attribute INIT_20 of inst : label is "0400000010000080001000008000100000000000000000C800C40040C800C000";
    attribute INIT_21 of inst : label is "720AD05C4927B0756ABEBEBEFBEBFEFBAE500000040005110084000111000400";
    attribute INIT_22 of inst : label is "DB8199D3407600525CA95AD852002C03B64A4F901A1C5AFC07E8F0019C01BBC9";
    attribute INIT_23 of inst : label is "807F24BAE2092C00058000F000160007C000D8000F00016000FC001D8002F6D3";
    attribute INIT_24 of inst : label is "91951991919197A3E0F6AEB446D77DD83DF5C760EFF6FF7002972B012972B012";
    attribute INIT_25 of inst : label is "E40F3BFBFABDDDF64151FF7C646464654664646465E8F83DABAD010547FDD991";
    attribute INIT_26 of inst : label is "9BF6D5AB766FDA7FB5766FDA46006BA209D993A2248332F323CE7E502F1B2483";
    attribute INIT_27 of inst : label is "285020EFF8A9ADE9962A5122EFF8A9ADE7B76DA6FDAB76DA9BF6ADD9BF6D6ADD";
    attribute INIT_28 of inst : label is "0C5B5E479768AC54560A668433893809F78F1E95AD9AC9A59289177FC54D6996";
    attribute INIT_29 of inst : label is "55DA6447056694A30809BDBB4809BDBB44A245FF9189082420428E9E9FE8BFED";
    attribute INIT_2A of inst : label is "E43196894B5EF5684921553569E130AED32255DA6447056694A309E130AED322";
    attribute INIT_2B of inst : label is "F7F6FF5CCE2C1FFFBFB7BA6C0DE24BF90C65A252D7BD5A1248754D59B037892F";
    attribute INIT_2C of inst : label is "001FF497F48007420217F48007420217F4A65BFE57A4EEFF9ADE6A6B99C583FF";
    attribute INIT_2D of inst : label is "95000A6A6F6E160CD80AA001F2924826000211483A4700A464C645721A400000";
    attribute INIT_2E of inst : label is "3BBDFFFA18919719487709645C648756914CCB8CA43BB09A665C64875492AAE5";
    attribute INIT_2F of inst : label is "429C439C55743103BCE6779CEBFA1881D89A7864F059805351924D35150CEE73";
    attribute INIT_30 of inst : label is "AF6D9DF7992465B9801354E943DD29B4C94BC92C4C029A2DD60C69CF39A12862";
    attribute INIT_31 of inst : label is "D2587CC209B64965B250D098053539817813944530026862E285B3840965236D";
    attribute INIT_32 of inst : label is "B466024D93B008CC069BB002EA64946DF99390003A522D603BDA3A487220D432";
    attribute INIT_33 of inst : label is "025C0492D99982B2466015B0DB9D804A164D798B7D3D24B92DD692A4B65B27FE";
    attribute INIT_34 of inst : label is "A32994C8C911A05697DE3AF914430C0A0010101B6D96DB2DB6DB6D058091012A";
    attribute INIT_35 of inst : label is "9B09677AEF6573DE127F443D95CF7949FE0961F8E50249B64D4D4D4D46A6E6A6";
    attribute INIT_36 of inst : label is "B1254C632490664D6B5AD0C1B3265B2F2F2F2F2864C21E3FFF11CC19B4B01CC1";
    attribute INIT_37 of inst : label is "3367365CAD92244893224C681A7A4C572B64891224C8ED7B26340C689172318C";
    attribute INIT_38 of inst : label is "F009A6D9D04FBE7F2B92B3F84C1095D9EE90E69399C583FFE6ECEEDCCE2C1FFF";
    attribute INIT_39 of inst : label is "919191951991919194A26097904C7F9D99191951991919194A2609790BC02642";
    attribute INIT_3A of inst : label is "2320000202000000000000033406200320020000000000000000000104C7F9F1";
    attribute INIT_3B of inst : label is "6ED1333D3592F4B17C583BE7CFCC3C383C380000000000000000000000022223";
    attribute INIT_3C of inst : label is "13989B479B3C9D765AE761A8EC1DDDA5E07817FFE6C47E2ABF0EB673F3437D67";
    attribute INIT_3D of inst : label is "9B387B3F6D1281C827774FB6DD9EDBD6BF93ACEE1D4751A8751A80D2EE1DDD91";
    attribute INIT_3E of inst : label is "DFB4875D96FE5E6BF04764EEEC2E1DF10C26CF18BFA1FFC60180671A5D733DB6";
    attribute INIT_3F of inst : label is "F78B598C7800027959B7D01A80B10ED01226D3E33CD3CD712F4BFDABB77ED2ED";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B8F75726584E0F09E0048401C746010854004139934811D543F94D7719E99B81";
    attribute INIT_01 of inst : label is "800510D2845071D000114811FB7C79C2820002FC22B6A024218000C0203B6B8C";
    attribute INIT_02 of inst : label is "2A292B42846424FCF6BF9ED7F3D8A152EA0C47A36880188F460052A966248202";
    attribute INIT_03 of inst : label is "60EFFB045144512414442082000000000012480110B30C2121A2480A5419935D";
    attribute INIT_04 of inst : label is "D461860008241C3A4003FE78330DF35123FE2DE597CFA22F0B45610AA7ACB45A";
    attribute INIT_05 of inst : label is "F00FFFDEFFFFFEFEE0000C0EFFF03C8E9A909B9D60A53A0400B34D58491B55CF";
    attribute INIT_06 of inst : label is "D63ACB588ECB3619D01067F31A5B1F55CAA80024807577908000001EF01FE00E";
    attribute INIT_07 of inst : label is "B3BE6CC9D9DB38C9CF0E747193931C48F2086461FDFC71891CFFB30DA91666B9";
    attribute INIT_08 of inst : label is "900A409034CC75B1A6EC938FDF3FEC3CB3872661AE8003419D25A52283F19836";
    attribute INIT_09 of inst : label is "6AC2F9291680484204C64A03C87588688FF71A4B6680E170540480168028C506";
    attribute INIT_0A of inst : label is "8892046E61E54100300061D404093ED548BB075AC06E902D0F2C4D2856094048";
    attribute INIT_0B of inst : label is "A5EF5BDA95BDAB6B52D6ADEF4B5EB7BD6B7B5694CD17ADAD4B5A95BDE2F3B396";
    attribute INIT_0C of inst : label is "A59343404BA84488D56040656D3124107260A0E08520695C11BAAFEEEFA392D6";
    attribute INIT_0D of inst : label is "A291000701A822D619B3FEB981BC044280B9E09284AB9521D8AABD008080A19E";
    attribute INIT_0E of inst : label is "161449841B2A22A6980B298EDAA17569F0131C9478E85188B622050B1A8C76ED";
    attribute INIT_0F of inst : label is "4198D72C09611AE1AF8CA8546547344AB3E8586B5A8A436569B86B8242A63309";
    attribute INIT_10 of inst : label is "031AE8576721213764DF967FDEA20151BF9FFF29F2CF935FE8B633A9B255FEB1";
    attribute INIT_11 of inst : label is "9B14A104D8B2CE8221402C277C04A929CEC91FDFF649FE21FFDFEF12002128A3";
    attribute INIT_12 of inst : label is "2BF966858010CE94842A7A1173AB0A4CA61540980191C461D1B6DBA1573D1B9B";
    attribute INIT_13 of inst : label is "33BDEFF090A7C6D22247BABEC6C25318F24CAB8B58C8D084A8A5CDDF9FB00001";
    attribute INIT_14 of inst : label is "8FFE80890CE7227FF0644EF62BB100CA4FF49B8BFE0677BDE33A7E93717FE08C";
    attribute INIT_15 of inst : label is "BF7EEE0307030735EA83550AF6AD6988E9EAB12068C3EDB2BC0422FB6CAF0118";
    attribute INIT_16 of inst : label is "544554544554544554544554544554544040004414104554544FFFFFFFF22243";
    attribute INIT_17 of inst : label is "5B6E924F249E8554544554544554544554544554544554544554544554544554";
    attribute INIT_18 of inst : label is "5DBDB28406492C9259249249152D925B24B64B6C9406DB6DB6DB6D96DB152DB7";
    attribute INIT_19 of inst : label is "3C000003EAAABF3333EAAABE2223FBBBBC0000BFFFEAAA20804925FFFFE4926D";
    attribute INIT_1A of inst : label is "3C000003E6667F3333E2223F3333EEEEFC000003E2223F3333E2223F3333E222";
    attribute INIT_1B of inst : label is "3C000003E6667F3333E2223F7777EAAABC000003E2223F3333E2223F3333E222";
    attribute INIT_1C of inst : label is "3C000003E6667FBBBBE6667E2223EEEEFC000003E2223F3333E2223F3333E222";
    attribute INIT_1D of inst : label is "8800000000000040000000004000000000000003E2223E2223E2223E2223E222";
    attribute INIT_1E of inst : label is "88000000080000400008000040000000000000000808804004000000C00C1908";
    attribute INIT_1F of inst : label is "44000000080000400008000000000400000000000808804004080000C0040808";
    attribute INIT_20 of inst : label is "88000000080000400008000140000000000000001D8044000018811000001D80";
    attribute INIT_21 of inst : label is "7927C93F9213735B811045111514000551444000080888400408088840040808";
    attribute INIT_22 of inst : label is "0649CB9724E502CE3918C63380A2980B0C300305024D9E6D739FB0268C161D08";
    attribute INIT_23 of inst : label is "417B6870FC309A0021400268004D000CA0019400368006D0010A003140046645";
    attribute INIT_24 of inst : label is "181AD83838181D2E83A15650B882BE9C3AE8A270D7E17E2801CE62811CE62806";
    attribute INIT_25 of inst : label is "0C007E198DC756AC41A1FEB00E0E0606B60E0E06074BA0E855942D0687FAC038";
    attribute INIT_26 of inst : label is "E01CBF780B8077550E0B807731978601FA21BA22A6E1BA89001F84550892AEEA";
    attribute INIT_27 of inst : label is "C7ABD7EAA1C6190300C7ABD7EAA1C6190880B97807780B97E01DE02E01CBDE02";
    attribute INIT_28 of inst : label is "A57A8304084711C388CC843192C72C610574119918B59B551D4E9F550AB2C300";
    attribute INIT_29 of inst : label is "174B930585C2EBCB807E10CB807E10CB8F57AFAA08109118908A04C4C1964002";
    attribute INIT_2A of inst : label is "162E084A19852A06EFB029C9C62CB8BA5C93174B930585C2EBCB862CB8BA5C93";
    attribute INIT_2B of inst : label is "E0284296E32E1FBF014254490970EC058B821286614A81BBEC0A72712425C3B0";
    attribute INIT_2C of inst : label is "00021B8A1B80080D480A1B800742020A1B8208BE028C662F82977B7ADC65C3F7";
    attribute INIT_2D of inst : label is "52EFF04675FBDF28842A2A15DAD999562428A1B2CAA7412479779710BA000000";
    attribute INIT_2E of inst : label is "9A94FBBE5CF17991475DF1B7E64475FBE3F6BCC8A3AEDF0FB5E64475FF1FEEF2";
    attribute INIT_2F of inst : label is "82D632D65D5CB9E196D33294EFBE5CF0B1BC8C7F18EDFF4201EDA422531E6B69";
    attribute INIT_30 of inst : label is "2DB6DB2C9249D0EDFF4210BBE14D24CDFDEA3FB66FFA1001C7322965ACB47973";
    attribute INIT_31 of inst : label is "1458684B2CB6CBFEFB732EDFF0202BCD450EDE613FE84232B7F8DA441DEFF649";
    attribute INIT_32 of inst : label is "4097FC0802F1212FFA10B1363B7B6A4FC33BD4895A957BCFDEF3BFEF789C8176";
    attribute INIT_33 of inst : label is "D92DB26D5E1E0234097FC1948917896D8494996A694C001A4012002D00C92500";
    attribute INIT_34 of inst : label is "D0381C1C1D912E615BF43FFC000000044000223924D249A4934927AAB64F6C96";
    attribute INIT_35 of inst : label is "5B4A62384F7972D94C7D023DE5CB6531F68459F0E1EDB5A6812121A1A090D0D0";
    attribute INIT_36 of inst : label is "154622309658100118463849A786C1403070307346BE943F7E504C85B4A504C8";
    attribute INIT_37 of inst : label is "0502506AD1BF36FCDB2E0291A8BE029AB46FCDBF36CB0D430148D4445A4B2E00";
    attribute INIT_38 of inst : label is "FA0FC45C2A47042A0B20A0F28C0F95814B714B72DC65C3F7E0A04A16E32E1FBF";
    attribute INIT_39 of inst : label is "3838181AD83838181D2E83A050607F8C038181AD83838181D2E83A0523E81F48";
    attribute INIT_3A of inst : label is "3034000000040004000400003C0420043004000000000000000000050607F8C0";
    attribute INIT_3B of inst : label is "78912645D71484A2BE9C38E3F3F43C3BC3C40000000400040004000400002024";
    attribute INIT_3C of inst : label is "9CECE017812420828875C141F0BE0885195618001ED17E0B9780A282E2224379";
    attribute INIT_3D of inst : label is "113E2E8780145BF54FD213DB566F6D581FA1AB4C6A1A8541A8142E8DF0BE083F";
    attribute INIT_3E of inst : label is "00CF0820A07E0E39786F85F044456AEB84970AC496A28025F940570A0C39BB56";
    attribute INIT_3F of inst : label is "F188C1CF380002621911FAB390B10A92121B656B20828A610A42A87058033816";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "B0F1468149470321F009248083040318D2002038000C11D7C8FE64D6D8F8F289";
    attribute INIT_01 of inst : label is "6C61B8C4E48CC28228E06211EA36CCC9084F22AC089242342118A4A6005BAB0A";
    attribute INIT_02 of inst : label is "A7B8330706E461BF56D7EADAFD58C21097A2ECEFF39344D956448D4C9324C302";
    attribute INIT_03 of inst : label is "D2EFE925390A400131800010000000000000000810D8453088CCE29A5A0C410A";
    attribute INIT_04 of inst : label is "90269A4020825C2A4012A18689B25533485F989D77A0AA4AC7B0FD233321ABCB";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000116411B104290294460A5145191FC321D";
    attribute INIT_06 of inst : label is "442D0FC18AA21060C0B047EA3C9216F10E8805397588092C0000000000000000";
    attribute INIT_07 of inst : label is "00D0401821200831C40E207063871C28FD5FDB096D651DDB429A80608F4D4011";
    attribute INIT_08 of inst : label is "232D82F9B7A05B43B7FAE5114452D0F008A61707860403690906842A8480020A";
    attribute INIT_09 of inst : label is "EB8B60215E8029B330C6AC7BE743A1FA1DF63A92422550674400250208B55B54";
    attribute INIT_0A of inst : label is "E1D7055E3018A220022046E400CD7D6881798C1B8E9829141C28DC28C2218071";
    attribute INIT_0B of inst : label is "EFBDCF7B3DFFF9EF77FFE7BDCF7FBFFF7BFFF7399BC5E7BDDFFFBCF7AFD5D55E";
    attribute INIT_0C of inst : label is "E011050259F9A247C52090C1CD2000004040803A2047EC3D44FBEBBBAAAD37FF";
    attribute INIT_0D of inst : label is "049B00C041A1264695FB5830D5E0E404C0D5C2D3250FA6352ACFB874A9252C9B";
    attribute INIT_0E of inst : label is "79C50FAEB4F34E36120FC40F9FE9754C8C42811310F2196EFF84856F4CD4D67F";
    attribute INIT_0F of inst : label is "4108C788486272C1EF934F15E760354A8BCD10CA54C397F56BB07BD26ABEBF5E";
    attribute INIT_10 of inst : label is "495AEF577509E9BFD6F9E2A784B45279F6294E0BC0230BDF8CA41B2C0095F822";
    attribute INIT_11 of inst : label is "9B1CB18541000A0A026044CAB08D000CDD125B9DE892D8878B5BD34221298B2B";
    attribute INIT_12 of inst : label is "2BFF8A178010D0020080F8E2BD8A319712021DC81A42867304B2CBE157FF9B1B";
    attribute INIT_13 of inst : label is "118C630DB5328802A474B4B6522618844120E5291CAC50142130322F9F800001";
    attribute INIT_14 of inst : label is "5DDB9C150AD292EEDC8088C220B5203C7600C9DADBA2318C755EC0593B5B4011";
    attribute INIT_15 of inst : label is "993E30A9E9ADEDA3A44788937CFC0782C12219847E0EEDEBBF90CDBB78EFC42B";
    attribute INIT_16 of inst : label is "1101001101001101001101001101001100004404045501001104444444411109";
    attribute INIT_17 of inst : label is "76D8C92192402544554100110100110100110100110100110100110100110100";
    attribute INIT_18 of inst : label is "58ADA310EF249E493C925924BFFB6DF6DBEDB7DB6FFB2496492C927924EABB6C";
    attribute INIT_19 of inst : label is "3C000003C0003C0003D1113C0003C0003C0014BFFFFFFE8209E492A4925D25A4";
    attribute INIT_1A of inst : label is "3C000003D1113C888BD1113C0003C0003C000003D1113C888BD1113C0003C000";
    attribute INIT_1B of inst : label is "3C000003D1113C888BD1113C0003C0003C000003C0003C888BD1113C0003C000";
    attribute INIT_1C of inst : label is "3C000003D1113C0003C888BD1113C0003C000003C0003C888BC0003C888BC000";
    attribute INIT_1D of inst : label is "2000000028000300002800020000380000000003C0003D999BC0003D999BC000";
    attribute INIT_1E of inst : label is "20000000240003000020000300002C000000000022222110102A22A110102222";
    attribute INIT_1F of inst : label is "2000000024000300002000034000280000000000222221101022022110103232";
    attribute INIT_20 of inst : label is "00000000240003800024000200002C0000000000222221101122222110112222";
    attribute INIT_21 of inst : label is "60AAC55C00471125014050140145554415400000332102222233023222223321";
    attribute INIT_22 of inst : label is "1A2909DF1474014018294A5A20612B1BBE008D831F557BEE41BC70A01C083917";
    attribute INIT_23 of inst : label is "007F0033E02A2800470005A000B40012800250004E0009C0003800170000B3C1";
    attribute INIT_24 of inst : label is "4F4F954D4D4D4C884216450E26181E39490638E505E42E6014062E004062E00A";
    attribute INIT_25 of inst : label is "7D702110B7478834B31C8A49D3D3D3D3E55353535322108591438ACC7229334F";
    attribute INIT_26 of inst : label is "907048D40E41CD88B20E41CDDB1E08228308D6BDD5355C157C0847AEC1FDD538";
    attribute INIT_27 of inst : label is "4B4183311041063F034B4183311041062940E0C41CD40E091073503907063503";
    attribute INIT_28 of inst : label is "E35463B4D84527E293C830A5268E68FD28D2224429F29D38FA1C398882187F03";
    attribute INIT_29 of inst : label is "789C627516271B9D18E4108518E41085168306110242044246377E9E91DEC007";
    attribute INIT_2A of inst : label is "D35B009DFAA086D0AEB062223E3DE1C4E308789C627516271B9D1E3DE1C4E308";
    attribute INIT_2B of inst : label is "E0E40C6ACDFCA7D7072063002043AD34D6C0277EA821B42BAC18888C00810EB4";
    attribute INIT_2C of inst : label is "4A2A5B2A5B000742022A5B000742022A5B36591E684A884790E5656559BF94FA";
    attribute INIT_2D of inst : label is "C67DA00896DD6E0A94AA821D9A5C93D897628EFBF867540E2872863220400F4F";
    attribute INIT_2E of inst : label is "CCC67EBA68875A953AB892BF6A53AB8D259FAD4A9D5C692CFD6A53AB892BAEB6";
    attribute INIT_2F of inst : label is "188718873D74D10CC53198C66EBA6886017A47968F2D6DC8756DF40447D33298";
    attribute INIT_30 of inst : label is "8E491EDB1DB69BC56D4854B7710C4C5F646164A32B6A4227131788718E7129A2";
    attribute INIT_31 of inst : label is "C9684EF4D1EDA49349316456D4050EC42E544C4D2DA10A1A3EC84AE40ECE4724";
    attribute INIT_32 of inst : label is "5DB5B52152C4B36B684204AB195B7A17C15D85A11462DADB56B17DFABEF81D2A";
    attribute INIT_33 of inst : label is "B6C76D801FE00E1A9B5B70C41F162567A006D4714E26490EDB39247B6C924800";
    attribute INIT_34 of inst : label is "BE9F4AB6A75D885671EC8B0C000000000000000C9239247248E49054EDB1DB63";
    attribute INIT_35 of inst : label is "4111C0A04E8C320A164A45BA30C828592888692AE6496FBEFB7B6AEA7D3D75F5";
    attribute INIT_36 of inst : label is "BAEAAEDBD75834F28425255D8B03593A9E9ADEDA606EEC8FAF865F64111865F6";
    attribute INIT_37 of inst : label is "076067A57949DBB64DAA6E111D8C66695E5276ED936ACA8337088D0F5A689B08";
    attribute INIT_38 of inst : label is "101C20A47E50823F5481407E8E20454D4B654B6559BF94FAE0EC0CEACDFCA7D7";
    attribute INIT_39 of inst : label is "4F4F4F4F954D4D4D4C8842176CC7229334F4F4F954D4D4D4C884217600405080";
    attribute INIT_3A of inst : label is "030400000004000400040003C4042807000400000000000000000006CC722927";
    attribute INIT_3B of inst : label is "8405C98A38E712981E394907FFFFC3C40000000000040004000400040000282F";
    attribute INIT_3C of inst : label is "33201BF71170D1469430C1CC8F11C154B51A1600019581843D2089186A700285";
    attribute INIT_3D of inst : label is "43A40606138DD90F6430E97FD1A5FF1717B187247E7B89C7B8DC4E1C8F11C155";
    attribute INIT_3E of inst : label is "83BA5451A45F89C3D2447C8E0C1E1DF40D26CE38BFA1FB46018067A84E989E2C";
    attribute INIT_3F of inst : label is "F0A00CA4A8000B207D435CE0D0B60A5612CFF6424514D328230C4590760EEC1D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "62098E904121202F40024A8187062529E410103A0A9055A908F96C444DEDBBA2";
    attribute INIT_01 of inst : label is "4001A09045090288AA014A55BB122288DC6BA364232480A842B2C0ECA20A4622";
    attribute INIT_02 of inst : label is "C41BBB0804B4EC0386E070DC0E18847926F97E2A21A1F3F4DE480BF9B5000004";
    attribute INIT_03 of inst : label is "0CA8214411104524100504800012012012010084A278083B8134E0C28F640010";
    attribute INIT_04 of inst : label is "544514524DB76AC78504AB2BE5E815350D00500658102A53BBEF770AB70B72D8";
    attribute INIT_05 of inst : label is "00000000000000000000000000000000EC826B328124009534B1441125A00243";
    attribute INIT_06 of inst : label is "2804A41499942515C0A14B66D1240202A528864000A200640000000000000000";
    attribute INIT_07 of inst : label is "A92D2A5B494A97F63CF1618FEC7F636F1AA0AAA0DCEFBB7E62A56904AD415881";
    attribute INIT_08 of inst : label is "0292411392CA09AA9C10B14911536AF8A11C0E502E024A050D1514A403694A54";
    attribute INIT_09 of inst : label is "7190A4A52401694262CE384C158781681FBE51248481D3E09445800C42C0890A";
    attribute INIT_0A of inst : label is "81F455CF12508520624485109CAB3EA08138948993D8449801418141900540C1";
    attribute INIT_0B of inst : label is "8C6318C690842108421084210846318C21084295134D8421084210843A15D550";
    attribute INIT_0C of inst : label is "341A02917445EEDC100843C099D04124894989788405243EEA05115451040631";
    attribute INIT_0D of inst : label is "0C6400640541A6DC53ACC2221600C80041B3CB19A70702418A0510628081E1D8";
    attribute INIT_0E of inst : label is "208CB114504184185868855A044788AD884BD5B398481EC100061D80286C2D22";
    attribute INIT_0F of inst : label is "052B521B2C802ACC448107597671B46C9C0C209290E34201EFB311094644502C";
    attribute INIT_10 of inst : label is "6539C68E1460E0E0859414A0C600C66328A9A323E284077F904803819247F943";
    attribute INIT_11 of inst : label is "1B1D1114A4820404082425267087840F3AC90B7AD648C98F53BCEB620CA82181";
    attribute INIT_12 of inst : label is "2BFD62192CD6F84300EAA8462220614412871A322F4F505601B6DB455F835B1B";
    attribute INIT_13 of inst : label is "339CE707C6B60E22A55913698A881D2925B62A8B199430182412C08F9F800001";
    attribute INIT_14 of inst : label is "33370815694ADB99BC60894A459720052C329B71B726739CE33506136E36F01D";
    attribute INIT_15 of inst : label is "3261048585C5C5B1844308A4963C858EE1C4510586099B0BED80E066C0FB6030";
    attribute INIT_16 of inst : label is "000111000111000111000111000111000455111051000111000EBEBEBEBF0F33";
    attribute INIT_17 of inst : label is "C002A497492EE555444111000111000111000111000111000111000111000111";
    attribute INIT_18 of inst : label is "3F9B63C0DA001C0028005000AEA001C0028007000EEA001C002A497492EEA001";
    attribute INIT_19 of inst : label is "FC000003D5557C4447C4447C4447C4447C00181555555402234003A492556C49";
    attribute INIT_1A of inst : label is "FC000003CCCCFC4447C4447C4447CCCCFC000003CCCCFC4447C4447C4447CCCC";
    attribute INIT_1B of inst : label is "FC000003EEEEFC4447C4447C4447CCCCFC000003DDDDFC4447CCCCFC4447CCCC";
    attribute INIT_1C of inst : label is "FC000003CCCCFE6667C4447E6667DDDDFC000003CCCCFC4447C4447C4447CCCC";
    attribute INIT_1D of inst : label is "0000000000000000001000000000000000000003CCCCFC4447CCCCFC4447CCCC";
    attribute INIT_1E of inst : label is "000000001000008000100000000000000000000011010282AA11010202220000";
    attribute INIT_1F of inst : label is "000000001000008000100000000000000000000000000282AA11010200200000";
    attribute INIT_20 of inst : label is "000000001000000000080001000000000000000000000282AA80000282AA8000";
    attribute INIT_21 of inst : label is "5A9614B39B39A010104411044401545044510000000001908900000190890000";
    attribute INIT_22 of inst : label is "53A4D038520FBED461DAD6B8F2009F802E52099013269D31340930910C111A40";
    attribute INIT_23 of inst : label is "EF790CC09C51DF003BE0037C006F800DF001BE0033C0067800CF0009E0073012";
    attribute INIT_24 of inst : label is "0C0AA40C0E0E088842148D2400110270410461C10C04A07DF69807DF69807DF6";
    attribute INIT_25 of inst : label is "E7362160149A0A164210084983830302A903038382221085234911084021320C";
    attribute INIT_26 of inst : label is "923088844648C808A04648CA4614492A21B8F638545D0639ED885BC2C3507418";
    attribute INIT_27 of inst : label is "C2A142811009246520C0A040811009246B4469448C84461112321119234A2111";
    attribute INIT_28 of inst : label is "0390CD95A340052002B820A5368168456082064023D23D20950A140884492520";
    attribute INIT_29 of inst : label is "588C4675063311C904403181044031810140819100000000000A809497850000";
    attribute INIT_2A of inst : label is "1111002C0804A4000D30262620CA30C4623A588C4675063311C900CA30C4623A";
    attribute INIT_2B of inst : label is "0464C6488B3820502326324A09630C0444400B02012900034C09898928258C30";
    attribute INIT_2C of inst : label is "020630863080074202063080074202063038E300C44310C030D440411167040A";
    attribute INIT_2D of inst : label is "82D3780E35B31C5B9955D5E89CDB6FA8D4E5380180E67615A37A362220C00742";
    attribute INIT_2E of inst : label is "808415414924B1912619B4B2C64261996D8618C8930CCB6C30C642619B4B1539";
    attribute INIT_2F of inst : label is "D0CEF08E1A229248041700841011493494D824125824DB8060DB1C064236020B";
    attribute INIT_30 of inst : label is "14003A087000E00CDBC066B7626C04F26D63CCA6E6DE03B5237C08E11C3BC524";
    attribute INIT_31 of inst : label is "544A4DC002A481BEDB67CFCDBC0644DC7940FC8F1B780C3A3EDACF843A552E00";
    attribute INIT_32 of inst : label is "A7E36E01D2C6A7C6DC0386BA3736C657CD51D7B160C7B9C6CE77B92619101062";
    attribute INIT_33 of inst : label is "0014003BA0000C1C7E36E0E4191635D036D911C34C740038005000E000924BFF";
    attribute INIT_34 of inst : label is "94140B1606118895103C430C0000000000000038005000E0014003BB8005000E";
    attribute INIT_35 of inst : label is "F1014AB044C29E69084C0F930A79A421301C51300DB69892512030A0289058D0";
    attribute INIT_36 of inst : label is "59294409671850138CE71B65AB8B4928585C5C5A48449C40A1409C8F101409C8";
    attribute INIT_37 of inst : label is "632E3286527DFBF6CCAC4881A11A6CA1949F7EFDB32B92242440D20F98099101";
    attribute INIT_38 of inst : label is "9E1820910048926A30A2400992A24150C610C6111167040A0C65C6488B382050";
    attribute INIT_39 of inst : label is "0E0C0C0AA40C0E0E088842151084021320C0C0AA40C0E0E088842150A2784028";
    attribute INIT_3A of inst : label is "101400004040808101020203FC06880410042000000080010002000108402126";
    attribute INIT_3B of inst : label is "A495894A28C6389102704107FFFFFFFFFFFFFFFFFFFBFFFBFFFBFFF800028A8C";
    attribute INIT_3C of inst : label is "49024A0716F0800335A4D51C85108364E50A160000D6614455A008912E7240A4";
    attribute INIT_3D of inst : label is "0306269E0900C10B2420494900A524426033874D68DA3D1DA391FC3C85108320";
    attribute INIT_3E of inst : label is "91940249CD80B1855A0428841C6F4ACB0CB70AC494E284ADFB405730DC50DC6C";
    attribute INIT_3F of inst : label is "F4D908DA2A0004225B031EBAA47204D49AA0016B0C304120611845023246408C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "710D8E1159292925059B6E920B0E2529740208B8A8A2D5FB5BFE82666BEB9FAB";
    attribute INIT_01 of inst : label is "534D821E5E482280A8F28ED5F70C22DAF86AA204AEB686A842F6C1BD80AF0716";
    attribute INIT_02 of inst : label is "84CD4A10C8293542A52854A50A9108D82288622AA9C510C456514AAB644934D0";
    attribute INIT_03 of inst : label is "AAA82189B66C9DB5B6DC24000010010010000005247160350C2943028A909803";
    attribute INIT_04 of inst : label is "4CE79E4924937060C077D24A219B1539AA40F446C8396E430B4667B541FA3E10";
    attribute INIT_05 of inst : label is "000000000000000000000000000000009AE4391089B484D49377DDB9B480132B";
    attribute INIT_06 of inst : label is "088090928884F492C2D94B2205B4C02391A93362AA2283320000000000000000";
    attribute INIT_07 of inst : label is "A534A92D272A500803009E0010008090100075D496A820440137E492F8009313";
    attribute INIT_08 of inst : label is "52120531526901E4B131172928577939E6144A4836124A855D9414A64BA5248E";
    attribute INIT_09 of inst : label is "418420A53049094222C48A441DA329B2949201B68E920042D09E924A1A684D8E";
    attribute INIT_0A of inst : label is "A9922457609485207244E55494895EACA93B04298278049661E061E0624504D9";
    attribute INIT_0B of inst : label is "84210842118C6318C6318C6318C210842318C21111450C6318C6118C72119110";
    attribute INIT_0C of inst : label is "2C379919400A55A81881498C81F00924C949C92C94A4253C4141440054664210";
    attribute INIT_0D of inst : label is "6E20005425492640528B9AFA75C49C16489141999366320DB9E4132392922431";
    attribute INIT_0E of inst : label is "2C8C99145E7967945928E5234C054950124B322139094A9104A64C922A5CC0B6";
    attribute INIT_0F of inst : label is "652BC21924C32A420439E45D656AB66EDBCDA6821EF94A49E79081094664502B";
    attribute INIT_10 of inst : label is "0D7B401A154DAD8988121EA8AEC25320242B97ACE798254AA0E9ABB1DF5CAA4F";
    attribute INIT_11 of inst : label is "5A31168046041A160320A52EF9B481A4060002D6B00080ACCAD6A204C4ADADB1";
    attribute INIT_12 of inst : label is "2BFD2E5C36D6C81ED49AA902F766295E96D7D903B941DD4519A69AE8DE055A5A";
    attribute INIT_13 of inst : label is "2AD6B5042140495AA59200008A9449CE0638209A513A1A964995FFF060000001";
    attribute INIT_14 of inst : label is "A2A452922BDE4B15229491CA6ED52003051B12A124C55AD6AAACA3225424AA9A";
    attribute INIT_15 of inst : label is "E541A98F8F8F8FE1C64BCC9C5514848FE6065624714952C5C8549254B1721524";
    attribute INIT_16 of inst : label is "000000000000000000000000000000000000000000000000000045104510FF12";
    attribute INIT_17 of inst : label is "D249A49149214000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "3D12441482924D249A493492542924D249A491492142924D249A491492142924";
    attribute INIT_19 of inst : label is "38000003A22238888BA22238888BA22238000BEAAAAAAA2000D248A49247246D";
    attribute INIT_1A of inst : label is "38000003A222391113A222391113A22238000003A222391113A222391113A222";
    attribute INIT_1B of inst : label is "380000038000391113AAAAB91113A22238000003A22239111380003911138000";
    attribute INIT_1C of inst : label is "38000003A222391113A222391113A22238000003A222391113AAAAB91113A222";
    attribute INIT_1D of inst : label is "080000001000000000000000000000000000000380003A222380003A22238000";
    attribute INIT_1E of inst : label is "0800000008000000000000000000080000000000080888000000000000000808";
    attribute INIT_1F of inst : label is "0800000028000000000000000000080000000000080888000008008000000808";
    attribute INIT_20 of inst : label is "0800000008000200000000020000180000000000080808000000000000000808";
    attribute INIT_21 of inst : label is "400200100003000EBEFAEBEFAFFBFFAAFAFE8000080808000008008800000808";
    attribute INIT_22 of inst : label is "0200003000043EC0005A529800000F802C000100060C08600008100004000800";
    attribute INIT_23 of inst : label is "0F7B0001800018001B000160002C00058000B000160002C00058000B00016000";
    attribute INIT_24 of inst : label is "5E57245E545E509E4D978B24CC912259998479664A24D061F000061F000061F6";
    attribute INIT_25 of inst : label is "57F2A935198F4C9F431D865F17951795C917951794279365E2C9310C76197C5C";
    attribute INIT_26 of inst : label is "12210CEC44488E4CB844488E442849321D9B925E45917595DCAA4EF2591645D6";
    attribute INIT_27 of inst : label is "CEE74EE99309252506CEE74EE993092529C4426488EC44219223B11122133B11";
    attribute INIT_28 of inst : label is "77924624814E2707131924A5379D79CD3CE253F13893892CB73A774C9C492506";
    attribute INIT_29 of inst : label is "5CBE66672F2F9DEB299339B3299339B32DCE9D9920000000001F489893E81FDF";
    attribute INIT_2A of inst : label is "E0FD2CEDE73DECD9CA20CF2F247032E5F3285CBE66672F2F9DEB247032E5F328";
    attribute INIT_2B of inst : label is "04CC8CDCCDCCC8E82264266E4DE4C8B83F4B3B79CF7B36728833CBC9B9379322";
    attribute INIT_2C of inst : label is "020F7DC73DC0074202073DC0074202073D40412044D600481E4A626399B9991D";
    attribute INIT_2D of inst : label is "00B2554D252A574A9BF5FFFF5092484009003B0436D64045AA5AA576C2C00742";
    attribute INIT_2E of inst : label is "08847FFEDDBD3135E4D12426C4DE4D104D14989AF2688268A4C4DE4D1242FEAD";
    attribute INIT_2F of inst : label is "B0F4A0B417DDBB58850210847FEEDDBCD3BB67A4CF48926A5892DAA7A0242281";
    attribute INIT_30 of inst : label is "5D24A8005492000892EA7AA5434D80A4484B88254495536B2A280B41682EBB76";
    attribute INIT_31 of inst : label is "555925524A80112492528A892AA6C889716896CE92554D23A292871C2A152E92";
    attribute INIT_32 of inst : label is "A0424BA9AA8048849553C0422224B757815DDC0272D62D64AB5A7A44D102902A";
    attribute INIT_33 of inst : label is "925D24ABFFFFF35F04249AFA95D402D036DD15DB657524BA497492A9252492AA";
    attribute INIT_34 of inst : label is "90B45A3E2ED59ED782209A88000000000000002A495492E925D24ABEA495492E";
    attribute INIT_35 of inst : label is "F72946F1D5CCD34F2A5826D7334D3CA9604E51610536D092432222A2219151D1";
    attribute INIT_36 of inst : label is "999DAAE2E59066D084A12555ABB24928E8E8E8ED29F3E091D14ACDAF7294ACDA";
    attribute INIT_37 of inst : label is "666C66C5AA76EDDA9590CAD03910C2F16A9DBB76A56452D465681F4993703D2D";
    attribute INIT_38 of inst : label is "9AD01491F758B2EA78B6E48A5331E0C9EFB9EFBB99B9991D0CCD8CDCCDCCC8E8";
    attribute INIT_39 of inst : label is "5E545E57245E545E519ECDB790CF61B7C5C5E57245E545E519ECDB792E6B604B";
    attribute INIT_3A of inst : label is "101000000000000000000000040008001000200000000000000000010CF61B7C";
    attribute INIT_3B of inst : label is "E6D7098F3CF696B322D99B8FFFFFFFFFFFFFFFFC000000000000000000000808";
    attribute INIT_3C of inst : label is "43A21B279324996718FDCB0AACD5A955C24E920000DE615E17B20813AA6B62E6";
    attribute INIT_3D of inst : label is "53C6EE4F8930E549952A4680119A00162833AF6CE85A1B0DA1F0DF9CACD5A9F4";
    attribute INIT_3E of inst : label is "913C0659C4A015217B3566AD4C1C3DF40D04CE38BFE1F94E0380673ACC7D993F";
    attribute INIT_3F of inst : label is "F0D90BDEAE0005664B537B0AB0A82EDE133249EF2492CB65295A65C22644F089";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "320E644450898C103269226D36B3180010480478000723A9E5FF46E2C9F9C9B8";
    attribute INIT_01 of inst : label is "3E321C4136A5B8A22A714323AA2CC8E54C2284C31200120C6392442482183327";
    attribute INIT_02 of inst : label is "D3892B0136C43442B6A856D50ADC834CE186258254D30C430504A6A40224C38D";
    attribute INIT_03 of inst : label is "38EC21B60982640208252000000200200201000E09208D9111E084582600111C";
    attribute INIT_04 of inst : label is "B2410424924913265491FF7E1880C19B48A0797CE01DC7090545A3ABA3AA1358";
    attribute INIT_05 of inst : label is "000000000000000000000000000000018849C910C40249C3BFE1060C9220B90C";
    attribute INIT_06 of inst : label is "0D4962ED88868B4D8D1431221C8624B86283690A2A2AA3D40000000000000000";
    attribute INIT_07 of inst : label is "58C316CDD9C588000000000000000000100001585CEC34C904801B6CA10E52C9";
    attribute INIT_08 of inst : label is "28DF619C1906921BE25E81DBC51586B698C3B135EC6920F01B40C211041AD830";
    attribute INIT_09 of inst : label is "D486621087046CE7984405303F390C20C4921C90C148810941B0492569026461";
    attribute INIT_0A of inst : label is "0C09E80FADFA61C03C23788867543C620CFD6C0C8E503248CF264F2659306204";
    attribute INIT_0B of inst : label is "318C6318C6318C6318C6318C6318C6318C6318C70105B18C6318C63180C80886";
    attribute INIT_0C of inst : label is "E69236341B38448AF316A482063524922424A4624251B29C04541005517298C6";
    attribute INIT_0D of inst : label is "199900C09034B2430C3881305B36254124914464491208310C10D89849489081";
    attribute INIT_0E of inst : label is "826265C30104104304831285B73027E8952114103474B18DB2312349858612DB";
    attribute INIT_0F of inst : label is "D0C64BC69208864336C410B04FC239D1883234C84906A1265A90CDE431170B84";
    attribute INIT_10 of inst : label is "18C61870C71B5B12F65964288D9B088CB68AC81ADA63D8CA878C436700B4A86A";
    attribute INIT_11 of inst : label is "0B94498189DB656AA0926FC22F6C0350CA925B5AD492D859539CEB13B2135B63";
    attribute INIT_12 of inst : label is "2BFF0331E58C483606003CF8201194854BAC35CE6941706F35B6DBB223410B0B";
    attribute INIT_13 of inst : label is "139CE70CB1A260D032708592616371F007C061499D8850C53048408810000001";
    attribute INIT_14 of inst : label is "4B3680C9C4A52059B0264CA112818000F304DB48B622739CF912E0DB6916C0C5";
    attribute INIT_15 of inst : label is "7761F8E5E5E5E5F33BB6B74768E739C4D9398DB2CA659B3388062566CCE20189";
    attribute INIT_16 of inst : label is "00000000000000000000000000000000000000000000000000005015054000FF";
    attribute INIT_17 of inst : label is "C001800300054000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "D08B72060600040008001000012000C001800300054600052488001492012000";
    attribute INIT_19 of inst : label is "3800000380003A222391113A2223911138002CAAAAAAAAAAAA4000A480040100";
    attribute INIT_1A of inst : label is "38000003911138888B911138888B911138000003911138888B911138888B9111";
    attribute INIT_1B of inst : label is "38000003BBBBB80003911138888B911138000003800038888BB33338888BB333";
    attribute INIT_1C of inst : label is "38000003911138888B911138888B911138000003911138000391113800039111";
    attribute INIT_1D of inst : label is "2000000020000080002000008000200000000003B33338888BB33338888BB333";
    attribute INIT_1E of inst : label is "0000000020000100002000010000200000000000222021100022202110002220";
    attribute INIT_1F of inst : label is "2000000000000100002800010000200000000000322121100000000110000000";
    attribute INIT_20 of inst : label is "000000002000010000200001000020000000000022202110102A28A110102220";
    attribute INIT_21 of inst : label is "3FF9FFCFFFFEFFE0150054055001555500554000000002222000000222200000";
    attribute INIT_22 of inst : label is "F9FFFFEFFFFBC1BFFFB5AD67FFFFF07FD3FFFEFFF9F3E7DFFFF7EFFFF3FFE7FF";
    attribute INIT_23 of inst : label is "F086FFFE7FFFF7FFE4FFFE9FFFD3FFFA7FFF4FFFE9FFFD3FFFA7FFF4FFFE9FFF";
    attribute INIT_24 of inst : label is "0F0A970F0F0F0F1FB7E8F3DB32CE23B95E9BA6E5723B519E0FFFFDE0FFFFDE0D";
    attribute INIT_25 of inst : label is "851C2CC9E270A168D36085B1C3C3C3C2A5C3C3C3C3C7EDFA3CF6CF4D8216E30F";
    attribute INIT_26 of inst : label is "CCD4DE139B3361B7479B3363B99734DDF3E8DDB1C0700E69670B308F4688E071";
    attribute INIT_27 of inst : label is "6118B196ECF4D2D7116118B196ECF4D2D639A9F336139A9BCCD84E6CCD4F84E6";
    attribute INIT_28 of inst : label is "8715B8175E219990CC46D65AD0E30E39D31DAD4D86DC6DC248C58CB767B6D711";
    attribute INIT_29 of inst : label is "AE071989C381C295DB6ED6CDDB6ED6CDD231636EC00000000000B2E2ED12F034";
    attribute INIT_2A of inst : label is "9213DB0C11E739B66DB1BB9B938DED7038C3AE071989C381C295D38DED7038C3";
    attribute INIT_2B of inst : label is "19BB5BAC533CA8E8CDDADD03A05A6F6484F6C30479CE6D9B6C6EE6E40E8169BD";
    attribute INIT_2C of inst : label is "023AD2BAD2800742023AD2000742023AD22514A13AC68928413626258A67951D";
    attribute INIT_2D of inst : label is "764B6062B1B3DE00C480820B5C5DB9982620EC92C187C122386387DDA5800742";
    attribute INIT_2E of inst : label is "C642155C2896C8F3F21D90BB234F21D921F72479F90EC90FBB234F21D90B10B6";
    attribute INIT_2F of inst : label is "184798071AB8510C40B18842000C28960D7C8C37186C5B03145B343017B71858";
    attribute INIT_30 of inst : label is "0D249800300002C45B4310B1782E6C496D762C8322DA18A4139384708E3030A2";
    attribute INIT_31 of inst : label is "086CBAD2498005B6DB692445B43112E6C6CC5C580B60609FBAC8C87688440600";
    attribute INIT_32 of inst : label is "0C916C0C02C13922DA1801311916CA05C011B489CDAD39D6CE733B721CC8CBA3";
    attribute INIT_33 of inst : label is "000C000140001018C916D0D0C1160965EDB2D306BACC00080010002001249000";
    attribute INIT_34 of inst : label is "BE170B9787199C5872349B8C0000000000000018003000200040014080010006";
    attribute INIT_35 of inst : label is "0194C47485D9FADA8F5A901767EB6A3D69231D6C125B2ECB397979F97CBCFCFC";
    attribute INIT_36 of inst : label is "5AC27705B6D8992631086041834B659E5E5E5E5F004A9491D1A62C60194A62C6";
    attribute INIT_37 of inst : label is "8992996E117DFBF6CE9F173DC5AF171B845F7EFDB3A70A028B9EE264DC8953D2";
    attribute INIT_38 of inst : label is "B926466E4820C7159AC9788E0BCF40E6525652558A67951D1132532C533CA8E8";
    attribute INIT_39 of inst : label is "0F0F0F0A970F0F0F0E1F37C874D0214E30F0F0A970F0F0F0E1F37C8752E499D4";
    attribute INIT_3A of inst : label is "232400038382020202000003F806A0072006000000020002000000034D0214C7";
    attribute INIT_3B of inst : label is "F00810379E4968CC23395C90000000000000000000000000000000000002A2A7";
    attribute INIT_3C of inst : label is "04E024BACC0A6699EB557070B0160EA619B4580001A3C1C6AF4C016C83101FF1";
    attribute INIT_3D of inst : label is "18302BB4F68F3160C583B2A4864A9249C84950C713A4E8764E874462B0160E9C";
    attribute INIT_3E of inst : label is "66C619A67B20646AF40580B0746A5FCF08A70ACD95C784A9FA40FFE5BFA992DA";
    attribute INIT_3F of inst : label is "F3BC60FA3A000C6334118AC2D106912224CB245ABAEB2CB296B5BA3CD99B0F36";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "080CC404540808802160040106138094B00002F80006A30091FE0391C8F8C091";
    attribute INIT_01 of inst : label is "2A05104216C5A402A07408A3220CD91155020DC10A00000C21A0002800396084";
    attribute INIT_02 of inst : label is "418D210096E42040228804510088814CE18320021ACB06400482C4040224828C";
    attribute INIT_03 of inst : label is "38CC01850145540104540000000040040040000D0431459008E0C258060880C9";
    attribute INIT_04 of inst : label is "8110410000003060C003FF7E0C81015958C06150901882090541A3A1008E1548";
    attribute INIT_05 of inst : label is "000000000000000000000000000000018041191050804983BFE2080A00001104";
    attribute INIT_06 of inst : label is "054902E18AA28841A48201220812A4B10380002A802AA9140000000000000000";
    attribute INIT_07 of inst : label is "40C0100C00040800000000000000000010004058484414C902800000210540D5";
    attribute INIT_08 of inst : label is "30DD618811009203825A8212451480A081800104AD2090601000800204420080";
    attribute INIT_09 of inst : label is "D0866000120068A510440628382108208492080251008101C000000600284544";
    attribute INIT_0A of inst : label is "0A8BE00400EC3101313061DE044414C408700C088E30290C0572057212A06008";
    attribute INIT_0B of inst : label is "318C6318C739CE739CE739CE6318C6318C6318C60104B18C6318C63190C88886";
    attribute INIT_0C of inst : label is "E25107101B3800025302800405649249521212420061A31C50514010512218C6";
    attribute INIT_0D of inst : label is "299B00C0487AAA420018000145250D22129150D0002210131020D91001008041";
    attribute INIT_0E of inst : label is "45400D820288288682032244B3206C405090040C2270C19DB628005B06091249";
    attribute INIT_0F of inst : label is "0802CB800049464336CA22944542654A8808144C6A88836D4090CDC020360B05";
    attribute INIT_10 of inst : label is "000008C045206012D6492228080A0104928A4C02820600EAA22462020004A828";
    attribute INIT_11 of inst : label is "19140501E5820E0E91094AC2280C0061C8924908449248691108490A20084207";
    attribute INIT_12 of inst : label is "2BFF0495A4854004050022A042221889ACB454DA288014C50492496011411919";
    attribute INIT_13 of inst : label is "1108420CB101505029718496C107460038006129CC980080A884200545400001";
    attribute INIT_14 of inst : label is "C99284A50294904C90252A94A201400013D2C9C8922221085916F859391240A1";
    attribute INIT_15 of inst : label is "D521B867676767734216C40369E42184816201A84854C92A888507324AA20149";
    attribute INIT_16 of inst : label is "000000000000000000000000000000000000000000000000000500155000000D";
    attribute INIT_17 of inst : label is "C001A49300054000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "10892A0506000C00180030005560004000800100001200052488001492002000";
    attribute INIT_19 of inst : label is "B80000038888B800038888B800038888B8003088888888000040008000040100";
    attribute INIT_1A of inst : label is "380000038888BA22238888BA22238888B80000038888BA22238888BA22238888";
    attribute INIT_1B of inst : label is "3800000380003AAAAB80003A22238888B800000380003A22238888BA22238000";
    attribute INIT_1C of inst : label is "B80000038888BA22238888BA22238888B800000380003AAAAB80003AAAAB8000";
    attribute INIT_1D of inst : label is "10000000000000000010000000001000000000038888B911138888B911138888";
    attribute INIT_1E of inst : label is "3000000010000080001000008000100000000000110010800891000080089100";
    attribute INIT_1F of inst : label is "100000003800000000100000800010000000000000000080089100008008B300";
    attribute INIT_20 of inst : label is "3000000010000080001000008000100000000000110010000011010000001100";
    attribute INIT_21 of inst : label is "80040020000200101555000555540000005540003320308008B320008008B320";
    attribute INIT_22 of inst : label is "0000002000080000000084200000000008000200040010000010000008001000";
    attribute INIT_23 of inst : label is "0000000100001000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "1B1A831B1B1B181E1784420372A8A02450620091420010000000000000000000";
    attribute INIT_25 of inst : label is "06202A110645C38880807410C6C6C6C6A0C6C6C6C60785E11080CE0201D0431B";
    attribute INIT_26 of inst : label is "21045D36208413C422208411B952821DF6015E0180200A89A80A840C08008062";
    attribute INIT_27 of inst : label is "9100815884420B17099301835884420B106208E84136208BA104D88210474D88";
    attribute INIT_28 of inst : label is "8516231458114088A0C81542020220710410B10D4ED0ED0448040AC422105709";
    attribute INIT_29 of inst : label is "3D0E800C0743A2161B2600461B2600461603068840000000000016828116C004";
    attribute INIT_2A of inst : label is "1222400831800000659023435225E1E874023D0E800C0743A2161225E1E87402";
    attribute INIT_2B of inst : label is "020020322812280810010100204264048890020C600000196408D0D400810990";
    attribute INIT_2C of inst : label is "022002A002800742022002800742022002A410202084880802211D1E45024501";
    attribute INIT_2D of inst : label is "6659205090994820A4AA000B4CCC99B81720A596C28440902922920026800742";
    attribute INIT_2E of inst : label is "CC42555C3042D8F3D248919B634D248B24936C79E92459249B634D2489194096";
    attribute INIT_2F of inst : label is "485398130AB860A4C0319842555C304201724812902449428449242806933018";
    attribute INIT_30 of inst : label is "0C001800300002444942959135284C49253A2582224A14A111938530A61030C1";
    attribute INIT_31 of inst : label is "0870A2C0018014924939244494293267464448280920509F9A48586708040600";
    attribute INIT_32 of inst : label is "0C91240A0240B922481400B111124A04A011148556B51092442131324CC8A9A2";
    attribute INIT_33 of inst : label is "000C000140001210C9124090A112056DA496D10AA34400080010002000000000";
    attribute INIT_34 of inst : label is "3E33199D8C311C24EA0211640000000000000008001000200040000080010006";
    attribute INIT_35 of inst : label is "0218C0280529CC120F520014A730483D48031D480259668A387878F87C3C7C7C";
    attribute INIT_36 of inst : label is "52C222209248102C6318C041020B451676767677008802101084684021884684";
    attribute INIT_37 of inst : label is "1001016A902F5EBC581C0A140DA4021AA40BD7AF16070040050A045448096240";
    attribute INIT_38 of inst : label is "282E452C480704151B01AA8601DF888400540056450245010200203228122808";
    attribute INIT_39 of inst : label is "1B1B1B1A831B1B1B181E1784E0201D0431B1B1A831B1B1B181E1784F40A099D0";
    attribute INIT_3A of inst : label is "000000000000000000000000000000000000000000000000000000020201D043";
    attribute INIT_3B of inst : label is "C80000434D118888A02450600000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0A20509AA11D504188510040A815080415C554000183BE8AAA000188828002C8";
    attribute INIT_3D of inst : label is "14080804408C3150C54228A48522924508056180322C8042C8040886A8950824";
    attribute INIT_3E of inst : label is "082214106020046AA00540A8443C39F00904CE31FFC1FD8E0380CFA6BA298310";
    attribute INIT_3F of inst : label is "F6B041762A000CD2A6195CE6F0974A9612D96C4AAAAA28CB18D6211104209C41";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
