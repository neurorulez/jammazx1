-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFF60C19552568AFFFFFFFFFFFF1652814B46C728D6F8D28905";
    attribute INIT_01 of inst : label is "FFFFFFFFA9D71659645D85FE819D4FA8FFFFFFFF0C142878B856995563665870";
    attribute INIT_02 of inst : label is "FFFFFFFF832752BBFFFFFFFFB62F4438FFFFFFFFFFFF284C8A22FBC0FFFF2120";
    attribute INIT_03 of inst : label is "CD45CEB9FFFF596A841EBF2E46745A7EFFFFFFFF93016D3EADFE155AAD9D5305";
    attribute INIT_04 of inst : label is "140E40E8CDAA02A29601A7078888888848888884888888488888844113114567";
    attribute INIT_05 of inst : label is "C140A40A40A40A14828AFC500930AE8CDAA02A29601AF074029D00AB4024069F";
    attribute INIT_06 of inst : label is "B02B02B20A28FDC02C42BAF16ED00A3402AD00902A3F503903A706AF00ADC06B";
    attribute INIT_07 of inst : label is "AE8A336ED00A28CD4029C18AE4028A3C6E4029C18AE4028AE8CDAB8029F02B02";
    attribute INIT_08 of inst : label is "0E88ABC1BB80280E88E9C1ABB900A28CD4029C18AE4028FD8AE4029C18AE40E8";
    attribute INIT_09 of inst : label is "078814068C1AA02A29601A7078A01ABB0AA469C288A88E88E8C5AA58069F80A8";
    attribute INIT_0A of inst : label is "AFC1AA58069F06A80A8A5806BC1C1AA02A29601A7078814068C1AA02A29601AF";
    attribute INIT_0B of inst : label is "0ABC02C02BC1D00AB402402BC1F00ABC02C02BC1D00AB402402BC1C12AE69601";
    attribute INIT_0C of inst : label is "7A8003BFFEAD503540FC143FA5AFFD7FFF5FEAAABAAAAEBD7FAF5FEE40A9C1F0";
    attribute INIT_0D of inst : label is "EDAFB48D24AA8FCBFE4929A3F2FE5928A3F2FE492BA3F2FF96FFC00033FBFD55";
    attribute INIT_0E of inst : label is "C6B0B3F510EDE8EB83A1FE50B22A91BFDE45DF2EF2AE1FFED904E815A5B7171B";
    attribute INIT_0F of inst : label is "268FCD8A051B82B2DBF3FED1141C9F04A8227932B581F1BD837ED896DBBD714A";
    attribute INIT_10 of inst : label is "3743030302C302C040403C3FFFFFFFFD75BA0A91982BB42BA1B50C62A15E06BE";
    attribute INIT_11 of inst : label is "EAA0200A00028182AAA0028000A0AA03C3FC444444444441541010100C100C00";
    attribute INIT_12 of inst : label is "A2A08028928982D5E28AD7A157BE8200AAAA80A8028A820092A0A02BABBAAAEE";
    attribute INIT_13 of inst : label is "BE2BE8022B78A82A8AA8ABF2A82AA8124B0982D7AF857BEF82B5C280A28028A2";
    attribute INIT_14 of inst : label is "0EC3555C5554B32CC9555555555CBC65768200A00A80A0028A8224980228A822";
    attribute INIT_15 of inst : label is "55555CB32CC555C5554B0EC35754153F33F335755C71CD5D573F33F315D5054B";
    attribute INIT_16 of inst : label is "EB91F5F9F548BA00F0F42C0FC1DD409DD73C0F01640000000000195D8BC95555";
    attribute INIT_17 of inst : label is "AFBAAEA8A80A2A04A800482A0AA2A002A8AAAA2A09501A28AE8B51782F0F40CB";
    attribute INIT_18 of inst : label is "A82A82A00A8A8200828982D5E2B55EFAA2BE8200AAA02A24A2A08828AD7A2A0A";
    attribute INIT_19 of inst : label is "A80A80228A82F888021578A822AAFBEBF2802AA8224A2A08AD7A17B557BED70A";
    attribute INIT_1A of inst : label is "D55539FE7D55755555FEFFFBF57F55555FBEFB5D5D55800A0A802A028A80AA04";
    attribute INIT_1B of inst : label is "5557EEFD5FBFFD55755555FF9FE7F575554FCCF54C5655C71C5655CF54CFCCD5";
    attribute INIT_1C of inst : label is "60180AEBBF97F5F9174A2A06C290A4380AA802202AAAFD31C0591757554EFBD5";
    attribute INIT_1D of inst : label is "7BEDEA0AAABE80A828A82A0092E0AAA8AAAAAB8AAA80504216808AF8AED74090";
    attribute INIT_1E of inst : label is "BE8AFA0002A028028A2A0891578A82FB57BEABE8028A8228028924A8228915E1";
    attribute INIT_1F of inst : label is "2A00A822498022608AF8AFA008ADED70AA2AA2AFCAA0A820492C26155EB5EB57";
    attribute INIT_20 of inst : label is "4FC3FC3575415B3B55C55554CE33B5573D5F4FFD155155555D6600200A00A80A";
    attribute INIT_21 of inst : label is "555557593FF4F57D3B55738C55554ED57B315D5054FC3FC3D5C555471CD5C555";
    attribute INIT_22 of inst : label is "AA03D20560AAEC80B710101C1705C26BBA757EABE0502409016CC00059480554";
    attribute INIT_23 of inst : label is "8A812A0A882AA2A0B5E4B157A0A02BAAE2BAE802A020022A0182AAA0008A80AA";
    attribute INIT_24 of inst : label is "00A82208260857BE15ED757B7A08028A80A820282A0892C90A82ABE17B55E2BE";
    attribute INIT_25 of inst : label is "72F195D56600028A80A80A8028A8122004A82F857BE802FB57A822A028ABF22A";
    attribute INIT_26 of inst : label is "45554ECEC5655FBEC5655CECECD5545554BC2F0D5D5555D50F7F0577F5525575";
    attribute INIT_27 of inst : label is "C008000000000000000006575592F25575715DFD54F7F0D5D5555D50BC2F0D55";
    attribute INIT_28 of inst : label is "0D58E141141D0768AEAA295100C10008108AE445DF9D542A80482304C02C509C";
    attribute INIT_29 of inst : label is "EEBB861151FFAA54318A266E4BDCD099BB56F07392AE145601EDA50541451527";
    attribute INIT_2A of inst : label is "268D55BFAD115155EC69896BBBAEEEBBBF288A3EE41515E68D43EEBB86115143";
    attribute INIT_2B of inst : label is "096952E0A63ACA2352F4BE045752EB95403FC02A58658987964B79AE198B3A86";
    attribute INIT_2C of inst : label is "A50EE659CB9672E59CB967045FA94F372243ACAEEFCEBAD69955156DA5522022";
    attribute INIT_2D of inst : label is "0242511067522919D0BA1E618A23821208BE9E6779EC9ECA742E87BBBBB36BC2";
    attribute INIT_2E of inst : label is "C018BE9D2113499134C442E879D1D91880444222088822222FB7A744869DDDD2";
    attribute INIT_2F of inst : label is "595D830402D1B2F0911F0667FFFFFF0E52B938A0A99841C49C2CBD2112321446";
    attribute INIT_30 of inst : label is "3743030302C302C040403C3FFFFFFFFD75BA0A91982BB42BA1B50C62A15E06BE";
    attribute INIT_31 of inst : label is "EAA0200A00028182AAA0028000A0AA03C3FC444444444441541010100C100C00";
    attribute INIT_32 of inst : label is "A2A08028928982D5E28AD7A157BE8200AAAA80A8028A820092A0A02BABBAAAEE";
    attribute INIT_33 of inst : label is "BE2BE8022B78A82A8AA8ABF2A82AA8124B0982D7AF857BEF82B5C280A28028A2";
    attribute INIT_34 of inst : label is "0EC3555C5554B32CC9555555555CBC65768200A00A80A0028A8224980228A822";
    attribute INIT_35 of inst : label is "55555CB32CC555C5554B0EC35754153F33F335755C71CD5D573F33F315D5054B";
    attribute INIT_36 of inst : label is "EB91F5F9F548BA00F0F42C0FC1DD409DD73C0F01640000000000195D8BC95555";
    attribute INIT_37 of inst : label is "AFBAAEA8A80A2A04A800482A0AA2A002A8AAAA2A09501A28AE8B51782F0F40CB";
    attribute INIT_38 of inst : label is "A82A82A00A8A8200828982D5E2B55EFAA2BE8200AAA02A24A2A08828AD7A2A0A";
    attribute INIT_39 of inst : label is "A80A80228A82F888021578A822AAFBEBF2802AA8224A2A08AD7A17B557BED70A";
    attribute INIT_3A of inst : label is "D55539FE7D55755555FEFFFBF57F55555FBEFB5D5D55800A0A802A028A80AA04";
    attribute INIT_3B of inst : label is "5557EEFD5FBFFD55755555FF9FE7F575554FCCF54C5655C71C5655CF54CFCCD5";
    attribute INIT_3C of inst : label is "60180AEBBF97F5F9174A2A06C290A4380AA802202AAAFD31C0591757554EFBD5";
    attribute INIT_3D of inst : label is "7BEDEA0AAABE80A828A82A0092E0AAA8AAAAAB8AAA80504216808AF8AED74090";
    attribute INIT_3E of inst : label is "BE8AFA0002A028028A2A0891578A82FB57BEABE8028A8228028924A8228915E1";
    attribute INIT_3F of inst : label is "2A00A822498022608AF8AFA008ADED70AA2AA2AFCAA0A820492C26155EB5EB57";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFF70074FE23C7FFFFFFFFFFFF07F202D30254262CDF279B02";
    attribute INIT_01 of inst : label is "FFFFFFFF4584CDCC9876F350EA5343CEFFFFFFFFA04ECD8E6F30274F9CBD3D00";
    attribute INIT_02 of inst : label is "FFFFFFFF330D7DC0FFFFFFFF381C0DCDFFFFFFFFFFFF3051F1BCA200FFFF0012";
    attribute INIT_03 of inst : label is "01763000FFFF3734D043D0F2698E3542FFFFFFFF3D830473725906FE7642D411";
    attribute INIT_04 of inst : label is "080C80C51C510118310014030500000060000007000000400000057677747666";
    attribute INIT_05 of inst : label is "006846846846841448710C1311301C71C51011831001C0380072001480480473";
    attribute INIT_06 of inst : label is "0A10A10221C73C04400071041CE0018800620120118F20320310418C002C0004";
    attribute INIT_07 of inst : label is "1C518710E011051C80041061C888614F1C88841061C88851C51C6340040A10A1";
    attribute INIT_08 of inst : label is "0C4887007340040C48C7006372011061C80071041C80863C51C80871061C8046";
    attribute INIT_09 of inst : label is "034008006005101183100140341001844854460C44474C48C60460C400634084";
    attribute INIT_0A of inst : label is "18C060C4006301440460C400700C05101183100140340080050051011831001C";
    attribute INIT_0B of inst : label is "218400400410D0218400400410C0218000000410C0218000000410C09C583100";
    attribute INIT_0C of inst : label is "355503FF555D557555C14170505FD7D7F5F5C3EBF0FAFC2AAB0AAADC800410D0";
    attribute INIT_0D of inst : label is "67259D876B87061FE5EAE1C18FE5EAE1C183E5EAE1C183F97AFDFFEAB3335550";
    attribute INIT_0E of inst : label is "3CCF115C30DF5A7C91FC63C0DA3FAC15438EA983DCBBCEE759C0DDC30B2F81C9";
    attribute INIT_0F of inst : label is "62CB53F0A2C3F0CC34D151F27E003DA32231CB1D6596491C5287AAEC34C7D8D3";
    attribute INIT_10 of inst : label is "3303030303C303C000003C3FFFFFFFFEC201F04F0C1C4E1C4F2D03C3205E70C8";
    attribute INIT_11 of inst : label is "492FAFF2FFFCBDB40003FCBFFF2D0033C3FC000000000000000000000C000C00";
    attribute INIT_12 of inst : label is "292ABE71D71EBCAA471CA8C5A924BC40C924AA4AA91CBC40D72F2A9201200048";
    attribute INIT_13 of inst : label is "24724BFC7291CBC91C91CC0C91324BD75E4DBCA8C9169249132ABCAA471691C7";
    attribute INIT_14 of inst : label is "D5350003000140501400000000014100000C5A45A4BFC5A91CBC75DBF075CBC7";
    attribute INIT_15 of inst : label is "00000140501000300014D53500034043443440300186100C004344344000D014";
    attribute INIT_16 of inst : label is "E391D579F558BA3FA7614AD2026680E668C0C202CC0000000000000014140000";
    attribute INIT_17 of inst : label is "49200491CAA472F5CBFF5E72D00B2FF4024000B2CB501A08AE8B51E42B06819B";
    attribute INIT_18 of inst : label is "4A8CA92AA31CAAF9F71DBCAA472AA4924724BC5A492A8C75C72F1F71CA8C72F2";
    attribute INIT_19 of inst : label is "CAA4BF075CBC91EBFC5A91CBC724924C0CAA924BC75C72F1CA8C592AA924AAF2";
    attribute INIT_1A of inst : label is "30004711C400000000051014400400000052050800004032A31032FF1CAA32F5";
    attribute INIT_1B of inst : label is "000015100144040000000004711C400C00100100010000155500001000100100";
    attribute INIT_1C of inst : label is "343F034BBF977579174228DF95C5FB4D066400302664212180B3420000220500";
    attribute INIT_1D of inst : label is "924A32F24924AA4A91CA92F9F76D000240000114000CD05214800AF8AED743F0";
    attribute INIT_1E of inst : label is "24A492DAA92A91691D72FDD5A91CBC92A924924AA91CBC71691D79CBC71D5A45";
    attribute INIT_1F of inst : label is "72AA4BC75DBF07AF1C91C92FF1CA4AAF247247303244CAAF5D7936DAA32A32A9";
    attribute INIT_20 of inst : label is "1035035000340B4B00100000110460004008502140040000000000C5A45A4BFC";
    attribute INIT_21 of inst : label is "000000004085002146000441000002C00B44000D010350350030001555003000";
    attribute INIT_22 of inst : label is "00335004608AAEA0A754108C1304C01BBA555EAAED4D715C75321210B3C00001";
    attribute INIT_23 of inst : label is "A4BD72A4A192476F2A39D5A92F2A920047204AA92FAFFC72FEB40003FF1CBD00";
    attribute INIT_24 of inst : label is "AA4BC79E7AF169245A4A869292F1691CAA4A869132F1D79D4CBC924592AA4724";
    attribute INIT_25 of inst : label is "15D400C00000691CAA4BFCAA91CBD7AFC9CBC916924BFC92A8CBC72A91CC0C72";
    attribute INIT_26 of inst : label is "30001050500001451000010505000300014D5350000000005050500500050010";
    attribute INIT_27 of inst : label is "131C000000000000000000030005D5001014014001050500000000054D535000";
    attribute INIT_28 of inst : label is "902EB8807D4D03688EB82B410D02709414ABE407D7955C2B8D55667D3D78B033";
    attribute INIT_29 of inst : label is "3084CB47DC0000001B549D938745C53DC88B6E4A0BE67D44CB6AD302C0DF6140";
    attribute INIT_2A of inst : label is "42EB804D5F27D857E2FACC024C093024C930DE69387DC520C9903084CB47DC90";
    attribute INIT_2B of inst : label is "08135F1F75EDBBBAD9959241F7143CBFEA955555FA550550E70741F240CD9C92";
    attribute INIT_2C of inst : label is "568B98C65431950C65431940C7C87CFB03B80A1331EFF1212121281751613231";
    attribute INIT_2D of inst : label is "414154051A855546A1800D1969AAA10101800D5428AA8AA940600155552595F9";
    attribute INIT_2E of inst : label is "6211800CA0007A95426546003684A441440001110444111060035A115068AA85";
    attribute INIT_2F of inst : label is "01C8CFF603E430C0153C3075FFFFFFD14E3D3FAE70E8CCC30A3CBD9111019005";
    attribute INIT_30 of inst : label is "3303030303C303C000003C3FFFFFFFFEC201F04F0C1C4E1C4F2D03C3205E70C8";
    attribute INIT_31 of inst : label is "492FAFF2FFFCBDB40003FCBFFF2D0033C3FC000000000000000000000C000C00";
    attribute INIT_32 of inst : label is "292ABE71D71EBCAA471CA8C5A924BC40C924AA4AA91CBC40D72F2A9201200048";
    attribute INIT_33 of inst : label is "24724BFC7291CBC91C91CC0C91324BD75E4DBCA8C9169249132ABCAA471691C7";
    attribute INIT_34 of inst : label is "D5350003000140501400000000014100000C5A45A4BFC5A91CBC75DBF075CBC7";
    attribute INIT_35 of inst : label is "00000140501000300014D53500034043443440300186100C004344344000D014";
    attribute INIT_36 of inst : label is "E391D579F558BA3FA7614AD2026680E668C0C202CC0000000000000014140000";
    attribute INIT_37 of inst : label is "49200491CAA472F5CBFF5E72D00B2FF4024000B2CB501A08AE8B51E42B06819B";
    attribute INIT_38 of inst : label is "4A8CA92AA31CAAF9F71DBCAA472AA4924724BC5A492A8C75C72F1F71CA8C72F2";
    attribute INIT_39 of inst : label is "CAA4BF075CBC91EBFC5A91CBC724924C0CAA924BC75C72F1CA8C592AA924AAF2";
    attribute INIT_3A of inst : label is "30004711C400000000051014400400000052050800004032A31032FF1CAA32F5";
    attribute INIT_3B of inst : label is "000015100144040000000004711C400C00100100010000155500001000100100";
    attribute INIT_3C of inst : label is "343F034BBF977579174228DF95C5FB4D066400302664212180B3420000220500";
    attribute INIT_3D of inst : label is "924A32F24924AA4A91CA92F9F76D000240000114000CD05214800AF8AED743F0";
    attribute INIT_3E of inst : label is "24A492DAA92A91691D72FDD5A91CBC92A924924AA91CBC71691D79CBC71D5A45";
    attribute INIT_3F of inst : label is "72AA4BC75DBF07AF1C91C92FF1CA4AAF247247303244CAAF5D7936DAA32A32A9";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFC702860B17CCFFFFFFFFFFFF1506801E89BC3F016D0C1808";
    attribute INIT_01 of inst : label is "FFFFFFFFBBA665E140F009514C0041CFFFFFFFFF10502F80C287A8600413B100";
    attribute INIT_02 of inst : label is "FFFFFFFFF21AD303FFFFFFFF20386983FFFFFFFFFFFF32600C4F1A51FFFF0010";
    attribute INIT_03 of inst : label is "31320121FFFF9487086084C730409041FFFFFFFF045088C020C215023030902A";
    attribute INIT_04 of inst : label is "30FF0FF1DFDD0DFB7D0CCF0F1011111121111110111111311111113030213202";
    attribute INIT_05 of inst : label is "C30F33F30F33F37077DCBCC2FC2FFB1DFDD0DFB6D0CCF0F0371CCFCB37307F1F";
    attribute INIT_06 of inst : label is "C0CCCCC2DF71FF07F07FECB8F7C0DCF33F0CFCC3FCFFC1FC1FC38F7C0CFF0333";
    attribute INIT_07 of inst : label is "FFECFFFBC1EF71FF0FB0D3DFF07BDC7FFF0BB0D3DFF07BEFF1FFDF4373C0CCCC";
    attribute INIT_08 of inst : label is "7F43B0E3EF47F47F43F0E3DFFC1EF73FF0FB1D3EFF0773FFEFF0F71D3EFF077D";
    attribute INIT_09 of inst : label is "0FFC30333C3DD0DFB7D0CCF0FED0CC743373343373343F43F1E3DEF4330F47F4";
    attribute INIT_0A of inst : label is "C3C3DEF4330F0F7437EDB4333C3C3DD0DFB7D0CCF0FFC70331C3DD0DFB6D0CCF";
    attribute INIT_0B of inst : label is "DCB07707F2D3CCECB07707F2D3CCFCB07707F2D3CCCCB07707F2D3C3F7FFAD0C";
    attribute INIT_0C of inst : label is "75555777AAAEAABAAAFFFFFFFFFEBEBFAFAFFE96BFA5AFD557F555FF07F0D3CC";
    attribute INIT_0D of inst : label is "087021C8B03F2036C20C0FC809C20C0FC80DC20C0FC80DB083CCEA957F775555";
    attribute INIT_0E of inst : label is "83E0D0063D660331F2C21023C430C0C023EF30A310A0ECC73F082F086459080C";
    attribute INIT_0F of inst : label is "450021C2080DC3E06650026A702A6F0427381C010410010012C3B4C166600E1F";
    attribute INIT_10 of inst : label is "3303030303C303C000003C3FFFFFFFFD0DC10C30CDCC1DCC1C5B4033205F7430";
    attribute INIT_11 of inst : label is "8A1D1FD1FFF474755557F47FFD1D5573C3FC000000000000000000000C000C00";
    attribute INIT_12 of inst : label is "2A2AF492492474AA8924AB4BAA2874804A28AA8AAA247480591D2AA256255589";
    attribute INIT_13 of inst : label is "289287F492A2474A24A24958A2128749248474AB4A2EA28A212AF4AA892EA249";
    attribute INIT_14 of inst : label is "000000000000040100000000000010001084BA8BA87F0BAA24749247FC924749";
    attribute INIT_15 of inst : label is "0000000401000000000000000000000000000000004100000000000000000000";
    attribute INIT_16 of inst : label is "E291DD797550BA013C8F62148044AA044040CB23660000000000000401000000";
    attribute INIT_17 of inst : label is "8A2558A24AA891D247FD2491D5551FF555555551CB501A08AE8B51481104411B";
    attribute INIT_18 of inst : label is "8AB4AA2AAD24ABD2492474AA892AA8A2892874BA8A2AB492491D24924AB491D2";
    attribute INIT_19 of inst : label is "4AA87FC92474A247F4BAA2474928A28958AAA287492495D24AB4BA2AAA28ABD2";
    attribute INIT_1A of inst : label is "000000000000000000000000000000000000000000008012AD2011FC24AAD1D2";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000001000100100041001000001001000";
    attribute INIT_1C of inst : label is "8410040ABF877D7857422814B62C44110446AA9A84441032C8D9C00000000000";
    attribute INIT_1D of inst : label is "A28AD1D28A28AA8AA24AA1D2491D555555555625555CD01294A02AFAAED74210";
    attribute INIT_1E of inst : label is "28A8A1FAAA2AA2EA2491D24BAA2474A2AA28A28AAA247492EA2492474924BA8B";
    attribute INIT_1F of inst : label is "92AA8749247FC91D24A24A1FD24A8ABD2892892562884ABD249211FAAD2AD2AA";
    attribute INIT_20 of inst : label is "0000000000000000000000010040000000000000000000000002004BA8BA87F0";
    attribute INIT_21 of inst : label is "0000000000000000000000100000100000000000000000000000000410000000";
    attribute INIT_22 of inst : label is "55737084688ABE200F4400982509425BFA555EAEE15F57D5C5610328D98C0000";
    attribute INIT_23 of inst : label is "A87492A8AFA2891D2AD24BAA1D2AA25589258AAA1D1FF491F4755557FD247D55";
    attribute INIT_24 of inst : label is "AA87492491D2EA28BA8ABEA2A1D2EA24AA8ABEA211D249248474A28BA2AA8928";
    attribute INIT_25 of inst : label is "000000000200EA24AA87F0AAA247491FF2474A2EA287F4A2AB47492AA2495892";
    attribute INIT_26 of inst : label is "0000010100100041001000101000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0328000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "6672200271ED416A8AB8AB450581505415ABA5175795DD2F835FE6C5815CD891";
    attribute INIT_29 of inst : label is "346228D71600000024171108002565CE1DD048820C3071E1948C1908C2DC5A98";
    attribute INIT_2A of inst : label is "4412326526A71E8CB12CDC54665199466B32CF499A716475233A352228D7163A";
    attribute INIT_2B of inst : label is "4C90891C370D03C8F71B2009C5AF31D5554015555946D568C6806DC7A0DCA0E8";
    attribute INIT_2C of inst : label is "546F048CC6233188CC6233005BC6D96033265359B82FF183818380985A08B3FE";
    attribute INIT_2D of inst : label is "5FDFFFEA8AAA82A2A3333C0AAAAAA444D3333D5FEBA0BA0000CCCD5555F55D35";
    attribute INIT_2E of inst : label is "AE63333F8D55CA88A88A8CCCFABC00EA8D13B44ED13B44ECCCCFAAFFF3A9AA95";
    attribute INIT_2F of inst : label is "AFAA2AA8A804450A45408100FFFFFF8120FCBC328E0F80181230FE8C4466AB9A";
    attribute INIT_30 of inst : label is "3303030303C303C000003C3FFFFFFFFD0DC10C30CDCC1DCC1C5B4033205F7430";
    attribute INIT_31 of inst : label is "8A1D1FD1FFF474755557F47FFD1D5573C3FC000000000000000000000C000C00";
    attribute INIT_32 of inst : label is "2A2AF492492474AA8924AB4BAA2874804A28AA8AAA247480591D2AA256255589";
    attribute INIT_33 of inst : label is "289287F492A2474A24A24958A2128749248474AB4A2EA28A212AF4AA892EA249";
    attribute INIT_34 of inst : label is "000000000000040100000000000010001084BA8BA87F0BAA24749247FC924749";
    attribute INIT_35 of inst : label is "0000000401000000000000000000000000000000004100000000000000000000";
    attribute INIT_36 of inst : label is "E291DD797550BA013C8F62148044AA044040CB23660000000000000401000000";
    attribute INIT_37 of inst : label is "8A2558A24AA891D247FD2491D5551FF555555551CB501A08AE8B51481104411B";
    attribute INIT_38 of inst : label is "8AB4AA2AAD24ABD2492474AA892AA8A2892874BA8A2AB492491D24924AB491D2";
    attribute INIT_39 of inst : label is "4AA87FC92474A247F4BAA2474928A28958AAA287492495D24AB4BA2AAA28ABD2";
    attribute INIT_3A of inst : label is "000000000000000000000000000000000000000000008012AD2011FC24AAD1D2";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000001000100100041001000001001000";
    attribute INIT_3C of inst : label is "8410040ABF877D7857422814B62C44110446AA9A84441032C8D9C00000000000";
    attribute INIT_3D of inst : label is "A28AD1D28A28AA8AA24AA1D2491D555555555625555CD01294A02AFAAED74210";
    attribute INIT_3E of inst : label is "28A8A1FAAA2AA2EA2491D24BAA2474A2AA28A28AAA247492EA2492474924BA8B";
    attribute INIT_3F of inst : label is "92AA8749247FC91D24A24A1FD24A8ABD2892892562884ABD249211FAAD2AD2AA";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFD9D079D01001FFFFFFFFFFFF49D0037210C301F771F12743";
    attribute INIT_01 of inst : label is "FFFFFFFF212BCE460C3073AF03BDAC0DFFFFFFFF8E840874F61C079DEBC036B4";
    attribute INIT_02 of inst : label is "FFFFFFFF02DE3071FFFFFFFF2C072EF4FFFFFFFFFFFF008D7018C511FFFF0000";
    attribute INIT_03 of inst : label is "BA9998A9FFFF3A1840AD2B100EF430BCFFFFFFFF70033D1DBF7E49D033AFE353";
    attribute INIT_04 of inst : label is "30F70F78DFCC0CF36C0CE70F98999999B999999B999999A999999A9ABB999998";
    attribute INIT_05 of inst : label is "C30F33F30F33F33037CE74C3DC3DF39DFCC0CF36C0CE70F0338CCCE33330378D";
    attribute INIT_06 of inst : label is "C0CCCCC3DF39DF037037CE78F7C0CE33339CFCC3DE37C0DC0DE78F7C0DC70339";
    attribute INIT_07 of inst : label is "F7CE33F7C2CF38EF0739D3CF70F7CE37F70379E3CF70F7CF78CFDF0339C0CCCC";
    attribute INIT_08 of inst : label is "37037AD3DF033037037AD3DFDC2CF38EF0738D3CF70F78DFCF70378E3CF70F7C";
    attribute INIT_09 of inst : label is "0FCFF0338C3CC0CF36C0CE70FCC0CEB033333033333037037AD3DDB033AF0330";
    attribute INIT_0A of inst : label is "EBC3DDB033AF0F3033CDB0339C3C3CC0CF36C0CE70FCFF0338C3CC0CF36C0CE7";
    attribute INIT_0B of inst : label is "CE70370379E3CCCE70370379E3CCCE70370379E3CCDE70370379E3C3F3F36C0C";
    attribute INIT_0C of inst : label is "30000333000C003AAAC0003F0F0EAAAB0000FFFFF5555EAAAB0000F70379E3CC";
    attribute INIT_0D of inst : label is "79C9E7398D0007B033434001E833434001E033434001E00CD0CCC00033330000";
    attribute INIT_0E of inst : label is "10443A68B23700340E509D0EE774350020C0CC20753D8335AC533451C1DF9152";
    attribute INIT_0F of inst : label is "8899BC1483501445747A9375AE007081447370000000000000F03CF7744BEC71";
    attribute INIT_10 of inst : label is "3303030303C303C000003C3FFFFFFFFCFCB340F4000CE40CE5DF0D00285F899A";
    attribute INIT_11 of inst : label is "CF3F3FF3FFFCFCFFFFFFFCFFFF3FFFF7C3FC000000000000000000000C000C00";
    attribute INIT_12 of inst : label is "3F3FFCF3CF3CFCFFCF3CFFCFFF3CFCFFCF3CFFCFFF3CFCFFCF3F3FF3FF3FFFCF";
    attribute INIT_13 of inst : label is "3CF3CFFCF3F3CFCF3CF3CFFCF3F3CFCF3CFCFCFFCF3FF3CF3F3FFCFFCF3FF3CF";
    attribute INIT_14 of inst : label is "00000000000000000000000000000000004CFFCFFCFFCFFF3CFCF3CFFCF3CFCF";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "F2D4DD7D7552AA849D27892240003F0005995444030000000000000000000000";
    attribute INIT_17 of inst : label is "CF3FFCF3CFFCF3F3CFFF3CF3FFFF3FFFFFFFFFF3DB501A8AAAAA55280A0280AB";
    attribute INIT_18 of inst : label is "CFFCFF3FFF3CFFF3CF3CFCFFCF3FFCF3CF3CFCFFCF3FFCF3CF3F3CF3CFFCF3F3";
    attribute INIT_19 of inst : label is "CFFCFFCF3CFCF3CFFCFFF3CFCF3CF3CFFCFFF3CFCF3CF3F3CFFCFF3FFF3CFFF3";
    attribute INIT_1A of inst : label is "000000000000000000000000000000000000000000004033FF3FF3FF3CFFF3F3";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "280A028AFFC57D7C4550A802709F24C9000000F0000166551100C00000000000";
    attribute INIT_1D of inst : label is "F3CFF3F3CF3CFFCFF3CFF3F3CF3FFFFFFFFFFF3FFFFDD01084A022FE2AF540A0";
    attribute INIT_1E of inst : label is "3CFCF3FFFF3FF3FF3CF3F3CFFF3CFCF3FF3CF3CFFF3CFCF3FF3CF3CFCF3CFFCF";
    attribute INIT_1F of inst : label is "F3FFCFCF3CFFCF3F3CF3CF3FF3CFCFFF3CF3CF3FF3CFCFFF3CF3F3FFFF3FF3FF";
    attribute INIT_20 of inst : label is "000000000000000000000000000000000000000000000000000100CFFCFFCFFC";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "FFF6748568AABA200D4400240902409AEA5D5FAEF12348D204866551001C0000";
    attribute INIT_23 of inst : label is "FCFCF3FCFFF3CF3F3FF3CFFF3F3FF3FFCF3FCFFF3F3FFCF3FCFFFFFFFF3CFFFF";
    attribute INIT_24 of inst : label is "FFCFCF3CF3F3FF3CFFCFFFF3F3F3FF3CFFCFFFF3F3F3CF3CFCFCF3CFF3FFCF3C";
    attribute INIT_25 of inst : label is "000000000100FF3CFFCFFCFFF3CFCF3FF3CFCF3FF3CFFCF3FFCFCF3FF3CFFCF3";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "655C000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "049AABD0AE49416A0ABAAB550240902409A3B51377D7DD2EA12348E208810106";
    attribute INIT_29 of inst : label is "0004550AE000000030EF33D101BECBCF42E220F3F904AE8EE2234340C0EBA320";
    attribute INIT_2A of inst : label is "8888FF47375AE4FD004383CF443D10F44D0094FD15AE0FB888F20004550AE0F2";
    attribute INIT_2B of inst : label is "63E7F1E33BCE336233F0E042BB033400000000000C3ACCCF4A01ACD03C0C240F";
    attribute INIT_2C of inst : label is "EBCB31C04C70131C04C701000A180C3D00F03D11110F740704070FE383F00D33";
    attribute INIT_2D of inst : label is "511115656555695953333EA555555AAA53333EA5555A55AA54CCCEAAAA4E2A46";
    attribute INIT_2E of inst : label is "5593333D66AA656656654CCCF956A8EA8E955A556955A554CCCFA55553565555";
    attribute INIT_2F of inst : label is "155541550155555055551555FFFFFF3E84300D009442C05100343D66AA995565";
    attribute INIT_30 of inst : label is "3303030303C303C000003C3FFFFFFFFCFCB340F4000CE40CE5DF0D00285F899A";
    attribute INIT_31 of inst : label is "CF3F3FF3FFFCFCFFFFFFFCFFFF3FFFF7C3FC000000000000000000000C000C00";
    attribute INIT_32 of inst : label is "3F3FFCF3CF3CFCFFCF3CFFCFFF3CFCFFCF3CFFCFFF3CFCFFCF3F3FF3FF3FFFCF";
    attribute INIT_33 of inst : label is "3CF3CFFCF3F3CFCF3CF3CFFCF3F3CFCF3CFCFCFFCF3FF3CF3F3FFCFFCF3FF3CF";
    attribute INIT_34 of inst : label is "00000000000000000000000000000000004CFFCFFCFFCFFF3CFCF3CFFCF3CFCF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "F2D4DD7D7552AA849D27892240003F0005995444030000000000000000000000";
    attribute INIT_37 of inst : label is "CF3FFCF3CFFCF3F3CFFF3CF3FFFF3FFFFFFFFFF3DB501A8AAAAA55280A0280AB";
    attribute INIT_38 of inst : label is "CFFCFF3FFF3CFFF3CF3CFCFFCF3FFCF3CF3CFCFFCF3FFCF3CF3F3CF3CFFCF3F3";
    attribute INIT_39 of inst : label is "CFFCFFCF3CFCF3CFFCFFF3CFCF3CF3CFFCFFF3CFCF3CF3F3CFFCFF3FFF3CFFF3";
    attribute INIT_3A of inst : label is "000000000000000000000000000000000000000000004033FF3FF3FF3CFFF3F3";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "280A028AFFC57D7C4550A802709F24C9000000F0000166551100C00000000000";
    attribute INIT_3D of inst : label is "F3CFF3F3CF3CFFCFF3CFF3F3CF3FFFFFFFFFFF3FFFFDD01084A022FE2AF540A0";
    attribute INIT_3E of inst : label is "3CFCF3FFFF3FF3FF3CF3F3CFFF3CFCF3FF3CF3CFFF3CFCF3FF3CF3CFCF3CFFCF";
    attribute INIT_3F of inst : label is "F3FFCFCF3CFFCF3F3CF3CF3FF3CFCFFF3CF3CF3FF3CFCFFF3CF3F3FFFF3FF3FF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
