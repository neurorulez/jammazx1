library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity berzerk_program1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of berzerk_program1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"40",X"3E",X"FF",X"32",X"5E",X"40",X"AF",X"32",X"66",X"40",X"01",X"0C",X"00",X"11",X"07",X"40",
		X"21",X"4D",X"10",X"ED",X"B0",X"CD",X"A5",X"1E",X"E1",X"F5",X"22",X"64",X"40",X"CD",X"39",X"10",
		X"CD",X"C2",X"20",X"11",X"5F",X"40",X"EB",X"CD",X"2E",X"10",X"F1",X"C3",X"29",X"05",X"06",X"03",
		X"7E",X"36",X"00",X"23",X"12",X"13",X"10",X"F8",X"C9",X"E5",X"2A",X"64",X"40",X"54",X"5D",X"29",
		X"19",X"29",X"19",X"11",X"53",X"31",X"19",X"22",X"64",X"40",X"7C",X"E1",X"C9",X"01",X"14",X"28",
		X"1E",X"74",X"01",X"08",X"01",X"20",X"04",X"00",X"08",X"01",X"8F",X"18",X"05",X"8F",X"1A",X"14",
		X"02",X"9F",X"1A",X"02",X"94",X"16",X"0A",X"92",X"16",X"02",X"BF",X"14",X"8F",X"09",X"9F",X"1A",
		X"8F",X"14",X"8F",X"09",X"BF",X"02",X"BF",X"14",X"8F",X"14",X"8F",X"0A",X"94",X"0A",X"9F",X"02",
		X"CF",X"14",X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"9F",X"12",
		X"04",X"9F",X"16",X"9F",X"14",X"00",X"FF",X"FF",X"FF",X"CD",X"1A",X"11",X"CD",X"50",X"0D",X"CD",
		X"A2",X"0C",X"CD",X"A2",X"20",X"CD",X"D5",X"30",X"CD",X"17",X"12",X"2E",X"12",X"57",X"12",X"41",
		X"12",X"6F",X"12",X"21",X"00",X"4B",X"CD",X"11",X"11",X"21",X"6E",X"40",X"3E",X"01",X"32",X"00",
		X"40",X"11",X"40",X"3F",X"D5",X"E5",X"7E",X"23",X"B6",X"23",X"B6",X"E1",X"E5",X"20",X"04",X"E1",
		X"D1",X"18",X"35",X"21",X"00",X"40",X"06",X"02",X"CD",X"53",X"2E",X"13",X"E1",X"06",X"06",X"CD",
		X"5D",X"2E",X"13",X"AF",X"4E",X"CD",X"EE",X"2D",X"13",X"23",X"4E",X"CD",X"EE",X"2D",X"13",X"23",
		X"4E",X"CD",X"EE",X"2D",X"23",X"D1",X"7A",X"C6",X"0C",X"57",X"3A",X"00",X"40",X"C6",X"01",X"27",
		X"32",X"00",X"40",X"FE",X"11",X"C2",X"C4",X"10",X"21",X"00",X"5B",X"CD",X"11",X"11",X"21",X"80",
		X"5D",X"3E",X"FF",X"06",X"40",X"77",X"23",X"10",X"FC",X"C9",X"21",X"00",X"81",X"01",X"00",X"07",
		X"CD",X"40",X"06",X"F3",X"ED",X"73",X"00",X"40",X"31",X"00",X"60",X"06",X"E0",X"11",X"00",X"00",
		X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",X"D5",
		X"10",X"EE",X"ED",X"7B",X"00",X"40",X"FB",X"DB",X"4A",X"CB",X"7F",X"20",X"0D",X"3A",X"07",X"40",
		X"FE",X"02",X"20",X"06",X"3E",X"08",X"32",X"22",X"40",X"C9",X"AF",X"32",X"22",X"40",X"C9",X"CD",
		X"8E",X"2D",X"90",X"0C",X"BE",X"1F",X"31",X"39",X"38",X"32",X"20",X"53",X"54",X"45",X"52",X"4E",
		X"20",X"45",X"6C",X"65",X"63",X"74",X"72",X"6F",X"6E",X"69",X"63",X"73",X"2C",X"20",X"49",X"6E",
		X"63",X"2E",X"00",X"C9",X"CD",X"07",X"12",X"CD",X"B5",X"0C",X"28",X"21",X"3D",X"28",X"0F",X"CD",
		X"C4",X"0D",X"CD",X"17",X"12",X"BE",X"12",X"08",X"13",X"E5",X"12",X"25",X"13",X"C9",X"CD",X"C4",
		X"0D",X"CD",X"17",X"12",X"7E",X"12",X"08",X"13",X"A0",X"12",X"25",X"13",X"C9",X"CD",X"BB",X"0D",
		X"CD",X"17",X"12",X"39",X"13",X"69",X"13",X"4C",X"13",X"80",X"13",X"21",X"A2",X"30",X"22",X"9A",
		X"F8",X"C9",X"CD",X"07",X"12",X"DB",X"60",X"E6",X"0F",X"28",X"26",X"47",X"E6",X"08",X"4F",X"78",
		X"E6",X"07",X"81",X"27",X"32",X"00",X"40",X"11",X"58",X"BE",X"21",X"00",X"40",X"06",X"02",X"CD",
		X"53",X"2E",X"CD",X"8E",X"2D",X"90",X"68",X"BE",X"30",X"30",X"30",X"20",X"3D",X"20",X"7E",X"00",
		X"C9",X"CD",X"8E",X"2D",X"90",X"48",X"BE",X"4E",X"6F",X"20",X"45",X"78",X"74",X"72",X"61",X"20",
		X"4C",X"69",X"76",X"65",X"73",X"00",X"C9",X"21",X"C0",X"5B",X"01",X"C0",X"02",X"AF",X"77",X"23",
		X"0D",X"C2",X"0E",X"12",X"10",X"F8",X"C9",X"E1",X"54",X"5D",X"01",X"08",X"00",X"09",X"E5",X"EB",
		X"DB",X"60",X"E6",X"C0",X"07",X"07",X"07",X"4F",X"09",X"7E",X"23",X"66",X"6F",X"E9",X"CD",X"8E",
		X"2D",X"90",X"50",X"2A",X"48",X"69",X"67",X"68",X"20",X"53",X"63",X"6F",X"72",X"65",X"73",X"00",
		X"C9",X"CD",X"8E",X"2D",X"90",X"44",X"2A",X"4D",X"65",X"69",X"6C",X"6C",X"65",X"75",X"72",X"20",
		X"53",X"63",X"6F",X"72",X"65",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"3C",X"2A",X"48",X"6F",X"65",
		X"63",X"68",X"73",X"74",X"65",X"72",X"20",X"47",X"65",X"62",X"6E",X"69",X"73",X"00",X"C9",X"CD",
		X"8E",X"2D",X"90",X"60",X"2A",X"52",X"65",X"63",X"6F",X"72",X"64",X"73",X"00",X"C9",X"CD",X"8E",
		X"2D",X"90",X"14",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",X"20",X"50",X"6C",X"61",X"79",X"65",
		X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"20",X"42",X"75",X"74",X"74",X"6F",X"6E",X"00",X"C9",
		X"CD",X"8E",X"2D",X"90",X"24",X"BE",X"50",X"6F",X"75",X"73",X"73",X"65",X"72",X"20",X"62",X"6F",
		X"75",X"74",X"6F",X"6E",X"20",X"73",X"74",X"61",X"72",X"74",X"20",X"31",X"00",X"C9",X"CD",X"8E",
		X"2D",X"90",X"04",X"BE",X"50",X"75",X"73",X"68",X"20",X"31",X"20",X"6F",X"72",X"20",X"32",X"20",
		X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"20",X"42",X"75",X"74",
		X"74",X"6F",X"6E",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"10",X"BE",X"50",X"6F",X"75",X"73",X"73",
		X"65",X"72",X"20",X"62",X"6F",X"75",X"74",X"6F",X"6E",X"20",X"73",X"74",X"61",X"72",X"74",X"20",
		X"31",X"20",X"6F",X"75",X"20",X"32",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"20",X"BE",X"53",X"74",
		X"61",X"72",X"74",X"6B",X"6E",X"6F",X"65",X"70",X"66",X"65",X"20",X"64",X"72",X"75",X"65",X"63",
		X"6B",X"65",X"6E",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"44",X"BE",X"50",X"75",X"6C",X"73",X"61",
		X"72",X"20",X"53",X"74",X"61",X"72",X"74",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"58",X"BE",X"49",
		X"6E",X"73",X"65",X"72",X"74",X"20",X"43",X"6F",X"69",X"6E",X"00",X"C9",X"CD",X"8E",X"2D",X"90",
		X"30",X"BE",X"49",X"6E",X"74",X"72",X"6F",X"64",X"75",X"69",X"72",X"65",X"20",X"6C",X"61",X"20",
		X"6D",X"6F",X"6E",X"6E",X"61",X"69",X"65",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"48",X"BE",X"4D",
		X"75",X"6E",X"7A",X"65",X"20",X"65",X"69",X"6E",X"77",X"65",X"72",X"66",X"65",X"6E",X"00",X"C9",
		X"CD",X"8E",X"2D",X"90",X"48",X"BE",X"50",X"6F",X"6E",X"67",X"61",X"20",X"6C",X"61",X"20",X"6D",
		X"6F",X"6E",X"65",X"64",X"61",X"00",X"C9",X"D3",X"4D",X"F3",X"F5",X"DB",X"4E",X"1F",X"38",X"6C",
		X"D3",X"4C",X"E5",X"C5",X"21",X"59",X"40",X"7E",X"23",X"46",X"A8",X"4F",X"DB",X"49",X"2F",X"77",
		X"2B",X"70",X"A1",X"E6",X"C0",X"2B",X"CB",X"7F",X"28",X"01",X"34",X"87",X"20",X"F7",X"21",X"A0",
		X"F8",X"CB",X"3E",X"21",X"C8",X"F8",X"35",X"F2",X"E3",X"13",X"36",X"3C",X"0E",X"08",X"CD",X"0F",
		X"08",X"3A",X"5E",X"40",X"B7",X"0E",X"07",X"CC",X"0F",X"08",X"21",X"A1",X"F8",X"7E",X"B7",X"28",
		X"02",X"3D",X"77",X"CD",X"B5",X"0C",X"2E",X"00",X"B7",X"28",X"08",X"FE",X"01",X"2E",X"01",X"28",
		X"02",X"2E",X"03",X"DB",X"49",X"2F",X"A5",X"6F",X"3A",X"56",X"40",X"B5",X"32",X"56",X"40",X"CA",
		X"07",X"14",X"CB",X"7F",X"CA",X"47",X"05",X"C1",X"E1",X"C3",X"A1",X"14",X"FD",X"E5",X"DD",X"E5",
		X"E5",X"D5",X"C5",X"08",X"F5",X"21",X"00",X"00",X"22",X"C1",X"F8",X"22",X"C3",X"F8",X"22",X"C5",
		X"F8",X"21",X"C7",X"F8",X"CB",X"06",X"06",X"03",X"2A",X"BF",X"F8",X"DA",X"47",X"14",X"21",X"AD",
		X"40",X"22",X"C5",X"F8",X"CD",X"B0",X"14",X"CD",X"0E",X"0F",X"21",X"AD",X"40",X"CB",X"66",X"C4",
		X"30",X"0F",X"2A",X"BF",X"F8",X"06",X"02",X"C5",X"CD",X"B0",X"14",X"C1",X"2A",X"BD",X"F8",X"EB",
		X"78",X"87",X"21",X"BF",X"F8",X"85",X"6F",X"7C",X"CE",X"00",X"67",X"73",X"23",X"72",X"EB",X"11",
		X"0E",X"00",X"19",X"11",X"FD",X"41",X"7D",X"BB",X"C2",X"70",X"14",X"7C",X"BA",X"CA",X"7A",X"14",
		X"7E",X"E6",X"80",X"28",X"EA",X"10",X"D0",X"C3",X"7D",X"14",X"21",X"BB",X"40",X"22",X"BF",X"F8",
		X"CD",X"99",X"09",X"2A",X"C5",X"F8",X"CD",X"25",X"15",X"2A",X"C3",X"F8",X"CD",X"25",X"15",X"2A",
		X"C1",X"F8",X"CD",X"25",X"15",X"CD",X"61",X"15",X"F1",X"08",X"C1",X"D1",X"E1",X"DD",X"E1",X"FD",
		X"E1",X"3E",X"01",X"D3",X"4F",X"D3",X"4C",X"3E",X"3F",X"ED",X"47",X"ED",X"5E",X"F1",X"FB",X"C9",
		X"22",X"BD",X"F8",X"FD",X"2A",X"BD",X"F8",X"CB",X"46",X"CA",X"D1",X"14",X"CB",X"86",X"23",X"7E",
		X"D3",X"4B",X"23",X"5E",X"23",X"56",X"23",X"7E",X"23",X"66",X"6F",X"CD",X"6F",X"15",X"2A",X"BD",
		X"F8",X"CB",X"4E",X"C8",X"CB",X"8E",X"11",X"09",X"00",X"19",X"5E",X"23",X"23",X"56",X"23",X"06",
		X"90",X"EB",X"CD",X"B6",X"2D",X"FD",X"77",X"01",X"EB",X"7E",X"23",X"66",X"6F",X"7E",X"23",X"66",
		X"6F",X"23",X"7E",X"2B",X"CB",X"7F",X"28",X"13",X"E6",X"7F",X"47",X"4E",X"23",X"23",X"EB",X"3A",
		X"22",X"40",X"B7",X"CA",X"09",X"15",X"ED",X"42",X"3E",X"09",X"EB",X"FD",X"75",X"04",X"FD",X"74",
		X"05",X"FD",X"73",X"02",X"FD",X"72",X"03",X"CD",X"6F",X"15",X"2A",X"BD",X"F8",X"DB",X"4E",X"CB",
		X"7F",X"C8",X"CB",X"EE",X"C9",X"22",X"BD",X"F8",X"CB",X"56",X"C8",X"E5",X"FD",X"E1",X"11",X"06",
		X"00",X"19",X"7E",X"23",X"35",X"C0",X"77",X"23",X"7E",X"23",X"86",X"77",X"23",X"7E",X"23",X"86",
		X"77",X"23",X"5E",X"23",X"56",X"13",X"13",X"EB",X"7E",X"23",X"B6",X"C2",X"54",X"15",X"23",X"7E",
		X"23",X"66",X"6F",X"3E",X"2B",X"EB",X"72",X"2B",X"73",X"3E",X"03",X"2A",X"BD",X"F8",X"B6",X"77",
		X"C9",X"21",X"03",X"80",X"06",X"18",X"7E",X"B7",X"28",X"01",X"35",X"23",X"10",X"F8",X"C9",X"06",
		X"00",X"7E",X"23",X"3D",X"CA",X"AB",X"15",X"3A",X"22",X"40",X"B7",X"7E",X"23",X"C2",X"95",X"15",
		X"01",X"1E",X"00",X"EB",X"08",X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"23",X"70",X"08",X"09",
		X"3D",X"C2",X"84",X"15",X"C9",X"01",X"E2",X"FF",X"EB",X"08",X"1A",X"13",X"77",X"2B",X"1A",X"13",
		X"77",X"2B",X"36",X"00",X"08",X"09",X"3D",X"C2",X"99",X"15",X"C9",X"3A",X"22",X"40",X"B7",X"7E",
		X"23",X"C2",X"C5",X"15",X"01",X"1F",X"00",X"EB",X"08",X"1A",X"13",X"77",X"23",X"70",X"08",X"09",
		X"3D",X"C2",X"B8",X"15",X"C9",X"01",X"E1",X"FF",X"EB",X"08",X"1A",X"13",X"77",X"2B",X"36",X"00",
		X"08",X"09",X"3D",X"C2",X"C9",X"15",X"C9",X"51",X"C5",X"D5",X"DD",X"6E",X"0C",X"DD",X"66",X"0D",
		X"5E",X"23",X"56",X"EB",X"57",X"23",X"7E",X"4F",X"CB",X"3F",X"C6",X"01",X"5F",X"DD",X"66",X"0B",
		X"DD",X"6E",X"09",X"CB",X"5A",X"CA",X"0E",X"16",X"E5",X"79",X"C6",X"03",X"84",X"67",X"D5",X"1E",
		X"05",X"CD",X"56",X"16",X"D1",X"E1",X"CA",X"25",X"16",X"CB",X"9A",X"C3",X"25",X"16",X"CB",X"52",
		X"CA",X"25",X"16",X"E5",X"3E",X"FD",X"84",X"67",X"D5",X"1E",X"05",X"CD",X"56",X"16",X"D1",X"E1",
		X"CA",X"25",X"16",X"CB",X"92",X"CB",X"4A",X"CA",X"3D",X"16",X"E5",X"3E",X"0B",X"85",X"6F",X"D5",
		X"CD",X"67",X"16",X"D1",X"E1",X"CA",X"52",X"16",X"CB",X"8A",X"C3",X"52",X"16",X"CB",X"42",X"CA",
		X"52",X"16",X"E5",X"3E",X"FD",X"85",X"6F",X"D5",X"CD",X"67",X"16",X"D1",X"E1",X"CA",X"52",X"16",
		X"CB",X"82",X"7A",X"D1",X"C1",X"C9",X"2D",X"1C",X"CD",X"78",X"16",X"C0",X"08",X"7D",X"C6",X"02",
		X"6F",X"08",X"1D",X"C2",X"58",X"16",X"C9",X"25",X"1C",X"CD",X"78",X"16",X"C0",X"08",X"7C",X"C6",
		X"02",X"67",X"08",X"1D",X"C2",X"69",X"16",X"C9",X"E5",X"CD",X"B4",X"2D",X"E6",X"0F",X"CB",X"5F",
		X"CA",X"85",X"16",X"EE",X"0F",X"EE",X"07",X"F3",X"D3",X"4B",X"CB",X"AC",X"7E",X"32",X"00",X"60",
		X"FB",X"3A",X"00",X"40",X"E6",X"01",X"E1",X"C9",X"7D",X"D6",X"08",X"1E",X"00",X"FE",X"30",X"38",
		X"0E",X"1E",X"06",X"FE",X"60",X"38",X"08",X"1E",X"0C",X"FE",X"90",X"38",X"02",X"1E",X"12",X"7C",
		X"D6",X"08",X"1D",X"D6",X"28",X"1C",X"30",X"FB",X"EB",X"01",X"26",X"40",X"26",X"00",X"09",X"7E",
		X"EB",X"C9",X"AF",X"32",X"A0",X"F8",X"21",X"FD",X"41",X"01",X"92",X"01",X"C3",X"40",X"06",X"FD",
		X"E5",X"DD",X"E5",X"E5",X"D5",X"C5",X"F5",X"CD",X"95",X"17",X"21",X"00",X"00",X"39",X"01",X"10",
		X"00",X"ED",X"B0",X"21",X"FD",X"41",X"46",X"23",X"7E",X"34",X"B8",X"20",X"02",X"36",X"00",X"7E",
		X"FE",X"01",X"28",X"F4",X"21",X"A0",X"F8",X"7E",X"B7",X"20",X"0D",X"36",X"01",X"3A",X"FD",X"41",
		X"B7",X"28",X"05",X"CD",X"8C",X"17",X"18",X"03",X"CD",X"95",X"17",X"21",X"70",X"F8",X"F9",X"EB",
		X"01",X"10",X"00",X"ED",X"B0",X"F1",X"C1",X"D1",X"E1",X"DD",X"E1",X"FD",X"E1",X"C9",X"FD",X"E5",
		X"DD",X"E5",X"E5",X"D5",X"C5",X"F5",X"CD",X"8C",X"17",X"21",X"00",X"00",X"39",X"01",X"10",X"00",
		X"ED",X"B0",X"C3",X"08",X"17",X"C5",X"FD",X"E5",X"DD",X"E5",X"E5",X"D5",X"C5",X"F5",X"21",X"FD",
		X"41",X"7E",X"FE",X"18",X"38",X"07",X"21",X"0E",X"00",X"39",X"F9",X"37",X"C9",X"34",X"CD",X"8F",
		X"17",X"21",X"00",X"00",X"39",X"01",X"10",X"00",X"ED",X"B0",X"F1",X"C1",X"D1",X"E1",X"DD",X"E1",
		X"FD",X"E1",X"C1",X"B7",X"C9",X"21",X"FD",X"41",X"7E",X"35",X"23",X"96",X"20",X"07",X"36",X"00",
		X"CD",X"95",X"17",X"18",X"96",X"CD",X"95",X"17",X"21",X"10",X"00",X"19",X"EB",X"E5",X"21",X"8F",
		X"43",X"B7",X"ED",X"52",X"44",X"4D",X"E1",X"EB",X"ED",X"B0",X"18",X"E4",X"0E",X"01",X"3E",X"4E",
		X"21",X"FF",X"41",X"18",X"05",X"21",X"FE",X"41",X"4E",X"23",X"06",X"00",X"EB",X"21",X"00",X"00",
		X"09",X"29",X"29",X"29",X"29",X"19",X"EB",X"C9",X"21",X"00",X"80",X"01",X"1B",X"00",X"C3",X"40",
		X"06",X"D5",X"C5",X"F5",X"21",X"00",X"80",X"01",X"00",X"03",X"7E",X"FE",X"FF",X"20",X"0B",X"3E",
		X"08",X"81",X"4F",X"23",X"10",X"F4",X"F1",X"37",X"18",X"16",X"06",X"01",X"57",X"A0",X"7A",X"28",
		X"05",X"0C",X"CB",X"00",X"18",X"F6",X"B0",X"77",X"06",X"00",X"21",X"03",X"80",X"09",X"F1",X"B7",
		X"C1",X"D1",X"C9",X"C5",X"F5",X"36",X"00",X"01",X"03",X"80",X"B7",X"ED",X"42",X"7D",X"FE",X"18",
		X"30",X"19",X"21",X"00",X"80",X"FE",X"08",X"38",X"05",X"23",X"D6",X"08",X"18",X"F7",X"06",X"FE",
		X"B7",X"28",X"05",X"CB",X"00",X"3D",X"20",X"FB",X"78",X"A6",X"77",X"F1",X"C1",X"C9",X"FD",X"E1",
		X"CD",X"B1",X"17",X"77",X"CD",X"CF",X"16",X"7E",X"B7",X"20",X"F9",X"CD",X"E3",X"17",X"FD",X"E9",
		X"CD",X"59",X"19",X"DD",X"36",X"00",X"96",X"01",X"FF",X"FF",X"CD",X"B1",X"17",X"EB",X"CD",X"1E",
		X"17",X"DD",X"CB",X"00",X"6E",X"C2",X"19",X"19",X"3A",X"5E",X"40",X"B7",X"28",X"18",X"1A",X"B7",
		X"28",X"03",X"79",X"18",X"18",X"2A",X"62",X"40",X"7E",X"23",X"22",X"62",X"40",X"CB",X"7F",X"28",
		X"08",X"CB",X"BF",X"12",X"18",X"D8",X"CD",X"8B",X"09",X"CB",X"67",X"20",X"0B",X"E6",X"0F",X"CD",
		X"D8",X"15",X"B9",X"C4",X"02",X"19",X"18",X"C6",X"47",X"1A",X"B7",X"20",X"14",X"AF",X"FD",X"21",
		X"1B",X"80",X"FD",X"B6",X"00",X"28",X"0E",X"FD",X"21",X"2A",X"80",X"AF",X"FD",X"B6",X"00",X"28",
		X"04",X"3E",X"00",X"18",X"D8",X"78",X"E6",X"0F",X"CA",X"2E",X"18",X"D5",X"CD",X"E6",X"1A",X"4F",
		X"06",X"00",X"50",X"21",X"A9",X"19",X"09",X"5E",X"21",X"CE",X"19",X"19",X"19",X"19",X"DD",X"36",
		X"08",X"00",X"DD",X"36",X"0A",X"00",X"7E",X"23",X"F3",X"DD",X"77",X"0C",X"7E",X"23",X"DD",X"77",
		X"0D",X"FB",X"DD",X"36",X"07",X"01",X"D1",X"EB",X"36",X"02",X"CD",X"1E",X"17",X"7E",X"B7",X"20",
		X"F9",X"EB",X"D5",X"46",X"23",X"4E",X"23",X"7E",X"F6",X"06",X"57",X"DD",X"7E",X"09",X"80",X"5F",
		X"DD",X"7E",X"0B",X"81",X"4F",X"FD",X"E5",X"E1",X"06",X"0F",X"AF",X"77",X"23",X"10",X"FC",X"F3",
		X"FD",X"72",X"00",X"FD",X"73",X"01",X"FD",X"71",X"02",X"FD",X"73",X"03",X"FD",X"71",X"04",X"FB",
		X"0E",X"00",X"E1",X"36",X"04",X"CD",X"1E",X"17",X"7E",X"B7",X"20",X"F9",X"36",X"0D",X"EB",X"C3",
		X"2E",X"18",X"E6",X"0F",X"D5",X"CD",X"20",X"30",X"21",X"BA",X"19",X"19",X"7E",X"23",X"66",X"F3",
		X"DD",X"77",X"0C",X"DD",X"74",X"0D",X"FB",X"D1",X"C9",X"CD",X"8B",X"1B",X"3E",X"10",X"CD",X"04",
		X"19",X"EB",X"36",X"96",X"CD",X"1E",X"17",X"3A",X"BC",X"F8",X"C6",X"55",X"F6",X"88",X"32",X"BC",
		X"F8",X"7E",X"B7",X"20",X"EF",X"DD",X"36",X"00",X"89",X"CD",X"1E",X"17",X"DD",X"CB",X"00",X"46",
		X"20",X"F7",X"36",X"1E",X"CD",X"1E",X"17",X"7E",X"B7",X"20",X"F9",X"DD",X"36",X"00",X"00",X"AF",
		X"32",X"A0",X"F8",X"CD",X"1E",X"17",X"C3",X"53",X"19",X"CD",X"89",X"19",X"3A",X"07",X"40",X"FE",
		X"01",X"3E",X"AA",X"28",X"02",X"3E",X"EE",X"32",X"BC",X"F8",X"2A",X"0A",X"40",X"DD",X"75",X"09",
		X"DD",X"74",X"0B",X"7D",X"6C",X"67",X"CD",X"98",X"16",X"EB",X"CB",X"F6",X"AF",X"CD",X"02",X"19",
		X"DD",X"36",X"06",X"01",X"DD",X"36",X"07",X"01",X"C9",X"21",X"AD",X"40",X"11",X"0E",X"00",X"06",
		X"18",X"CB",X"7E",X"28",X"05",X"19",X"10",X"F9",X"37",X"C9",X"E5",X"01",X"0E",X"00",X"CD",X"40",
		X"06",X"DD",X"E1",X"DD",X"CB",X"00",X"FE",X"B7",X"C9",X"00",X"0C",X"04",X"00",X"10",X"0E",X"02",
		X"10",X"08",X"0A",X"06",X"08",X"00",X"0C",X"04",X"00",X"12",X"8F",X"39",X"97",X"39",X"97",X"39",
		X"97",X"39",X"97",X"39",X"A7",X"39",X"A7",X"39",X"A7",X"39",X"97",X"39",X"B7",X"39",X"8F",X"39",
		X"00",X"00",X"00",X"00",X"C3",X"39",X"08",X"02",X"60",X"00",X"CB",X"39",X"08",X"03",X"20",X"00",
		X"D3",X"39",X"07",X"07",X"A0",X"00",X"DB",X"39",X"06",X"08",X"80",X"00",X"E3",X"39",X"FF",X"07",
		X"90",X"00",X"EB",X"39",X"FF",X"03",X"10",X"00",X"F3",X"39",X"FF",X"FF",X"50",X"00",X"FB",X"39",
		X"07",X"01",X"40",X"00",X"C5",X"D5",X"E5",X"CD",X"81",X"09",X"C2",X"84",X"07",X"3A",X"5E",X"40",
		X"B7",X"28",X"08",X"3E",X"01",X"32",X"80",X"F8",X"C3",X"1E",X"1A",X"CD",X"95",X"1A",X"CD",X"53",
		X"1A",X"3A",X"5E",X"40",X"B7",X"20",X"1E",X"2A",X"9A",X"F8",X"7C",X"B5",X"28",X"1A",X"DB",X"44",
		X"E6",X"C0",X"FE",X"40",X"20",X"12",X"7E",X"CB",X"7F",X"20",X"0A",X"23",X"D3",X"44",X"CB",X"77",
		X"28",X"06",X"C3",X"2A",X"1A",X"21",X"00",X"00",X"22",X"9A",X"F8",X"E1",X"D1",X"C1",X"F1",X"D3",
		X"4C",X"ED",X"45",X"21",X"80",X"F8",X"46",X"23",X"56",X"23",X"5E",X"23",X"0E",X"41",X"CB",X"80",
		X"CB",X"C2",X"ED",X"51",X"0D",X"ED",X"41",X"0C",X"CB",X"82",X"ED",X"51",X"0D",X"ED",X"59",X"0C",
		X"0C",X"06",X"03",X"79",X"0C",X"51",X"5E",X"23",X"4F",X"7E",X"23",X"ED",X"79",X"79",X"4A",X"ED",
		X"59",X"14",X"14",X"10",X"F1",X"0D",X"3E",X"00",X"06",X"04",X"B6",X"23",X"ED",X"79",X"E6",X"C0",
		X"C6",X"40",X"10",X"F6",X"C9",X"3A",X"91",X"F8",X"B7",X"C4",X"B9",X"1D",X"3A",X"90",X"F8",X"B7",
		X"C4",X"37",X"1E",X"2A",X"8D",X"F8",X"7C",X"B5",X"C8",X"E9",X"21",X"00",X"00",X"22",X"8D",X"F8",
		X"C9",X"E1",X"22",X"8D",X"F8",X"C9",X"F5",X"E5",X"21",X"00",X"00",X"AF",X"22",X"80",X"F8",X"32",
		X"82",X"F8",X"22",X"89",X"F8",X"22",X"8B",X"F8",X"AF",X"32",X"8F",X"F8",X"E1",X"F1",X"C9",X"21",
		X"00",X"00",X"AF",X"22",X"80",X"F8",X"32",X"82",X"F8",X"22",X"89",X"F8",X"22",X"8B",X"F8",X"AF",
		X"32",X"8F",X"F8",X"C3",X"AA",X"1A",X"F5",X"3A",X"8F",X"F8",X"FE",X"0A",X"DA",X"F4",X"1A",X"CA",
		X"F4",X"1A",X"F1",X"C9",X"3E",X"0A",X"32",X"8F",X"F8",X"E5",X"21",X"03",X"1B",X"22",X"8D",X"F8",
		X"E1",X"F1",X"C9",X"21",X"80",X"F8",X"36",X"92",X"23",X"36",X"92",X"23",X"36",X"92",X"21",X"89",
		X"F8",X"36",X"00",X"23",X"36",X"05",X"23",X"36",X"06",X"23",X"36",X"06",X"21",X"32",X"00",X"22",
		X"83",X"F8",X"21",X"32",X"00",X"22",X"85",X"F8",X"21",X"32",X"00",X"22",X"87",X"F8",X"3E",X"32",
		X"32",X"92",X"F8",X"CD",X"B1",X"1A",X"2A",X"83",X"F8",X"11",X"0F",X"00",X"19",X"22",X"83",X"F8",
		X"2A",X"85",X"F8",X"11",X"11",X"00",X"19",X"22",X"85",X"F8",X"2A",X"87",X"F8",X"11",X"10",X"00",
		X"19",X"22",X"87",X"F8",X"21",X"92",X"F8",X"35",X"C2",X"33",X"1B",X"3E",X"32",X"32",X"92",X"F8",
		X"CD",X"B1",X"1A",X"2A",X"83",X"F8",X"11",X"0A",X"00",X"19",X"22",X"83",X"F8",X"2A",X"85",X"F8",
		X"11",X"0D",X"00",X"19",X"22",X"85",X"F8",X"2A",X"87",X"F8",X"11",X"0F",X"00",X"19",X"22",X"87",
		X"F8",X"21",X"92",X"F8",X"35",X"C2",X"60",X"1B",X"C3",X"CF",X"1A",X"F5",X"3A",X"8F",X"F8",X"FE",
		X"0D",X"DA",X"99",X"1B",X"CA",X"99",X"1B",X"F1",X"C9",X"3E",X"0D",X"32",X"8F",X"F8",X"E5",X"21",
		X"A8",X"1B",X"22",X"8D",X"F8",X"E1",X"F1",X"C9",X"21",X"80",X"F8",X"36",X"90",X"23",X"36",X"90",
		X"23",X"36",X"90",X"21",X"89",X"F8",X"36",X"00",X"23",X"36",X"06",X"23",X"36",X"07",X"23",X"36",
		X"07",X"3E",X"10",X"32",X"92",X"F8",X"21",X"E6",X"00",X"22",X"83",X"F8",X"21",X"14",X"00",X"2A",
		X"85",X"F8",X"21",X"0A",X"00",X"2A",X"86",X"F8",X"3E",X"14",X"32",X"94",X"F8",X"CD",X"B1",X"1A",
		X"21",X"85",X"F8",X"7E",X"C6",X"05",X"77",X"21",X"87",X"F8",X"7E",X"C6",X"1E",X"77",X"21",X"94",
		X"F8",X"35",X"C2",X"DD",X"1B",X"21",X"83",X"F8",X"7E",X"C6",X"FC",X"77",X"21",X"92",X"F8",X"35",
		X"C2",X"CC",X"1B",X"C3",X"CF",X"1A",X"F5",X"3A",X"8F",X"F8",X"FE",X"0B",X"DA",X"14",X"1C",X"CA",
		X"14",X"1C",X"F1",X"C9",X"3E",X"0B",X"32",X"8F",X"F8",X"E5",X"21",X"23",X"1C",X"22",X"8D",X"F8",
		X"E1",X"F1",X"C9",X"21",X"80",X"F8",X"36",X"82",X"23",X"36",X"80",X"23",X"36",X"80",X"21",X"89",
		X"F8",X"36",X"03",X"23",X"36",X"07",X"23",X"36",X"07",X"23",X"36",X"07",X"21",X"01",X"00",X"22",
		X"83",X"F8",X"21",X"01",X"00",X"22",X"85",X"F8",X"21",X"05",X"00",X"22",X"87",X"F8",X"CD",X"B1",
		X"1A",X"21",X"80",X"F8",X"36",X"92",X"23",X"36",X"90",X"23",X"36",X"90",X"3E",X"37",X"32",X"94",
		X"F8",X"3E",X"06",X"32",X"92",X"F8",X"CD",X"B1",X"1A",X"21",X"92",X"F8",X"35",X"C2",X"66",X"1C",
		X"2A",X"83",X"F8",X"11",X"01",X"00",X"19",X"22",X"83",X"F8",X"21",X"94",X"F8",X"35",X"C2",X"61",
		X"1C",X"C3",X"CF",X"1A",X"F5",X"3A",X"8F",X"F8",X"FE",X"0B",X"DA",X"92",X"1C",X"CA",X"92",X"1C",
		X"F1",X"C9",X"3E",X"0B",X"32",X"8F",X"F8",X"E5",X"21",X"A1",X"1C",X"22",X"8D",X"F8",X"E1",X"F1",
		X"C9",X"21",X"80",X"F8",X"36",X"92",X"23",X"36",X"92",X"23",X"36",X"92",X"21",X"89",X"F8",X"36",
		X"00",X"23",X"36",X"06",X"23",X"36",X"06",X"23",X"36",X"07",X"21",X"14",X"00",X"22",X"83",X"F8",
		X"21",X"2D",X"00",X"22",X"85",X"F8",X"21",X"5A",X"00",X"22",X"87",X"F8",X"3E",X"04",X"32",X"94",
		X"F8",X"3E",X"50",X"32",X"92",X"F8",X"CD",X"B1",X"1A",X"2A",X"83",X"F8",X"11",X"08",X"00",X"19",
		X"22",X"83",X"F8",X"2A",X"85",X"F8",X"11",X"11",X"00",X"19",X"22",X"85",X"F8",X"2A",X"87",X"F8",
		X"11",X"2F",X"00",X"19",X"22",X"87",X"F8",X"21",X"92",X"F8",X"35",X"C2",X"D6",X"1C",X"21",X"94",
		X"F8",X"35",X"C2",X"D1",X"1C",X"C3",X"CF",X"1A",X"F5",X"3A",X"8F",X"F8",X"FE",X"0C",X"DA",X"16",
		X"1D",X"CA",X"16",X"1D",X"F1",X"C9",X"3E",X"0C",X"32",X"8F",X"F8",X"E5",X"21",X"25",X"1D",X"22",
		X"8D",X"F8",X"E1",X"F1",X"C9",X"21",X"80",X"F8",X"36",X"92",X"23",X"36",X"92",X"23",X"36",X"92",
		X"21",X"89",X"F8",X"36",X"00",X"23",X"36",X"07",X"23",X"36",X"07",X"23",X"36",X"07",X"21",X"C8",
		X"00",X"22",X"83",X"F8",X"21",X"3C",X"00",X"22",X"85",X"F8",X"21",X"28",X"00",X"22",X"87",X"F8",
		X"3E",X"14",X"32",X"94",X"F8",X"3E",X"14",X"32",X"92",X"F8",X"CD",X"B1",X"1A",X"2A",X"83",X"F8",
		X"11",X"14",X"00",X"19",X"22",X"83",X"F8",X"2A",X"85",X"F8",X"11",X"06",X"00",X"19",X"22",X"85",
		X"F8",X"2A",X"87",X"F8",X"11",X"04",X"00",X"19",X"22",X"87",X"F8",X"21",X"92",X"F8",X"35",X"C2",
		X"5A",X"1D",X"3E",X"14",X"32",X"92",X"F8",X"CD",X"B1",X"1A",X"2A",X"83",X"F8",X"11",X"EC",X"FF",
		X"19",X"22",X"83",X"F8",X"2A",X"85",X"F8",X"11",X"FA",X"FF",X"19",X"22",X"85",X"F8",X"2A",X"87",
		X"F8",X"11",X"FC",X"FF",X"19",X"22",X"87",X"F8",X"21",X"92",X"F8",X"35",X"C2",X"87",X"1D",X"21",
		X"94",X"F8",X"35",X"C2",X"55",X"1D",X"C3",X"CF",X"1A",X"AF",X"32",X"91",X"F8",X"32",X"90",X"F8",
		X"3A",X"8F",X"F8",X"FE",X"0B",X"DA",X"CC",X"1D",X"CA",X"CC",X"1D",X"C9",X"3E",X"0B",X"32",X"8F",
		X"F8",X"21",X"80",X"F8",X"36",X"92",X"23",X"36",X"92",X"23",X"36",X"92",X"21",X"89",X"F8",X"36",
		X"00",X"23",X"36",X"07",X"23",X"36",X"07",X"23",X"36",X"07",X"21",X"30",X"00",X"22",X"83",X"F8",
		X"21",X"38",X"00",X"22",X"85",X"F8",X"21",X"40",X"00",X"22",X"87",X"F8",X"ED",X"5F",X"E6",X"1F",
		X"32",X"94",X"F8",X"CD",X"B1",X"1A",X"3A",X"94",X"F8",X"E6",X"07",X"C2",X"18",X"1E",X"21",X"8A",
		X"F8",X"7E",X"3D",X"77",X"23",X"77",X"23",X"77",X"21",X"83",X"F8",X"7E",X"C6",X"06",X"77",X"21",
		X"85",X"F8",X"7E",X"C6",X"07",X"77",X"21",X"87",X"F8",X"7E",X"C6",X"08",X"77",X"21",X"94",X"F8",
		X"35",X"C2",X"03",X"1E",X"C3",X"CF",X"1A",X"AF",X"32",X"90",X"F8",X"3A",X"8F",X"F8",X"FE",X"0A",
		X"DA",X"47",X"1E",X"CA",X"47",X"1E",X"C9",X"3E",X"0A",X"32",X"8F",X"F8",X"21",X"80",X"F8",X"36",
		X"82",X"23",X"36",X"80",X"23",X"36",X"80",X"21",X"89",X"F8",X"36",X"03",X"23",X"36",X"07",X"23",
		X"36",X"07",X"23",X"36",X"07",X"21",X"01",X"00",X"22",X"83",X"F8",X"21",X"01",X"00",X"22",X"85",
		X"F8",X"21",X"02",X"00",X"22",X"87",X"F8",X"CD",X"B1",X"1A",X"21",X"80",X"F8",X"36",X"92",X"23",
		X"36",X"90",X"23",X"36",X"90",X"3E",X"37",X"32",X"94",X"F8",X"CD",X"B1",X"1A",X"21",X"85",X"F8",
		X"7E",X"C6",X"01",X"77",X"21",X"87",X"F8",X"7E",X"C6",X"01",X"77",X"21",X"94",X"F8",X"35",X"C2",
		X"8A",X"1E",X"C3",X"CF",X"1A",X"E1",X"22",X"05",X"40",X"CD",X"1A",X"11",X"CD",X"20",X"24",X"3A",
		X"5E",X"40",X"B7",X"20",X"20",X"CD",X"59",X"19",X"01",X"12",X"10",X"3A",X"21",X"40",X"FE",X"02",
		X"28",X"02",X"06",X"06",X"DD",X"71",X"00",X"3E",X"0A",X"CD",X"0E",X"18",X"3E",X"1B",X"A9",X"4F",
		X"10",X"F2",X"CD",X"77",X"20",X"FB",X"AF",X"32",X"23",X"40",X"32",X"66",X"40",X"3E",X"5A",X"32",
		X"A1",X"F8",X"3A",X"0D",X"40",X"C6",X"06",X"FE",X"17",X"38",X"08",X"D6",X"16",X"FE",X"07",X"38",
		X"F4",X"18",X"F4",X"32",X"0D",X"40",X"32",X"9E",X"F8",X"01",X"20",X"18",X"CD",X"35",X"17",X"01",
		X"9F",X"2E",X"CD",X"35",X"17",X"3A",X"12",X"40",X"B7",X"28",X"0A",X"E6",X"03",X"20",X"06",X"01",
		X"9B",X"31",X"CD",X"35",X"17",X"AF",X"32",X"1F",X"40",X"01",X"A1",X"21",X"CD",X"35",X"17",X"21",
		X"0D",X"40",X"35",X"20",X"F4",X"3A",X"9E",X"F8",X"32",X"0D",X"40",X"CD",X"CF",X"16",X"DD",X"21",
		X"AD",X"40",X"DD",X"CB",X"00",X"56",X"CA",X"8D",X"1F",X"DD",X"7E",X"0B",X"32",X"0B",X"40",X"47",
		X"DD",X"7E",X"09",X"32",X"0A",X"40",X"DD",X"CB",X"00",X"6E",X"C2",X"67",X"1F",X"11",X"D5",X"1E",
		X"D5",X"FE",X"05",X"DA",X"3D",X"20",X"FE",X"F6",X"D2",X"04",X"20",X"78",X"FE",X"05",X"DA",X"CC",
		X"1F",X"FE",X"BE",X"D2",X"94",X"1F",X"D1",X"CD",X"CF",X"20",X"3A",X"67",X"40",X"B7",X"C4",X"A2",
		X"20",X"3A",X"A1",X"F8",X"B7",X"20",X"0A",X"3D",X"32",X"A1",X"F8",X"01",X"E5",X"2E",X"CD",X"35",
		X"17",X"3A",X"5E",X"40",X"B7",X"28",X"03",X"CD",X"27",X"0D",X"C3",X"2B",X"1F",X"CD",X"B6",X"1A",
		X"2A",X"05",X"40",X"E9",X"3E",X"0A",X"32",X"0B",X"40",X"21",X"09",X"40",X"34",X"21",X"F3",X"23",
		X"E5",X"CD",X"74",X"20",X"28",X"06",X"11",X"DF",X"5F",X"C3",X"E7",X"1F",X"11",X"00",X"44",X"3E",
		X"1B",X"21",X"00",X"01",X"19",X"01",X"00",X"19",X"D5",X"ED",X"B0",X"D1",X"01",X"00",X"01",X"2B",
		X"36",X"00",X"0D",X"C2",X"BF",X"1F",X"10",X"F7",X"3D",X"20",X"E6",X"C9",X"3E",X"B2",X"32",X"0B",
		X"40",X"21",X"09",X"40",X"35",X"21",X"C6",X"23",X"E5",X"CD",X"74",X"20",X"28",X"06",X"11",X"00",
		X"46",X"C3",X"AF",X"1F",X"11",X"FF",X"5D",X"3E",X"1A",X"01",X"00",X"19",X"21",X"00",X"FF",X"19",
		X"D5",X"ED",X"B8",X"D1",X"01",X"00",X"01",X"23",X"36",X"00",X"0D",X"C2",X"F7",X"1F",X"10",X"F7",
		X"3D",X"20",X"E6",X"C9",X"3E",X"13",X"32",X"0A",X"40",X"21",X"08",X"40",X"34",X"21",X"7C",X"23",
		X"E5",X"CD",X"74",X"20",X"28",X"06",X"11",X"E0",X"5F",X"C3",X"58",X"20",X"11",X"00",X"44",X"3E",
		X"20",X"01",X"FF",X"19",X"21",X"01",X"00",X"19",X"D5",X"ED",X"B0",X"06",X"D0",X"11",X"E1",X"FF",
		X"36",X"00",X"2B",X"36",X"00",X"19",X"10",X"F8",X"D1",X"3D",X"20",X"E5",X"C9",X"3E",X"E4",X"32",
		X"0A",X"40",X"21",X"08",X"40",X"35",X"21",X"A1",X"23",X"E5",X"CD",X"74",X"20",X"28",X"06",X"11",
		X"00",X"46",X"C3",X"1F",X"20",X"11",X"00",X"5E",X"3E",X"20",X"01",X"00",X"1A",X"21",X"FF",X"FF",
		X"19",X"D5",X"ED",X"B8",X"11",X"1F",X"00",X"36",X"00",X"23",X"36",X"00",X"19",X"10",X"F8",X"D1",
		X"3D",X"20",X"E7",X"C9",X"CD",X"01",X"0E",X"F3",X"CD",X"98",X"20",X"21",X"BB",X"40",X"22",X"BF",
		X"F8",X"21",X"AD",X"40",X"22",X"BD",X"F8",X"01",X"50",X"01",X"CD",X"40",X"06",X"CD",X"C2",X"16",
		X"CD",X"A8",X"17",X"3A",X"22",X"40",X"B7",X"C9",X"21",X"1B",X"80",X"01",X"69",X"00",X"CD",X"40",
		X"06",X"C9",X"AF",X"32",X"67",X"40",X"11",X"00",X"D5",X"21",X"68",X"40",X"06",X"06",X"CD",X"53",
		X"2E",X"3A",X"21",X"40",X"FE",X"02",X"C0",X"11",X"B0",X"D5",X"21",X"6B",X"40",X"06",X"06",X"C3",
		X"53",X"2E",X"3A",X"07",X"40",X"FE",X"02",X"21",X"6B",X"40",X"C8",X"21",X"68",X"40",X"C9",X"21",
		X"66",X"40",X"7E",X"B7",X"C8",X"4F",X"ED",X"44",X"F3",X"86",X"77",X"FB",X"79",X"F5",X"0F",X"0F",
		X"0F",X"0F",X"06",X"01",X"CD",X"EA",X"20",X"F1",X"06",X"00",X"E6",X"0F",X"4F",X"3A",X"B9",X"F8",
		X"F5",X"C5",X"CD",X"FB",X"20",X"C1",X"F1",X"3D",X"20",X"F6",X"C9",X"3E",X"FF",X"32",X"67",X"40",
		X"1E",X"04",X"CD",X"C2",X"20",X"23",X"23",X"23",X"CB",X"38",X"08",X"04",X"2B",X"1D",X"10",X"FC",
		X"08",X"30",X"08",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"7B",X"FE",X"02",X"28",X"0D",
		X"79",X"86",X"27",X"77",X"30",X"06",X"2B",X"0E",X"01",X"1D",X"20",X"EF",X"C9",X"7E",X"47",X"81",
		X"27",X"77",X"0E",X"02",X"38",X"01",X"0D",X"E6",X"F0",X"08",X"78",X"E6",X"F0",X"47",X"08",X"90",
		X"27",X"28",X"13",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"11",X"40",X"B7",X"28",X"08",X"90",X"38",
		X"0C",X"28",X"0A",X"32",X"11",X"40",X"0D",X"CA",X"2C",X"21",X"C3",X"26",X"21",X"47",X"DB",X"60",
		X"E6",X"0F",X"90",X"32",X"11",X"40",X"C5",X"D5",X"E5",X"21",X"0C",X"40",X"34",X"CD",X"08",X"1D",
		X"CD",X"40",X"24",X"E1",X"D1",X"C1",X"C3",X"56",X"21",X"CD",X"89",X"19",X"DA",X"65",X"17",X"ED",
		X"5F",X"0F",X"38",X"05",X"CD",X"73",X"30",X"18",X"03",X"CD",X"7F",X"30",X"DD",X"36",X"09",X"92",
		X"DD",X"36",X"0B",X"68",X"21",X"F1",X"38",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"0E",X"00",X"18",
		X"1E",X"ED",X"5F",X"E6",X"01",X"C2",X"11",X"37",X"21",X"1F",X"40",X"34",X"7E",X"32",X"20",X"40",
		X"CD",X"89",X"19",X"DA",X"65",X"17",X"CD",X"FB",X"22",X"AF",X"0E",X"FF",X"CD",X"2E",X"22",X"DD",
		X"36",X"06",X"02",X"DD",X"36",X"07",X"01",X"DD",X"36",X"00",X"86",X"CD",X"B1",X"17",X"3A",X"0F",
		X"40",X"FE",X"28",X"30",X"02",X"3E",X"28",X"47",X"CD",X"39",X"10",X"E6",X"F8",X"0F",X"0F",X"0F",
		X"80",X"77",X"CD",X"CF",X"16",X"DD",X"CB",X"00",X"6E",X"20",X"04",X"7E",X"B7",X"20",X"F3",X"0E",
		X"00",X"FD",X"21",X"AD",X"40",X"C5",X"FD",X"7E",X"09",X"DD",X"96",X"09",X"57",X"01",X"00",X"00",
		X"28",X"06",X"06",X"01",X"38",X"02",X"06",X"02",X"FD",X"7E",X"0B",X"C6",X"02",X"DD",X"96",X"0B",
		X"5F",X"28",X"06",X"0E",X"04",X"38",X"02",X"0E",X"08",X"78",X"81",X"C1",X"CD",X"81",X"2C",X"CD",
		X"2E",X"22",X"CD",X"CF",X"16",X"DD",X"CB",X"00",X"6E",X"CA",X"F1",X"21",X"18",X"2C",X"E5",X"21",
		X"23",X"40",X"CB",X"4E",X"28",X"03",X"AF",X"18",X"09",X"E6",X"0F",X"28",X"05",X"CB",X"46",X"CC",
		X"D8",X"15",X"B9",X"28",X"13",X"4F",X"CD",X"20",X"30",X"21",X"69",X"23",X"19",X"7E",X"23",X"66",
		X"F3",X"DD",X"77",X"0C",X"DD",X"74",X"0D",X"FB",X"E1",X"C9",X"CD",X"E3",X"17",X"DD",X"E5",X"CD",
		X"06",X"1C",X"E1",X"11",X"08",X"00",X"19",X"F3",X"72",X"23",X"7E",X"D6",X"04",X"77",X"23",X"72",
		X"23",X"7E",X"D6",X"06",X"77",X"23",X"01",X"4B",X"39",X"71",X"23",X"70",X"FB",X"DD",X"36",X"07",
		X"01",X"DD",X"36",X"06",X"01",X"DD",X"E5",X"01",X"05",X"01",X"CD",X"FB",X"20",X"21",X"1F",X"40",
		X"7E",X"B7",X"CA",X"D9",X"22",X"35",X"32",X"10",X"40",X"20",X"3E",X"3A",X"20",X"40",X"F5",X"01",
		X"01",X"01",X"CD",X"FB",X"20",X"F1",X"3D",X"20",X"F5",X"CD",X"8E",X"2D",X"00",X"60",X"D5",X"42",
		X"4F",X"4E",X"55",X"53",X"00",X"F5",X"3A",X"20",X"40",X"47",X"AF",X"C6",X"01",X"27",X"10",X"FB",
		X"0F",X"0F",X"0F",X"0F",X"6F",X"E6",X"F0",X"67",X"3E",X"0F",X"A5",X"6F",X"F1",X"E5",X"21",X"00",
		X"00",X"39",X"08",X"06",X"04",X"CD",X"5D",X"2E",X"E1",X"DD",X"E1",X"3E",X"1E",X"CD",X"0E",X"18",
		X"21",X"82",X"C1",X"DD",X"7E",X"04",X"BD",X"20",X"06",X"DD",X"7E",X"05",X"BC",X"28",X"05",X"CD",
		X"CF",X"16",X"18",X"EC",X"DD",X"36",X"00",X"00",X"C3",X"65",X"17",X"CD",X"39",X"10",X"D6",X"18",
		X"30",X"FC",X"C6",X"18",X"06",X"00",X"4F",X"21",X"26",X"40",X"09",X"7E",X"E6",X"F0",X"28",X"04",
		X"79",X"3C",X"18",X"EA",X"CB",X"FE",X"21",X"39",X"23",X"09",X"09",X"56",X"23",X"5E",X"CD",X"2D",
		X"23",X"82",X"DD",X"77",X"09",X"CD",X"2D",X"23",X"83",X"DD",X"77",X"0B",X"C9",X"D5",X"CD",X"39",
		X"10",X"D1",X"D6",X"1A",X"30",X"FC",X"C6",X"1A",X"C9",X"0C",X"08",X"34",X"08",X"5C",X"08",X"84",
		X"08",X"AC",X"08",X"D4",X"08",X"0C",X"38",X"34",X"38",X"5C",X"38",X"84",X"38",X"AC",X"38",X"D4",
		X"38",X"0C",X"68",X"34",X"68",X"5C",X"68",X"84",X"68",X"AC",X"68",X"D4",X"68",X"0C",X"98",X"34",
		X"98",X"5C",X"98",X"84",X"98",X"AC",X"98",X"D4",X"98",X"05",X"39",X"23",X"39",X"23",X"39",X"23",
		X"39",X"2D",X"39",X"37",X"39",X"37",X"39",X"37",X"39",X"41",X"39",X"6B",X"CD",X"4B",X"26",X"DD",
		X"CB",X"18",X"C6",X"DD",X"CB",X"1E",X"C6",X"DD",X"CB",X"24",X"C6",X"DD",X"CB",X"2A",X"C6",X"2A",
		X"0A",X"40",X"6C",X"26",X"F0",X"CD",X"98",X"16",X"21",X"18",X"00",X"19",X"CB",X"CE",X"C3",X"27",
		X"24",X"CD",X"4B",X"26",X"DD",X"CB",X"1D",X"CE",X"DD",X"CB",X"23",X"CE",X"DD",X"CB",X"29",X"CE",
		X"DD",X"CB",X"2F",X"CE",X"2A",X"0A",X"40",X"6C",X"26",X"10",X"CD",X"98",X"16",X"21",X"18",X"00",
		X"19",X"CB",X"C6",X"C3",X"27",X"24",X"CD",X"4B",X"26",X"DD",X"CB",X"2A",X"DE",X"DD",X"CB",X"2B",
		X"DE",X"DD",X"CB",X"2C",X"DE",X"DD",X"CB",X"2D",X"DE",X"DD",X"CB",X"2E",X"DE",X"DD",X"CB",X"2F",
		X"DE",X"2A",X"0A",X"40",X"65",X"2E",X"10",X"CD",X"98",X"16",X"21",X"18",X"00",X"19",X"CB",X"D6",
		X"C3",X"27",X"24",X"CD",X"4B",X"26",X"DD",X"CB",X"18",X"D6",X"DD",X"CB",X"19",X"D6",X"DD",X"CB",
		X"1A",X"D6",X"DD",X"CB",X"1B",X"D6",X"DD",X"CB",X"1C",X"D6",X"DD",X"CB",X"1D",X"D6",X"2A",X"0A",
		X"40",X"65",X"2E",X"B4",X"CD",X"98",X"16",X"21",X"18",X"00",X"19",X"CB",X"DE",X"C3",X"27",X"24",
		X"21",X"12",X"40",X"35",X"CD",X"4B",X"26",X"DD",X"21",X"26",X"40",X"CD",X"77",X"24",X"CD",X"77",
		X"24",X"CD",X"77",X"24",X"CD",X"F1",X"24",X"CD",X"52",X"0E",X"CD",X"F3",X"26",X"CD",X"A2",X"20",
		X"3A",X"07",X"40",X"FE",X"02",X"21",X"38",X"D5",X"20",X"02",X"2E",X"E8",X"06",X"00",X"CD",X"B6",
		X"2D",X"EB",X"08",X"3A",X"0C",X"40",X"47",X"08",X"05",X"28",X"14",X"C5",X"0E",X"80",X"CD",X"EE",
		X"2D",X"13",X"08",X"3A",X"22",X"40",X"B7",X"28",X"02",X"1B",X"1B",X"08",X"C1",X"10",X"EC",X"3A",
		X"5E",X"40",X"B7",X"C4",X"A2",X"0C",X"C9",X"06",X"05",X"C5",X"CD",X"39",X"10",X"01",X"91",X"24",
		X"C5",X"E6",X"03",X"CA",X"AF",X"24",X"3D",X"CA",X"99",X"24",X"3D",X"CA",X"C5",X"24",X"C3",X"DB",
		X"24",X"C1",X"DD",X"23",X"10",X"E3",X"DD",X"23",X"C9",X"DD",X"CB",X"06",X"CE",X"DD",X"CB",X"07",
		X"C6",X"3A",X"64",X"40",X"07",X"D0",X"DD",X"CB",X"1E",X"CE",X"DD",X"CB",X"1F",X"C6",X"C9",X"DD",
		X"CB",X"00",X"CE",X"DD",X"CB",X"01",X"C6",X"3A",X"64",X"40",X"07",X"D0",X"DD",X"CB",X"18",X"CE",
		X"DD",X"CB",X"19",X"C6",X"C9",X"DD",X"CB",X"01",X"DE",X"DD",X"CB",X"07",X"D6",X"3A",X"64",X"40",
		X"07",X"D0",X"DD",X"CB",X"19",X"DE",X"DD",X"CB",X"1F",X"D6",X"C9",X"DD",X"CB",X"00",X"DE",X"DD",
		X"CB",X"06",X"D6",X"3A",X"64",X"40",X"07",X"D0",X"DD",X"CB",X"18",X"DE",X"DD",X"CB",X"1E",X"D6",
		X"C9",X"26",X"04",X"DD",X"21",X"26",X"40",X"01",X"04",X"04",X"CD",X"26",X"25",X"3E",X"30",X"84",
		X"67",X"10",X"F7",X"DD",X"21",X"38",X"40",X"0E",X"08",X"CD",X"26",X"25",X"DD",X"21",X"26",X"40",
		X"01",X"01",X"06",X"2E",X"08",X"CD",X"58",X"25",X"3E",X"28",X"85",X"6F",X"10",X"F7",X"DD",X"2B",
		X"0E",X"02",X"CD",X"58",X"25",X"C9",X"C5",X"2E",X"08",X"06",X"06",X"E5",X"C5",X"DD",X"7E",X"18",
		X"A1",X"28",X"10",X"DD",X"7E",X"00",X"A1",X"28",X"05",X"CD",X"BE",X"25",X"18",X"0E",X"CD",X"A8",
		X"25",X"18",X"09",X"DD",X"7E",X"00",X"A1",X"28",X"03",X"CD",X"92",X"25",X"C1",X"E1",X"DD",X"23",
		X"3E",X"28",X"85",X"6F",X"10",X"D5",X"C1",X"C9",X"C5",X"26",X"04",X"06",X"04",X"E5",X"C5",X"DD",
		X"7E",X"18",X"A1",X"28",X"10",X"DD",X"7E",X"00",X"A1",X"28",X"05",X"CD",X"17",X"26",X"18",X"0E",
		X"CD",X"01",X"26",X"18",X"09",X"DD",X"7E",X"00",X"A1",X"28",X"03",X"CD",X"EB",X"25",X"C1",X"E1",
		X"11",X"06",X"00",X"DD",X"19",X"3E",X"30",X"84",X"67",X"10",X"D2",X"11",X"E9",X"FF",X"DD",X"19",
		X"C1",X"C9",X"06",X"0B",X"C5",X"E5",X"CD",X"44",X"26",X"21",X"AB",X"27",X"CD",X"6F",X"15",X"E1",
		X"C1",X"3E",X"04",X"85",X"6F",X"10",X"ED",X"C9",X"06",X"0B",X"C5",X"E5",X"CD",X"44",X"26",X"21",
		X"A5",X"27",X"CD",X"6F",X"15",X"E1",X"C1",X"3E",X"04",X"85",X"6F",X"10",X"ED",X"C9",X"E5",X"CD",
		X"44",X"26",X"21",X"C9",X"27",X"CD",X"6F",X"15",X"E1",X"3E",X"04",X"85",X"6F",X"06",X"09",X"C5",
		X"E5",X"CD",X"44",X"26",X"21",X"C3",X"27",X"CD",X"6F",X"15",X"E1",X"C1",X"3E",X"04",X"85",X"6F",
		X"10",X"ED",X"CD",X"44",X"26",X"21",X"CF",X"27",X"C3",X"6F",X"15",X"06",X"0D",X"C5",X"E5",X"CD",
		X"44",X"26",X"21",X"AB",X"27",X"CD",X"6F",X"15",X"E1",X"C1",X"3E",X"04",X"84",X"67",X"10",X"ED",
		X"C9",X"06",X"0D",X"C5",X"E5",X"CD",X"44",X"26",X"21",X"A5",X"27",X"CD",X"6F",X"15",X"E1",X"C1",
		X"3E",X"04",X"84",X"67",X"10",X"ED",X"C9",X"E5",X"CD",X"44",X"26",X"21",X"B7",X"27",X"CD",X"6F",
		X"15",X"E1",X"3E",X"04",X"84",X"67",X"06",X"0B",X"C5",X"E5",X"CD",X"44",X"26",X"21",X"B1",X"27",
		X"CD",X"6F",X"15",X"E1",X"C1",X"3E",X"04",X"84",X"67",X"10",X"ED",X"CD",X"44",X"26",X"21",X"BD",
		X"27",X"C3",X"6F",X"15",X"06",X"10",X"CD",X"B6",X"2D",X"EB",X"C9",X"2A",X"08",X"40",X"22",X"64",
		X"40",X"3A",X"22",X"40",X"B7",X"20",X"05",X"21",X"6A",X"5E",X"18",X"03",X"21",X"4A",X"44",X"11",
		X"14",X"00",X"AF",X"0E",X"0C",X"06",X"0C",X"77",X"23",X"10",X"FC",X"19",X"0D",X"20",X"F6",X"01",
		X"30",X"00",X"11",X"26",X"40",X"21",X"4C",X"27",X"ED",X"B0",X"DD",X"21",X"26",X"40",X"2A",X"08",
		X"40",X"7D",X"E6",X"03",X"5F",X"16",X"00",X"62",X"6B",X"29",X"19",X"29",X"EB",X"DD",X"19",X"DD",
		X"CB",X"00",X"86",X"DD",X"21",X"26",X"40",X"2A",X"08",X"40",X"7D",X"3C",X"E6",X"03",X"5F",X"16",
		X"00",X"62",X"6B",X"29",X"19",X"29",X"EB",X"DD",X"19",X"DD",X"CB",X"05",X"8E",X"DD",X"21",X"26",
		X"40",X"2A",X"08",X"40",X"7C",X"E6",X"03",X"3C",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"CB",X"00",
		X"96",X"DD",X"21",X"26",X"40",X"2A",X"08",X"40",X"7C",X"3C",X"E6",X"03",X"3C",X"5F",X"16",X"00",
		X"DD",X"19",X"DD",X"CB",X"12",X"9E",X"21",X"12",X"40",X"34",X"7E",X"FE",X"21",X"38",X"06",X"FE",
		X"FF",X"28",X"02",X"36",X"13",X"7E",X"B7",X"28",X"05",X"E6",X"03",X"CC",X"84",X"35",X"DD",X"21",
		X"26",X"40",X"C9",X"21",X"7C",X"27",X"7E",X"B7",X"C8",X"4F",X"23",X"46",X"23",X"E5",X"CD",X"05",
		X"27",X"E1",X"C3",X"F6",X"26",X"C5",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"19",X"CB",X"38",
		X"CB",X"19",X"CB",X"38",X"CB",X"19",X"08",X"3A",X"22",X"40",X"B7",X"CA",X"29",X"27",X"21",X"FF",
		X"87",X"ED",X"42",X"C1",X"08",X"3F",X"C3",X"2F",X"27",X"21",X"00",X"81",X"09",X"C1",X"08",X"CB",
		X"51",X"11",X"F0",X"0F",X"28",X"03",X"11",X"0F",X"F0",X"3A",X"22",X"40",X"B7",X"28",X"03",X"7A",
		X"53",X"5F",X"7E",X"A2",X"57",X"3A",X"A2",X"F8",X"A3",X"B2",X"77",X"C9",X"05",X"04",X"04",X"04",
		X"04",X"06",X"01",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"02",X"09",X"08",
		X"08",X"08",X"08",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"08",X"34",
		X"08",X"64",X"08",X"94",X"08",X"C4",X"F8",X"04",X"F8",X"34",X"F8",X"64",X"F8",X"94",X"F8",X"C4",
		X"30",X"04",X"58",X"04",X"80",X"04",X"A8",X"04",X"D0",X"04",X"30",X"C4",X"58",X"C4",X"80",X"C4",
		X"A8",X"C4",X"D0",X"C4",X"00",X"01",X"04",X"F0",X"90",X"90",X"F0",X"01",X"04",X"60",X"F0",X"F0",
		X"60",X"01",X"04",X"60",X"60",X"60",X"60",X"01",X"04",X"00",X"60",X"60",X"60",X"01",X"04",X"60",
		X"60",X"60",X"00",X"01",X"04",X"00",X"F0",X"F0",X"00",X"01",X"04",X"00",X"70",X"70",X"00",X"01",
		X"04",X"00",X"E0",X"E0",X"00",X"CD",X"C2",X"20",X"E5",X"23",X"23",X"0E",X"06",X"EB",X"D5",X"CD",
		X"34",X"08",X"58",X"16",X"00",X"1D",X"19",X"D1",X"0E",X"00",X"1A",X"1B",X"CD",X"68",X"29",X"1A",
		X"1B",X"CD",X"68",X"29",X"1A",X"1B",X"CD",X"68",X"29",X"06",X"03",X"AF",X"CD",X"68",X"29",X"10",
		X"FA",X"0E",X"06",X"CD",X"34",X"08",X"E5",X"0E",X"00",X"7E",X"E6",X"F0",X"81",X"4F",X"23",X"10",
		X"F8",X"E1",X"2B",X"71",X"0E",X"0A",X"11",X"6E",X"40",X"E1",X"E5",X"D5",X"06",X"03",X"1A",X"BE",
		X"38",X"11",X"20",X"04",X"13",X"23",X"10",X"F6",X"D1",X"21",X"06",X"00",X"19",X"EB",X"E1",X"0D",
		X"20",X"E8",X"C9",X"D1",X"D5",X"06",X"00",X"0D",X"28",X"14",X"21",X"00",X"00",X"09",X"29",X"09",
		X"29",X"E5",X"19",X"2B",X"54",X"5D",X"01",X"06",X"00",X"09",X"EB",X"C1",X"ED",X"B8",X"D1",X"E1",
		X"06",X"03",X"7E",X"23",X"12",X"13",X"10",X"FA",X"EB",X"E5",X"CD",X"1A",X"11",X"CD",X"CD",X"0D",
		X"CD",X"A2",X"20",X"CD",X"17",X"12",X"85",X"29",X"C4",X"29",X"A4",X"29",X"E0",X"29",X"08",X"06",
		X"01",X"21",X"07",X"40",X"CD",X"5D",X"2E",X"CD",X"17",X"12",X"FF",X"29",X"BD",X"2A",X"60",X"2A",
		X"17",X"2B",X"CD",X"8E",X"2D",X"90",X"78",X"62",X"5F",X"5F",X"5F",X"00",X"CD",X"17",X"12",X"67",
		X"2B",X"67",X"2B",X"AD",X"2B",X"08",X"2C",X"CD",X"B1",X"17",X"E5",X"FD",X"E1",X"06",X"00",X"21",
		X"78",X"60",X"CD",X"B6",X"2D",X"EB",X"E1",X"E5",X"06",X"03",X"36",X"20",X"23",X"10",X"FB",X"E1",
		X"3E",X"1E",X"32",X"0C",X"40",X"06",X"03",X"0E",X"41",X"C5",X"3A",X"22",X"40",X"CD",X"EE",X"2D",
		X"C1",X"FD",X"36",X"00",X"0F",X"CD",X"CF",X"16",X"FD",X"7E",X"00",X"B7",X"20",X"F7",X"FD",X"36",
		X"00",X"3C",X"FD",X"7E",X"00",X"B7",X"20",X"0B",X"3A",X"0C",X"40",X"3D",X"32",X"0C",X"40",X"28",
		X"3A",X"18",X"EB",X"CD",X"8B",X"09",X"CB",X"67",X"28",X"54",X"71",X"C5",X"3A",X"22",X"40",X"B7",
		X"01",X"40",X"00",X"28",X"03",X"01",X"C0",X"FF",X"D5",X"EB",X"09",X"EB",X"3A",X"22",X"40",X"F6",
		X"90",X"0E",X"5F",X"CD",X"EE",X"2D",X"D1",X"C1",X"23",X"3A",X"22",X"40",X"B7",X"13",X"28",X"02",
		X"1B",X"1B",X"CD",X"8B",X"09",X"CB",X"67",X"20",X"F9",X"10",X"9E",X"21",X"6E",X"40",X"11",X"1B",
		X"F9",X"01",X"00",X"1E",X"7E",X"E6",X"F0",X"12",X"13",X"81",X"4F",X"7E",X"23",X"07",X"07",X"07",
		X"07",X"E6",X"F0",X"12",X"13",X"81",X"4F",X"10",X"EB",X"79",X"32",X"1A",X"F9",X"C9",X"CB",X"47",
		X"20",X"0F",X"CB",X"5F",X"20",X"0B",X"CB",X"4F",X"20",X"0B",X"CB",X"57",X"20",X"07",X"C3",X"D2",
		X"28",X"3E",X"FF",X"18",X"02",X"3E",X"01",X"81",X"FE",X"40",X"20",X"02",X"3E",X"5A",X"FE",X"5B",
		X"20",X"02",X"3E",X"41",X"4F",X"C3",X"B9",X"28",X"F5",X"07",X"07",X"07",X"07",X"CD",X"71",X"29",
		X"F1",X"E6",X"F0",X"08",X"7E",X"E6",X"F0",X"81",X"27",X"77",X"08",X"86",X"27",X"77",X"2B",X"0E",
		X"00",X"D0",X"0E",X"10",X"C9",X"CD",X"8E",X"2D",X"90",X"20",X"08",X"43",X"6F",X"6E",X"67",X"72",
		X"61",X"74",X"75",X"6C",X"61",X"74",X"69",X"6F",X"6E",X"73",X"20",X"50",X"6C",X"61",X"79",X"65",
		X"72",X"20",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"10",X"08",X"46",X"65",X"6C",X"69",X"63",X"69",
		X"74",X"61",X"74",X"69",X"6F",X"6E",X"73",X"20",X"61",X"75",X"20",X"6A",X"6F",X"75",X"65",X"75",
		X"72",X"20",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"20",X"08",X"47",X"72",X"61",X"74",X"75",X"6C",
		X"69",X"65",X"72",X"65",X"2C",X"20",X"53",X"70",X"69",X"65",X"6C",X"65",X"72",X"20",X"00",X"C9",
		X"CD",X"8E",X"2D",X"90",X"20",X"08",X"46",X"65",X"6C",X"69",X"63",X"69",X"74",X"61",X"63",X"69",
		X"6F",X"6E",X"65",X"73",X"20",X"6A",X"75",X"67",X"61",X"64",X"6F",X"72",X"20",X"00",X"C9",X"CD",
		X"8E",X"2D",X"90",X"08",X"20",X"59",X"6F",X"75",X"20",X"68",X"61",X"76",X"65",X"20",X"6A",X"6F",
		X"69",X"6E",X"65",X"64",X"20",X"74",X"68",X"65",X"20",X"69",X"6D",X"6D",X"6F",X"72",X"74",X"61",
		X"6C",X"73",X"00",X"CD",X"8E",X"2D",X"90",X"10",X"30",X"69",X"6E",X"20",X"74",X"68",X"65",X"20",
		X"46",X"52",X"45",X"4E",X"5A",X"59",X"20",X"68",X"61",X"6C",X"6C",X"20",X"6F",X"66",X"20",X"66",
		X"61",X"6D",X"65",X"00",X"CD",X"8E",X"2D",X"90",X"18",X"50",X"45",X"6E",X"74",X"65",X"72",X"20",
		X"79",X"6F",X"75",X"72",X"20",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"73",X"3A",X"00",X"C9",
		X"CD",X"8E",X"2D",X"90",X"08",X"20",X"56",X"6F",X"75",X"73",X"20",X"61",X"76",X"65",X"7A",X"20",
		X"6A",X"6F",X"69",X"6E",X"74",X"20",X"6C",X"65",X"73",X"20",X"69",X"6D",X"6D",X"6F",X"72",X"74",
		X"65",X"6C",X"73",X"00",X"CD",X"8E",X"2D",X"90",X"18",X"30",X"64",X"75",X"20",X"70",X"61",X"6E",
		X"74",X"68",X"65",X"6F",X"6E",X"20",X"46",X"52",X"45",X"4E",X"5A",X"59",X"2E",X"00",X"CD",X"8E",
		X"2D",X"90",X"08",X"50",X"49",X"6E",X"73",X"63",X"72",X"69",X"72",X"65",X"20",X"76",X"6F",X"73",
		X"20",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"73",X"3A",X"00",X"C9",X"CD",X"8E",X"2D",
		X"90",X"08",X"20",X"44",X"61",X"73",X"20",X"57",X"61",X"72",X"20",X"65",X"69",X"6E",X"20",X"52",
		X"75",X"68",X"6D",X"76",X"6F",X"6C",X"6C",X"65",X"72",X"20",X"53",X"69",X"65",X"67",X"21",X"00",
		X"CD",X"8E",X"2D",X"90",X"08",X"40",X"54",X"72",X"61",X"67",X"20",X"44",X"65",X"69",X"6E",X"65",
		X"6E",X"20",X"4E",X"61",X"6D",X"65",X"6E",X"20",X"69",X"6E",X"20",X"64",X"69",X"65",X"00",X"CD",
		X"8E",X"2D",X"90",X"10",X"50",X"48",X"65",X"6C",X"64",X"65",X"6E",X"6C",X"69",X"73",X"74",X"65",
		X"20",X"65",X"69",X"6E",X"21",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"04",X"20",X"53",X"65",X"20",
		X"70",X"75",X"6E",X"74",X"61",X"6A",X"65",X"20",X"65",X"73",X"74",X"61",X"20",X"65",X"6E",X"74",
		X"72",X"65",X"20",X"6C",X"6F",X"73",X"20",X"64",X"69",X"65",X"7A",X"00",X"CD",X"8E",X"2D",X"90",
		X"08",X"30",X"6D",X"65",X"6A",X"6F",X"72",X"65",X"73",X"2E",X"00",X"CD",X"8E",X"2D",X"90",X"18",
		X"50",X"45",X"6E",X"74",X"72",X"65",X"20",X"73",X"75",X"73",X"20",X"69",X"6E",X"69",X"63",X"69",
		X"61",X"6C",X"65",X"73",X"3A",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"08",X"80",X"4D",X"6F",X"76",
		X"65",X"20",X"73",X"74",X"69",X"63",X"6B",X"20",X"74",X"6F",X"20",X"63",X"68",X"61",X"6E",X"67",
		X"65",X"20",X"6C",X"65",X"74",X"74",X"65",X"72",X"00",X"CD",X"8E",X"2D",X"90",X"08",X"90",X"74",
		X"68",X"65",X"6E",X"20",X"70",X"72",X"65",X"73",X"73",X"20",X"46",X"49",X"52",X"45",X"20",X"74",
		X"6F",X"20",X"73",X"74",X"6F",X"72",X"65",X"20",X"69",X"74",X"2E",X"00",X"C9",X"CD",X"8E",X"2D",
		X"90",X"04",X"80",X"50",X"6F",X"75",X"73",X"73",X"65",X"7A",X"20",X"62",X"61",X"74",X"6F",X"6E",
		X"6E",X"65",X"74",X"20",X"70",X"6F",X"75",X"72",X"20",X"76",X"6F",X"73",X"00",X"CD",X"8E",X"2D",
		X"90",X"04",X"90",X"69",X"6E",X"69",X"74",X"69",X"61",X"6C",X"65",X"73",X"2E",X"20",X"50",X"6F",
		X"75",X"73",X"73",X"65",X"7A",X"20",X"46",X"49",X"52",X"45",X"20",X"71",X"75",X"61",X"6E",X"64",
		X"00",X"CD",X"8E",X"2D",X"90",X"04",X"A0",X"6C",X"65",X"74",X"74",X"72",X"65",X"20",X"63",X"6F",
		X"72",X"72",X"65",X"63",X"74",X"65",X"00",X"C9",X"CD",X"8E",X"2D",X"90",X"04",X"80",X"4D",X"6F",
		X"76",X"69",X"65",X"6E",X"64",X"6F",X"20",X"6C",X"61",X"20",X"70",X"61",X"6C",X"61",X"6E",X"63",
		X"61",X"20",X"70",X"61",X"72",X"61",X"00",X"CD",X"8E",X"2D",X"90",X"04",X"90",X"63",X"61",X"6D",
		X"62",X"69",X"61",X"72",X"20",X"6C",X"61",X"73",X"20",X"6C",X"65",X"74",X"72",X"61",X"73",X"2C",
		X"20",X"6C",X"75",X"65",X"67",X"6F",X"00",X"CD",X"8E",X"2D",X"90",X"04",X"A0",X"61",X"70",X"6C",
		X"61",X"73",X"74",X"65",X"20",X"65",X"6C",X"20",X"62",X"6F",X"74",X"6F",X"6E",X"20",X"64",X"65",
		X"20",X"64",X"69",X"73",X"70",X"61",X"72",X"6F",X"00",X"CD",X"8E",X"2D",X"90",X"04",X"B0",X"70",
		X"61",X"72",X"61",X"20",X"72",X"65",X"74",X"65",X"6E",X"65",X"72",X"6C",X"61",X"73",X"2E",X"00",
		X"C9",X"E5",X"C5",X"F5",X"4F",X"7E",X"B7",X"20",X"1D",X"3A",X"23",X"40",X"CB",X"57",X"20",X"16",
		X"3A",X"0E",X"40",X"B7",X"28",X"10",X"47",X"21",X"39",X"80",X"D5",X"11",X"0F",X"00",X"7E",X"B7",
		X"28",X"08",X"19",X"10",X"F9",X"D1",X"F1",X"C1",X"E1",X"C9",X"D1",X"7A",X"FE",X"FE",X"D2",X"DF",
		X"2C",X"FE",X"08",X"38",X"2A",X"7B",X"FE",X"F6",X"30",X"1F",X"FE",X"05",X"38",X"1B",X"7A",X"CB",
		X"41",X"28",X"03",X"ED",X"44",X"57",X"7B",X"CB",X"51",X"28",X"03",X"ED",X"44",X"5F",X"92",X"FE",
		X"F6",X"30",X"12",X"FE",X"06",X"30",X"CF",X"18",X"0C",X"79",X"E6",X"03",X"4F",X"18",X"06",X"79",
		X"E6",X"0C",X"4F",X"18",X"00",X"E5",X"06",X"0F",X"AF",X"77",X"23",X"10",X"FC",X"CD",X"84",X"1C",
		X"21",X"A9",X"19",X"09",X"4E",X"21",X"58",X"2D",X"09",X"09",X"09",X"DD",X"70",X"08",X"DD",X"70",
		X"0A",X"7E",X"23",X"F3",X"DD",X"77",X"0C",X"7E",X"DD",X"77",X"0D",X"FB",X"23",X"DD",X"36",X"07",
		X"01",X"46",X"23",X"4E",X"23",X"56",X"DD",X"7E",X"09",X"80",X"47",X"DD",X"7E",X"0B",X"81",X"4F",
		X"E1",X"7A",X"F6",X"03",X"F3",X"77",X"23",X"70",X"23",X"71",X"23",X"70",X"23",X"71",X"FB",X"F1",
		X"C1",X"E1",X"36",X"0A",X"CD",X"CF",X"16",X"DD",X"CB",X"00",X"6E",X"20",X"04",X"7E",X"B7",X"20",
		X"F3",X"3A",X"1F",X"40",X"87",X"87",X"C6",X"05",X"4F",X"3A",X"0F",X"40",X"CB",X"3F",X"B9",X"38",
		X"01",X"79",X"77",X"0E",X"10",X"C3",X"25",X"22",X"05",X"39",X"00",X"00",X"00",X"00",X"05",X"39",
		X"07",X"01",X"60",X"00",X"05",X"39",X"08",X"02",X"20",X"00",X"05",X"39",X"08",X"04",X"A0",X"00",
		X"05",X"39",X"06",X"0B",X"80",X"00",X"05",X"39",X"FF",X"04",X"90",X"00",X"05",X"39",X"FF",X"02",
		X"10",X"00",X"05",X"39",X"00",X"01",X"50",X"00",X"05",X"39",X"06",X"00",X"40",X"00",X"E1",X"46",
		X"23",X"5E",X"23",X"56",X"23",X"EB",X"CD",X"B6",X"2D",X"EB",X"4E",X"CB",X"B9",X"CD",X"EE",X"2D",
		X"47",X"3A",X"22",X"40",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"23",X"7E",X"B7",X"78",X"C2",
		X"9A",X"2D",X"23",X"E9",X"06",X"90",X"3A",X"22",X"40",X"B7",X"3E",X"07",X"20",X"15",X"A5",X"B0",
		X"D3",X"4B",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"01",X"00",
		X"64",X"09",X"C9",X"A5",X"B0",X"CB",X"DF",X"D3",X"4B",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",
		X"1D",X"CB",X"3C",X"CB",X"1D",X"44",X"4D",X"21",X"FF",X"7F",X"B7",X"ED",X"42",X"C9",X"E5",X"21",
		X"00",X"00",X"06",X"00",X"09",X"29",X"29",X"29",X"09",X"01",X"E1",X"C2",X"09",X"D5",X"F5",X"EB",
		X"3A",X"22",X"40",X"B7",X"1A",X"20",X"26",X"B7",X"F2",X"0F",X"2E",X"01",X"60",X"00",X"09",X"3E",
		X"09",X"01",X"1F",X"00",X"08",X"F1",X"F5",X"F3",X"D3",X"4B",X"1A",X"E6",X"7F",X"13",X"77",X"23",
		X"36",X"00",X"FB",X"09",X"08",X"3D",X"C2",X"14",X"2E",X"F1",X"D1",X"E1",X"C9",X"B7",X"F2",X"35",
		X"2E",X"01",X"A0",X"FF",X"09",X"3E",X"09",X"01",X"E1",X"FF",X"08",X"F1",X"F5",X"F3",X"D3",X"4B",
		X"1A",X"E6",X"7F",X"13",X"77",X"2B",X"36",X"00",X"FB",X"09",X"08",X"3D",X"C2",X"3A",X"2E",X"F1",
		X"D1",X"E1",X"C9",X"C5",X"06",X"00",X"EB",X"CD",X"B6",X"2D",X"EB",X"08",X"C1",X"CB",X"81",X"78",
		X"3D",X"20",X"02",X"CB",X"C1",X"7E",X"CB",X"40",X"20",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"2B",X"23",X"E6",X"0F",X"20",X"08",X"CB",X"41",X"20",X"06",X"3E",X"20",X"18",X"08",
		X"CB",X"C1",X"C6",X"90",X"27",X"C6",X"40",X"27",X"E5",X"C5",X"4F",X"08",X"CD",X"EE",X"2D",X"08",
		X"C1",X"E1",X"3A",X"22",X"40",X"B7",X"20",X"03",X"13",X"18",X"01",X"1B",X"10",X"C1",X"C9",X"AF",
		X"32",X"5C",X"40",X"2A",X"0A",X"40",X"7D",X"FE",X"20",X"30",X"04",X"2E",X"02",X"18",X"06",X"FE",
		X"F0",X"38",X"02",X"2E",X"F8",X"7C",X"FE",X"B4",X"38",X"02",X"26",X"A0",X"22",X"24",X"40",X"3A",
		X"20",X"40",X"47",X"3A",X"0F",X"40",X"0F",X"0F",X"E6",X"07",X"80",X"32",X"10",X"40",X"1E",X"00",
		X"3E",X"28",X"CD",X"0E",X"18",X"21",X"10",X"40",X"35",X"20",X"F5",X"2A",X"24",X"40",X"3E",X"1E",
		X"32",X"A1",X"F8",X"18",X"07",X"11",X"80",X"54",X"EB",X"11",X"02",X"00",X"D5",X"E5",X"CD",X"89",
		X"19",X"E1",X"D1",X"DA",X"65",X"17",X"7B",X"B7",X"20",X"0E",X"D5",X"E5",X"CD",X"60",X"30",X"C1",
		X"D1",X"3E",X"3C",X"CD",X"0E",X"18",X"60",X"69",X"DD",X"75",X"09",X"DD",X"74",X"0B",X"AF",X"DD",
		X"77",X"08",X"DD",X"77",X"0A",X"21",X"03",X"3A",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",
		X"07",X"01",X"DD",X"36",X"06",X"02",X"16",X"00",X"DD",X"36",X"00",X"86",X"AF",X"CD",X"E0",X"2F",
		X"3E",X"3C",X"CD",X"0E",X"18",X"DD",X"CB",X"00",X"B6",X"FD",X"21",X"AD",X"40",X"D5",X"FD",X"7E",
		X"09",X"DD",X"96",X"09",X"06",X"00",X"28",X"08",X"06",X"02",X"30",X"04",X"06",X"01",X"ED",X"44",
		X"57",X"FD",X"7E",X"0B",X"83",X"5A",X"C6",X"01",X"FE",X"B0",X"DA",X"5F",X"2F",X"3E",X"AF",X"DD",
		X"96",X"0B",X"0E",X"00",X"28",X"08",X"0E",X"08",X"30",X"04",X"0E",X"04",X"ED",X"44",X"57",X"78",
		X"81",X"42",X"4B",X"D1",X"CD",X"E0",X"2F",X"DD",X"CB",X"00",X"76",X"28",X"29",X"DD",X"CB",X"00",
		X"B6",X"CD",X"06",X"1C",X"14",X"D5",X"21",X"23",X"3A",X"15",X"CA",X"90",X"2F",X"21",X"37",X"3A",
		X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"07",X"01",X"01",X"02",X"01",X"CD",X"FB",X"20",
		X"D1",X"7A",X"FE",X"03",X"28",X"05",X"CD",X"CF",X"16",X"18",X"8E",X"AF",X"DD",X"77",X"08",X"DD",
		X"77",X"0A",X"2F",X"32",X"5C",X"40",X"CD",X"68",X"30",X"21",X"4B",X"3A",X"DD",X"75",X"0C",X"DD",
		X"74",X"0D",X"DD",X"36",X"06",X"04",X"3E",X"3C",X"CD",X"0E",X"18",X"DD",X"36",X"00",X"81",X"3E",
		X"0A",X"CD",X"0E",X"18",X"7B",X"FE",X"07",X"30",X"01",X"1C",X"2A",X"24",X"40",X"C3",X"08",X"2F",
		X"E6",X"0F",X"C2",X"EB",X"2F",X"01",X"00",X"00",X"C3",X"19",X"30",X"C5",X"08",X"21",X"4B",X"30",
		X"06",X"00",X"4B",X"09",X"09",X"7E",X"DD",X"77",X"06",X"23",X"7E",X"C1",X"B8",X"30",X"01",X"47",
		X"B9",X"30",X"01",X"4F",X"08",X"CB",X"57",X"28",X"06",X"08",X"78",X"ED",X"44",X"47",X"08",X"CB",
		X"47",X"28",X"06",X"08",X"79",X"ED",X"44",X"4F",X"08",X"DD",X"71",X"08",X"DD",X"70",X"0A",X"C9",
		X"4F",X"06",X"00",X"21",X"A9",X"19",X"09",X"5E",X"50",X"21",X"37",X"30",X"19",X"7E",X"DD",X"77",
		X"08",X"23",X"7E",X"DD",X"77",X"0A",X"C9",X"00",X"00",X"01",X"FF",X"01",X"00",X"01",X"01",X"00",
		X"01",X"FF",X"01",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"03",X"01",X"01",X"01",X"01",
		X"03",X"01",X"04",X"01",X"06",X"01",X"08",X"01",X"0A",X"01",X"0C",X"E1",X"22",X"9A",X"F8",X"C9",
		X"CD",X"5B",X"30",X"7D",X"1C",X"02",X"47",X"FF",X"CD",X"5B",X"30",X"7E",X"03",X"02",X"05",X"01",
		X"15",X"47",X"FF",X"CD",X"5B",X"30",X"7C",X"1B",X"1C",X"07",X"17",X"1B",X"18",X"47",X"FF",X"CD",
		X"5B",X"30",X"7C",X"1B",X"1C",X"16",X"06",X"0A",X"0F",X"47",X"FF",X"CD",X"5B",X"30",X"7E",X"0A",
		X"0F",X"16",X"17",X"15",X"0A",X"1C",X"47",X"FF",X"CD",X"5B",X"30",X"7B",X"0E",X"07",X"0A",X"0F",
		X"47",X"FF",X"7D",X"10",X"09",X"0B",X"11",X"45",X"FF",X"CD",X"1A",X"11",X"CD",X"99",X"0D",X"CD",
		X"5F",X"11",X"FD",X"21",X"84",X"31",X"DD",X"21",X"35",X"31",X"21",X"10",X"0C",X"11",X"04",X"05",
		X"CD",X"EB",X"30",X"FD",X"21",X"8A",X"31",X"DD",X"21",X"58",X"31",X"21",X"10",X"54",X"11",X"05",
		X"08",X"CD",X"E7",X"30",X"C9",X"FD",X"21",X"95",X"31",X"DD",X"21",X"58",X"31",X"21",X"3D",X"02",
		X"11",X"03",X"04",X"CD",X"EB",X"30",X"C9",X"06",X"FF",X"18",X"02",X"06",X"00",X"0E",X"01",X"E5",
		X"DD",X"E5",X"DD",X"7E",X"00",X"A1",X"CA",X"1B",X"31",X"C5",X"D5",X"E5",X"CD",X"B4",X"2D",X"EB",
		X"FD",X"E5",X"E1",X"CD",X"6F",X"15",X"E1",X"D1",X"C1",X"78",X"B7",X"CA",X"1B",X"31",X"06",X"00",
		X"DD",X"E3",X"DD",X"E3",X"DD",X"E3",X"DD",X"E3",X"10",X"F6",X"47",X"7D",X"83",X"6F",X"DD",X"23",
		X"DD",X"7E",X"00",X"DD",X"B6",X"FF",X"C2",X"F2",X"30",X"DD",X"E1",X"E1",X"7C",X"82",X"67",X"CB",
		X"21",X"C2",X"EF",X"30",X"C9",X"CE",X"DB",X"DB",X"FB",X"73",X"00",X"03",X"03",X"FF",X"FF",X"03",
		X"03",X"00",X"FF",X"FF",X"DB",X"DB",X"C3",X"00",X"FF",X"FF",X"1B",X"1B",X"FF",X"EE",X"00",X"FF",
		X"FF",X"0E",X"1C",X"38",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"1B",X"1B",X"03",X"03",X"00",X"FF",
		X"FF",X"1B",X"1B",X"FF",X"EE",X"00",X"FF",X"FF",X"DB",X"DB",X"C3",X"C3",X"00",X"FF",X"FF",X"0E",
		X"1C",X"38",X"FF",X"FF",X"00",X"E3",X"F3",X"FB",X"DF",X"CF",X"C7",X"00",X"07",X"0F",X"FC",X"FC",
		X"0F",X"07",X"00",X"00",X"01",X"04",X"40",X"E0",X"E0",X"40",X"01",X"09",X"7C",X"84",X"84",X"84",
		X"FC",X"84",X"84",X"84",X"F8",X"01",X"04",X"C0",X"C0",X"C0",X"00",X"3A",X"12",X"40",X"CB",X"5F",
		X"CA",X"AB",X"31",X"CB",X"57",X"CA",X"10",X"33",X"C3",X"BD",X"33",X"CB",X"57",X"C2",X"46",X"32",
		X"21",X"E5",X"35",X"CD",X"0F",X"35",X"11",X"94",X"C8",X"21",X"83",X"3B",X"CD",X"56",X"35",X"11",
		X"15",X"C9",X"21",X"84",X"4A",X"CD",X"56",X"35",X"11",X"2E",X"C9",X"21",X"8C",X"48",X"CD",X"56",
		X"35",X"21",X"71",X"3A",X"11",X"88",X"40",X"CD",X"60",X"35",X"21",X"8D",X"3A",X"11",X"9C",X"58",
		X"CD",X"60",X"35",X"21",X"B1",X"3A",X"11",X"8E",X"55",X"CD",X"60",X"35",X"DD",X"36",X"06",X"01",
		X"21",X"95",X"3A",X"11",X"93",X"5C",X"CD",X"60",X"35",X"DD",X"36",X"06",X"01",X"C1",X"C1",X"D1",
		X"DD",X"E1",X"CD",X"CF",X"16",X"3A",X"1F",X"40",X"B7",X"FA",X"10",X"32",X"FE",X"0D",X"30",X"F2",
		X"21",X"63",X"3A",X"CD",X"4D",X"35",X"3E",X"32",X"CD",X"0E",X"18",X"D5",X"DD",X"E3",X"D1",X"21",
		X"79",X"3A",X"CD",X"4D",X"35",X"3E",X"3C",X"CD",X"0E",X"18",X"01",X"79",X"21",X"CD",X"35",X"17",
		X"3E",X"5A",X"CD",X"0E",X"18",X"21",X"8D",X"3A",X"CD",X"4D",X"35",X"D5",X"DD",X"E3",X"D1",X"3E",
		X"1E",X"CD",X"0E",X"18",X"18",X"BC",X"CD",X"8B",X"30",X"21",X"21",X"36",X"CD",X"0F",X"35",X"11",
		X"6A",X"C7",X"21",X"84",X"3C",X"CD",X"56",X"35",X"11",X"BC",X"C7",X"21",X"94",X"3C",X"CD",X"56",
		X"35",X"CD",X"F4",X"32",X"CD",X"CF",X"16",X"3A",X"5C",X"40",X"B7",X"20",X"0C",X"3A",X"AD",X"40",
		X"CB",X"6F",X"28",X"F0",X"CD",X"06",X"33",X"18",X"37",X"CD",X"F4",X"32",X"CD",X"C9",X"32",X"11",
		X"6E",X"52",X"01",X"E8",X"2E",X"CD",X"35",X"17",X"11",X"AA",X"52",X"01",X"E8",X"2E",X"CD",X"35",
		X"17",X"11",X"94",X"28",X"01",X"E8",X"2E",X"CD",X"35",X"17",X"11",X"94",X"5A",X"01",X"E8",X"2E",
		X"CD",X"35",X"17",X"CD",X"CF",X"16",X"3A",X"AD",X"40",X"CB",X"6F",X"28",X"F6",X"CD",X"E1",X"32",
		X"CD",X"B6",X"32",X"C3",X"65",X"17",X"11",X"4A",X"C8",X"21",X"84",X"56",X"CD",X"56",X"35",X"11",
		X"5A",X"C8",X"21",X"94",X"56",X"CD",X"56",X"35",X"C9",X"11",X"0E",X"C8",X"21",X"8B",X"41",X"CD",
		X"56",X"35",X"11",X"1C",X"C8",X"21",X"95",X"41",X"CD",X"56",X"35",X"21",X"5D",X"36",X"CD",X"0F",
		X"35",X"11",X"2A",X"C8",X"21",X"84",X"56",X"CD",X"56",X"35",X"11",X"3A",X"C8",X"21",X"94",X"56",
		X"CD",X"56",X"35",X"C9",X"11",X"70",X"C8",X"21",X"84",X"45",X"CD",X"56",X"35",X"11",X"82",X"C8",
		X"21",X"94",X"45",X"CD",X"56",X"35",X"11",X"6A",X"C8",X"21",X"8C",X"56",X"CD",X"56",X"35",X"C9",
		X"21",X"D5",X"36",X"CD",X"0F",X"35",X"CD",X"72",X"34",X"11",X"E3",X"CC",X"21",X"88",X"3C",X"CD",
		X"56",X"35",X"11",X"E3",X"CC",X"21",X"88",X"4C",X"CD",X"56",X"35",X"11",X"E3",X"CC",X"21",X"9C",
		X"44",X"CD",X"56",X"35",X"11",X"F5",X"CC",X"21",X"9C",X"54",X"CD",X"56",X"35",X"11",X"C5",X"CD",
		X"21",X"83",X"5C",X"CD",X"56",X"35",X"11",X"CB",X"CD",X"21",X"90",X"5C",X"CD",X"56",X"35",X"11",
		X"C5",X"CD",X"21",X"9C",X"5C",X"CD",X"56",X"35",X"21",X"0F",X"3B",X"11",X"8C",X"3F",X"CD",X"60",
		X"35",X"DD",X"36",X"06",X"01",X"21",X"25",X"3B",X"11",X"8C",X"48",X"CD",X"60",X"35",X"DD",X"36",
		X"06",X"01",X"21",X"B1",X"3A",X"11",X"88",X"5E",X"CD",X"60",X"35",X"DD",X"36",X"06",X"01",X"21",
		X"95",X"3A",X"11",X"9C",X"5E",X"CD",X"60",X"35",X"DD",X"36",X"06",X"01",X"C1",X"D1",X"E1",X"DD",
		X"E1",X"CD",X"CF",X"16",X"CD",X"4D",X"34",X"28",X"F8",X"F3",X"0A",X"CB",X"97",X"02",X"1A",X"CB",
		X"97",X"12",X"7E",X"E6",X"F9",X"77",X"DD",X"7E",X"00",X"E6",X"F9",X"DD",X"77",X"00",X"FB",X"3E",
		X"02",X"32",X"23",X"40",X"01",X"01",X"02",X"CD",X"FB",X"20",X"C3",X"65",X"17",X"21",X"99",X"36",
		X"CD",X"0F",X"35",X"CD",X"72",X"34",X"11",X"0B",X"CB",X"21",X"84",X"44",X"CD",X"56",X"35",X"11",
		X"49",X"CB",X"21",X"98",X"44",X"CD",X"56",X"35",X"11",X"87",X"CB",X"21",X"92",X"47",X"CD",X"56",
		X"35",X"21",X"D9",X"3A",X"11",X"90",X"3A",X"CD",X"60",X"35",X"DD",X"36",X"06",X"01",X"21",X"FF",
		X"3A",X"11",X"8C",X"54",X"CD",X"60",X"35",X"21",X"CD",X"3A",X"11",X"84",X"3C",X"CD",X"60",X"35",
		X"DD",X"36",X"06",X"01",X"21",X"CD",X"3A",X"11",X"9E",X"3C",X"CD",X"60",X"35",X"DD",X"36",X"06",
		X"01",X"DD",X"E1",X"E1",X"D1",X"C1",X"CD",X"CF",X"16",X"CD",X"4D",X"34",X"28",X"F8",X"F3",X"0A",
		X"E6",X"FB",X"02",X"7E",X"E6",X"FB",X"77",X"DD",X"7E",X"00",X"E6",X"FB",X"DD",X"77",X"00",X"D5",
		X"DD",X"E1",X"21",X"ED",X"3A",X"DD",X"74",X"0D",X"DD",X"75",X"0C",X"FB",X"3E",X"05",X"32",X"23",
		X"40",X"01",X"01",X"02",X"CD",X"FB",X"20",X"CD",X"98",X"30",X"C3",X"65",X"17",X"FD",X"21",X"1B",
		X"80",X"CD",X"5D",X"34",X"FD",X"21",X"2A",X"80",X"CD",X"5D",X"34",X"AF",X"C9",X"FD",X"7E",X"01",
		X"FE",X"80",X"D8",X"FE",X"A8",X"D0",X"FD",X"7E",X"02",X"FE",X"38",X"D8",X"FE",X"66",X"D0",X"33",
		X"33",X"C9",X"3A",X"22",X"40",X"B7",X"20",X"2C",X"DD",X"21",X"B0",X"82",X"11",X"20",X"00",X"CD",
		X"B9",X"34",X"06",X"0B",X"CD",X"C7",X"34",X"CD",X"B9",X"34",X"F3",X"21",X"80",X"34",X"E5",X"CD",
		X"92",X"25",X"E1",X"CD",X"EB",X"25",X"21",X"A8",X"34",X"CD",X"EB",X"25",X"21",X"80",X"64",X"CD",
		X"92",X"25",X"FB",X"C9",X"DD",X"21",X"4F",X"86",X"11",X"E0",X"FF",X"CD",X"E4",X"34",X"06",X"0B",
		X"CD",X"F2",X"34",X"CD",X"E4",X"34",X"C3",X"8A",X"34",X"06",X"05",X"DD",X"E5",X"E1",X"3A",X"BA",
		X"F8",X"77",X"23",X"10",X"FC",X"06",X"01",X"3A",X"BA",X"F8",X"E6",X"F0",X"4F",X"DD",X"7E",X"00",
		X"E6",X"0F",X"B1",X"DD",X"77",X"00",X"DD",X"7E",X"05",X"E6",X"0F",X"B1",X"DD",X"77",X"05",X"DD",
		X"19",X"10",X"EA",X"C9",X"06",X"05",X"DD",X"E5",X"E1",X"3A",X"BA",X"F8",X"77",X"2B",X"10",X"FC",
		X"06",X"01",X"3A",X"BA",X"F8",X"E6",X"0F",X"4F",X"DD",X"7E",X"00",X"E6",X"F0",X"B1",X"DD",X"77",
		X"00",X"DD",X"7E",X"FB",X"E6",X"F0",X"B1",X"DD",X"77",X"FB",X"DD",X"19",X"10",X"EA",X"C9",X"3A",
		X"22",X"40",X"B7",X"20",X"1A",X"DD",X"21",X"B0",X"82",X"11",X"1B",X"00",X"0E",X"0C",X"06",X"05",
		X"7E",X"23",X"DD",X"77",X"00",X"DD",X"23",X"10",X"F7",X"DD",X"19",X"0D",X"20",X"F0",X"C9",X"DD",
		X"21",X"4F",X"86",X"11",X"E5",X"FF",X"0E",X"0C",X"06",X"05",X"7E",X"23",X"07",X"07",X"07",X"07",
		X"DD",X"77",X"00",X"DD",X"2B",X"10",X"F3",X"DD",X"19",X"0D",X"20",X"EC",X"C9",X"F3",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"FB",X"C9",X"F3",X"CD",X"B4",X"2D",X"EB",X"CD",X"6F",X"15",X"FB",X"C9",
		X"D5",X"E5",X"CD",X"89",X"19",X"E1",X"D1",X"D8",X"DD",X"73",X"09",X"DD",X"72",X"0B",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"07",X"01",X"DD",X"36",X"06",X"02",X"DD",X"36",X"00",X"86",
		X"E1",X"DD",X"E5",X"E9",X"DD",X"21",X"26",X"40",X"DD",X"CB",X"21",X"DE",X"DD",X"CB",X"21",X"D6",
		X"DD",X"CB",X"21",X"CE",X"DD",X"CB",X"21",X"C6",X"DD",X"CB",X"1B",X"DE",X"DD",X"CB",X"27",X"D6",
		X"DD",X"CB",X"20",X"CE",X"DD",X"CB",X"22",X"C6",X"DD",X"CB",X"09",X"DE",X"DD",X"CB",X"09",X"D6",
		X"DD",X"CB",X"09",X"CE",X"DD",X"CB",X"09",X"C6",X"DD",X"CB",X"03",X"DE",X"DD",X"CB",X"0F",X"D6",
		X"DD",X"CB",X"08",X"CE",X"DD",X"CB",X"0A",X"C6",X"DD",X"CB",X"09",X"FE",X"DD",X"CB",X"27",X"9E",
		X"DD",X"CB",X"2D",X"96",X"DD",X"CB",X"26",X"8E",X"DD",X"CB",X"27",X"86",X"DD",X"CB",X"27",X"8E",
		X"DD",X"CB",X"28",X"86",X"C9",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"55",X"55",X"55",X"77",X"77",X"55",X"55",X"55",X"77",X"77",X"55",X"55",X"55",X"77",X"74",X"41",
		X"11",X"13",X"33",X"74",X"46",X"66",X"63",X"33",X"74",X"46",X"66",X"63",X"33",X"74",X"46",X"66",
		X"63",X"33",X"74",X"46",X"66",X"63",X"33",X"74",X"46",X"66",X"63",X"33",X"74",X"46",X"66",X"63",
		X"33",X"77",X"77",X"77",X"77",X"77",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",
		X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",
		X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",
		X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"77",X"77",X"77",
		X"77",X"77",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",
		X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"31",X"33",X"13",X"33",X"73",X"33",X"33",X"33",X"33",
		X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"73",
		X"33",X"33",X"33",X"33",X"73",X"33",X"33",X"33",X"33",X"77",X"77",X"77",X"77",X"77",X"76",X"66",
		X"22",X"26",X"66",X"76",X"66",X"22",X"26",X"66",X"76",X"66",X"22",X"26",X"66",X"76",X"66",X"CC",
		X"C6",X"66",X"7C",X"3C",X"33",X"3C",X"3C",X"7C",X"3C",X"33",X"3C",X"3C",X"7C",X"3C",X"11",X"1C",
		X"3C",X"7C",X"3C",X"11",X"1C",X"3C",X"7C",X"3C",X"11",X"1C",X"3C",X"7C",X"3C",X"11",X"1C",X"3C",
		X"7C",X"CC",X"11",X"1C",X"CC",X"77",X"77",X"77",X"77",X"77",X"73",X"33",X"33",X"33",X"33",X"73",
		X"33",X"55",X"53",X"33",X"73",X"33",X"55",X"53",X"33",X"73",X"66",X"55",X"53",X"33",X"73",X"66",
		X"55",X"53",X"33",X"73",X"33",X"55",X"56",X"63",X"73",X"33",X"55",X"56",X"63",X"73",X"66",X"55",
		X"56",X"63",X"73",X"66",X"55",X"56",X"63",X"77",X"77",X"77",X"77",X"77",X"73",X"33",X"33",X"33",
		X"33",X"21",X"1F",X"40",X"34",X"7E",X"32",X"20",X"40",X"CD",X"89",X"19",X"DA",X"65",X"17",X"CD",
		X"FB",X"22",X"AF",X"0E",X"FF",X"CD",X"BD",X"37",X"DD",X"36",X"06",X"02",X"DD",X"36",X"07",X"01",
		X"DD",X"36",X"00",X"86",X"CD",X"B1",X"17",X"3A",X"0F",X"40",X"FE",X"2D",X"30",X"02",X"3E",X"2D",
		X"47",X"CD",X"39",X"10",X"E6",X"F8",X"0F",X"0F",X"0F",X"80",X"77",X"CD",X"CF",X"16",X"DD",X"CB",
		X"00",X"6E",X"20",X"04",X"7E",X"B7",X"20",X"F3",X"0E",X"00",X"FD",X"21",X"AD",X"40",X"C5",X"FD",
		X"7E",X"09",X"D6",X"01",X"DD",X"96",X"09",X"57",X"01",X"00",X"00",X"28",X"06",X"06",X"01",X"38",
		X"02",X"06",X"02",X"FD",X"7E",X"0B",X"C6",X"02",X"DD",X"96",X"0B",X"5F",X"28",X"06",X"0E",X"04",
		X"38",X"02",X"0E",X"08",X"78",X"81",X"C1",X"CD",X"E4",X"37",X"E5",X"E6",X"0F",X"28",X"19",X"21",
		X"23",X"40",X"CB",X"4E",X"28",X"03",X"AF",X"18",X"0F",X"CB",X"46",X"CC",X"D8",X"15",X"CB",X"47",
		X"20",X"04",X"CB",X"4F",X"28",X"02",X"E6",X"03",X"B9",X"E1",X"28",X"04",X"4F",X"CD",X"BD",X"37",
		X"CD",X"CF",X"16",X"DD",X"CB",X"00",X"6E",X"CA",X"5A",X"37",X"C3",X"5A",X"22",X"E5",X"CD",X"20",
		X"30",X"21",X"D2",X"37",X"19",X"7E",X"23",X"66",X"F3",X"DD",X"77",X"0C",X"DD",X"74",X"0D",X"FB",
		X"E1",X"C9",X"57",X"39",X"5F",X"39",X"5F",X"39",X"5F",X"39",X"6B",X"39",X"77",X"39",X"77",X"39",
		X"77",X"39",X"83",X"39",X"E5",X"C5",X"F5",X"4F",X"7E",X"B7",X"20",X"1D",X"3A",X"23",X"40",X"CB",
		X"57",X"20",X"16",X"3A",X"0E",X"40",X"B7",X"28",X"10",X"47",X"21",X"39",X"80",X"D5",X"11",X"0F",
		X"00",X"7E",X"B7",X"28",X"08",X"19",X"10",X"F9",X"D1",X"F1",X"C1",X"E1",X"C9",X"D1",X"7A",X"FE",
		X"FE",X"D2",X"42",X"38",X"FE",X"06",X"38",X"2A",X"7B",X"FE",X"F6",X"30",X"1F",X"FE",X"02",X"38",
		X"1B",X"7A",X"CB",X"41",X"28",X"03",X"ED",X"44",X"57",X"7B",X"CB",X"51",X"28",X"03",X"ED",X"44",
		X"5F",X"92",X"FE",X"F6",X"30",X"12",X"FE",X"06",X"30",X"CF",X"18",X"0C",X"79",X"E6",X"03",X"4F",
		X"18",X"06",X"79",X"E6",X"0C",X"4F",X"18",X"00",X"E5",X"06",X"0F",X"AF",X"77",X"23",X"10",X"FC",
		X"CD",X"84",X"1C",X"21",X"A9",X"19",X"09",X"4E",X"21",X"BB",X"38",X"09",X"09",X"09",X"DD",X"70",
		X"08",X"DD",X"70",X"0A",X"7E",X"23",X"F3",X"DD",X"77",X"0C",X"7E",X"DD",X"77",X"0D",X"FB",X"23",
		X"DD",X"36",X"07",X"01",X"46",X"23",X"4E",X"23",X"56",X"DD",X"7E",X"09",X"80",X"47",X"DD",X"7E",
		X"0B",X"81",X"4F",X"E1",X"7A",X"F6",X"03",X"F3",X"77",X"23",X"70",X"23",X"71",X"23",X"70",X"23",
		X"71",X"FB",X"F1",X"C1",X"E1",X"36",X"0A",X"CD",X"CF",X"16",X"DD",X"CB",X"00",X"6E",X"20",X"04",
		X"7E",X"B7",X"20",X"F3",X"3A",X"1F",X"40",X"87",X"87",X"C6",X"05",X"4F",X"3A",X"0F",X"40",X"CB",
		X"3F",X"B9",X"38",X"01",X"79",X"77",X"0E",X"10",X"C3",X"B3",X"37",X"57",X"39",X"00",X"00",X"00",
		X"00",X"57",X"39",X"05",X"00",X"60",X"00",X"57",X"39",X"06",X"01",X"20",X"00",X"57",X"39",X"06",
		X"02",X"A0",X"00",X"57",X"39",X"06",X"0A",X"80",X"00",X"57",X"39",X"00",X"02",X"90",X"00",X"57",
		X"39",X"00",X"01",X"10",X"00",X"57",X"39",X"00",X"00",X"50",X"00",X"57",X"39",X"05",X"00",X"40",
		X"00",X"E8",X"C9",X"EB",X"C9",X"EF",X"C9",X"F4",X"C9",X"FA",X"C9",X"01",X"CA",X"09",X"CA",X"12",
		X"CA",X"1C",X"CA",X"27",X"CA",X"01",X"C0",X"0E",X"C0",X"1B",X"C0",X"28",X"C0",X"35",X"C0",X"42",
		X"C0",X"42",X"C0",X"42",X"C0",X"42",X"C0",X"42",X"C0",X"4F",X"C0",X"5C",X"C0",X"69",X"C0",X"00",
		X"00",X"05",X"39",X"76",X"C0",X"83",X"C0",X"90",X"C0",X"00",X"00",X"23",X"39",X"EB",X"C0",X"F8",
		X"C0",X"05",X"C1",X"00",X"00",X"2D",X"39",X"9D",X"C0",X"AA",X"C0",X"B7",X"C0",X"00",X"00",X"37",
		X"39",X"C4",X"C0",X"D1",X"C0",X"DE",X"C0",X"00",X"00",X"41",X"39",X"12",X"C1",X"36",X"C1",X"5A",
		X"C1",X"82",X"C1",X"00",X"00",X"51",X"39",X"33",X"CA",X"33",X"CA",X"00",X"00",X"57",X"39",X"9F",
		X"CA",X"B1",X"CA",X"9F",X"CA",X"C3",X"CA",X"00",X"00",X"5F",X"39",X"45",X"CA",X"33",X"CA",X"45",
		X"CA",X"57",X"CA",X"00",X"00",X"6B",X"39",X"D5",X"CA",X"E7",X"CA",X"D5",X"CA",X"F9",X"CA",X"00",
		X"00",X"77",X"39",X"69",X"CA",X"7B",X"CA",X"69",X"CA",X"8D",X"CA",X"00",X"00",X"83",X"39",X"A7",
		X"C2",X"A7",X"C2",X"00",X"00",X"8F",X"39",X"DD",X"C2",X"DD",X"C2",X"B9",X"C2",X"B9",X"C2",X"CB",
		X"C2",X"CB",X"C2",X"00",X"00",X"97",X"39",X"13",X"C3",X"13",X"C3",X"EF",X"C2",X"EF",X"C2",X"01",
		X"C3",X"01",X"C3",X"00",X"00",X"A7",X"39",X"37",X"C3",X"25",X"C3",X"4A",X"C3",X"5D",X"C3",X"00",
		X"00",X"B7",X"39",X"70",X"C3",X"70",X"C3",X"00",X"00",X"C3",X"39",X"81",X"C3",X"81",X"C3",X"00",
		X"00",X"CB",X"39",X"92",X"C3",X"92",X"C3",X"00",X"00",X"D3",X"39",X"A3",X"C3",X"A3",X"C3",X"00",
		X"00",X"DB",X"39",X"B4",X"C3",X"B4",X"C3",X"00",X"00",X"E3",X"39",X"C5",X"C3",X"C5",X"C3",X"00",
		X"00",X"EB",X"39",X"D6",X"C3",X"D6",X"C3",X"00",X"00",X"F3",X"39",X"E7",X"C3",X"E7",X"C3",X"00",
		X"00",X"FB",X"39",X"85",X"C1",X"8B",X"C1",X"92",X"C1",X"9A",X"C1",X"A3",X"C1",X"AD",X"C1",X"FA",
		X"C1",X"C4",X"C1",X"D2",X"C1",X"E0",X"C1",X"EE",X"C1",X"E0",X"C1",X"D2",X"C1",X"C4",X"C1",X"00",
		X"00",X"0F",X"3A",X"FA",X"C1",X"07",X"C2",X"15",X"C2",X"23",X"C2",X"31",X"C2",X"23",X"C2",X"15",
		X"C2",X"07",X"C2",X"00",X"00",X"23",X"3A",X"FA",X"C1",X"3D",X"C2",X"4B",X"C2",X"59",X"C2",X"67",
		X"C2",X"59",X"C2",X"4B",X"C2",X"3D",X"C2",X"00",X"00",X"37",X"3A",X"59",X"C2",X"67",X"C2",X"59",
		X"C2",X"4B",X"C2",X"3D",X"C2",X"73",X"C2",X"80",X"C2",X"8D",X"C2",X"9A",X"C2",X"82",X"C1",X"00",
		X"00",X"5D",X"3A",X"A1",X"C8",X"AF",X"C8",X"BD",X"C8",X"CB",X"C8",X"D9",X"C8",X"E7",X"C8",X"F5",
		X"C8",X"07",X"C9",X"A1",X"C8",X"00",X"00",X"71",X"3A",X"6A",X"C9",X"75",X"C9",X"7F",X"C9",X"86",
		X"C9",X"8D",X"C9",X"86",X"C9",X"7F",X"C9",X"75",X"C9",X"00",X"00",X"79",X"3A",X"6A",X"C9",X"6A",
		X"C9",X"00",X"00",X"8D",X"3A",X"94",X"C9",X"9B",X"C9",X"A2",X"C9",X"A9",X"C9",X"B0",X"C9",X"B7",
		X"C9",X"BE",X"C9",X"C5",X"C9",X"CC",X"C9",X"D3",X"C9",X"DA",X"C9",X"E1",X"C9",X"00",X"00",X"95",
		X"3A",X"E1",X"C9",X"DA",X"C9",X"D3",X"C9",X"CC",X"C9",X"C5",X"C9",X"BE",X"C9",X"B7",X"C9",X"B0",
		X"C9",X"A9",X"C9",X"A2",X"C9",X"9B",X"C9",X"94",X"C9",X"00",X"00",X"B1",X"3A",X"33",X"CC",X"4D",
		X"CC",X"67",X"CC",X"81",X"CC",X"00",X"00",X"CD",X"3A",X"AD",X"CC",X"BF",X"CC",X"D1",X"CC",X"9B",
		X"CC",X"D1",X"CC",X"AD",X"CC",X"BF",X"CC",X"9B",X"CC",X"00",X"00",X"D9",X"3A",X"9B",X"CB",X"A5",
		X"CB",X"B3",X"CB",X"C5",X"CB",X"DB",X"CB",X"F5",X"CB",X"13",X"CC",X"00",X"00",X"F9",X"3A",X"91",
		X"CB",X"9B",X"CB",X"A5",X"CB",X"B3",X"CB",X"A5",X"CB",X"9B",X"CB",X"00",X"00",X"FF",X"3A",X"FF",
		X"CC",X"82",X"C1",X"82",X"C1",X"11",X"CD",X"82",X"C1",X"23",X"CD",X"35",X"CD",X"47",X"CD",X"82",
		X"C1",X"00",X"00",X"0F",X"3B",X"82",X"C1",X"59",X"CD",X"6B",X"CD",X"7D",X"CD",X"82",X"C1",X"82",
		X"C1",X"82",X"C1",X"8F",X"CD",X"A1",X"CD",X"B3",X"CD",X"82",X"C1",X"00",X"00",X"25",X"3B",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"97",X"13",X"D7",X"00",
		X"07",X"01",X"0B",X"3C",X"7E",X"C7",X"D7",X"C7",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",
		X"3C",X"7E",X"E3",X"EB",X"E3",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",
		X"F5",X"F1",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F8",X"FA",X"F8",X"7E",
		X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"FC",X"FD",X"FC",X"7E",X"3C",X"DB",X"7E",
		X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",
		X"0B",X"3C",X"7E",X"3F",X"BF",X"3F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",
		X"1F",X"5F",X"1F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",X"8F",
		X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"DB",
		X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"6D",X"FF",X"FE",X"36",
		X"01",X"0B",X"3C",X"7E",X"F1",X"F5",X"F1",X"7E",X"3C",X"B6",X"FF",X"7F",X"6C",X"01",X"0B",X"3C",
		X"7E",X"8F",X"AF",X"8F",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",
		X"8F",X"7E",X"3C",X"B6",X"FF",X"7F",X"6C",X"01",X"0B",X"3C",X"7E",X"8F",X"AF",X"8F",X"7E",X"3C",
		X"6D",X"FF",X"FE",X"36",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"FF",X"1F",X"F8",
		X"E7",X"01",X"0B",X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"1F",X"F8",X"FF",X"07",X"01",X"0B",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"7E",X"3C",X"F8",X"FF",X"1F",X"E0",X"01",X"0B",X"3C",X"7E",X"FF",
		X"C7",X"D7",X"46",X"3C",X"FF",X"1F",X"F8",X"E7",X"01",X"0B",X"3C",X"7E",X"FF",X"C7",X"D7",X"46",
		X"3C",X"F8",X"FF",X"1F",X"E0",X"01",X"0B",X"3C",X"7E",X"FF",X"C7",X"D7",X"46",X"3C",X"1F",X"F8",
		X"FF",X"07",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"07",X"E0",X"0F",X"78",X"13",X"C8",X"0A",X"D0",X"03",X"40",X"33",X"CC",X"09",X"F0",
		X"02",X"48",X"1E",X"78",X"06",X"60",X"02",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"C0",X"06",X"60",X"12",X"48",X"08",X"90",X"10",X"08",X"22",X"44",X"24",X"48",X"0A",X"90",
		X"13",X"60",X"08",X"18",X"14",X"20",X"02",X"40",X"06",X"60",X"02",X"13",X"00",X"00",X"02",X"00",
		X"00",X"20",X"01",X"08",X"10",X"00",X"02",X"40",X"20",X"12",X"08",X"01",X"80",X"20",X"08",X"82",
		X"40",X"02",X"04",X"10",X"21",X"00",X"08",X"04",X"20",X"02",X"04",X"08",X"20",X"20",X"10",X"08",
		X"18",X"0C",X"01",X"01",X"00",X"00",X"82",X"01",X"02",X"18",X"18",X"00",X"82",X"01",X"03",X"10",
		X"38",X"10",X"00",X"82",X"01",X"04",X"10",X"38",X"38",X"10",X"00",X"82",X"01",X"05",X"18",X"3C",
		X"3C",X"3C",X"18",X"00",X"82",X"01",X"06",X"38",X"7C",X"7C",X"7C",X"7C",X"38",X"00",X"82",X"01",
		X"07",X"38",X"7C",X"FE",X"FE",X"FE",X"7C",X"1C",X"00",X"82",X"01",X"08",X"18",X"7E",X"5A",X"FF",
		X"FF",X"7E",X"7E",X"18",X"00",X"81",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",
		X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",
		X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",X"01",X"0A",
		X"18",X"7E",X"7E",X"DB",X"FF",X"BD",X"DB",X"66",X"7E",X"18",X"00",X"82",X"01",X"09",X"00",X"00",
		X"00",X"3C",X"5A",X"FF",X"FF",X"C3",X"7E",X"00",X"81",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",
		X"FF",X"C3",X"7E",X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",
		X"7E",X"7E",X"18",X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",X"7E",X"7E",
		X"18",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"C3",X"7E",X"7E",X"18",X"00",X"81",X"01",
		X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"80",X"80",X"01",X"0A",X"18",
		X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"40",X"80",X"01",X"0A",X"18",X"7E",X"7E",
		X"DB",X"FF",X"FF",X"E7",X"5A",X"7E",X"18",X"01",X"0A",X"18",X"7E",X"7E",X"DB",X"FF",X"FF",X"E7",
		X"5A",X"7E",X"18",X"00",X"82",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"3C",X"5A",X"C3",X"FF",
		X"00",X"82",X"01",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"5A",X"FF",X"00",X"82",X"01",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"FF",X"00",X"82",X"01",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"18",X"01",X"10",X"18",X"18",X"00",X"3C",X"5A",
		X"9A",X"59",X"18",X"18",X"24",X"22",X"41",X"41",X"81",X"81",X"C0",X"01",X"10",X"00",X"18",X"18",
		X"00",X"3C",X"5C",X"5A",X"3A",X"18",X"18",X"14",X"12",X"F2",X"82",X"02",X"03",X"01",X"10",X"18",
		X"18",X"00",X"3C",X"3C",X"3C",X"1A",X"18",X"18",X"0C",X"0A",X"0F",X"78",X"48",X"08",X"0C",X"01",
		X"10",X"18",X"18",X"00",X"3C",X"5A",X"59",X"9A",X"18",X"18",X"24",X"44",X"82",X"82",X"81",X"81",
		X"03",X"01",X"10",X"00",X"18",X"18",X"00",X"3C",X"3A",X"3A",X"DC",X"18",X"18",X"28",X"48",X"4F",
		X"41",X"40",X"80",X"01",X"10",X"18",X"18",X"00",X"3C",X"3C",X"3C",X"58",X"18",X"18",X"30",X"50",
		X"F0",X"1E",X"12",X"10",X"30",X"01",X"10",X"00",X"18",X"18",X"00",X"3C",X"5A",X"5A",X"5A",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"3C",X"01",X"11",X"18",X"24",X"24",X"42",X"81",X"81",X"81",
		X"81",X"81",X"42",X"24",X"24",X"24",X"24",X"24",X"42",X"3C",X"01",X"11",X"18",X"24",X"24",X"7E",
		X"C3",X"A5",X"A5",X"A5",X"E7",X"66",X"24",X"24",X"24",X"24",X"66",X"42",X"3C",X"01",X"11",X"3C",
		X"3C",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"3C",X"3C",X"3C",X"7E",X"7E",X"7E",
		X"01",X"0F",X"18",X"19",X"02",X"1C",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"1C",X"01",X"0F",X"18",X"18",X"00",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"18",X"18",X"1C",X"1A",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"3C",X"3C",X"3A",X"3A",X"3A",X"18",X"18",X"18",
		X"18",X"18",X"18",X"1C",X"01",X"0F",X"18",X"18",X"00",X"3C",X"3C",X"5C",X"9C",X"1C",X"18",X"18",
		X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"18",X"18",X"00",X"F8",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"98",X"58",X"20",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"38",X"01",X"0F",X"18",X"18",X"00",X"1D",X"1B",X"19",X"18",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1C",X"00",X"3E",X"41",X"5D",X"51",X"5D",X"41",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"00",X"10",X"14",X"14",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"14",X"14",X"7F",
		X"14",X"7F",X"14",X"14",X"14",X"14",X"7F",X"54",X"54",X"7F",X"15",X"15",X"7F",X"14",X"20",X"51",
		X"22",X"04",X"08",X"10",X"22",X"45",X"02",X"00",X"18",X"24",X"28",X"10",X"29",X"46",X"46",X"39",
		X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"08",X"10",X"10",X"10",X"10",X"10",
		X"08",X"04",X"10",X"08",X"04",X"04",X"04",X"04",X"04",X"08",X"10",X"00",X"00",X"08",X"2A",X"1C",
		X"1C",X"2A",X"08",X"00",X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"00",X"80",X"00",X"00",
		X"00",X"18",X"18",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"20",
		X"40",X"1C",X"22",X"41",X"41",X"41",X"41",X"41",X"22",X"1C",X"08",X"18",X"08",X"08",X"08",X"08",
		X"08",X"08",X"1C",X"3E",X"41",X"01",X"01",X"3E",X"40",X"40",X"40",X"7F",X"3E",X"41",X"01",X"01",
		X"1E",X"01",X"01",X"41",X"3E",X"02",X"06",X"0A",X"12",X"22",X"7F",X"02",X"02",X"02",X"7F",X"40",
		X"40",X"40",X"7E",X"01",X"01",X"41",X"3E",X"3E",X"41",X"40",X"40",X"7E",X"41",X"41",X"41",X"3E",
		X"7F",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"08",X"3E",X"41",X"41",X"41",X"3E",X"41",X"41",
		X"41",X"3E",X"3E",X"41",X"41",X"41",X"3F",X"01",X"01",X"41",X"3E",X"00",X"00",X"00",X"18",X"18",
		X"00",X"00",X"18",X"18",X"98",X"18",X"00",X"00",X"18",X"18",X"08",X"10",X"00",X"02",X"04",X"08",
		X"10",X"20",X"10",X"08",X"04",X"02",X"00",X"00",X"00",X"3E",X"00",X"3E",X"00",X"00",X"00",X"20",
		X"10",X"08",X"04",X"02",X"04",X"08",X"10",X"20",X"1C",X"22",X"02",X"02",X"04",X"08",X"08",X"00",
		X"08",X"3E",X"41",X"4F",X"49",X"49",X"4F",X"40",X"40",X"3F",X"3E",X"41",X"41",X"41",X"7F",X"41",
		X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"41",X"41",X"41",X"7E",X"3E",X"41",X"40",X"40",
		X"40",X"40",X"40",X"41",X"3E",X"7E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"7E",X"7F",X"40",
		X"40",X"40",X"7C",X"40",X"40",X"40",X"7F",X"7F",X"40",X"40",X"40",X"7C",X"40",X"40",X"40",X"40",
		X"3E",X"41",X"40",X"40",X"47",X"41",X"41",X"41",X"3F",X"41",X"41",X"41",X"41",X"7F",X"41",X"41",
		X"41",X"41",X"1C",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"1C",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"41",X"3E",X"41",X"42",X"44",X"48",X"50",X"68",X"44",X"42",X"41",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"7F",X"41",X"63",X"55",X"49",X"41",X"41",X"41",X"41",X"41",X"41",
		X"61",X"51",X"49",X"45",X"43",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"41",X"41",X"41",X"41",
		X"3E",X"7E",X"41",X"41",X"41",X"7E",X"40",X"40",X"40",X"40",X"3E",X"41",X"41",X"41",X"41",X"41",
		X"45",X"42",X"3D",X"7E",X"41",X"41",X"41",X"7E",X"48",X"44",X"42",X"41",X"3E",X"41",X"40",X"40",
		X"3E",X"01",X"01",X"41",X"3E",X"7F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"41",X"41",
		X"41",X"41",X"41",X"41",X"41",X"41",X"3E",X"41",X"41",X"41",X"22",X"22",X"14",X"14",X"08",X"08",
		X"41",X"41",X"41",X"41",X"41",X"49",X"55",X"63",X"41",X"41",X"41",X"22",X"14",X"08",X"14",X"22",
		X"41",X"41",X"41",X"41",X"22",X"14",X"08",X"08",X"08",X"08",X"08",X"7F",X"01",X"02",X"04",X"08",
		X"10",X"20",X"40",X"7F",X"3C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"3C",X"00",X"00",X"40",
		X"20",X"10",X"08",X"04",X"02",X"01",X"3C",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"3C",X"08",
		X"14",X"22",X"41",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"18",X"18",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"46",X"42",
		X"42",X"46",X"3A",X"40",X"40",X"40",X"5C",X"62",X"42",X"42",X"62",X"5C",X"00",X"00",X"00",X"3C",
		X"42",X"40",X"40",X"42",X"3C",X"02",X"02",X"02",X"3A",X"46",X"42",X"42",X"46",X"3A",X"00",X"00",
		X"00",X"3C",X"42",X"7E",X"40",X"40",X"3C",X"0C",X"12",X"10",X"10",X"38",X"10",X"10",X"10",X"10",
		X"BA",X"46",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",X"40",X"40",X"40",X"7C",X"42",X"42",X"42",
		X"42",X"42",X"00",X"08",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"84",X"04",X"04",X"04",X"04",
		X"04",X"04",X"44",X"38",X"40",X"40",X"40",X"44",X"48",X"50",X"70",X"48",X"44",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"76",X"49",X"49",X"49",X"49",X"49",X"00",
		X"00",X"00",X"7C",X"42",X"42",X"42",X"42",X"42",X"00",X"00",X"00",X"3C",X"42",X"42",X"42",X"42",
		X"3C",X"DC",X"62",X"42",X"42",X"62",X"5C",X"40",X"40",X"40",X"BA",X"46",X"42",X"42",X"46",X"3A",
		X"02",X"02",X"02",X"00",X"00",X"00",X"5C",X"62",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"3C",
		X"42",X"30",X"0C",X"42",X"3C",X"00",X"10",X"10",X"7C",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"42",X"42",X"42",X"42",X"42",X"3C",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"28",X"10",
		X"00",X"00",X"00",X"41",X"41",X"41",X"49",X"49",X"36",X"00",X"00",X"00",X"42",X"24",X"18",X"18",
		X"24",X"42",X"C2",X"42",X"42",X"42",X"46",X"3A",X"02",X"42",X"3C",X"00",X"00",X"00",X"7E",X"04",
		X"08",X"10",X"20",X"7E",X"0C",X"10",X"10",X"10",X"20",X"10",X"10",X"10",X"0C",X"08",X"08",X"08",
		X"00",X"00",X"08",X"08",X"08",X"00",X"18",X"04",X"04",X"04",X"02",X"04",X"04",X"04",X"18",X"08",
		X"00",X"1C",X"2A",X"08",X"08",X"14",X"22",X"00",X"55",X"2A",X"55",X"2A",X"55",X"2A",X"55",X"2A",
		X"55",X"08",X"00",X"1C",X"2A",X"08",X"08",X"14",X"22",X"00",X"02",X"28",X"00",X"0F",X"00",X"3F",
		X"00",X"FF",X"01",X"FF",X"03",X"FF",X"07",X"FF",X"0F",X"FF",X"1F",X"FF",X"1F",X"FF",X"3F",X"FF",
		X"3F",X"FF",X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"7F",X"FF",X"7F",X"FF",X"3F",X"FF",X"3F",X"FF",X"1F",X"FF",X"1F",X"FF",X"0F",X"FF",
		X"07",X"FF",X"03",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"3F",X"00",X"0F",X"02",X"28",X"F0",X"00",
		X"FC",X"00",X"FF",X"00",X"FF",X"80",X"FF",X"C0",X"FF",X"E0",X"FF",X"F0",X"FF",X"F8",X"FF",X"F8",
		X"FF",X"FC",X"FF",X"FC",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FC",X"FF",X"FC",X"FF",X"F8",X"FF",X"F8",
		X"FF",X"F0",X"FF",X"E0",X"FF",X"C0",X"FF",X"80",X"FF",X"00",X"FC",X"00",X"F0",X"00",X"01",X"0C",
		X"20",X"30",X"18",X"0C",X"06",X"03",X"70",X"F8",X"C8",X"C8",X"F8",X"70",X"01",X"0C",X"04",X"0C",
		X"18",X"30",X"60",X"C0",X"0E",X"1F",X"13",X"13",X"1F",X"0E",X"02",X"07",X"00",X"03",X"00",X"1F",
		X"00",X"3C",X"00",X"60",X"00",X"C0",X"01",X"80",X"01",X"00",X"02",X"07",X"C0",X"00",X"F8",X"00",
		X"3C",X"00",X"06",X"00",X"03",X"00",X"01",X"80",X"00",X"80",X"02",X"07",X"01",X"00",X"01",X"80",
		X"00",X"C0",X"00",X"60",X"00",X"3C",X"00",X"1F",X"00",X"03",X"02",X"07",X"00",X"80",X"01",X"80",
		X"03",X"00",X"06",X"00",X"3C",X"00",X"F8",X"00",X"C0",X"00",X"02",X"02",X"FF",X"FF",X"FF",X"FF",
		X"02",X"08",X"00",X"30",X"00",X"78",X"00",X"CC",X"01",X"86",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"F0",X"02",X"08",X"0C",X"00",X"1E",X"00",X"33",X"00",X"61",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"C0",X"01",X"0B",X"F8",X"F8",X"98",X"68",X"68",X"08",X"68",X"68",X"68",X"F8",
		X"F8",X"02",X"06",X"00",X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",X"80",X"FF",X"00",X"02",
		X"06",X"60",X"00",X"FF",X"00",X"05",X"80",X"02",X"80",X"05",X"80",X"FF",X"00",X"02",X"06",X"06",
		X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",
		X"60",X"05",X"B0",X"02",X"80",X"05",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",X"00",X"02",
		X"B0",X"07",X"98",X"02",X"80",X"FF",X"00",X"02",X"06",X"00",X"00",X"FF",X"00",X"05",X"80",X"02",
		X"80",X"05",X"98",X"FF",X"0C",X"02",X"08",X"00",X"00",X"FF",X"00",X"02",X"80",X"07",X"80",X"02",
		X"80",X"FF",X"00",X"00",X"0C",X"00",X"06",X"02",X"06",X"00",X"00",X"FF",X"00",X"05",X"80",X"02",
		X"80",X"05",X"80",X"FF",X"00",X"01",X"17",X"30",X"78",X"FC",X"FC",X"FC",X"8C",X"B4",X"B4",X"8C",
		X"B4",X"B4",X"8C",X"FC",X"FC",X"78",X"30",X"30",X"78",X"30",X"34",X"3F",X"1F",X"04",X"02",X"1D",
		X"3F",X"FC",X"1F",X"F8",X"0F",X"F0",X"07",X"E0",X"FF",X"FF",X"80",X"01",X"93",X"29",X"AA",X"B9",
		X"BB",X"39",X"AA",X"A9",X"AA",X"A9",X"80",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"09",X"00",X"00",X"00",X"00",
		X"C0",X"40",X"40",X"40",X"78",X"01",X"08",X"00",X"00",X"00",X"00",X"C0",X"40",X"40",X"78",X"01",
		X"05",X"00",X"00",X"00",X"00",X"F8",X"01",X"05",X"00",X"78",X"40",X"40",X"C0",X"01",X"05",X"78",
		X"40",X"40",X"40",X"C0",X"01",X"05",X"04",X"04",X"FC",X"04",X"04",X"01",X"05",X"02",X"0C",X"74",
		X"84",X"08",X"01",X"05",X"02",X"1A",X"24",X"C8",X"08",X"01",X"05",X"09",X"12",X"24",X"48",X"90",
		X"01",X"05",X"10",X"13",X"24",X"58",X"40",X"01",X"05",X"10",X"21",X"2E",X"30",X"40",X"01",X"05",
		X"20",X"20",X"3F",X"20",X"20",X"01",X"05",X"40",X"30",X"2E",X"21",X"10",X"01",X"05",X"40",X"58",
		X"24",X"13",X"10",X"01",X"05",X"90",X"48",X"24",X"12",X"09",X"01",X"05",X"08",X"C8",X"24",X"1A",
		X"02",X"01",X"05",X"08",X"84",X"74",X"0C",X"02",X"01",X"01",X"5A",X"01",X"02",X"FF",X"5A",X"01",
		X"03",X"7E",X"FF",X"5A",X"01",X"04",X"DB",X"7E",X"FF",X"5A",X"01",X"05",X"3C",X"DB",X"7E",X"FF",
		X"5A",X"01",X"06",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"07",X"FF",X"7E",X"3C",X"DB",X"7E",
		X"FF",X"5A",X"01",X"08",X"EF",X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"09",X"FF",X"EF",
		X"FF",X"7E",X"3C",X"DB",X"7E",X"FF",X"5A",X"01",X"0A",X"7E",X"FF",X"EF",X"FF",X"7E",X"3C",X"DB",
		X"7E",X"FF",X"5A",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",
		X"10",X"38",X"28",X"28",X"6C",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",X"92",X"BA",
		X"90",X"38",X"10",X"38",X"28",X"68",X"0C",X"01",X"10",X"38",X"54",X"7C",X"28",X"38",X"10",X"7C",
		X"92",X"BA",X"12",X"38",X"10",X"38",X"28",X"2C",X"60",X"01",X"10",X"38",X"7C",X"7C",X"38",X"38",
		X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"38",X"28",X"28",X"6C",X"01",X"10",X"38",X"7C",X"7C",
		X"38",X"38",X"10",X"7C",X"92",X"BA",X"12",X"38",X"10",X"38",X"28",X"2C",X"60",X"01",X"10",X"38",
		X"7C",X"7C",X"38",X"38",X"10",X"7C",X"92",X"BA",X"90",X"38",X"10",X"38",X"28",X"68",X"0C",X"01",
		X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"38",X"28",X"28",
		X"3C",X"01",X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"7C",
		X"44",X"44",X"66",X"01",X"10",X"38",X"74",X"7C",X"30",X"38",X"10",X"7C",X"92",X"BA",X"92",X"38",
		X"10",X"10",X"10",X"10",X"18",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",X"10",X"7C",X"92",X"BA",
		X"92",X"38",X"10",X"38",X"28",X"28",X"78",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",X"10",X"7C",
		X"92",X"BA",X"92",X"38",X"10",X"7C",X"44",X"44",X"CC",X"01",X"10",X"38",X"5C",X"7C",X"18",X"38",
		X"10",X"7C",X"92",X"BA",X"92",X"38",X"10",X"10",X"10",X"10",X"30",X"02",X"1E",X"80",X"00",X"80",
		X"00",X"80",X"00",X"80",X"07",X"80",X"08",X"80",X"10",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
		X"20",X"40",X"40",X"40",X"40",X"20",X"80",X"1F",X"00",X"02",X"1E",X"00",X"01",X"00",X"01",X"00",
		X"01",X"E0",X"01",X"10",X"01",X"08",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",
		X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",
		X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"04",X"01",X"02",
		X"02",X"02",X"02",X"01",X"04",X"00",X"F8",X"01",X"08",X"3C",X"00",X"FF",X"FF",X"FF",X"7E",X"7E",
		X"3C",X"02",X"04",X"0F",X"FF",X"08",X"01",X"08",X"01",X"0F",X"FF",X"02",X"04",X"0F",X"FF",X"08",
		X"01",X"09",X"F9",X"0F",X"FF",X"02",X"06",X"0F",X"FF",X"08",X"01",X"0B",X"FD",X"0F",X"FF",X"01",
		X"F8",X"00",X"F0",X"02",X"08",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"03",X"FC",X"03",
		X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0A",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",
		X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0C",X"0F",X"FF",X"08",
		X"01",X"0F",X"BF",X"0F",X"BF",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",
		X"FC",X"01",X"F8",X"00",X"F0",X"02",X"0E",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",
		X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",
		X"F8",X"00",X"F0",X"02",X"0F",X"0F",X"FF",X"08",X"01",X"0F",X"BF",X"0F",X"BF",X"07",X"BE",X"07",
		X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"07",X"BE",X"03",X"FC",X"03",X"FC",X"01",
		X"F8",X"00",X"F0",X"02",X"0C",X"1E",X"00",X"33",X"00",X"73",X"80",X"73",X"80",X"F3",X"C0",X"FF",
		X"C0",X"FF",X"C0",X"F3",X"C0",X"73",X"80",X"73",X"80",X"33",X"00",X"1E",X"00",X"02",X"0C",X"1E",
		X"00",X"3F",X"00",X"4F",X"80",X"67",X"80",X"E7",X"C0",X"FF",X"C0",X"FF",X"C0",X"F9",X"C0",X"79",
		X"80",X"7C",X"80",X"3F",X"00",X"1E",X"00",X"02",X"0C",X"1E",X"00",X"3F",X"00",X"7F",X"80",X"7F",
		X"80",X"FF",X"C0",X"8C",X"40",X"8C",X"40",X"FF",X"C0",X"7F",X"80",X"7F",X"80",X"3F",X"00",X"1E",
		X"00",X"02",X"0C",X"1E",X"00",X"3F",X"00",X"7C",X"80",X"79",X"80",X"F9",X"C0",X"FF",X"C0",X"FF",
		X"C0",X"E7",X"C0",X"67",X"80",X"4F",X"80",X"3F",X"00",X"1E",X"00",X"02",X"08",X"FF",X"F0",X"CF",
		X"30",X"B6",X"D0",X"BE",X"D0",X"A6",X"D0",X"B6",X"D0",X"C7",X"30",X"FF",X"F0",X"02",X"08",X"FF",
		X"F0",X"CE",X"30",X"B7",X"70",X"BF",X"70",X"A7",X"70",X"B7",X"70",X"C6",X"30",X"FF",X"F0",X"02",
		X"08",X"FF",X"F0",X"BB",X"B0",X"D7",X"30",X"EF",X"B0",X"EF",X"B0",X"D7",X"B0",X"BB",X"10",X"FF",
		X"F0",X"02",X"08",X"FF",X"F0",X"BA",X"10",X"D6",X"F0",X"EE",X"30",X"EF",X"D0",X"EF",X"D0",X"EE",
		X"30",X"FF",X"F0",X"01",X"10",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"18",X"18",X"3C",
		X"18",X"18",X"3C",X"18",X"18",X"01",X"08",X"3C",X"18",X"18",X"3C",X"18",X"18",X"3C",X"18",X"02",
		X"08",X"0E",X"00",X"01",X"C0",X"00",X"30",X"00",X"20",X"00",X"40",X"00",X"30",X"00",X"0C",X"00",
		X"03",X"02",X"08",X"0E",X"00",X"01",X"C0",X"00",X"30",X"00",X"70",X"00",X"C0",X"00",X"30",X"00",
		X"0C",X"00",X"03",X"02",X"08",X"00",X"00",X"0F",X"80",X"00",X"60",X"00",X"80",X"01",X"80",X"00",
		X"60",X"00",X"18",X"00",X"07",X"02",X"08",X"00",X"00",X"00",X"00",X"0E",X"00",X"01",X"C0",X"00",
		X"60",X"00",X"E0",X"00",X"1C",X"00",X"07",X"02",X"08",X"00",X"00",X"0C",X"00",X"03",X"80",X"00",
		X"70",X"00",X"20",X"00",X"40",X"00",X"38",X"00",X"07",X"02",X"08",X"00",X"00",X"00",X"01",X"00",
		X"C6",X"00",X"A8",X"01",X"30",X"02",X"00",X"04",X"00",X"08",X"00",X"02",X"08",X"00",X"01",X"00",
		X"02",X"00",X"64",X"00",X"98",X"01",X"00",X"02",X"00",X"04",X"00",X"08",X"00",X"02",X"08",X"00",
		X"00",X"00",X"03",X"00",X"0C",X"00",X"10",X"00",X"E0",X"03",X"00",X"04",X"00",X"08",X"00",X"02",
		X"08",X"00",X"03",X"00",X"0C",X"00",X"30",X"00",X"80",X"00",X"30",X"01",X"C0",X"0E",X"00",X"00",
		X"00",X"02",X"08",X"00",X"03",X"00",X"0E",X"00",X"18",X"00",X"D0",X"01",X"B0",X"02",X"00",X"04",
		X"00",X"08",X"00",X"02",X"08",X"00",X"00",X"00",X"07",X"00",X"8C",X"00",X"C8",X"01",X"B0",X"02",
		X"10",X"04",X"00",X"08",X"00",X"02",X"02",X"FF",X"F8",X"FF",X"F8",X"02",X"02",X"FF",X"F0",X"FF",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
