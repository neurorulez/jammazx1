-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "3604059C9964FAD6B8D2579D8A7FFABB731D296D2C9AD4E6BB9EAB93270C72A1";
    attribute INIT_01 of inst : label is "356C9D5AD4BE693F9E44FE1650DFF1453689B63AD8C898644C3B2B24D116A56D";
    attribute INIT_02 of inst : label is "2A62797EB49340AC35D98100027B810C67DC16CFB0C93473D39F4D9826212481";
    attribute INIT_03 of inst : label is "44070EA18BBB0B30216CAB3A27DB3C9ED5599718E621C6208C8E6990650A508D";
    attribute INIT_04 of inst : label is "09B8750C644F206A77EAA679A56797EB413745614D4F6E9F556B831D111721C7";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF7ECB0254DEA666796AD4CF27B6A7184CCB81D8E10ABC0E384";
    attribute INIT_06 of inst : label is "CC2876AC742F3BE29FFF78E98A4FF3D8F1CA7E3C9AD4E6BB773A51941042E30D";
    attribute INIT_07 of inst : label is "190D2B45D7D77AF349371569B469BFEFEA8CBEA765133E74819CA32C0C12720C";
    attribute INIT_08 of inst : label is "FEFB53ABF9F776345D7DFF922234B878CFF648A2E654695F32C8442C94063FFB";
    attribute INIT_09 of inst : label is "02088808820000000000000AAAA7DD813E04EE11B70E5C21DD6C4A23DD72DD7D";
    attribute INIT_0A of inst : label is "0031981453486210000808020202088A88020082088A82088088020880000882";
    attribute INIT_0B of inst : label is "DB64594000000026A6800000002E2E35F65D4D378A760E9AAAF5A7AED20B2800";
    attribute INIT_0C of inst : label is "F36DCEF20F571FB8EFFD3BFFF623977A8A80A8082D04EE3B85B11A924AEFFF7F";
    attribute INIT_0D of inst : label is "230B18B26FDEF8EE4DA4CFDC86DEF6C4EE4DAE677FF985001443BBBF86B7D951";
    attribute INIT_0E of inst : label is "FF00EFA00F6A69976BF17D4AD824CC000000AEB776C000001800001ADC08E622";
    attribute INIT_0F of inst : label is "00A44C3023D8D936F037CC58B9DB99B733B98FD9E8FB3C97EEBF19BCE9ACE73C";
    attribute INIT_10 of inst : label is "BDF881498676CF4D9668B9B03DE74CC8E7F1CDC9FDBD7F6F7D7DCD8275F5FE62";
    attribute INIT_11 of inst : label is "3EC4875080B0419300040EA6A869B76774910410C2040042083002AB675C1334";
    attribute INIT_12 of inst : label is "6FF926494FF5269E77ECEF23306022BF02536629630A2FCA527380FEF67FC7FF";
    attribute INIT_13 of inst : label is "88661B130D8986C4C36269B130D8B8644C222EB3B21DDDDDDDD5924EC83B7F4F";
    attribute INIT_14 of inst : label is "01369D925E49F3C964C2E5DE7BFB000008BB77FE5DBCBF3279EDCB0A7CCF3D22";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFE806CEB3C8251A88CFF3CE7FDDBFF2ECBF3275CAE49AC012";
    attribute INIT_16 of inst : label is "75750E96C3FD754A35291AFCD33AE7AB36B747EECD747CF729F3F5057036C31D";
    attribute INIT_17 of inst : label is "0004404004004000444004000400AAAA80AAFFFFED0B03ECB88E40F7914FFFAE";
    attribute INIT_18 of inst : label is "F033C3330CC0F03C0C00000000000A8000000000000000000000440440040000";
    attribute INIT_19 of inst : label is "444A25128888C444688891188D1111A22244447BBBB8002AAAAAA0000C30FC30";
    attribute INIT_1A of inst : label is "911EEEE4A231188D1188D11A251288D111111223446894462344A2311A234444";
    attribute INIT_1B of inst : label is "111111111111156A88C46231188C47BBAAD5AD5AD7BBA2344A2446894488C468";
    attribute INIT_1C of inst : label is "A855AAC807B3D45EA00BC050EFA0FFFFFE888888888888888888888D11111111";
    attribute INIT_1D of inst : label is "3555555555BCEAF48E429C1FD567AD4A5295295EB52B52B52B52B57918801FFC";
    attribute INIT_1E of inst : label is "03FD0EC1D52C237B6D6A56A56A56A56AA356AE24FFAADFABFCAFFAA109C6B220";
    attribute INIT_1F of inst : label is "D9FD5495FD7FD52A8D9EE524924B65ADDFD54D7F54AFFEFFAAACA1B9A12DBAF0";
    attribute INIT_20 of inst : label is "D395B4E57FFFFFFFFFFFFFFFBFF9999BB2FAF7EB7FFFFFFFD7B7FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "4B6DB24924A492492DB2DED24B6D96DB6DB2492DB6DB64B65B6DB6D94DDB4E56";
    attribute INIT_22 of inst : label is "B972A55B972A55B976E5DB972A55B976E5DB972A55B976E5D6DB6D9249492492";
    attribute INIT_23 of inst : label is "2B75CA674D9CB24B2C924965B2C965B65B24965B2C924965B2C965B65B64B65C";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFEC76246FFB6592CF696DB65A9592DD6D6D6D6D6D6CB60DD28460";
    attribute INIT_25 of inst : label is "020225AF61A9FF32BE9CD09E4D3F59DBF594DA65B4D948ECB47D25FE4C27252D";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF98842A904A42A904A457A915CA457A915CA10202";
    attribute INIT_27 of inst : label is "E73F8D8621FE6B1B3F5DB75AC29639A58EEEDBA9F0D236C1636B813A261B920D";
    attribute INIT_28 of inst : label is "0CC37BBFFE46EFF3BD9F359DF97C4DC30F04C28268A77DA7671C3AD57DE716F1";
    attribute INIT_29 of inst : label is "319400A40E7600C41600C43300620100221A00482C51D03F8A0E89421120771E";
    attribute INIT_2A of inst : label is "801008318000208E0000200000008D2020000A8836510D3400ABC04444ECEAE7";
    attribute INIT_2B of inst : label is "8018801200AAB960AA76C150ED82A9DB3B80808118060208E002020060080823";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF937DA4B4";
    attribute INIT_2D of inst : label is "92C9B583C4860E26BCF259CF9CCF24FE38EF137D3F3D9A24D5133EA39938F509";
    attribute INIT_2E of inst : label is "E98F9FBCF9CFFBBFF2D9A61303FFFE7ECD29BA94431A74DBB1CE4DDF3498884D";
    attribute INIT_2F of inst : label is "FFFFEDA6DCD79A79B9CF39D7F5DE78E9A71D269AA764FF12C40927DAAABAAEA4";
    attribute INIT_30 of inst : label is "D395B4E57FFFFFFFFFFFFFFFBFF9999BB2FAF7EB7FFFFFFFD7B7FFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "4B6DB24924A492492DB2DED24B6D96DB6DB2492DB6DB64B65B6DB6D94DDB4E56";
    attribute INIT_32 of inst : label is "B972A55B972A55B976E5DB972A55B976E5DB972A55B976E5D6DB6D9249492492";
    attribute INIT_33 of inst : label is "2B75CA674D9CB24B2C924965B2C965B65B24965B2C924965B2C965B65B64B65C";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFEC76246FFB6592CF696DB65A9592DD6D6D6D6D6D6CB60DD28460";
    attribute INIT_35 of inst : label is "020225AF61A9FF32BE9CD09E4D3F59DBF594DA65B4D948ECB47D25FE4C27252D";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF98842A904A42A904A457A915CA457A915CA10202";
    attribute INIT_37 of inst : label is "E73F8D8621FE6B1B3F5DB75AC29639A58EEEDBA9F0D236C1636B813A261B920D";
    attribute INIT_38 of inst : label is "0CC37BBFFE46EFF3BD9F359DF97C4DC30F04C28268A77DA7671C3AD57DE716F1";
    attribute INIT_39 of inst : label is "319400A40E7600C41600C43300620100221A00482C51D03F8A0E89421120771E";
    attribute INIT_3A of inst : label is "801008318000208E0000200000008D2020000A8836510D3400ABC04444ECEAE7";
    attribute INIT_3B of inst : label is "8018801200AAB960AA76C150ED82A9DB3B80808118060208E002020060080823";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF937DA4B4";
    attribute INIT_3D of inst : label is "92C9B583C4860E26BCF259CF9CCF24FE38EF137D3F3D9A24D5133EA39938F509";
    attribute INIT_3E of inst : label is "E98F9FBCF9CFFBBFF2D9A61303FFFE7ECD29BA94431A74DBB1CE4DDF3498884D";
    attribute INIT_3F of inst : label is "FFFFEDA6DCD79A79B9CF39D7F5DE78E9A71D269AA764FF12C40927DAAABAAEA4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1EC14284EBC034CA486CD8001038804121A440C81919BF165045E468D16716DC";
    attribute INIT_01 of inst : label is "C3C166A70B087783413D44CBE2E45CBE3AFA4EA13ABFA34FD1A6DC432E21D092";
    attribute INIT_02 of inst : label is "C56422CBE7858003D24632FFFD9076F0B8A1A0208296C90820413251D543483E";
    attribute INIT_03 of inst : label is "9220739558E051444AA65C5450461040299547EAB3D57A2F55F7FEB5F265E5D4";
    attribute INIT_04 of inst : label is "DE039CAAA88412BF5C94D42098822CBE78593266A9A05909FFC2D4524C846E54";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF8154EDAA90454B42A69A8410055438AB5E8DA290B42572A62";
    attribute INIT_06 of inst : label is "C6969112C6D040C40F11840A128AECFD141020A019BD06544C97EA9889B47954";
    attribute INIT_07 of inst : label is "6A3EC68C6A0E4DB7B744DEDD4B6645905FD7471FEFD04A915A72D85BB62DC310";
    attribute INIT_08 of inst : label is "100CBAD40E280268C6B060C3F57272A9680080140B88A220A75A9DD5B9EB8003";
    attribute INIT_09 of inst : label is "080A0A0A028AAAAAAAAAAAA0000140F67DDB88990A942A5A8684B17754AC8684";
    attribute INIT_0A of inst : label is "105C199920332DE0080A000808080A00000802080A08880A0A00080A08080A08";
    attribute INIT_0B of inst : label is "C2AF670000000037F3800000003773182AF7CCAD549AD303CD1240926C056334";
    attribute INIT_0C of inst : label is "02AE9557D4D19DE9830760C0584548A93B1693E6B12D54554E5FAAF5BA3B078F";
    attribute INIT_0D of inst : label is "032289D700025180365286003B2266E700364F2C1834327898B55557FB60909A";
    attribute INIT_0E of inst : label is "FF0005063197440324AAABB1A25E840000015361D1BBBFFFF7FFFFED83B72802";
    attribute INIT_0F of inst : label is "367AAFAF55460A0AE2959148B29B250542AAA2327A464091179012A03645481D";
    attribute INIT_10 of inst : label is "827993B27C1691B1A5640205C618B6EB00342009440151010546149090054C7D";
    attribute INIT_11 of inst : label is "BEC9ADA4229B32B762B32487EE6E182188E8041002001000040082002A218D1B";
    attribute INIT_12 of inst : label is "7BB2128483E60304FDF83D7DE9D35F8CED88ABB7254F0205C004A9FE10AAC955";
    attribute INIT_13 of inst : label is "62CC41E620F31079883C4C1E220F3B879CC3C463E375F5F5F5E637029E63DBCC";
    attribute INIT_14 of inst : label is "A2C90A07E08604373A5642000950A008220C51FED5AD0000808A0B5745EF3FFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFCC0151548C5D990A2084012A608FF62D0040025C43710A0C";
    attribute INIT_16 of inst : label is "C5B2AB5558901FB7DDD2B401554C19704B2DF90216DF9110400C92F7C35B79C4";
    attribute INIT_17 of inst : label is "1115515115115111555115111515FFFFD5BBFFFFA298BC15CED56D00220788A2";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFF41044401111111111111111111111551551151111";
    attribute INIT_19 of inst : label is "AAA82D428022D4012228105A841154A2A85504554117EAD406F11FFFFFFFFFFF";
    attribute INIT_1A of inst : label is "B41AFAFAA0B50A0C5082C14A8452A0C16BBBFE83052831420B14A0B14A8305BB";
    attribute INIT_1B of inst : label is "545454545454556A8A41629058A417EBE2448D18D3BBE0B05A8416290582D420";
    attribute INIT_1C of inst : label is "C09866108282101B850ABFFB4005FFFFFE080808080808080808080C54545454";
    attribute INIT_1D of inst : label is "A4CCCCCC6681E60DC541B4C499A49B26C9B364C60366C06C9909931ACC0AA551";
    attribute INIT_1E of inst : label is "07370498F5188C292C06CD80D9321326773198AEBBBA7BBAF6EBBA633880F3C4";
    attribute INIT_1F of inst : label is "8222206220AA2200082318010080401862220688224001005404238BD073C310";
    attribute INIT_20 of inst : label is "428490A138B6EEEDBBBB6EEEFFFE1E1A30FAFFA6FFFFFFFFB16EDFFFFFFFFAFF";
    attribute INIT_21 of inst : label is "B4926DB493926DB6DA693DE9269B6DA6DB6D249B4D36DA6D369A6DF8DC090A12";
    attribute INIT_22 of inst : label is "56AC10356AC10356AD5AB56AC10356AD5AB56AC10356AD5ABDA69B692724DB6D";
    attribute INIT_23 of inst : label is "79600062614B6D34DA6934DB69A4DB6DB6D36934DA6934DB69A4DB6DB6936903";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFC8240D2406DB69A494D34DB31B024A9292929292919CC7F080C2";
    attribute INIT_25 of inst : label is "CAE845183204A017C361070032408260E4B3892CD0CB3C058A056A15D8AA6FE0";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFAC440090064189026424090906424890926ACAE8";
    attribute INIT_27 of inst : label is "75202C0045A8C98A0191364447E118F846E342FAF1807B05076F63130039809C";
    attribute INIT_28 of inst : label is "6D1380DFFE973FF4C06F47E6419CC05B5522379039D18115E5C8B27201004A80";
    attribute INIT_29 of inst : label is "D0A699301624E0981EE1D812F05C12704C19C030089BCD10916041C96A0E0485";
    attribute INIT_2A of inst : label is "38085C03A8465088E0007000A0014BB3AEDFE18FF090FA2E3F0842505068E222";
    attribute INIT_2B of inst : label is "CC1410042018DA201AB04035608062C13AC085C13A8065088E001704EA019402";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0832802E";
    attribute INIT_2D of inst : label is "EF2E99B3D879B9D96EFCA1F320061900F5DCE5B6DCBE0DDB26604360254E2FE4";
    attribute INIT_2E of inst : label is "AAE0E0800025448FF75A940DA6000180164641208A299944DD91B2E4386D67B2";
    attribute INIT_2F of inst : label is "FFFFCDD34AEA4C0DC411405C00401300A9C46CF9F58305A16A52DC59AAB6A1EA";
    attribute INIT_30 of inst : label is "428490A138B6EEEDBBBB6EEEFFFE1E1A30FAFFA6FFFFFFFFB16EDFFFFFFFFAFF";
    attribute INIT_31 of inst : label is "B4926DB493926DB6DA693DE9269B6DA6DB6D249B4D36DA6D369A6DF8DC090A12";
    attribute INIT_32 of inst : label is "56AC10356AC10356AD5AB56AC10356AD5AB56AC10356AD5ABDA69B692724DB6D";
    attribute INIT_33 of inst : label is "79600062614B6D34DA6934DB69A4DB6DB6D36934DA6934DB69A4DB6DB6936903";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFC8240D2406DB69A494D34DB31B024A9292929292919CC7F080C2";
    attribute INIT_35 of inst : label is "CAE845183204A017C361070032408260E4B3892CD0CB3C058A056A15D8AA6FE0";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFAC440090064189026424090906424890926ACAE8";
    attribute INIT_37 of inst : label is "75202C0045A8C98A0191364447E118F846E342FAF1807B05076F63130039809C";
    attribute INIT_38 of inst : label is "6D1380DFFE973FF4C06F47E6419CC05B5522379039D18115E5C8B27201004A80";
    attribute INIT_39 of inst : label is "D0A699301624E0981EE1D812F05C12704C19C030089BCD10916041C96A0E0485";
    attribute INIT_3A of inst : label is "38085C03A8465088E0007000A0014BB3AEDFE18FF090FA2E3F0842505068E222";
    attribute INIT_3B of inst : label is "CC1410042018DA201AB04035608062C13AC085C13A8065088E001704EA019402";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0832802E";
    attribute INIT_3D of inst : label is "EF2E99B3D879B9D96EFCA1F320061900F5DCE5B6DCBE0DDB26604360254E2FE4";
    attribute INIT_3E of inst : label is "AAE0E0800025448FF75A940DA6000180164641208A299944DD91B2E4386D67B2";
    attribute INIT_3F of inst : label is "FFFFCDD34AEA4C0DC411405C00401300A9C46CF9F58305A16A52DC59AAB6A1EA";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "1AC321886BE00E83F1FE84851A83355435B86A014150AD742A8D7F3163455444";
    attribute INIT_01 of inst : label is "729FB3B3CF6F7A6F3615F68FF0F778FF3D2B3890E252B9315C916E6C2B3F6CCD";
    attribute INIT_02 of inst : label is "EA49D92D573EC4001FBAA233004FE600FBECF7DBEA7B6C46D1371B4972727DB8";
    attribute INIT_03 of inst : label is "C2325FE4D7725156EB8EBF766DC1EC362FDCD5B27F64EC81DADA23B4274C3BD9";
    attribute INIT_04 of inst : label is "9312FFA68CFB03D5EE17F3D83D5D92D573EC754AE7C964F6AABB574B0CCA6BD2";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF015DCC2E5C672F7AC63E7B0D837322E5DF836250E6555C943";
    attribute INIT_06 of inst : label is "9A6845AC64694A06A066CCEB3ADFBDDDE4528FA550AF6415557505AD8C84F1C4";
    attribute INIT_07 of inst : label is "03C36AF2AFD31250DE868937A143D369757A201822C944C7CBD6295D3B375199";
    attribute INIT_08 of inst : label is "1FBFEF5C6EFB35AF2AE7CFFB77A09F99A2B2006ABDCECF5583DBD13DAD2D17FA";
    attribute INIT_09 of inst : label is "00041404490555555555555555213822AE88CC227939E6EA7AC0D000889B7AC0";
    attribute INIT_0A of inst : label is "545A44CB229A8420000405014151044551004811044A50040010000400000450";
    attribute INIT_0B of inst : label is "33AE708000000011110000000019190DBAFAA879D7C85D73EF8DA26E36055669";
    attribute INIT_0C of inst : label is "7BD2532893CAD7FE3E7E8F9EE6F48B9383A43864B959324CDE23B468A95E7DF0";
    attribute INIT_0D of inst : label is "0120C3FD9F12133F1FE2A07E6FF224213F1FF3D1F3E7A70D9D34CCCFF89F3DCF";
    attribute INIT_0E of inst : label is "FF00012A87FDECC4DB3ACEDAB6C284000001509EEF115FFFEFFFFFE27D118800";
    attribute INIT_0F of inst : label is "5460A0E344D44B0CDA275C100BD2B097693BABABD0757085DD9D0BA55B65AC01";
    attribute INIT_10 of inst : label is "78D387A3F4B4957D2141031DD55C9622021FA885F5107C457125D812D481FC05";
    attribute INIT_11 of inst : label is "3817ADA423BF231D4BE335B54E2E16257CEA040082040002082080007AA09CBA";
    attribute INIT_12 of inst : label is "7EF802444416108CDFBC557941B303754403AF30254C1D4C5004ADD5DED56EAA";
    attribute INIT_13 of inst : label is "F721AE00D7006B8035C092E04D700EB8065C01AC05D20200AA7827169C1BFF83";
    attribute INIT_14 of inst : label is "B2668F87BF9862C7CBB4E71218ADD5555DED8F54F139EF1C206A1275E5C71F6E";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFCF615A570E41D0CE9F9242156C7AA709EF1C29760C73CB31";
    attribute INIT_16 of inst : label is "108A33EF585FEADEC5FFD6CDD67AA35154D2A3D2512A3D514A75F022F606F1D4";
    attribute INIT_17 of inst : label is "0000000000000000000000000001AEBAD5AFFFFF9C171FD5C30E4694A350338E";
    attribute INIT_18 of inst : label is "F3FFFFFFFFFFFFFFFFFFFFF54050511040000000000000000000000000000000";
    attribute INIT_19 of inst : label is "05080402000040002000100804000080004000015414051550550CC0CCFFFF3F";
    attribute INIT_1A of inst : label is "1005005580100804008040080402004014141601002010020100801008010014";
    attribute INIT_1B of inst : label is "0000000000000AD1804020100804015420408408410520100804020100804020";
    attribute INIT_1C of inst : label is "E2E1E04A72A42BF0550EFEAAAFBBFFFFFE000000000000000000000400000000";
    attribute INIT_1D of inst : label is "8C3C03C180BCB496954214D8E02480013FB0003E009FC003F9006F618C23130C";
    attribute INIT_1E of inst : label is "443604C8F015A7292C013F8007F200DEE20F82875005F0055E1500F69C8266AE";
    attribute INIT_1F of inst : label is "B0A00A002A0A014ABB0A009A4936D27B4A00240A80155000000F7948CC713215";
    attribute INIT_20 of inst : label is "46AC91AB7EB6EEEDBBBB6EEFFFEAB54860BAF7A03FEFFEA68FFCDFFFFFF6FEFF";
    attribute INIT_21 of inst : label is "400000025C4B402028001484B80904800010924900126124920024828D891AB2";
    attribute INIT_22 of inst : label is "00010A100010A1000400100010A1000400100010A100040016808044B8968040";
    attribute INIT_23 of inst : label is "11540A32400AA480000402002482002002480000000402002482002002482480";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFCC2618C52249241D2000049C6149080000000000061C47A15A40";
    attribute INIT_25 of inst : label is "8AEE248ECC645555ADBCA506C36ECADDF1E50979521E506F2A3DC6CF89C77B44";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF9A7228C823221C847219848661219148645CDABE";
    attribute INIT_27 of inst : label is "A427AAC0465E428A0B5791126094102504D6EFD090D03667230E41290212008C";
    attribute INIT_28 of inst : label is "C9D15F5554BA9AA6AFAAE1358C3444B25D0F2787B8AB47C3231B88D005A376A0";
    attribute INIT_29 of inst : label is "A1C80A40142200400F01E00A01400F80F002004056774C28302041C0090E0009";
    attribute INIT_2A of inst : label is "80118824804D00120000200000000738014016047301869C10D3465500768604";
    attribute INIT_2B of inst : label is "E050C8199160510160A202C144058288054098804804D0092002620120034024";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5376A01C";
    attribute INIT_2D of inst : label is "79EF3D0A81A3356DF8AFBDBED00061FCEDBBBEFF67B7350DB7773C408F746BC4";
    attribute INIT_2E of inst : label is "4B47ADA52862AE7AA713D330B57FE6CDFB5B79ECDBBE9DFCE95EDB77BD87C6DB";
    attribute INIT_2F of inst : label is "FFFFD6C3C0770E20F441220BCFB63ADB2E8976FD5B0C3FB3EC711D90FFFFA342";
    attribute INIT_30 of inst : label is "46AC91AB7EB6EEEDBBBB6EEFFFEAB54860BAF7A03FEFFEA68FFCDFFFFFF6FEFF";
    attribute INIT_31 of inst : label is "400000025C4B402028001484B80904800010924900126124920024828D891AB2";
    attribute INIT_32 of inst : label is "00010A100010A1000400100010A1000400100010A100040016808044B8968040";
    attribute INIT_33 of inst : label is "11540A32400AA480000402002482002002480000000402002482002002482480";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFCC2618C52249241D2000049C6149080000000000061C47A15A40";
    attribute INIT_35 of inst : label is "8AEE248ECC645555ADBCA506C36ECADDF1E50979521E506F2A3DC6CF89C77B44";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF9A7228C823221C847219848661219148645CDABE";
    attribute INIT_37 of inst : label is "A427AAC0465E428A0B5791126094102504D6EFD090D03667230E41290212008C";
    attribute INIT_38 of inst : label is "C9D15F5554BA9AA6AFAAE1358C3444B25D0F2787B8AB47C3231B88D005A376A0";
    attribute INIT_39 of inst : label is "A1C80A40142200400F01E00A01400F80F002004056774C28302041C0090E0009";
    attribute INIT_3A of inst : label is "80118824804D00120000200000000738014016047301869C10D3465500768604";
    attribute INIT_3B of inst : label is "E050C8199160510160A202C144058288054098804804D0092002620120034024";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5376A01C";
    attribute INIT_3D of inst : label is "79EF3D0A81A3356DF8AFBDBED00061FCEDBBBEFF67B7350DB7773C408F746BC4";
    attribute INIT_3E of inst : label is "4B47ADA52862AE7AA713D330B57FE6CDFB5B79ECDBBE9DFCE95EDB77BD87C6DB";
    attribute INIT_3F of inst : label is "FFFFD6C3C0770E20F441220BCFB63ADB2E8976FD5B0C3FB3EC711D90FFFFA342";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "DEB8E1E3797804EEDEDE818C0A01100125362899120D8E3B5CCC6D993326947C";
    attribute INIT_01 of inst : label is "73D9911CAF3298275A03938D153928D10C0769B5A6D074603A39322C3B12265D";
    attribute INIT_02 of inst : label is "5F7F6DB44FDBD00176DAEFFCFE4BABD47184BA49B6D9BCE27092CBDB762A2DA8";
    attribute INIT_03 of inst : label is "1A231AADCB3C11A26E4BE222B6C9B45A046DBF3EE67DCED589989B129F178999";
    attribute INIT_04 of inst : label is "1398D56E456D025927A237682BF6DB44FDBE5F7C4C49B6DAA0A906D86E872336";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF02C557C6C73267144546ED168A37AC6DCBCC06CE943C19B3A";
    attribute INIT_06 of inst : label is "ACB6457A62A3580280237B5714F561298CD2046C0D8C2B65D9B19962F3F6E934";
    attribute INIT_07 of inst : label is "B18DF9E88FF57B6B7842ADA4EA77FA4D34497201548354454B2443451B34901C";
    attribute INIT_08 of inst : label is "A496491EBC611DDF88E54AD367FBACB1AEB680CF84444EF5ADC4F7DC4F2C9555";
    attribute INIT_09 of inst : label is "00000101404EEEEEEEEEEEEEEEAA5E2B67BFCCFF9B5E6F7AD8E2DCAA89B258E3";
    attribute INIT_0A of inst : label is "5564A2AFA30387C0040104050505014540040005014401004040000004040140";
    attribute INIT_0B of inst : label is "0DE2BF800000003ABA800000003A3A37DE1C9E9886515A1A69C4E12597CF22B5";
    attribute INIT_0C of inst : label is "D5E4E67186E24E3D2A570A94B4B5AEBDD5DC5D745EAA6799E9EB3976DC4E75D0";
    attribute INIT_0D of inst : label is "012187A0CF2E45A81B3A46502D9C69BD281B336152A56BAE8EB9999FE497AF6F";
    attribute INIT_0E of inst : label is "FF00E474D2C9340D6D10D77E79788400000176D67795BF9E780000125F7F1C00";
    attribute INIT_0F of inst : label is "05F2ED7E57D359016CE65F77E99CB8B67133EB8B547161E5C55CAB8C197DA731";
    attribute INIT_10 of inst : label is "B87E9353452EB5C3E87663D517C2DC0FA10269A58D34624D48A50B1CF5918F69";
    attribute INIT_11 of inst : label is "31BF93F3317C3B3A3AC2B9AC5FBF94F55EAA000000000000000000464C489135";
    attribute INIT_12 of inst : label is "8EFCC146700BCAE2576F062AE899C9B1DFC2655E333DCC67D1B391FEF4AAA555";
    attribute INIT_13 of inst : label is "6820A0005000280014000A0005000A80044000A001500000AA8086D543B56E76";
    attribute INIT_14 of inst : label is "F26EE2632C5836435A9F299618AB0A0008B217FE519D82DC3ED3D7493C12CF6E";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFF38FC97231FA9D5AEEAAC21590BFF28D821DB4640C3E88B0";
    attribute INIT_16 of inst : label is "7F5931A3C54DAB797DEF4F7A8E27331B56DA32F2D1232F134829622A7339C9A4";
    attribute INIT_17 of inst : label is "644446646466464644644446446B50152E11FFFFEEBBA02C1C4E2831A140115D";
    attribute INIT_18 of inst : label is "FF3FFFFFFFFFFCFFFFFFFFFEBABBEAFEC4E6C646464646446444444444444444";
    attribute INIT_19 of inst : label is "EBB804024004620020441008048008801142203BFBEBEAFEFAFEB3FFFF33FFF3";
    attribute INIT_1A of inst : label is "100BBBEE80100C4488C44008048A4448AEFBAF112224522311229118891122AE";
    attribute INIT_1B of inst : label is "AAA88A88888AABBBC46231188C4622EEE040840842BBE0100804020100804020";
    attribute INIT_1C of inst : label is "84001E18431C0504114AABAFEFBFFFFFFF5444445445555444455544AAA8888A";
    attribute INIT_1D of inst : label is "8403C03C07B0CB492C4E143081C37F00004F600D9000360006C000E1084C20C1";
    attribute INIT_1E of inst : label is "0E2C8EA1993884300B20006C000D8001E2007DC40500C5000C0050E310D16201";
    attribute INIT_1F of inst : label is "800A00028020A000180050000000011800A000A002000555000E210D11610F10";
    attribute INIT_20 of inst : label is "00000000710000000000000140B54008259500DFC00013D8030360006C000DCE";
    attribute INIT_21 of inst : label is "224920000200000011208000064000124928000024801000004900500C400000";
    attribute INIT_22 of inst : label is "1020000102000010204081020000102040810200001020408D12490004000000";
    attribute INIT_23 of inst : label is "91C1008242880002080000410000410410000012080000410000410410000008";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFC8642045B000000D2049200801020A929292929295150D128070";
    attribute INIT_25 of inst : label is "57330614004CF719E8B58782C36508F1EA243889B1A24AD12972AA23CAE96324";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF980001000400100040430810C20430810C221766";
    attribute INIT_27 of inst : label is "9CC252E076F7AA0E03F6B490628418A10657ADAC00D03D5EA20A41A3001A008C";
    attribute INIT_28 of inst : label is "4D2DD39FFE040FF0E9CF818769ACCD936535769AA9F3F6876718A4C344E13589";
    attribute INIT_29 of inst : label is "000204101C08C1182AC1582560AC10E01C11803040330D8851A147480B0A349A";
    attribute INIT_2A of inst : label is "1802040018043000600010006000C331BFDFE807D520F18C3F61070000602821";
    attribute INIT_2B of inst : label is "C6280C081880700080E00101C00203802EC02040018043000600810006010C00";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9973B00C";
    attribute INIT_2D of inst : label is "1C5339C96DE16D6C9DF2CADE94006300DB77B649615BBF0D91130E51A86263A4";
    attribute INIT_2E of inst : label is "6325C52D3862B6BFF23BD6B0F12504C9991B2BB56DFED7F6ABF8D9194D8C46D9";
    attribute INIT_2F of inst : label is "FFFFE9B6C2D45A0CACD52A4C0C920A490C49FFDA472C123C8DDB0C8DAAAAAAB0";
    attribute INIT_30 of inst : label is "00000000710000000000000140B54008259500DFC00013D8030360006C000DCE";
    attribute INIT_31 of inst : label is "224920000200000011208000064000124928000024801000004900500C400000";
    attribute INIT_32 of inst : label is "1020000102000010204081020000102040810200001020408D12490004000000";
    attribute INIT_33 of inst : label is "91C1008242880002080000410000410410000012080000410000410410000008";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFC8642045B000000D2049200801020A929292929295150D128070";
    attribute INIT_35 of inst : label is "57330614004CF719E8B58782C36508F1EA243889B1A24AD12972AA23CAE96324";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF980001000400100040430810C20430810C221766";
    attribute INIT_37 of inst : label is "9CC252E076F7AA0E03F6B490628418A10657ADAC00D03D5EA20A41A3001A008C";
    attribute INIT_38 of inst : label is "4D2DD39FFE040FF0E9CF818769ACCD936535769AA9F3F6876718A4C344E13589";
    attribute INIT_39 of inst : label is "000204101C08C1182AC1582560AC10E01C11803040330D8851A147480B0A349A";
    attribute INIT_3A of inst : label is "1802040018043000600010006000C331BFDFE807D520F18C3F61070000602821";
    attribute INIT_3B of inst : label is "C6280C081880700080E00101C00203802EC02040018043000600810006010C00";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9973B00C";
    attribute INIT_3D of inst : label is "1C5339C96DE16D6C9DF2CADE94006300DB77B649615BBF0D91130E51A86263A4";
    attribute INIT_3E of inst : label is "6325C52D3862B6BFF23BD6B0F12504C9991B2BB56DFED7F6ABF8D9194D8C46D9";
    attribute INIT_3F of inst : label is "FFFFE9B6C2D45A0CACD52A4C0C920A490C49FFDA472C123C8DDB0C8DAAAAAAB0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "0AA2702261408C89B19210A41C3D11446036704600C18820408C5B0502001549";
    attribute INIT_01 of inst : label is "C2A09BB18F66586F3605B78F3CB378F3AD0B48152040B128589006786E376EE4";
    attribute INIT_02 of inst : label is "4444DB6D573255514DB2AA4300DEAA50C104B6DC12492616E336894D726E6E38";
    attribute INIT_03 of inst : label is "2BEB0B84C6200E39620246766DC06C362CD8B436407C8DA59A1BBB98BB148918";
    attribute INIT_04 of inst : label is "F3585C260CDB1A55C41662D8088DB6D57B241246E4DB6DB6A81B47C8AA836172";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF00D554AC4D67273EF70C5B0D8772F0E5EA812E42B41D0B90A";
    attribute INIT_06 of inst : label is "5960E314D4A33907003A02CBDAC565519A44241CC18A3052111133CAEA912081";
    attribute INIT_07 of inst : label is "231B6AC30E12A6E6DA86AB77034400DB6570552ACEA720C10B05072F1E341059";
    attribute INIT_08 of inst : label is "8DC246186041342C30EAD58146A29211B4BE40242CCCC2257DECCCDECC2C155A";
    attribute INIT_09 of inst : label is "0441110104550505050505050541B22A66A93300399CE47270C0D1557696F0C2";
    attribute INIT_0A of inst : label is "5450A22C28C094A0040101044454010011044514010114010511044115054114";
    attribute INIT_0B of inst : label is "03EAB2B5AD6CFB510014ED14CD0091813E92A8B9E7A85C4061ADC66D122752A5";
    attribute INIT_0C of inst : label is "32C4422082CC642856AA15AB6260F111999519571D2C324CA8423026B18A8CA0";
    attribute INIT_0D of inst : label is "592087A4DAA59390312AFAA83895ACA554312A02B568AB2AECA0CCCF99BC9CCB";
    attribute INIT_0E of inst : label is "FF6679249848D2041B3CCE4AB148840AA22829BC4C15206197FFFFE6F55215D1";
    attribute INIT_0F of inst : label is "B15E1A8A1083F1255F095BC14912B6E96D4BC10B5F21653085C82BBCD928A565";
    attribute INIT_10 of inst : label is "6C505A1644A08689060536141220934766A283364066911881AAB110C31A48D0";
    attribute INIT_11 of inst : label is "E5B105B43F69FBF7DE9BF13C0FAEC858890A000000000000000000E99880C0C1";
    attribute INIT_12 of inst : label is "4AB0CD9A98170936D52801CF9A85136D54EC6D53940F1B74841413D441801402";
    attribute INIT_13 of inst : label is "7562855142A8A15450AA2855142A8215400AA2855042ADDD770025CCD3925A72";
    attribute INIT_14 of inst : label is "A3D31E0B303028468B378E0214AEF55D7743ED553139E2102E48E605CD124FFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFC24BDF37B54A91A03B98CB951D6AA909E2102C6510651DE1";
    attribute INIT_16 of inst : label is "A092B1E7DCDB6A4C49C9D6C1966C23172DB6A321CB6A330B30A198AA4A4B2081";
    attribute INIT_17 of inst : label is "31339331393B1393933B1933B1AAFBFAEBEBFFFF98D6200D861C4E3393801D8A";
    attribute INIT_18 of inst : label is "F0F3C3330CC0F33C0C00000FEAEBABBFB919391BB19313B31193111131111339";
    attribute INIT_19 of inst : label is "FBE9148B545562A2A545588C46A8AAD1516A2A2AEBBAAFBFFEEABC000CFCFC3C";
    attribute INIT_1A of inst : label is "100BEBAFC0500D562091602806AA11623AEBEF112220180A012291100C0500BA";
    attribute INIT_1B of inst : label is "0222000220202BAA9140201009148BAFB44AD62D6BEBE0100804020100804020";
    attribute INIT_1C of inst : label is "D30101A843861104550BBBAEFABEFFFFFF010110001110111000100402000222";
    attribute INIT_1D of inst : label is "84003FF3F998FFDFF9DB181081C9FF0000009FF46FFFF600003FFFA10F3FDFC2";
    attribute INIT_1E of inst : label is "F6241482FF50863B68DFFFEC00007FFF63FFF887FFAB7FAAB6AAAE4310E0C398";
    attribute INIT_1F of inst : label is "FFFF56B7FFD55FFFEFBFFDB6DB6DBECFFFF56FFFFFFFFFFFAAA6218999B1E21F";
    attribute INIT_20 of inst : label is "B1916C643E5B9D36E74DB9D279FFFFF038D1EFFFFFE81227FDFFFDA46BFFFBFF";
    attribute INIT_21 of inst : label is "6FFFFB6DB6B6DB6DBFFBFFDB6FFFFFFFFFFB6DBFFFFFFFFFFFFFFF900F96C645";
    attribute INIT_22 of inst : label is "BD7AB56BD7AB56BD7AF5EBD7AB56BD7AF5EBD7AB56BD7AF5E7FFFFDB6D6DB6DB";
    attribute INIT_23 of inst : label is "51C2A102C08EDB6FF7FFFFBEDF7FBEDBEDB6FFEFF7FFFFBEDF7FBEDBEDB6DB5E";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFDC2E00477FFFFFF7EDFFFFF211FC0D6D6D6D6D6D681C17F48469";
    attribute INIT_25 of inst : label is "35155910184657310896079383642A85F8807A203708078407D10A8092C8E201";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF8007601DC07701DC076C11DB0476C11DB0442404";
    attribute INIT_27 of inst : label is "763301604F51B8410A140004076101D8400828001D414056B422FA8B83A8C0D1";
    attribute INIT_28 of inst : label is "59041E55547A2AAB0F2A3B1888A2BB5640A90654A50204048497803215E5F20F";
    attribute INIT_29 of inst : label is "D16F8B7C0037F0FE34F09E38F91F1C788F1FE0FC7A8C49D112264C2DAC0E08F4";
    attribute INIT_2A of inst : label is "01F983F387C20F9C0000000000000C00155FF103A4807A300F380155541AF240";
    attribute INIT_2B of inst : label is "00458001011282111204222408444810815F983F387E20F9C07E60FCE1F883E7";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF59320030";
    attribute INIT_2D of inst : label is "34CB18128B2125C4B8A6999A0030C101C932E25B4333651893369A5C81606281";
    attribute INIT_2E of inst : label is "4B05050CB972A96AA91312E0A825058A096129ACEBB4C9A6495989332F044F89";
    attribute INIT_2F of inst : label is "FFFFD6DC530A70460640006811B81ADBAC08F6D9481818370F7418D144050343";
    attribute INIT_30 of inst : label is "B1916C643E5B9D36E74DB9D279FFFFF038D1EFFFFFE81227FDFFFDA46BFFFBFF";
    attribute INIT_31 of inst : label is "6FFFFB6DB6B6DB6DBFFBFFDB6FFFFFFFFFFB6DBFFFFFFFFFFFFFFF900F96C645";
    attribute INIT_32 of inst : label is "BD7AB56BD7AB56BD7AF5EBD7AB56BD7AF5EBD7AB56BD7AF5E7FFFFDB6D6DB6DB";
    attribute INIT_33 of inst : label is "51C2A102C08EDB6FF7FFFFBEDF7FBEDBEDB6FFEFF7FFFFBEDF7FBEDBEDB6DB5E";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFDC2E00477FFFFFF7EDFFFFF211FC0D6D6D6D6D6D681C17F48469";
    attribute INIT_35 of inst : label is "35155910184657310896079383642A85F8807A203708078407D10A8092C8E201";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF8007601DC07701DC076C11DB0476C11DB0442404";
    attribute INIT_37 of inst : label is "763301604F51B8410A140004076101D8400828001D414056B422FA8B83A8C0D1";
    attribute INIT_38 of inst : label is "59041E55547A2AAB0F2A3B1888A2BB5640A90654A50204048497803215E5F20F";
    attribute INIT_39 of inst : label is "D16F8B7C0037F0FE34F09E38F91F1C788F1FE0FC7A8C49D112264C2DAC0E08F4";
    attribute INIT_3A of inst : label is "01F983F387C20F9C0000000000000C00155FF103A4807A300F380155541AF240";
    attribute INIT_3B of inst : label is "00458001011282111204222408444810815F983F387E20F9C07E60FCE1F883E7";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF59320030";
    attribute INIT_3D of inst : label is "34CB18128B2125C4B8A6999A0030C101C932E25B4333651893369A5C81606281";
    attribute INIT_3E of inst : label is "4B05050CB972A96AA91312E0A825058A096129ACEBB4C9A6495989332F044F89";
    attribute INIT_3F of inst : label is "FFFFD6DC530A70460640006811B81ADBAC08F6D9481818370F7418D144050343";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "53CCFDAD61AC0589BBB690801603E40452B45823046198D8511CDBA346883D5B";
    attribute INIT_01 of inst : label is "0E1522A1A946D86FB645B5AB31B35AB36C0B41990640B1285890466018244895";
    attribute INIT_02 of inst : label is "58CCDB6EAFF6D5540DC3AAFCFCD8AAC88718A69236522496D136DB49526A6820";
    attribute INIT_03 of inst : label is "2BEE563CC8532A31420286746DD06CB668DCC8A25544A9441852AA48AB158958";
    attribute INIT_04 of inst : label is "B272B1E60CDB2A3A0AD472D90B0DB6EAFF6C144EA4DB6DB7D55B5748ABB20A92";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF000755AA4D472D329D0E5B2D9753ECE5058D3A46AD905493A";
    attribute INIT_06 of inst : label is "FD6DE165ADA100E58FE490DB56C55315D4461C046198D84827137782C2B1260B";
    attribute INIT_07 of inst : label is "231922C52C8206CE48B68B6816C400DB6AC2DF039D2900C12B1D390D5AB47DDF";
    attribute INIT_08 of inst : label is "4DA6D05961C630AD52D0240456221295A1C2004CECCCC2CEFD04D5504D2C7BBE";
    attribute INIT_09 of inst : label is "0140500044155005500550055060412AC2ABFFFF39DCE57642DAD6AAAA96C2D8";
    attribute INIT_0A of inst : label is "4513D82CB008D5B0000005014151004555014451004011004055014051014051";
    attribute INIT_0B of inst : label is "0382B6D150DAA4C888B161B268998888382D58BDF62D5CA165ADA26DB6140AAD";
    attribute INIT_0C of inst : label is "36C65322A294C25081202048606C80959591D9015B2233CCAAD2B0A292952220";
    attribute INIT_0D of inst : label is "09081575A2F615C40372E38C21B625ADC603680409100B202C88CCCFE1B05CCB";
    attribute INIT_0E of inst : label is "FF42416594DA13001BBEEED8B0588422288029B0B0D57F9E68000006C556C680";
    attribute INIT_0F of inst : label is "2058241A01024F404255952B507325254AAA31107A22039887087060124C41EC";
    attribute INIT_10 of inst : label is "8BD192B8064CCA0900C408201804969608F3B16D662D598AA7C0335499555520";
    attribute INIT_11 of inst : label is "B9BCA5A19078EBA21A1FF5B6AF6E80701B83000000000000000000049BB2830B";
    attribute INIT_12 of inst : label is "D449264757EE6EAC1AB5E9DB2FEF6B8755C40556EC1C61D580C3BB54D4D576A8";
    attribute INIT_13 of inst : label is "402A0005000280014000A0005000280015000A000500020A28002F058716A4E2";
    attribute INIT_14 of inst : label is "2F0AAF326800C18102041260295BAA082AB611559B31B4704D58C602000007FB";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFC1B20D82E158B18022C8042BB28AAC59B420E06C60133E00";
    attribute INIT_16 of inst : label is "0F042DA706DB76DA5BDB56D1B6644F390DB74E1A4374E19118670DAAAAD9060B";
    attribute INIT_17 of inst : label is "C66C6C6E464EE464EEC46EEC46D454151101FFFFA19860002C3AD80082C7F200";
    attribute INIT_18 of inst : label is "FF3FFFFFFFFFFCFFFFFFFFF55501540024E46CE646CCE64E4E6E46EEE46EE6C6";
    attribute INIT_19 of inst : label is "54080403410462083044100804820A841142209454155555004013FFFF33FFF3";
    attribute INIT_1A of inst : label is "5881540595100C4602804A88048B01400054060180B1188A4500C0522C458840";
    attribute INIT_1B of inst : label is "00202220000225148048A452291401502568D48D4154355AAD56AA45AAD56AB5";
    attribute INIT_1C of inst : label is "EC01001023883EEFABE411504540FFFFFF100001110100000111011620222000";
    attribute INIT_1D of inst : label is "07FFFFF10120802005051028FE0BFF000000000FFFFFF600000000508EC01FC1";
    attribute INIT_1E of inst : label is "0A3FEC8590A840292FFFFFEC00000000A3FFF947FFABFFAABEAAAA8108D18389";
    attribute INIT_1F of inst : label is "B4AA0202AAAAAA955A4002DB6DB6DB7B4AA024AAAB555555000A008EEEC1E410";
    attribute INIT_20 of inst : label is "008000207180080002000081863FFFFC3BEF18FFC000000003FF6000000007D2";
    attribute INIT_21 of inst : label is "26DB6924929249249B69BDC926DB6DB6DB69249B6DB6DB6DB6DB6DF18C600200";
    attribute INIT_22 of inst : label is "162C183162C183162C58B162C183162C58B162C183162C58BDB6DB4925249249";
    attribute INIT_23 of inst : label is "F1E510E2430B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D8B";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFC9E4F0C5B6DB6DBDA4DB6DBC3103880000000000071FEF0B0870";
    attribute INIT_25 of inst : label is "9DD900000044A91315B8030C01787B0AF488CCA21AA88C94465309CC9ACE660B";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF8000F003C00F003C008000200008000200088CC8";
    attribute INIT_27 of inst : label is "2CEC92075EAD2D0E242A08200608018200D054D191E06297C79463D7063D8219";
    attribute INIT_28 of inst : label is "184820F554D2EAAF107A7338F344C9460339CF9C79142A0C1C1981002902F7B9";
    attribute INIT_29 of inst : label is "01028817E000EE1C00EE1C00760E00770E01DF380100080850A146C928C85694";
    attribute INIT_2A of inst : label is "11FC8BF917F22FE447FE2FFC5FF8B0413FDFE00B880170402F0405FFFC012040";
    attribute INIT_2B of inst : label is "040208E010070602070C040E18081C302EDFC8BF917F22FE447F22FE45FC8BF9";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7DB20081";
    attribute INIT_2D of inst : label is "38DB0B168801650DB9A69B9E806701A04B3206DB73730101B3371C688D61E61B";
    attribute INIT_2E of inst : label is "DB1F1FC460A5748AAEB3A3002CCB0A3D5BD379ACCBBCB1E58B5E1B336C00561B";
    attribute INIT_2F of inst : label is "FFFFC4536AE64C8DC44180D209B59ADBEC3874D0A1C060B12C400721EEBFF746";
    attribute INIT_30 of inst : label is "008000207180080002000081863FFFFC3BEF18FFC000000003FF6000000007D2";
    attribute INIT_31 of inst : label is "26DB6924929249249B69BDC926DB6DB6DB69249B6DB6DB6DB6DB6DF18C600200";
    attribute INIT_32 of inst : label is "162C183162C183162C58B162C183162C58B162C183162C58BDB6DB4925249249";
    attribute INIT_33 of inst : label is "F1E510E2430B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D8B";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFC9E4F0C5B6DB6DBDA4DB6DBC3103880000000000071FEF0B0870";
    attribute INIT_35 of inst : label is "9DD900000044A91315B8030C01787B0AF488CCA21AA88C94465309CC9ACE660B";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF8000F003C00F003C008000200008000200088CC8";
    attribute INIT_37 of inst : label is "2CEC92075EAD2D0E242A08200608018200D054D191E06297C79463D7063D8219";
    attribute INIT_38 of inst : label is "184820F554D2EAAF107A7338F344C9460339CF9C79142A0C1C1981002902F7B9";
    attribute INIT_39 of inst : label is "01028817E000EE1C00EE1C00760E00770E01DF380100080850A146C928C85694";
    attribute INIT_3A of inst : label is "11FC8BF917F22FE447FE2FFC5FF8B0413FDFE00B880170402F0405FFFC012040";
    attribute INIT_3B of inst : label is "040208E010070602070C040E18081C302EDFC8BF917F22FE447F22FE45FC8BF9";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7DB20081";
    attribute INIT_3D of inst : label is "38DB0B168801650DB9A69B9E806701A04B3206DB73730101B3371C688D61E61B";
    attribute INIT_3E of inst : label is "DB1F1FC460A5748AAEB3A3002CCB0A3D5BD379ACCBBCB1E58B5E1B336C00561B";
    attribute INIT_3F of inst : label is "FFFFC4536AE64C8DC44180D209B59ADBEC3874D0A1C060B12C400721EEBFF746";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "CF58176869F810E5B0B65A840A07745130B82899135C84E70ECC1B193324D866";
    attribute INIT_01 of inst : label is "274DB91884321B6F36199604103960410CB364B992DB336D99B9222C41162C5F";
    attribute INIT_02 of inst : label is "0272DB6D4716D1156DC8033302D90304679EB2D9F2DB6E76F1B61B9D76262C80";
    attribute INIT_03 of inst : label is "10261EE5C9700B74245922222DC96C36045DD6B0DD65AC19895913BF1306055B";
    attribute INIT_04 of inst : label is "5330F72E445B065D2E2236D8606DB6D4716EC9F06C5B6DB6AA8B5658419E23C6";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF03400644E63764986E46DB0D8636206DD78082C01CF41E300";
    attribute INIT_06 of inst : label is "08B22C0E6235082280EEC84310D53065E5421E645C84E721D9709888C8C1C934";
    attribute INIT_07 of inst : label is "912B6CC8AED996C2D9460374A87192DB754B15068699046C8B24C90E0C109138";
    attribute INIT_08 of inst : label is "2D96E95839E7964C8AE9D3B05678CBB093E200B28464581F01FAD99FEDAC9FFB";
    attribute INIT_09 of inst : label is "05414101005000055550000555A24803240C00009B8E4C32CAD045555536CAC0";
    attribute INIT_0A of inst : label is "0034C00C33088620040100040404010004050144010105014545054155054105";
    attribute INIT_0B of inst : label is "0BA0288A06010111110A96499340002DBA3E8E39B6605C1D75EDE36C360D0030";
    attribute INIT_0C of inst : label is "90DCF76C1662CF794E98D3A766259330E0E08E0008C1675D8B8AB70ECC5EBC10";
    attribute INIT_0D of inst : label is "0189C17DA4BE61DE0B7165BC05BE4000DE0B66DA74EB81C007059DDFFDB2186B";
    attribute INIT_0E of inst : label is "FF42E61862DD3286DB36CEDB39608488AA082DB2F2819FFFFFFFFFF6C8180000";
    attribute INIT_0F of inst : label is "2018609A0290CF04BA075D00EB9CBCB7793B258BC2B17852CCAF0B145B71AF24";
    attribute INIT_10 of inst : label is "90AD4AC90D2726CFC872499023864A00C3F7E5E1FCBC7F2EFCBBD010F1F1FB04";
    attribute INIT_11 of inst : label is "881C8363121067B744063DB55F3FAF92E00600000000000000000052EC48932C";
    attribute INIT_12 of inst : label is "1EFC36C5F402C7E84F7F575B7BA785900657A018210CC50611A89AABFC2AED55";
    attribute INIT_13 of inst : label is "8020000000000000000000000000000000000000000002A02A80D1000720FEE4";
    attribute INIT_14 of inst : label is "032FE7E20658F7C060C0238AB2A800A2801712ABD1B5AFD13C81C10D34020DB3";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFC3FF445024601CD564A55755BA955E0DAF91B6C2A4008E30";
    attribute INIT_16 of inst : label is "9069A1B744DB6ADB61DB66488633B3090DB6B2C6436B2D7508F96A02E324E934";
    attribute INIT_17 of inst : label is "1B1B31931B1131B13193B3193B0055401401FFFFE659803450C621508140772C";
    attribute INIT_18 of inst : label is "F3FFFFFFFFFFFFFFFFFFFFF5555400003B99333B193BBB913BB33933339331B3";
    attribute INIT_19 of inst : label is "000D56AA0101400830001AAD56020084004000950015555555554CC0CCFFFF3F";
    attribute INIT_1A of inst : label is "12240005801AA914A8D5400D5622546A950007552A3552A355AA951AA951AA55";
    attribute INIT_1B of inst : label is "00202222222000559148A45229140000254AD628415560100804031100804020";
    attribute INIT_1C of inst : label is "86FEFF90224A0505414015505005FFFFFE011111110100000111100402222000";
    attribute INIT_1D of inst : label is "0400000EFE48800002241B21FFD200FFFFFFFFF4000009FFFFFFFF90086FE039";
    attribute INIT_1E of inst : label is "CA3BCF79EF284236D8000013FFFFFFFF22000144005440554555552000A90271";
    attribute INIT_1F of inst : label is "CB55FDFD5555556AACB5AD249249248CB55FDB5554AAAAAAFFF000080001041F";
    attribute INIT_20 of inst : label is "FF7FFFDFA97FF7FFFDFFFF7EF9E000006195EF803FFFFFFFFD009FFFFFFFFAFF";
    attribute INIT_21 of inst : label is "D92496DB6D6DB6DB64964236D92492492496DB6492492492492492021A5FFDFF";
    attribute INIT_22 of inst : label is "E9D3E7CE9D3E7CE9D3A74E9D3E7CE9D3A74E9D3E7CE9D3A7464924B6DADB6DB6";
    attribute INIT_23 of inst : label is "9329D4A3129C9249249249249249249249249249249249249249249249249274";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFE2712806492492465B24924011FC9FFFFFFFFFFFF813CCF20054";
    attribute INIT_25 of inst : label is "40007F2554895D103DBD802EC37E2E95F2804C201A0804C40660269240A12124";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFBCC7031C0C7031C0C77F31DFCC77F31DFCC01555";
    attribute INIT_27 of inst : label is "A00F8CC2C65668001244B7DCC1F7307DCC2489FC3641844EB8E62C8112C88866";
    attribute INIT_28 of inst : label is "04C6794AABCF95573CA578B9A8BA4DC1088E1F67942254F3E3D5BEE47DA35C39";
    attribute INIT_29 of inst : label is "F37D13E81E4F11E26F11E26F89F13788F13620C4DEFF9158102044A48301339C";
    attribute INIT_2A of inst : label is "30031806300C6018C0006000C0018FB304401F9077F20FBE40FBC800009EDCC7";
    attribute INIT_2B of inst : label is "CC7D981F31F8F861F8F0C3F1E187E3C3104031806300C6018C00C6018C031806";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC931223E";
    attribute INIT_2D of inst : label is "124361C3E5802C2DB4F24859296960F0197616D9090BB005B112CB6A82726124";
    attribute INIT_2E of inst : label is "43279F146ACABA955C1B063001FF8E7CDB0B7C846B322D91619E5B190D81065B";
    attribute INIT_2F of inst : label is "FFFFEF31E63DC634794650CF05B29CD90E4B349B52AC72B1AC0B039C11400EF2";
    attribute INIT_30 of inst : label is "FF7FFFDFA97FF7FFFDFFFF7EF9E000006195EF803FFFFFFFFD009FFFFFFFFAFF";
    attribute INIT_31 of inst : label is "D92496DB6D6DB6DB64964236D92492492496DB6492492492492492021A5FFDFF";
    attribute INIT_32 of inst : label is "E9D3E7CE9D3E7CE9D3A74E9D3E7CE9D3A74E9D3E7CE9D3A7464924B6DADB6DB6";
    attribute INIT_33 of inst : label is "9329D4A3129C9249249249249249249249249249249249249249249249249274";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFE2712806492492465B24924011FC9FFFFFFFFFFFF813CCF20054";
    attribute INIT_35 of inst : label is "40007F2554895D103DBD802EC37E2E95F2804C201A0804C40660269240A12124";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFBCC7031C0C7031C0C77F31DFCC77F31DFCC01555";
    attribute INIT_37 of inst : label is "A00F8CC2C65668001244B7DCC1F7307DCC2489FC3641844EB8E62C8112C88866";
    attribute INIT_38 of inst : label is "04C6794AABCF95573CA578B9A8BA4DC1088E1F67942254F3E3D5BEE47DA35C39";
    attribute INIT_39 of inst : label is "F37D13E81E4F11E26F11E26F89F13788F13620C4DEFF9158102044A48301339C";
    attribute INIT_3A of inst : label is "30031806300C6018C0006000C0018FB304401F9077F20FBE40FBC800009EDCC7";
    attribute INIT_3B of inst : label is "CC7D981F31F8F861F8F0C3F1E187E3C3104031806300C6018C00C6018C031806";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC931223E";
    attribute INIT_3D of inst : label is "124361C3E5802C2DB4F24859296960F0197616D9090BB005B112CB6A82726124";
    attribute INIT_3E of inst : label is "43279F146ACABA955C1B063001FF8E7CDB0B7C846B322D91619E5B190D81065B";
    attribute INIT_3F of inst : label is "FFFFEF31E63DC634794650CF05B29CD90E4B349B52AC72B1AC0B039C11400EF2";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "1E4055A840A0504491136A840E077BABFC9C3803004884E2388C0971E3041052";
    attribute INIT_01 of inst : label is "A5FC91188C324D27122C920C109920C127D9BC3AF0FD9E76CF3FE23405122479";
    attribute INIT_02 of inst : label is "062249240622450424EE02BFFE4D02B4679E924F20C92772519209DF36222680";
    attribute INIT_03 of inst : label is "58240E218D500A546049622224CF2412044DD292D525A4208F4FF92C79051549";
    attribute INIT_04 of inst : label is "5920710C444902C8AAA2364820E4924062264BA06C49249200097359619401D6";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFF020C0546E6326E986EC6C9048236304C958ECAC25CA00EB09";
    attribute INIT_06 of inst : label is "92C0241C2455082380EFE849127FFCB4F5461E044884E21711F00088C8A2C100";
    attribute INIT_07 of inst : label is "11B13E6EA57DD2444F0201228022DA49202A301C085914668906890418301111";
    attribute INIT_08 of inst : label is "24F2454E39E79F66EA5FBF7053D1EF319BF200B70444483F24966EC966A45FF1";
    attribute INIT_09 of inst : label is "05455404051FFFFAAAAAAAAFFFE16E82980A0C0C9B9A6C60EA60C80809B26A61";
    attribute INIT_0A of inst : label is "002840083E898560000401004050040015014550040154050515054551014415";
    attribute INIT_0B of inst : label is "09002580000000333B00000000333B3F902C0410D3784F5D34E4A32412082020";
    attribute INIT_0C of inst : label is "926AF676063ACA55FDF97F7F36259BB181809800190076598AAA9B94A755DA70";
    attribute INIT_0D of inst : label is "01810145359A617E2931A7FC149A4484FE293DEFEFDF83000C01DD9FFC9B0869";
    attribute INIT_0E of inst : label is "FF42A6208E48A68F491E444F9950840000A3D49ABB011FFFF7FFFFF268150800";
    attribute INIT_0F of inst : label is "B03C60BB22F2C6047A0A4D01A90E9CDA3951A689CAD131D34CB52934493CA740";
    attribute INIT_10 of inst : label is "D4AD2AAD042287CE80200D5017464E02C3C5E6E2BCDCAF377D3FD11072F2B704";
    attribute INIT_11 of inst : label is "94840740123062844D062A541D3DBEF3E180000000000000000000AB4228F3AA";
    attribute INIT_12 of inst : label is "554AB255540406AC2A5442503B265ED8055F0015200C170554201E2AA62A8955";
    attribute INIT_13 of inst : label is "1560000000000000000000000000000000000000000007FFD50097008522A4A4";
    attribute INIT_14 of inst : label is "43BC8D8A1668FBC1E1C8E5CA3AAEFFFFFFF5DAAAA09CCF10B4894108B0CD3522";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFC3FC0701A45008D555354755ACD55584CF503EC2B4118A50";
    attribute INIT_16 of inst : label is "D2FBF0F20C49204F5189F268923A2309049203664120367518F1B002A216C100";
    attribute INIT_17 of inst : label is "E8E2AAA8E2EA8E6A8A2A28A6E2AAFFFFEAFEFFFFF45D00208B82475081C077BE";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFEAA68484A6A6846AAA48A2A88A6A8A6A";
    attribute INIT_19 of inst : label is "AAA804020000480020101008040000800440803FFFEBFABFABAAAFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "100AAAAF8010080400804008040200403FFFFA010020100201008010080100AA";
    attribute INIT_1B of inst : label is "2202000000000ABF8040201008048BFFE040848D6AAAA0100804020100804020";
    attribute INIT_1C of inst : label is "C7010018E20E7AAFEEAABEAAFFEFFFFFFE000000001011111000000400000222";
    attribute INIT_1D of inst : label is "8C0000010079800007273939801200000000000C00000000000000630C701001";
    attribute INIT_1E of inst : label is "0E640C819039C63B6800000000000000C702018EAAAAEAAAAEAAAAC610C9C601";
    attribute INIT_1F of inst : label is "EB5556B55555556ABEB5ADB6DB6DB6DEB5556B5556AAAAAAAAAE710800630630";
    attribute INIT_20 of inst : label is "9111244471C9111244449111CEA0000E71C672800000000003008000000006F7";
    attribute INIT_21 of inst : label is "6DB6DB6DB6B6DB6DB6DB6B5B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB630C724444";
    attribute INIT_22 of inst : label is "AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56F6DB6DB6D6DB6DB";
    attribute INIT_23 of inst : label is "F3C9E4E7D39EDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB56";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFA7D39C76DB6DB6F6DB6DB6E61931C2424242424263C0F031864";
    attribute INIT_25 of inst : label is "99990010004D5D10BC9E800F413E6ADDF2004C001A00054006A100DA08852102";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF80400100040010004000100004000100004CD999";
    attribute INIT_27 of inst : label is "884F96D24C5F288C0B6680000000000000F6EDE8B2C0B7452B6525820258002A";
    attribute INIT_28 of inst : label is "04CB7D8AABCC1557BEC570BDE9A95681005C550EB0B36680000680027CAB473A";
    attribute INIT_29 of inst : label is "01000000000000002000002000001000001000004000010810204480050033A8";
    attribute INIT_2A of inst : label is "000000000000000000000000000000002F800008000100002000040000000000";
    attribute INIT_2B of inst : label is "000000000000002000004000008000013F800000000000000000000000000000";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC931A000";
    attribute INIT_2D of inst : label is "1A49208346800CA49CD649CFE869A2F05966524B3939D01491134F6A8B316110";
    attribute INIT_2E of inst : label is "49179F9468EABED55609965043FF8F7FC9393D84691E34F1A08F491926810549";
    attribute INIT_2F of inst : label is "FFFFFB33E677CE34FD47D0CF1C9E8849262926DA0B347E92A48D0788AAA6AFA2";
    attribute INIT_30 of inst : label is "9111244471C9111244449111CEA0000E71C672800000000003008000000006F7";
    attribute INIT_31 of inst : label is "6DB6DB6DB6B6DB6DB6DB6B5B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB630C724444";
    attribute INIT_32 of inst : label is "AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56AD5AB56F6DB6DB6D6DB6DB";
    attribute INIT_33 of inst : label is "F3C9E4E7D39EDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB56";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFA7D39C76DB6DB6F6DB6DB6E61931C2424242424263C0F031864";
    attribute INIT_35 of inst : label is "99990010004D5D10BC9E800F413E6ADDF2004C001A00054006A100DA08852102";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF80400100040010004000100004000100004CD999";
    attribute INIT_37 of inst : label is "884F96D24C5F288C0B6680000000000000F6EDE8B2C0B7452B6525820258002A";
    attribute INIT_38 of inst : label is "04CB7D8AABCC1557BEC570BDE9A95681005C550EB0B36680000680027CAB473A";
    attribute INIT_39 of inst : label is "01000000000000002000002000001000001000004000010810204480050033A8";
    attribute INIT_3A of inst : label is "000000000000000000000000000000002F800008000100002000040000000000";
    attribute INIT_3B of inst : label is "000000000000002000004000008000013F800000000000000000000000000000";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC931A000";
    attribute INIT_3D of inst : label is "1A49208346800CA49CD649CFE869A2F05966524B3939D01491134F6A8B316110";
    attribute INIT_3E of inst : label is "49179F9468EABED55609965043FF8F7FC9393D84691E34F1A08F491926810549";
    attribute INIT_3F of inst : label is "FFFFFB33E677CE34FD47D0CF1C9E8849262926DA0B347E92A48D0788AAA6AFA2";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
