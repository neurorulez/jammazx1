-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_8E is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(11 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_8E is

	signal rom_addr : std_logic_vector(11 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(11 downto 0) <= ADDR;
	end process;

	ROM_8E_0 : RAMB16_S4
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"0000CEEC0008CC08EEC000000CC80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_02 => x"FFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFF00000033FFFFFFFF",
		INIT_03 => x"33000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFF",
		INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => x"000000000660000000000000000000000000000000000000026C800000008C62",
		INIT_06 => x"000EE0000CE222EC046222EC08888EE8046222EC06EEAA22022EE22008C622C8",
		INIT_07 => x"00AA00000EE0000000000000EE00AAEE0C2EAA2C0C2AAA2C002226C80CE222EC",
		INIT_08 => x"08C622EE0EE000000EE222200EE226C808C622640EE222EC0EE888EE00000000",
		INIT_09 => x"0CE222EC0EE08CEE0EE080EE0EE222200EE8CE62046222EC022EE2200EE000EE",
		INIT_0A => x"0CEC8CEC008CEC800CE222EC000EE000046222EC0EE8CE620CE2AECA0EE88880",
		INIT_0B => x"F1111111F00000001111111F0000000F0000000006EEA222000EE00006EC8CE6",
		INIT_0C => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_0D => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_0E => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_0F => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_10 => x"0000000000000377000000007730000000000008000003488000000000100000",
		INIT_11 => x"008CE7777FF80000777EC80000008FF7000008CC0037FC88CC80000088CF7300",
		INIT_12 => x"000CEECC000133579126C0003730000000000EFF00000FFFFFE00000FFF00000",
		INIT_13 => x"00000000000000000000000000000000000CEECC0001337F9126C000F7300000",
		INIT_14 => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_15 => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_16 => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_17 => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_18 => x"33333333000000003333FFFF0000FFFFFFFF3333FFFF00003333333300000000",
		INIT_19 => x"33333333000000003333FFFF0000FFFF33333333000000003333FFFF0000FFFF",
		INIT_1A => x"33333333000000003333FFFF0000FFFF33333333000000003333FFFF0000FFFF",
		INIT_1B => x"FFFFFFFFFFFFFF00FFFF0000FF00000000000000FFFFFFFFFFFFFF00FFFF0000",
		INIT_1C => x"00000000FFFFFFFF00FFFFFF0000FFFF00000000000000000000000000000000",
		INIT_1D => x"00000000000000000000000000000000FFFFFFFF00FFFFFF0000FFFF000000FF",
		INIT_1E => x"0000000000000000000000000FFFF0000000FFFFEFF73000EEEEEEEE000037FF",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"00000000000000008044666E000000000000000000000008C800000000000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"FFFFFFFFFFFFFFFF000000FF000000FF33333333FFFFFFFF33333333FFFFFFFF",
		INIT_23 => x"FF000000FF000000FFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFF00000000",
		INIT_24 => x"AAAAAAAAFFFFFFFFAAAAAAAAFFFFFFFF008C42AA0F0FFFFFAAAAAAAAFFFFFFFF",
		INIT_25 => x"AAAAAAAAFFFFFFFFAAAAAAAAFFFFFFFFAAAAAAAAFFFFFFFFAAAAAAAAFFFFFFFF",
		INIT_26 => x"AAAA222237FFFE8022222222017FFFC0AAAAAAAAFFFFFFFFAAAAAAAAFFF73100",
		INIT_27 => x"AAAAAAAAF710008EAAAAAAAA88800000222222AA0FFF000CAAAAAAAA8000007F",
		INIT_28 => x"22222AAA310000002222222200000000AAAAAAAA00008C28AAAAA222EFFFF773",
		INIT_29 => x"22222AAA18AF8CEFAA24C800EC8FF0F02AAAAAAA001F71CFA2222222FFFFBBB0",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_2D => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_2E => x"FFFFF000FFFFF000EFFFF000FFFFF00088888888888888888888888888888888",
		INIT_2F => x"888888889BFFF88889BFF000FFFFF88888888000FEC8888889BFF000FFFFF888",
		INIT_30 => x"00000000000037FF00000000FF73000000000000005773770000000073777300",
		INIT_31 => x"008CE7777FF80000777EC80000008FF7000008CC0037FC88CC80000088CF7300",
		INIT_32 => x"00004A4A00EFFDEF04EEE000FFEFFF0000004A4A00EFFDEF0CEEA000FFEFFF00",
		INIT_33 => x"00004A4A00EFFDEF04EEE000FFEFFF0000004A4A00EFFDEF008CE000FFEFFF00",
		INIT_34 => x"F1111F1FF1F33F1FF1333F1FF1D5F51FCCCCCCCCCCCCCCCCCCCCCC00FECCCCCC",
		INIT_35 => x"F1F1111FF1F3331FF1F33F1FF1F3371FF1F33F1FF1F11F1FF1333F1FF1F33F1F",
		INIT_36 => x"00000E0000E22E0000222E0000C4E40000622E0000EAAA000002E20000E22E00",
		INIT_37 => x"00E0000000E2220000E22E0000E2260000E22E0000E00E0000222E0000E22E00",
		INIT_38 => x"00008CCA0000133724C800007330000000000EFF00000FFFFFE00000FFF00000",
		INIT_39 => x"000CEECC000133779126C00037300000000CEECC000133779126C00077300000",
		INIT_3A => x"0000CEEF0000011FFEEC000031100000000000CC00087077EEECC000FFF77000",
		INIT_3B => x"0000CEEF0000011FFEEC0000311000000000CEEF0000011FFEEC000031100000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0000",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8E_1 : RAMB16_S4
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"004EF737007337FF37FE4000F7337000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_02 => x"FFFFFFFFFFFFFFFFFFFFFFFF000000CCFFFFFFFFFFFFFFFF00000000FFFFFFFF",
		INIT_03 => x"00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC000000FFFFFFFFFFFFFFFF",
		INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => x"00000000000000000111111000000000000000000000000008C73000000037C8",
		INIT_06 => x"0CC89BEC037D99900EEAAAB90136CFF00089BFD804C99BF6004FF00003788C73",
		INIT_07 => x"00FFF00007755702000CE00077203322078BAB87078BAA8706F999F706F999F6",
		INIT_08 => x"037C89990FF999980FF999800FF88C73037C88C40FF999F6037C8C7300000000",
		INIT_09 => x"07F888F70FF731FF0FF737FF0FF000000FF136C8000000FF088FF8800FF111FF",
		INIT_0A => x"0FF131FF0FF101FF0FF000FF088FF88006F999D40FF889F707F888F70FF88887",
		INIT_0B => x"F0000000F88888880000000F8888888F000000000889BFEC0CF11FC00CE737EC",
		INIT_0C => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_0D => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_0E => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_0F => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_10 => x"00000CEE00000000EEC000000000000000002C010000000012E2000000000000",
		INIT_11 => x"EFF1000000137EEE00001FFEEEE7310000CEF31100000133113FEC0033100000",
		INIT_12 => x"007FFFFF00000000FFC013000000000000000FFF00000001FFF0000010000000",
		INIT_13 => x"00000000000000000000000000000000007FFFFF00000001FFC0130010000000",
		INIT_14 => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_15 => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_16 => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_17 => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_18 => x"00000000CCCCCCCC0000FFFFCCCCFFFFFFFF0000FFFFCCCC00000000CCCCCCCC",
		INIT_19 => x"00000000CCCCCCCC0000FFFFCCCCFFFF00000000CCCCCCCC0000FFFFCCCCFFFF",
		INIT_1A => x"00000000CCCCCCCC0000FFFFCCCCFFFF00000000CCCCCCCC0000FFFFCCCCFFFF",
		INIT_1B => x"FFFFFFFFFFFFFF00FFFF0000FF00000000000000FFFFFFFFFFFFFF00FFFF0000",
		INIT_1C => x"00000000FFFFFFFF00FFFFFF0000FFFF00000000000000000000000000000000",
		INIT_1D => x"00000000000000000000000000000000FFFFFFFF00FFFFFF0000FFFF000000FF",
		INIT_1E => x"FFEC8000FFFFFFFF00008CEF0FFFF0000000FFFF110000001111111100000001",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"0000000000000000100000000000000000000000CCC66331013264CC00000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"FFFFFFFFFFFFFFFF000000FF000000FF00000000FFFFFFFF00000000FFFFFFFF",
		INIT_23 => x"FF000000FF000000FFFFFFFFFFFFFFFFFFFFFFFFCCCCCCCCFFFFFFFFCCCCCCCC",
		INIT_24 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0E1CEFFF0F0FFFFFFFFFFFFFFFFFFFFF",
		INIT_25 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_26 => x"398C000080017FFF6EEEE800C001BBB2FFFFFFFFFFFFFFFFFFFFFFF7F70EFFEC",
		INIT_27 => x"8880000010004677003FFF33310000080CC8000007FF000F13733008F7080001",
		INIT_28 => x"CC88000100000800000000004CEEEFFF00000000CEFFF0630088CCCC31100000",
		INIT_29 => x"C4000F73FFFFFFFF7F1EC1E0FFFFF0F001FFFF710001CFFF1888CCC0FFFF718C",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_2D => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_2E => x"FFFFF000FFFFF000FFFFF0007FFFF000FFFFFFFFFFFFFFFFFFFFFFF77FFFFFFF",
		INIT_2F => x"FFFFF137FFFFFFFFFFFFF000FFFFF37FFFFFF000FFFFF137FFFFFEC8FFFFFFFF",
		INIT_30 => x"0000CEFF00000000FFEC00000000000000CEEACE00000000EECEEE0000000000",
		INIT_31 => x"EFF1000000137EEE00001FFEEEE7310000CEF31100000133113FEC0033100000",
		INIT_32 => x"0000101000233133057730003133310000001010002331330577300031333100",
		INIT_33 => x"0000101000233133077720003133310000001010002331330737300031333100",
		INIT_34 => x"F8CCCF8FF8FDDD8FF8FDDD8FF8F8988FFFFFFFFFFFFFFFFFFFFFFFC8FFFFFFFF",
		INIT_35 => x"F8FDDC8FF8FDDC8FF8999F8FF8FCCE8FF8F9998FF8FDDF8FF8FDDF8FF8FDDF8F",
		INIT_36 => x"0044470000755500007555000070100000645700006447000002700000744700",
		INIT_37 => x"0075540000755400001117000074460000711100007557000075570000755700",
		INIT_38 => x"0006FFFF00000000FC8160000000000000000FFF00000017FFF0000071000000",
		INIT_39 => x"007FFFFF00000000FFC0130000000000007FFFFF00000000FFC0130000000000",
		INIT_3A => x"0003FFFF00000000FFFF300012000000000800AA00034888AAAAA00043000000",
		INIT_3B => x"0003FFFF00000000FFFF3000120000000003FFFF00000000FFFF300012000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0000",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
