library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity eprom_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of eprom_1 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"ED",X"56",X"00",X"00",X"C3",X"A7",X"17",X"E5",X"26",X"C0",X"6F",X"36",X"00",X"E1",X"C9",
		X"E5",X"26",X"C0",X"6F",X"36",X"01",X"E1",X"C9",X"C5",X"D5",X"E5",X"C3",X"11",X"01",X"00",X"00",
		X"C5",X"D5",X"E5",X"3E",X"01",X"C3",X"11",X"01",X"21",X"00",X"C0",X"06",X"0A",X"C3",X"0B",X"01",
		X"6F",X"26",X"C0",X"36",X"01",X"C3",X"D8",X"00",X"32",X"10",X"D0",X"F5",X"3A",X"E0",X"C3",X"A7",
		X"28",X"3F",X"CD",X"BE",X"15",X"CD",X"B5",X"23",X"CD",X"22",X"02",X"CD",X"D6",X"02",X"CD",X"92",
		X"67",X"21",X"E0",X"C3",X"36",X"00",X"FB",X"CD",X"A9",X"00",X"F3",X"ED",X"73",X"27",X"C4",X"2A",
		X"27",X"C4",X"11",X"00",X"C0",X"ED",X"52",X"7C",X"FE",X"08",X"D2",X"AB",X"24",X"3E",X"01",X"32",
		X"E0",X"C3",X"F1",X"E1",X"E5",X"F5",X"11",X"00",X"C0",X"ED",X"52",X"D2",X"B0",X"24",X"F1",X"FB",
		X"C9",X"ED",X"73",X"23",X"C4",X"31",X"21",X"C4",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",
		X"22",X"02",X"CD",X"D6",X"02",X"CD",X"92",X"67",X"CD",X"BE",X"15",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"ED",X"7B",X"23",X"C4",X"F1",X"FB",X"C9",X"21",X"00",X"C0",X"7E",X"A7",X"28",X"21",
		X"35",X"20",X"1E",X"22",X"DE",X"C3",X"CB",X"25",X"3E",X"0A",X"85",X"6F",X"ED",X"73",X"21",X"C4",
		X"5E",X"23",X"56",X"EB",X"F9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"D9",X"E1",X"D1",X"C1",
		X"C9",X"2C",X"7D",X"FE",X"0A",X"20",X"D5",X"C9",X"1E",X"00",X"CB",X"3F",X"CB",X"1B",X"1F",X"CB",
		X"1B",X"1F",X"CB",X"1B",X"57",X"E5",X"21",X"2C",X"C0",X"19",X"EB",X"E1",X"CB",X"25",X"4D",X"3E",
		X"0A",X"85",X"6F",X"73",X"23",X"72",X"3E",X"10",X"83",X"5F",X"30",X"01",X"14",X"21",X"30",X"03",
		X"06",X"00",X"09",X"4E",X"23",X"46",X"EB",X"71",X"23",X"70",X"C9",X"36",X"00",X"23",X"10",X"FB",
		X"C9",X"D9",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"2A",X"DE",X"C3",X"77",X"CB",X"25",X"3E",
		X"0A",X"85",X"6F",X"ED",X"73",X"25",X"C4",X"ED",X"5B",X"25",X"C4",X"73",X"23",X"72",X"ED",X"7B",
		X"21",X"C4",X"2A",X"DE",X"C3",X"18",X"9A",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"09",X"0D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"09",X"0D",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"05",X"09",X"0D",X"11",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"06",X"09",X"0D",X"11",X"15",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"09",
		X"0D",X"11",X"15",X"19",X"1E",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"09",X"0E",X"11",X"15",
		X"19",X"1D",X"01",X"00",X"00",X"00",X"00",X"01",X"05",X"09",X"0D",X"11",X"15",X"19",X"1D",X"01",
		X"05",X"00",X"00",X"00",X"01",X"05",X"09",X"0E",X"11",X"16",X"19",X"1D",X"01",X"05",X"09",X"00",
		X"00",X"01",X"05",X"09",X"0D",X"11",X"15",X"19",X"1D",X"01",X"05",X"09",X"0D",X"00",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"12",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CD",X"2C",X"02",X"CD",X"51",X"02",X"CD",X"96",X"02",X"C9",X"DD",X"21",X"2B",X"C4",
		X"3A",X"0C",X"D0",X"CB",X"67",X"CD",X"41",X"02",X"DD",X"21",X"2D",X"C4",X"3A",X"0C",X"D0",X"CB",
		X"6F",X"3E",X"FF",X"20",X"08",X"AF",X"DD",X"BE",X"00",X"C8",X"DD",X"34",X"01",X"DD",X"77",X"00",
		X"C9",X"DD",X"21",X"2B",X"C4",X"3A",X"C1",X"C4",X"07",X"07",X"07",X"CD",X"68",X"02",X"DD",X"21",
		X"2D",X"C4",X"3A",X"C1",X"C4",X"07",X"07",X"07",X"E6",X"06",X"16",X"00",X"5F",X"21",X"20",X"03",
		X"3A",X"FF",X"BF",X"FE",X"76",X"28",X"03",X"21",X"28",X"03",X"19",X"DD",X"7E",X"01",X"96",X"D8",
		X"DD",X"77",X"01",X"3E",X"EF",X"CD",X"AE",X"67",X"3E",X"05",X"CD",X"AE",X"67",X"23",X"3A",X"32",
		X"C4",X"86",X"32",X"32",X"C4",X"C9",X"3A",X"31",X"C4",X"A7",X"20",X"0B",X"3A",X"32",X"C4",X"FE",
		X"09",X"30",X"04",X"CD",X"2C",X"20",X"C9",X"CD",X"38",X"20",X"C9",X"3A",X"32",X"C4",X"FE",X"09",
		X"D0",X"DD",X"21",X"2F",X"C4",X"3A",X"0C",X"D0",X"CB",X"57",X"CD",X"41",X"02",X"DD",X"7E",X"01",
		X"A7",X"C8",X"21",X"32",X"C4",X"86",X"77",X"DD",X"36",X"01",X"00",X"3E",X"EF",X"CD",X"AE",X"67",
		X"3E",X"05",X"CD",X"AE",X"67",X"C9",X"3A",X"31",X"C4",X"A7",X"C0",X"CD",X"AB",X"02",X"3A",X"0C",
		X"D0",X"CB",X"5F",X"28",X"05",X"AF",X"32",X"31",X"C4",X"C9",X"F3",X"CD",X"BF",X"95",X"3E",X"0E",
		X"32",X"FF",X"C7",X"CD",X"38",X"20",X"CD",X"17",X"21",X"CD",X"D0",X"21",X"3E",X"FF",X"32",X"31",
		X"C4",X"11",X"1B",X"03",X"21",X"60",X"E4",X"AF",X"CD",X"F1",X"21",X"11",X"00",X"00",X"06",X"03",
		X"32",X"10",X"D0",X"1B",X"7B",X"B2",X"20",X"F8",X"10",X"F6",X"C7",X"04",X"54",X"49",X"4C",X"54",
		X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"06",X"02",X"01",X"01",X"02",X"01",X"01",
		X"92",X"91",X"F7",X"30",X"00",X"00",X"23",X"36",X"B5",X"05",X"82",X"80",X"EA",X"4E",X"E2",X"76",
		X"3A",X"0C",X"D0",X"CB",X"77",X"28",X"F9",X"AF",X"32",X"18",X"D0",X"32",X"10",X"D0",X"21",X"00",
		X"00",X"3A",X"0C",X"D0",X"CB",X"77",X"28",X"F9",X"7E",X"32",X"18",X"D0",X"32",X"10",X"D0",X"3A",
		X"0C",X"D0",X"CB",X"77",X"28",X"F9",X"23",X"7D",X"FE",X"FF",X"20",X"E5",X"CD",X"90",X"04",X"7C",
		X"FE",X"BF",X"20",X"DD",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"CD",X"17",X"21",X"3A",X"18",
		X"D0",X"FE",X"55",X"20",X"13",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"CD",X"D0",X"21",X"3A",
		X"18",X"D0",X"32",X"8A",X"ED",X"A7",X"28",X"23",X"32",X"35",X"C4",X"AF",X"21",X"20",X"E5",X"11",
		X"AA",X"03",X"CD",X"D2",X"03",X"32",X"10",X"D0",X"18",X"FB",X"10",X"42",X"41",X"44",X"20",X"48",
		X"41",X"52",X"44",X"57",X"41",X"52",X"45",X"20",X"20",X"20",X"20",X"3E",X"00",X"F7",X"CD",X"59",
		X"04",X"CD",X"2C",X"20",X"FB",X"3A",X"35",X"C4",X"A7",X"28",X"FA",X"18",X"FD",X"CD",X"92",X"67",
		X"18",X"F3",X"C5",X"F5",X"F5",X"1A",X"47",X"0E",X"FF",X"F1",X"07",X"07",X"07",X"13",X"EB",X"12",
		X"13",X"ED",X"A0",X"1B",X"CD",X"0D",X"21",X"10",X"F6",X"F1",X"C1",X"C9",X"21",X"00",X"00",X"3A",
		X"0C",X"D0",X"CB",X"77",X"28",X"F9",X"7E",X"32",X"18",X"D0",X"32",X"10",X"D0",X"3A",X"0C",X"D0",
		X"CB",X"77",X"28",X"F9",X"23",X"7D",X"FE",X"FF",X"20",X"E5",X"CD",X"90",X"04",X"7C",X"FE",X"BF",
		X"20",X"DD",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"CD",X"17",X"21",X"3A",X"18",X"D0",X"FE",
		X"55",X"20",X"13",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"CD",X"D0",X"21",X"3A",X"18",X"D0",
		X"32",X"8A",X"ED",X"A7",X"28",X"23",X"32",X"35",X"C4",X"AF",X"21",X"20",X"E5",X"11",X"AA",X"03",
		X"CD",X"D2",X"03",X"32",X"10",X"D0",X"18",X"FB",X"10",X"42",X"41",X"44",X"20",X"48",X"41",X"52",
		X"44",X"57",X"41",X"52",X"45",X"20",X"20",X"20",X"20",X"E5",X"D5",X"C5",X"7B",X"E5",X"7A",X"57",
		X"84",X"65",X"6B",X"5F",X"30",X"01",X"14",X"C1",X"09",X"13",X"21",X"4E",X"03",X"11",X"EC",X"03",
		X"01",X"6D",X"00",X"1A",X"ED",X"A1",X"20",X"07",X"13",X"78",X"B1",X"20",X"F6",X"18",X"0D",X"ED",
		X"5F",X"32",X"32",X"C4",X"32",X"33",X"C4",X"32",X"34",X"C4",X"ED",X"47",X"C1",X"D1",X"E1",X"C9",
		X"E5",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"1E",X"21",X"B3",X"04",X"CD",X"50",X"20",
		X"7E",X"32",X"2B",X"E3",X"AF",X"32",X"2A",X"E3",X"23",X"7E",X"32",X"EB",X"E2",X"AF",X"32",X"EA",
		X"E2",X"E1",X"C9",X"31",X"31",X"31",X"30",X"20",X"39",X"20",X"38",X"20",X"37",X"20",X"36",X"20",
		X"35",X"20",X"34",X"20",X"33",X"20",X"32",X"20",X"31",X"20",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"09",X"0D",X"03",X"15",X"00",X"1E",X"01",X"06",X"09",X"0D",X"00",X"00",X"09",X"0D",X"03",
		X"15",X"19",X"00",X"01",X"05",X"0A",X"0D",X"03",X"00",X"00",X"0D",X"03",X"16",X"19",X"1D",X"00",
		X"05",X"09",X"0D",X"03",X"16",X"00",X"00",X"03",X"15",X"19",X"1D",X"01",X"00",X"09",X"0D",X"03",
		X"15",X"19",X"00",X"00",X"15",X"19",X"1D",X"01",X"05",X"00",X"0D",X"03",X"15",X"19",X"1D",X"00",
		X"00",X"19",X"1D",X"01",X"05",X"09",X"00",X"03",X"15",X"19",X"1D",X"01",X"00",X"00",X"1E",X"01",
		X"05",X"09",X"0D",X"00",X"15",X"1A",X"1D",X"01",X"05",X"00",X"00",X"01",X"05",X"09",X"0D",X"03",
		X"00",X"19",X"1D",X"01",X"05",X"0A",X"00",X"00",X"05",X"09",X"0E",X"03",X"15",X"00",X"1D",X"01",
		X"05",X"09",X"0D",X"00",X"00",X"09",X"0D",X"03",X"16",X"19",X"00",X"01",X"05",X"09",X"0D",X"03",
		X"00",X"00",X"0D",X"03",X"15",X"19",X"1D",X"00",X"05",X"09",X"0D",X"03",X"15",X"00",X"00",X"03",
		X"15",X"19",X"1D",X"02",X"00",X"0A",X"0E",X"03",X"15",X"19",X"00",X"00",X"15",X"19",X"1D",X"01",
		X"05",X"00",X"0D",X"03",X"15",X"19",X"1D",X"00",X"00",X"19",X"1D",X"01",X"05",X"09",X"00",X"03",
		X"15",X"19",X"1D",X"02",X"00",X"E7",X"AF",X"32",X"36",X"C4",X"21",X"00",X"20",X"01",X"00",X"10",
		X"3A",X"36",X"C4",X"86",X"32",X"36",X"C4",X"23",X"0B",X"78",X"B1",X"20",X"F3",X"3A",X"36",X"C4",
		X"21",X"46",X"35",X"BE",X"28",X"08",X"32",X"75",X"EE",X"32",X"6C",X"C6",X"ED",X"5E",X"AF",X"32",
		X"74",X"C4",X"32",X"C4",X"C4",X"21",X"FE",X"C4",X"06",X"09",X"77",X"23",X"10",X"FC",X"3E",X"01",
		X"32",X"D5",X"C4",X"CD",X"82",X"54",X"CD",X"2F",X"21",X"21",X"63",X"C4",X"11",X"64",X"C4",X"01",
		X"0A",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"72",X"ED",X"FE",X"20",X"32",X"83",X"ED",X"28",X"2F",
		X"E7",X"21",X"83",X"06",X"11",X"6E",X"07",X"06",X"20",X"1A",X"BE",X"20",X"06",X"23",X"13",X"10",
		X"F8",X"18",X"08",X"3E",X"EE",X"CD",X"AE",X"67",X"32",X"CE",X"C4",X"3A",X"7B",X"C4",X"CB",X"B7",
		X"32",X"7B",X"C4",X"3A",X"72",X"ED",X"E6",X"03",X"CD",X"75",X"55",X"E7",X"CD",X"70",X"22",X"CD",
		X"4E",X"21",X"3E",X"48",X"32",X"39",X"C4",X"DD",X"21",X"6B",X"C4",X"DD",X"36",X"00",X"01",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"21",X"3D",X"C4",X"DD",X"36",X"03",X"04",X"DD",
		X"36",X"04",X"01",X"DD",X"36",X"10",X"01",X"DD",X"36",X"1C",X"01",X"3A",X"72",X"ED",X"FE",X"20",
		X"28",X"54",X"3A",X"66",X"EF",X"A7",X"20",X"4E",X"CD",X"D0",X"21",X"3E",X"0B",X"CD",X"AE",X"67",
		X"CD",X"0E",X"28",X"06",X"1E",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",
		X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",
		X"E7",X"10",X"E6",X"CD",X"62",X"28",X"06",X"32",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",
		X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",
		X"32",X"18",X"D0",X"E7",X"10",X"E6",X"11",X"86",X"19",X"3E",X"80",X"32",X"3A",X"C4",X"47",X"3A",
		X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"78",X"86",X"E1",
		X"21",X"0D",X"D0",X"2B",X"CB",X"76",X"28",X"FC",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"21",
		X"92",X"B6",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"19",X"CD",X"D0",X"21",X"7E",X"32",X"62",
		X"C4",X"22",X"71",X"C4",X"3E",X"03",X"F7",X"3E",X"06",X"F7",X"CD",X"4A",X"0E",X"E7",X"3A",X"66",
		X"EF",X"A7",X"28",X"03",X"CD",X"2B",X"29",X"21",X"48",X"0E",X"11",X"A7",X"C4",X"01",X"02",X"00",
		X"ED",X"B0",X"21",X"A5",X"C4",X"36",X"E4",X"23",X"3A",X"3A",X"C4",X"77",X"32",X"61",X"C4",X"AF",
		X"32",X"63",X"EF",X"32",X"70",X"C4",X"32",X"73",X"C4",X"32",X"7A",X"C4",X"3E",X"78",X"32",X"48",
		X"C4",X"E7",X"3E",X"FF",X"32",X"C4",X"C4",X"E7",X"3A",X"66",X"EF",X"A7",X"20",X"06",X"3A",X"7C",
		X"C4",X"32",X"61",X"C4",X"CD",X"A8",X"0C",X"3A",X"3A",X"C4",X"DD",X"96",X"08",X"21",X"00",X"00",
		X"22",X"78",X"C4",X"22",X"76",X"C4",X"22",X"65",X"C6",X"22",X"67",X"C6",X"18",X"20",X"06",X"1E",
		X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",
		X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"E7",X"10",X"E6",X"3A",X"8A",
		X"ED",X"67",X"3A",X"75",X"EE",X"B4",X"20",X"FD",X"3A",X"C4",X"C4",X"32",X"75",X"C4",X"AF",X"32",
		X"C4",X"C4",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",
		X"3E",X"92",X"86",X"E1",X"21",X"0D",X"D0",X"2B",X"CB",X"76",X"28",X"FC",X"32",X"18",X"D0",X"CB",
		X"76",X"28",X"FC",X"3A",X"83",X"ED",X"32",X"18",X"D0",X"2A",X"74",X"ED",X"23",X"22",X"74",X"ED",
		X"3A",X"64",X"EF",X"2A",X"74",X"ED",X"11",X"00",X"07",X"ED",X"52",X"38",X"21",X"20",X"03",X"3C",
		X"18",X"1C",X"2A",X"74",X"ED",X"11",X"00",X"0E",X"ED",X"52",X"38",X"12",X"20",X"03",X"3C",X"18",
		X"0D",X"2A",X"74",X"ED",X"11",X"00",X"15",X"ED",X"52",X"38",X"03",X"20",X"01",X"3C",X"FE",X"03",
		X"38",X"02",X"3E",X"03",X"32",X"64",X"EF",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"2A",X"78",
		X"C4",X"23",X"22",X"78",X"C4",X"11",X"18",X"15",X"A7",X"ED",X"52",X"20",X"05",X"3E",X"01",X"32",
		X"CE",X"C4",X"2A",X"71",X"C4",X"7E",X"A7",X"20",X"11",X"32",X"62",X"EF",X"3E",X"03",X"CF",X"3E",
		X"06",X"CF",X"3E",X"00",X"D7",X"AF",X"DF",X"3E",X"03",X"DF",X"3A",X"62",X"EF",X"A7",X"28",X"16",
		X"3E",X"FF",X"32",X"C4",X"C4",X"CD",X"E4",X"0E",X"3A",X"86",X"ED",X"32",X"C4",X"C4",X"3E",X"00",
		X"D7",X"AF",X"DF",X"3E",X"03",X"DF",X"3A",X"75",X"C4",X"32",X"C4",X"C4",X"21",X"6A",X"C4",X"7E",
		X"2B",X"BE",X"C4",X"BF",X"09",X"FE",X"02",X"20",X"10",X"21",X"6C",X"C4",X"7E",X"23",X"B6",X"20",
		X"08",X"3E",X"00",X"32",X"69",X"C4",X"32",X"6A",X"C4",X"3A",X"37",X"C4",X"3C",X"32",X"37",X"C4",
		X"FE",X"0C",X"CC",X"16",X"0E",X"CD",X"2C",X"51",X"3A",X"6D",X"C4",X"A7",X"28",X"17",X"DD",X"21",
		X"55",X"C4",X"3A",X"62",X"C4",X"DD",X"77",X"02",X"21",X"AD",X"C4",X"CD",X"CA",X"10",X"FD",X"21",
		X"AD",X"C4",X"CD",X"C0",X"56",X"3A",X"6C",X"C4",X"A7",X"28",X"19",X"DD",X"21",X"49",X"C4",X"3A",
		X"62",X"C4",X"DD",X"77",X"02",X"21",X"A9",X"C4",X"CD",X"CA",X"10",X"FD",X"21",X"A9",X"C4",X"CD",
		X"C0",X"56",X"18",X"2C",X"3A",X"6D",X"C4",X"A7",X"28",X"26",X"21",X"AD",X"C4",X"11",X"A9",X"C4",
		X"01",X"04",X"00",X"ED",X"B0",X"21",X"AD",X"C4",X"CD",X"2F",X"0B",X"21",X"55",X"C4",X"11",X"49",
		X"C4",X"01",X"0C",X"00",X"ED",X"B0",X"3A",X"6D",X"C4",X"32",X"6C",X"C4",X"AF",X"32",X"6D",X"C4",
		X"3A",X"6B",X"C4",X"A7",X"28",X"75",X"DD",X"21",X"3D",X"C4",X"3A",X"62",X"C4",X"DD",X"77",X"02",
		X"3A",X"62",X"C4",X"21",X"4C",X"09",X"CD",X"50",X"20",X"3A",X"63",X"EF",X"BE",X"38",X"4D",X"DD",
		X"7E",X"03",X"FE",X"08",X"38",X"04",X"FE",X"18",X"38",X"42",X"AF",X"32",X"63",X"EF",X"3A",X"62",
		X"C4",X"FE",X"0E",X"30",X"04",X"3C",X"32",X"62",X"C4",X"DD",X"7E",X"03",X"E6",X"07",X"CB",X"57",
		X"28",X"03",X"3D",X"18",X"01",X"3C",X"47",X"DD",X"7E",X"03",X"E6",X"18",X"B0",X"DD",X"77",X"03",
		X"18",X"1A",X"09",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"00",X"19",X"19",X"23",
		X"23",X"2D",X"3C",X"50",X"78",X"8C",X"A0",X"B4",X"C8",X"DC",X"F0",X"FF",X"21",X"A5",X"C4",X"CD",
		X"CA",X"10",X"FD",X"21",X"A5",X"C4",X"CD",X"C0",X"56",X"18",X"2C",X"3A",X"6C",X"C4",X"A7",X"28",
		X"26",X"21",X"A9",X"C4",X"11",X"A5",X"C4",X"01",X"04",X"00",X"ED",X"B0",X"21",X"49",X"C4",X"11",
		X"3D",X"C4",X"01",X"0C",X"00",X"ED",X"B0",X"21",X"A9",X"C4",X"CD",X"2F",X"0B",X"3A",X"6C",X"C4",
		X"32",X"6B",X"C4",X"AF",X"32",X"6C",X"C4",X"CD",X"34",X"0B",X"CD",X"6A",X"0A",X"CD",X"A8",X"0C",
		X"E7",X"C3",X"8E",X"07",X"2A",X"88",X"ED",X"06",X"EA",X"3A",X"6A",X"C6",X"BE",X"20",X"05",X"23",
		X"10",X"FA",X"A7",X"C9",X"3D",X"BE",X"20",X"05",X"3A",X"6C",X"C6",X"18",X"F2",X"37",X"C9",X"FE",
		X"02",X"C8",X"F5",X"3A",X"69",X"C4",X"32",X"6A",X"C4",X"FE",X"02",X"28",X"4C",X"FE",X"01",X"28",
		X"1F",X"3E",X"01",X"32",X"41",X"C4",X"21",X"48",X"0E",X"11",X"A7",X"C4",X"ED",X"A0",X"ED",X"A0",
		X"21",X"A9",X"C4",X"11",X"AA",X"C4",X"01",X"07",X"00",X"36",X"00",X"ED",X"B0",X"C3",X"68",X"0A",
		X"3E",X"02",X"32",X"41",X"C4",X"21",X"A5",X"C4",X"11",X"A9",X"C4",X"7E",X"C6",X"08",X"12",X"23",
		X"13",X"ED",X"A0",X"D9",X"21",X"90",X"1B",X"CD",X"BA",X"20",X"3E",X"A8",X"B4",X"D9",X"77",X"D9",
		X"7D",X"D9",X"ED",X"A0",X"77",X"3C",X"12",X"18",X"4F",X"21",X"48",X"0E",X"11",X"A7",X"C4",X"ED",
		X"A0",X"ED",X"A0",X"DD",X"21",X"3D",X"C4",X"DD",X"36",X"04",X"01",X"21",X"3D",X"C4",X"11",X"49",
		X"C4",X"01",X"18",X"00",X"ED",X"B0",X"DD",X"7E",X"03",X"47",X"3D",X"4F",X"E6",X"07",X"20",X"02",
		X"0C",X"0C",X"DD",X"71",X"0F",X"78",X"3C",X"4F",X"E6",X"07",X"20",X"02",X"0D",X"0D",X"DD",X"71",
		X"1B",X"21",X"A5",X"C4",X"11",X"A9",X"C4",X"01",X"08",X"00",X"ED",X"B0",X"DD",X"21",X"6B",X"C4",
		X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"01",X"F1",X"C9",X"3A",X"6B",X"C4",X"A7",X"28",X"10",
		X"3A",X"A5",X"C4",X"FE",X"F8",X"38",X"09",X"21",X"A5",X"C4",X"CD",X"2F",X"0B",X"32",X"6B",X"C4",
		X"3A",X"6C",X"C4",X"A7",X"28",X"10",X"3A",X"A9",X"C4",X"FE",X"F8",X"38",X"09",X"21",X"A9",X"C4",
		X"CD",X"2F",X"0B",X"32",X"6C",X"C4",X"3A",X"6D",X"C4",X"A7",X"28",X"10",X"3A",X"AD",X"C4",X"FE",
		X"F8",X"38",X"09",X"21",X"AD",X"C4",X"CD",X"2F",X"0B",X"32",X"6D",X"C4",X"21",X"6B",X"C4",X"06",
		X"03",X"AF",X"BE",X"20",X"09",X"23",X"10",X"FA",X"3E",X"FF",X"32",X"62",X"EF",X"C9",X"21",X"FE",
		X"C4",X"CB",X"46",X"28",X"1E",X"23",X"23",X"7E",X"FE",X"D9",X"38",X"17",X"FE",X"F0",X"30",X"13",
		X"2B",X"3A",X"3A",X"C4",X"D6",X"20",X"BE",X"30",X"0A",X"C6",X"20",X"BE",X"38",X"05",X"2B",X"CB",
		X"E6",X"CB",X"F6",X"21",X"01",X"C5",X"CB",X"46",X"28",X"1E",X"23",X"23",X"7E",X"FE",X"D9",X"38",
		X"17",X"FE",X"F0",X"30",X"13",X"2B",X"3A",X"3A",X"C4",X"D6",X"20",X"BE",X"30",X"0A",X"C6",X"20",
		X"BE",X"38",X"05",X"2B",X"CB",X"E6",X"CB",X"F6",X"21",X"04",X"C5",X"CB",X"46",X"28",X"1E",X"23",
		X"23",X"7E",X"FE",X"D9",X"38",X"17",X"FE",X"F0",X"30",X"13",X"2B",X"3A",X"3A",X"C4",X"D6",X"20",
		X"BE",X"30",X"0A",X"C6",X"20",X"BE",X"38",X"05",X"2B",X"CB",X"E6",X"CB",X"F6",X"A7",X"C9",X"AF",
		X"77",X"23",X"77",X"C9",X"DD",X"21",X"B1",X"C4",X"21",X"63",X"C4",X"CB",X"7E",X"20",X"5C",X"3A",
		X"65",X"C4",X"BE",X"20",X"20",X"C5",X"3A",X"39",X"C4",X"47",X"DD",X"7E",X"02",X"E6",X"07",X"B0",
		X"DD",X"77",X"02",X"DD",X"77",X"06",X"47",X"3A",X"65",X"C4",X"FE",X"02",X"20",X"03",X"DD",X"70",
		X"0A",X"C1",X"C3",X"82",X"0C",X"A7",X"20",X"14",X"7E",X"32",X"64",X"C4",X"FE",X"02",X"20",X"07",
		X"F5",X"3E",X"09",X"CD",X"AE",X"67",X"F1",X"CB",X"FF",X"77",X"18",X"08",X"CB",X"FE",X"3A",X"8A",
		X"ED",X"32",X"64",X"C4",X"CD",X"91",X"0C",X"11",X"83",X"0C",X"CD",X"4A",X"20",X"1A",X"32",X"66",
		X"C4",X"32",X"68",X"C4",X"AF",X"32",X"67",X"C4",X"C3",X"82",X"0C",X"3A",X"68",X"C4",X"A7",X"28",
		X"07",X"3D",X"32",X"68",X"C4",X"C3",X"82",X"0C",X"3A",X"66",X"C4",X"32",X"68",X"C4",X"CD",X"91",
		X"0C",X"CB",X"27",X"21",X"87",X"0C",X"CD",X"56",X"20",X"EB",X"E9",X"21",X"20",X"0F",X"CD",X"BA",
		X"20",X"3A",X"64",X"C4",X"A7",X"3A",X"67",X"C4",X"20",X"04",X"47",X"3E",X"09",X"90",X"CB",X"27",
		X"0E",X"48",X"FE",X"0E",X"20",X"02",X"0E",X"60",X"CD",X"50",X"20",X"7C",X"B1",X"67",X"3A",X"67",
		X"C4",X"3C",X"32",X"67",X"C4",X"FE",X"0A",X"20",X"03",X"CD",X"9A",X"0C",X"DD",X"75",X"03",X"DD",
		X"74",X"02",X"23",X"DD",X"75",X"07",X"DD",X"74",X"06",X"C3",X"82",X"0C",X"DD",X"21",X"B1",X"C4",
		X"21",X"D0",X"0B",X"CD",X"BA",X"20",X"23",X"3E",X"48",X"B4",X"DD",X"77",X"0A",X"DD",X"75",X"0B",
		X"3A",X"64",X"C4",X"A7",X"3A",X"67",X"C4",X"20",X"1A",X"FE",X"07",X"20",X"0D",X"AF",X"DD",X"77",
		X"09",X"DD",X"77",X"08",X"32",X"86",X"C4",X"32",X"85",X"C4",X"DD",X"35",X"01",X"DD",X"34",X"05",
		X"C3",X"6E",X"0C",X"A7",X"20",X"0C",X"DD",X"7E",X"01",X"D6",X"08",X"DD",X"77",X"09",X"DD",X"36",
		X"08",X"E8",X"DD",X"34",X"01",X"DD",X"35",X"05",X"DD",X"7E",X"01",X"FE",X"D9",X"30",X"09",X"DD",
		X"7E",X"05",X"FE",X"16",X"38",X"0D",X"18",X"16",X"DD",X"35",X"01",X"DD",X"35",X"05",X"DD",X"35",
		X"09",X"18",X"0B",X"DD",X"34",X"01",X"DD",X"34",X"05",X"DD",X"34",X"09",X"18",X"00",X"3A",X"67",
		X"C4",X"3C",X"32",X"67",X"C4",X"FE",X"08",X"20",X"09",X"CD",X"9A",X"0C",X"C3",X"82",X"0C",X"CD",
		X"9A",X"0C",X"C9",X"00",X"03",X"01",X"00",X"00",X"00",X"BB",X"0B",X"FC",X"0B",X"7F",X"0C",X"00",
		X"00",X"3A",X"64",X"C4",X"47",X"3A",X"65",X"C4",X"B0",X"C9",X"3A",X"64",X"C4",X"32",X"65",X"C4",
		X"3A",X"63",X"C4",X"CB",X"BF",X"32",X"63",X"C4",X"DD",X"21",X"B1",X"C4",X"E5",X"21",X"61",X"C4",
		X"3A",X"66",X"EF",X"A7",X"28",X"05",X"3A",X"A6",X"C4",X"18",X"03",X"3A",X"7C",X"C4",X"47",X"96",
		X"70",X"47",X"DD",X"7E",X"01",X"80",X"30",X"15",X"CB",X"78",X"28",X"1B",X"DD",X"7E",X"05",X"80",
		X"FE",X"16",X"DA",X"B7",X"0D",X"FE",X"D9",X"D2",X"B7",X"0D",X"C3",X"E0",X"0D",X"CB",X"78",X"C2",
		X"B7",X"0D",X"FE",X"D9",X"DA",X"E0",X"0D",X"3E",X"D9",X"DD",X"96",X"01",X"47",X"DD",X"36",X"01",
		X"D9",X"DD",X"86",X"05",X"DD",X"77",X"05",X"3A",X"65",X"C4",X"FE",X"02",X"28",X"09",X"3A",X"63",
		X"C4",X"E6",X"0F",X"FE",X"02",X"20",X"07",X"78",X"DD",X"86",X"09",X"DD",X"77",X"09",X"3A",X"CE",
		X"C4",X"A7",X"CA",X"05",X"0E",X"3E",X"18",X"CD",X"AE",X"67",X"3E",X"03",X"CF",X"21",X"89",X"C4",
		X"11",X"8A",X"C4",X"01",X"27",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"65",X"C4",X"E6",X"0F",X"FE",
		X"02",X"28",X"15",X"3A",X"63",X"C4",X"E6",X"0F",X"FE",X"02",X"28",X"0C",X"21",X"B9",X"C4",X"CD",
		X"34",X"0E",X"21",X"85",X"C4",X"CD",X"34",X"0E",X"DD",X"21",X"6B",X"C4",X"DD",X"36",X"00",X"00",
		X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"21",X"B1",X"C4",X"DD",X"7E",X"01",X"FE",
		X"F8",X"28",X"03",X"DD",X"34",X"01",X"DD",X"7E",X"05",X"FE",X"F8",X"28",X"03",X"DD",X"34",X"05",
		X"3A",X"65",X"C4",X"E6",X"0F",X"FE",X"02",X"28",X"09",X"3A",X"63",X"C4",X"E6",X"0F",X"FE",X"02",
		X"20",X"0A",X"DD",X"7E",X"09",X"FE",X"F8",X"28",X"03",X"DD",X"34",X"09",X"E1",X"E5",X"CD",X"AB",
		X"0E",X"E7",X"DD",X"7E",X"01",X"FE",X"F8",X"20",X"C3",X"DD",X"7E",X"05",X"FE",X"F8",X"20",X"BC",
		X"E1",X"06",X"64",X"11",X"10",X"00",X"CD",X"23",X"27",X"E7",X"10",X"F7",X"AF",X"32",X"83",X"ED",
		X"32",X"62",X"EF",X"32",X"CE",X"C4",X"C9",X"3E",X"16",X"DD",X"96",X"05",X"47",X"DD",X"36",X"05",
		X"16",X"DD",X"86",X"01",X"DD",X"77",X"01",X"3A",X"65",X"C4",X"FE",X"02",X"28",X"09",X"3A",X"63",
		X"C4",X"E6",X"0F",X"FE",X"02",X"20",X"2E",X"78",X"DD",X"86",X"09",X"DD",X"77",X"09",X"18",X"25",
		X"78",X"DD",X"86",X"01",X"DD",X"77",X"01",X"78",X"DD",X"86",X"05",X"DD",X"77",X"05",X"3A",X"65",
		X"C4",X"FE",X"02",X"28",X"09",X"3A",X"63",X"C4",X"E6",X"0F",X"FE",X"02",X"20",X"07",X"78",X"DD",
		X"86",X"09",X"DD",X"77",X"09",X"E1",X"CD",X"AB",X"0E",X"DD",X"7E",X"01",X"32",X"3A",X"C4",X"DD",
		X"7E",X"05",X"32",X"3B",X"C4",X"C9",X"AF",X"32",X"37",X"C4",X"3A",X"38",X"C4",X"3C",X"32",X"38",
		X"C4",X"FE",X"06",X"20",X"04",X"AF",X"32",X"38",X"C4",X"21",X"40",X"0E",X"CD",X"50",X"20",X"7E",
		X"32",X"39",X"C4",X"C9",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"C9",
		X"48",X"50",X"58",X"60",X"58",X"50",X"E0",X"80",X"61",X"B8",X"06",X"06",X"78",X"FE",X"02",X"CC",
		X"AB",X"0E",X"21",X"6F",X"0E",X"78",X"3D",X"CB",X"27",X"CD",X"56",X"20",X"EB",X"11",X"7B",X"0E",
		X"78",X"3D",X"CD",X"4A",X"20",X"1A",X"CD",X"81",X"0E",X"3E",X"05",X"DF",X"10",X"DE",X"C9",X"20",
		X"0F",X"00",X"0F",X"E0",X"0E",X"C0",X"0E",X"A0",X"0E",X"80",X"0E",X"50",X"50",X"58",X"60",X"48",
		X"48",X"CD",X"BA",X"20",X"DD",X"21",X"B1",X"C4",X"DD",X"75",X"03",X"B4",X"67",X"DD",X"74",X"02",
		X"23",X"DD",X"75",X"07",X"DD",X"74",X"06",X"3E",X"E8",X"DD",X"77",X"00",X"DD",X"77",X"04",X"3A",
		X"3A",X"C4",X"DD",X"77",X"01",X"D6",X"10",X"DD",X"77",X"05",X"C9",X"E5",X"D5",X"C5",X"21",X"B1",
		X"C4",X"11",X"7D",X"C4",X"06",X"02",X"3A",X"65",X"C4",X"FE",X"02",X"28",X"09",X"3A",X"63",X"C4",
		X"E6",X"0F",X"FE",X"02",X"20",X"01",X"04",X"7E",X"C6",X"04",X"12",X"13",X"23",X"7E",X"C6",X"04",
		X"12",X"13",X"23",X"7E",X"E6",X"07",X"F6",X"40",X"12",X"13",X"23",X"ED",X"A0",X"03",X"10",X"E7",
		X"C1",X"D1",X"E1",X"C9",X"3E",X"1A",X"CD",X"AE",X"67",X"21",X"7D",X"C4",X"11",X"7E",X"C4",X"01",
		X"3F",X"00",X"36",X"00",X"ED",X"B0",X"21",X"20",X"0F",X"3E",X"50",X"CD",X"81",X"0E",X"CD",X"AB",
		X"0E",X"3E",X"03",X"CF",X"3E",X"0A",X"DF",X"21",X"60",X"10",X"3E",X"48",X"CD",X"81",X"0E",X"3E",
		X"05",X"DF",X"21",X"80",X"10",X"3E",X"60",X"CD",X"81",X"0E",X"3E",X"0A",X"DF",X"21",X"B1",X"C4",
		X"11",X"B2",X"C4",X"01",X"0B",X"00",X"36",X"00",X"ED",X"B0",X"21",X"7D",X"C4",X"11",X"7E",X"C4",
		X"01",X"07",X"00",X"36",X"00",X"ED",X"B0",X"3E",X"00",X"32",X"38",X"C4",X"21",X"A0",X"10",X"CD",
		X"BA",X"20",X"4D",X"7C",X"32",X"6E",X"C4",X"21",X"A3",X"0F",X"3A",X"38",X"C4",X"CB",X"27",X"CD",
		X"56",X"20",X"1A",X"47",X"21",X"7D",X"C4",X"CD",X"83",X"0F",X"21",X"AB",X"0F",X"3A",X"38",X"C4",
		X"CD",X"50",X"20",X"46",X"E7",X"10",X"FD",X"3A",X"38",X"C4",X"3C",X"32",X"38",X"C4",X"FE",X"04",
		X"20",X"D5",X"21",X"7D",X"C4",X"11",X"7E",X"C4",X"01",X"40",X"00",X"36",X"00",X"ED",X"B0",X"3E",
		X"3C",X"DF",X"C9",X"C5",X"13",X"1A",X"4F",X"13",X"1A",X"C6",X"E8",X"77",X"23",X"79",X"47",X"3A",
		X"3A",X"C4",X"80",X"77",X"23",X"3A",X"6E",X"C4",X"F6",X"48",X"77",X"23",X"C1",X"71",X"23",X"0C",
		X"10",X"E1",X"C9",X"AF",X"0F",X"BC",X"0F",X"BC",X"0F",X"CF",X"0F",X"06",X"08",X"0A",X"0C",X"06",
		X"F0",X"F8",X"F0",X"00",X"F0",X"08",X"00",X"F8",X"00",X"00",X"00",X"08",X"09",X"E8",X"F8",X"E8",
		X"00",X"E8",X"08",X"F8",X"F8",X"F8",X"00",X"F8",X"08",X"08",X"F8",X"08",X"00",X"08",X"08",X"08",
		X"E8",X"F8",X"E8",X"00",X"E8",X"08",X"F8",X"F8",X"F8",X"08",X"08",X"F8",X"08",X"00",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"00",
		X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"12",X"03",X"03",X"03",
		X"12",X"03",X"03",X"00",X"00",X"00",X"00",X"03",X"03",X"12",X"03",X"03",X"03",X"12",X"03",X"03",
		X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"03",X"00",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"E5",X"DD",X"7E",X"03",X"E6",X"0F",
		X"FE",X"06",X"38",X"12",X"FE",X"0B",X"30",X"0E",X"DD",X"7E",X"02",X"C6",X"02",X"FE",X"0F",X"38",
		X"02",X"3E",X"0E",X"DD",X"77",X"02",X"DD",X"7E",X"0B",X"A7",X"28",X"56",X"DD",X"35",X"0B",X"20",
		X"05",X"3E",X"03",X"CD",X"AE",X"67",X"E5",X"3A",X"7A",X"C4",X"47",X"3A",X"3A",X"C4",X"90",X"23",
		X"77",X"2B",X"E1",X"3A",X"6F",X"ED",X"CB",X"4F",X"28",X"1B",X"3A",X"FF",X"BF",X"FE",X"76",X"20",
		X"14",X"3A",X"C1",X"C4",X"CB",X"7F",X"28",X"0D",X"3A",X"C0",X"C4",X"CB",X"57",X"20",X"1F",X"CB",
		X"D7",X"CB",X"87",X"18",X"0B",X"3A",X"C0",X"C4",X"CB",X"47",X"20",X"12",X"CB",X"C7",X"CB",X"97",
		X"32",X"C0",X"C4",X"AF",X"DD",X"77",X"0B",X"3E",X"03",X"CD",X"AE",X"67",X"18",X"04",X"AF",X"DD",
		X"77",X"02",X"CD",X"4A",X"11",X"CD",X"7E",X"12",X"E1",X"C9",X"E5",X"DD",X"7E",X"03",X"D5",X"E5",
		X"DD",X"E5",X"D1",X"CD",X"4F",X"12",X"E1",X"D1",X"DD",X"7E",X"01",X"CD",X"BF",X"11",X"DD",X"CB",
		X"00",X"4E",X"28",X"02",X"2F",X"3C",X"23",X"F5",X"86",X"DD",X"77",X"08",X"F1",X"CD",X"AD",X"11",
		X"DD",X"7E",X"01",X"0F",X"0F",X"0F",X"0F",X"CD",X"BF",X"11",X"DD",X"CB",X"00",X"46",X"28",X"02",
		X"2F",X"3C",X"2B",X"F5",X"86",X"DD",X"77",X"07",X"F1",X"CD",X"AD",X"11",X"DD",X"34",X"05",X"3E",
		X"01",X"DD",X"BE",X"02",X"20",X"06",X"DD",X"CB",X"05",X"46",X"28",X"0F",X"DD",X"7E",X"06",X"47",
		X"3C",X"E6",X"0F",X"4F",X"78",X"E6",X"F0",X"B1",X"DD",X"77",X"06",X"E1",X"C9",X"D5",X"E5",X"11",
		X"04",X"00",X"DD",X"46",X"04",X"4F",X"79",X"86",X"77",X"19",X"10",X"FA",X"E1",X"D1",X"C9",X"E6",
		X"0F",X"28",X"5E",X"FE",X"01",X"20",X"05",X"11",X"27",X"12",X"18",X"15",X"FE",X"05",X"20",X"05",
		X"11",X"31",X"12",X"18",X"0C",X"FE",X"07",X"20",X"05",X"11",X"3B",X"12",X"18",X"03",X"11",X"45",
		X"12",X"DD",X"7E",X"02",X"CB",X"3F",X"30",X"07",X"DD",X"CB",X"05",X"46",X"28",X"01",X"3C",X"A7",
		X"28",X"2F",X"D5",X"4F",X"3D",X"E6",X"03",X"CB",X"3F",X"28",X"01",X"13",X"1A",X"38",X"04",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"47",X"D1",X"79",X"3C",X"CD",X"4A",X"20",X"1A",X"81",X"4F",X"DD",
		X"7E",X"06",X"E6",X"03",X"11",X"23",X"12",X"CD",X"4A",X"20",X"1A",X"A0",X"79",X"20",X"01",X"3D",
		X"C9",X"AF",X"C9",X"01",X"02",X"04",X"08",X"15",X"7F",X"00",X"FF",X"FE",X"FD",X"FD",X"FC",X"FB",
		X"FA",X"5F",X"5F",X"00",X"FF",X"FF",X"FE",X"FE",X"FD",X"FD",X"FC",X"75",X"1F",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"7A",X"12",X"CD",X"50",X"20",X"ED",X"A0",X"F1",X"E6",
		X"0F",X"21",X"6A",X"12",X"CD",X"50",X"20",X"ED",X"A0",X"C9",X"F0",X"F1",X"F5",X"F7",X"FF",X"7F",
		X"5F",X"1F",X"0F",X"1F",X"5F",X"7F",X"FF",X"F7",X"F5",X"F1",X"01",X"00",X"02",X"03",X"E5",X"CD",
		X"18",X"13",X"E1",X"CD",X"87",X"12",X"C9",X"FD",X"21",X"FE",X"C4",X"FD",X"7E",X"00",X"CB",X"47",
		X"28",X"10",X"CB",X"67",X"20",X"0C",X"FD",X"56",X"01",X"FD",X"5E",X"02",X"CD",X"D1",X"12",X"FD",
		X"77",X"00",X"FD",X"7E",X"03",X"CB",X"47",X"28",X"10",X"CB",X"67",X"20",X"0C",X"FD",X"56",X"04",
		X"FD",X"5E",X"05",X"CD",X"D1",X"12",X"FD",X"77",X"03",X"FD",X"7E",X"06",X"CB",X"47",X"28",X"10",
		X"CB",X"67",X"20",X"0C",X"FD",X"56",X"07",X"FD",X"5E",X"08",X"CD",X"D1",X"12",X"FD",X"77",X"06",
		X"C9",X"E5",X"F5",X"23",X"7E",X"D6",X"12",X"BA",X"30",X"3B",X"C6",X"0E",X"BA",X"38",X"36",X"2B",
		X"7E",X"D6",X"08",X"BB",X"30",X"2F",X"C6",X"0C",X"BB",X"38",X"2A",X"D6",X"03",X"BB",X"38",X"14",
		X"D6",X"06",X"BB",X"30",X"0F",X"CD",X"BA",X"14",X"CB",X"67",X"20",X"04",X"CB",X"DF",X"18",X"07",
		X"CB",X"9F",X"18",X"03",X"CD",X"BA",X"14",X"DD",X"77",X"03",X"DD",X"CB",X"06",X"BE",X"F1",X"CB",
		X"E7",X"CB",X"EF",X"E1",X"C9",X"F1",X"E1",X"C9",X"7E",X"23",X"DD",X"CB",X"06",X"7E",X"C2",X"1B",
		X"14",X"FE",X"E4",X"DA",X"1B",X"14",X"FE",X"EC",X"D2",X"1B",X"14",X"3A",X"3A",X"C4",X"C6",X"0C",
		X"96",X"DA",X"1B",X"14",X"47",X"3A",X"3B",X"C4",X"D6",X"04",X"96",X"D2",X"1B",X"14",X"2F",X"3C",
		X"B8",X"38",X"08",X"11",X"15",X"14",X"0E",X"01",X"78",X"18",X"05",X"11",X"0F",X"14",X"0E",X"00",
		X"E5",X"06",X"03",X"21",X"0C",X"14",X"BE",X"38",X"05",X"23",X"10",X"FA",X"18",X"FE",X"3A",X"73",
		X"C4",X"A7",X"28",X"05",X"3E",X"03",X"CD",X"AE",X"67",X"ED",X"5F",X"F6",X"80",X"32",X"73",X"C4",
		X"78",X"3D",X"CB",X"27",X"EB",X"CD",X"56",X"20",X"DD",X"CB",X"06",X"FE",X"21",X"00",X"00",X"22",
		X"78",X"C4",X"2A",X"76",X"C4",X"23",X"22",X"76",X"C4",X"18",X"0F",X"7C",X"A7",X"20",X"0B",X"7D",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"04",X"38",X"02",X"3E",X"04",X"CD",X"4A",X"20",X"1A",
		X"DD",X"77",X"03",X"21",X"61",X"C4",X"3A",X"7C",X"C4",X"96",X"CB",X"7F",X"47",X"28",X"01",X"2F",
		X"FE",X"10",X"E1",X"38",X"0C",X"CB",X"78",X"20",X"05",X"34",X"34",X"34",X"18",X"03",X"35",X"35",
		X"35",X"3A",X"59",X"C6",X"FE",X"03",X"C0",X"DD",X"7E",X"0B",X"A7",X"C0",X"3E",X"78",X"DD",X"77",
		X"0B",X"3A",X"3A",X"C4",X"96",X"32",X"7A",X"C4",X"3E",X"19",X"CD",X"AE",X"67",X"AF",X"B9",X"28",
		X"05",X"35",X"35",X"35",X"18",X"03",X"34",X"34",X"34",X"2B",X"36",X"E4",X"23",X"C9",X"1C",X"19",
		X"1F",X"1B",X"1A",X"1C",X"19",X"1F",X"1B",X"1B",X"1E",X"19",X"1F",X"1D",X"1E",X"02",X"07",X"01",
		X"03",X"02",X"04",X"07",X"01",X"05",X"05",X"04",X"07",X"01",X"05",X"06",X"03",X"08",X"1E",X"F8",
		X"13",X"F3",X"13",X"EE",X"13",X"FD",X"13",X"02",X"14",X"07",X"14",X"56",X"2B",X"5E",X"3E",X"1C",
		X"BA",X"38",X"0D",X"DD",X"CB",X"03",X"66",X"28",X"19",X"CD",X"BA",X"14",X"CB",X"A7",X"18",X"77",
		X"3E",X"E0",X"BA",X"30",X"0D",X"DD",X"CB",X"03",X"66",X"20",X"07",X"CD",X"BA",X"14",X"CB",X"E7",
		X"18",X"65",X"3E",X"1C",X"BB",X"38",X"72",X"3A",X"70",X"C4",X"A7",X"20",X"37",X"21",X"62",X"14",
		X"3A",X"72",X"ED",X"CD",X"50",X"20",X"3A",X"62",X"C4",X"BE",X"30",X"28",X"7E",X"32",X"62",X"C4",
		X"18",X"22",X"07",X"07",X"08",X"00",X"07",X"07",X"07",X"00",X"07",X"05",X"07",X"07",X"08",X"06",
		X"07",X"05",X"07",X"07",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"07",X"08",X"07",X"00",X"07",
		X"00",X"00",X"00",X"00",X"DD",X"7E",X"03",X"E6",X"18",X"28",X"04",X"FE",X"18",X"20",X"2A",X"CD",
		X"BA",X"14",X"CB",X"67",X"20",X"06",X"CB",X"DF",X"CB",X"A7",X"18",X"0B",X"CB",X"9F",X"18",X"07",
		X"3E",X"F0",X"BB",X"30",X"14",X"18",X"12",X"DD",X"77",X"03",X"DD",X"CB",X"06",X"BE",X"3A",X"63",
		X"EF",X"3C",X"32",X"63",X"EF",X"DD",X"36",X"0B",X"00",X"C9",X"DD",X"7E",X"03",X"4F",X"2F",X"3C",
		X"E6",X"07",X"47",X"79",X"E6",X"18",X"B0",X"CB",X"5F",X"20",X"04",X"CB",X"DF",X"18",X"02",X"CB",
		X"9F",X"C9",X"C9",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"00",X"11",X"00",X"0D",X"00",X"09",X"00",
		X"0D",X"00",X"11",X"00",X"15",X"16",X"00",X"12",X"00",X"0E",X"00",X"0A",X"00",X"0E",X"00",X"12",
		X"00",X"16",X"15",X"00",X"11",X"00",X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"15",X"15",
		X"00",X"11",X"00",X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"15",X"15",X"00",X"11",X"00",
		X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"15",X"16",X"00",X"FF",X"06",X"FF",X"06",X"FF",
		X"06",X"FF",X"06",X"FF",X"00",X"16",X"15",X"00",X"11",X"00",X"0D",X"00",X"0A",X"00",X"0D",X"00",
		X"12",X"00",X"15",X"15",X"00",X"11",X"00",X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"16",
		X"15",X"00",X"11",X"00",X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"15",X"15",X"00",X"11",
		X"00",X"0D",X"00",X"09",X"00",X"0D",X"00",X"11",X"00",X"15",X"06",X"00",X"06",X"00",X"FF",X"00",
		X"06",X"00",X"FF",X"00",X"06",X"00",X"06",X"15",X"00",X"11",X"00",X"0D",X"00",X"09",X"00",X"0D",
		X"00",X"11",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"C4",
		X"C4",X"A7",X"CA",X"3C",X"16",X"21",X"0C",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"BE",X"C4",X"C6",
		X"16",X"47",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",
		X"78",X"86",X"E1",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"7C",X"C4",X"32",X"18",X"D0",
		X"CB",X"76",X"28",X"FC",X"CB",X"7E",X"20",X"FC",X"11",X"7C",X"C4",X"1A",X"32",X"C6",X"C4",X"3A",
		X"BE",X"C4",X"CD",X"4A",X"20",X"E5",X"D5",X"21",X"7D",X"C4",X"11",X"00",X"E8",X"01",X"40",X"00",
		X"ED",X"B0",X"D1",X"E1",X"3A",X"18",X"D0",X"12",X"E5",X"21",X"C6",X"C4",X"96",X"32",X"C5",X"C4",
		X"E1",X"CB",X"7E",X"20",X"FC",X"3E",X"0E",X"32",X"00",X"D0",X"3A",X"01",X"D0",X"32",X"BD",X"C4",
		X"D5",X"CD",X"4A",X"20",X"E1",X"3A",X"18",X"D0",X"86",X"77",X"18",X"16",X"21",X"7D",X"C4",X"11",
		X"00",X"E8",X"01",X"40",X"00",X"ED",X"B0",X"3E",X"0E",X"32",X"00",X"D0",X"3A",X"01",X"D0",X"32",
		X"BD",X"C4",X"3A",X"66",X"EF",X"A7",X"3E",X"FF",X"20",X"0A",X"3A",X"BF",X"C4",X"47",X"3A",X"10",
		X"D0",X"B8",X"28",X"06",X"32",X"BF",X"C4",X"32",X"C0",X"C4",X"3A",X"7B",X"C4",X"32",X"08",X"D0",
		X"21",X"BE",X"15",X"11",X"95",X"16",X"01",X"28",X"00",X"1A",X"ED",X"A1",X"20",X"07",X"13",X"78",
		X"B1",X"20",X"F6",X"18",X"0F",X"ED",X"5F",X"32",X"71",X"ED",X"32",X"BE",X"C4",X"32",X"18",X"D0",
		X"3E",X"ED",X"ED",X"47",X"C9",X"3A",X"C4",X"C4",X"A7",X"CA",X"3C",X"16",X"21",X"0C",X"D0",X"CB",
		X"76",X"28",X"FC",X"3A",X"BE",X"C4",X"C6",X"16",X"47",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",
		X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"78",X"86",X"E1",X"32",X"18",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"1D",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1D",X"1D",X"19",X"19",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"1D",
		X"19",X"19",X"15",X"15",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"19",X"19",X"15",X"15",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"1D",X"19",X"1A",X"15",X"16",X"11",X"12",X"0D",X"0D",
		X"00",X"00",X"00",X"00",X"19",X"19",X"15",X"15",X"11",X"11",X"0D",X"0D",X"09",X"00",X"00",X"00",
		X"00",X"19",X"15",X"15",X"11",X"12",X"0D",X"0D",X"09",X"09",X"00",X"00",X"00",X"00",X"15",X"15",
		X"11",X"11",X"0D",X"0D",X"09",X"09",X"05",X"00",X"00",X"00",X"00",X"15",X"11",X"11",X"0D",X"0E",
		X"09",X"09",X"05",X"05",X"00",X"00",X"00",X"00",X"11",X"11",X"0E",X"0D",X"0A",X"09",X"06",X"05",
		X"01",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"09",X"09",X"05",X"05",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"09",X"09",X"05",X"05",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"05",X"05",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"21",X"AD",X"17",X"C3",X"D3",X"2D",X"3E",X"00",X"32",
		X"7B",X"C4",X"32",X"08",X"D0",X"F3",X"21",X"00",X"C0",X"11",X"01",X"C0",X"01",X"FF",X"07",X"36",
		X"00",X"ED",X"B0",X"21",X"00",X"E0",X"11",X"01",X"E0",X"01",X"FF",X"0F",X"36",X"00",X"ED",X"B0",
		X"3A",X"7B",X"C4",X"CB",X"FF",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"3A",X"18",X"D0",X"31",X"FE",
		X"C7",X"CD",X"DB",X"67",X"06",X"00",X"3A",X"0C",X"D0",X"CB",X"7F",X"28",X"05",X"10",X"F7",X"C3",
		X"98",X"03",X"CD",X"C9",X"9E",X"CD",X"06",X"27",X"ED",X"5F",X"28",X"EA",X"21",X"E6",X"17",X"3A",
		X"18",X"D0",X"CD",X"17",X"21",X"CD",X"55",X"18",X"CD",X"38",X"20",X"3E",X"0F",X"32",X"00",X"D0",
		X"3A",X"01",X"D0",X"32",X"C1",X"C4",X"CD",X"BF",X"95",X"AF",X"21",X"9E",X"E5",X"11",X"8B",X"18",
		X"CD",X"F1",X"21",X"AF",X"21",X"64",X"E7",X"11",X"9A",X"18",X"CD",X"F1",X"21",X"AF",X"21",X"2A",
		X"E5",X"11",X"B7",X"18",X"CD",X"F1",X"21",X"3E",X"0F",X"32",X"00",X"D0",X"3A",X"01",X"D0",X"32",
		X"C1",X"C4",X"3E",X"0F",X"32",X"00",X"D0",X"3A",X"01",X"D0",X"32",X"C1",X"C4",X"3E",X"01",X"32",
		X"E0",X"C3",X"C3",X"40",X"03",X"CD",X"2C",X"20",X"CD",X"73",X"18",X"3A",X"0C",X"D0",X"E6",X"30",
		X"C8",X"CD",X"38",X"20",X"AF",X"21",X"20",X"E5",X"11",X"80",X"18",X"CD",X"F1",X"21",X"32",X"10",
		X"D0",X"18",X"FB",X"06",X"00",X"DD",X"21",X"00",X"00",X"DD",X"21",X"00",X"00",X"10",X"F6",X"C9",
		X"0A",X"49",X"2E",X"4F",X"20",X"45",X"52",X"52",X"4F",X"52",X"2E",X"0E",X"48",X"41",X"52",X"44",
		X"57",X"41",X"52",X"45",X"20",X"43",X"48",X"45",X"43",X"4B",X"1C",X"57",X"41",X"49",X"54",X"20",
		X"55",X"4E",X"54",X"49",X"4C",X"20",X"54",X"49",X"4D",X"45",X"52",X"20",X"52",X"45",X"41",X"43",
		X"48",X"45",X"53",X"20",X"27",X"30",X"27",X"07",X"54",X"49",X"4D",X"45",X"52",X"20",X"3A",X"AF",
		X"32",X"08",X"D0",X"06",X"00",X"11",X"00",X"80",X"78",X"2F",X"3C",X"F5",X"21",X"09",X"19",X"CD",
		X"50",X"20",X"4E",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"F1",X"F5",X"21",X"09",X"1B",
		X"CD",X"50",X"20",X"7E",X"B1",X"12",X"13",X"F1",X"21",X"09",X"1D",X"CD",X"50",X"20",X"7E",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"12",X"13",X"10",X"CD",X"AF",X"CB",X"F7",X"32",X"08",
		X"D0",X"CD",X"09",X"1F",X"AF",X"32",X"08",X"D0",X"C9",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"0F",X"0B",X"0B",X"00",X"00",X"00",X"0B",X"00",X"0F",X"07",X"07",X"00",X"00",X"00",
		X"07",X"00",X"00",X"04",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",
		X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",
		X"00",X"00",X"0F",X"0F",X"0B",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"0B",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"0B",X"00",X"00",X"0F",X"0F",X"0C",X"09",X"0F",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"0A",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0A",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0D",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"0C",X"00",X"00",X"0F",X"0D",X"0B",X"08",X"05",
		X"0F",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",X"0F",X"00",X"00",X"0E",X"0F",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0C",X"09",X"08",X"00",X"00",X"0F",X"0F",X"0C",X"0A",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0D",X"0B",X"09",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"05",X"0D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"08",X"00",X"00",X"05",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"0F",X"08",X"0A",X"00",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"0A",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"0A",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"0A",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"0A",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"0A",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",
		X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",X"00",X"00",X"00",X"0F",X"0F",X"0B",X"08",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0A",X"07",X"00",X"00",X"00",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"0A",X"00",X"00",X"0F",X"0F",X"0C",X"0A",X"08",X"07",X"00",X"00",X"0F",X"0B",X"09",X"08",X"0F",
		X"00",X"00",X"0F",X"05",X"05",X"05",X"02",X"0C",X"09",X"00",X"0F",X"06",X"06",X"06",X"04",X"0D",
		X"0A",X"00",X"0F",X"07",X"07",X"07",X"06",X"0E",X"0B",X"00",X"0F",X"08",X"08",X"08",X"08",X"0F",
		X"0C",X"00",X"0F",X"00",X"00",X"00",X"00",X"0B",X"08",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"08",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"07",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",
		X"06",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0B",X"08",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0D",X"0B",X"09",X"07",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"00",
		X"0F",X"00",X"00",X"00",X"0B",X"0B",X"0B",X"00",X"0B",X"00",X"0F",X"00",X"07",X"07",X"07",X"00",
		X"07",X"00",X"0F",X"00",X"04",X"04",X"04",X"00",X"04",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"05",X"03",X"03",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",
		X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",X"08",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",
		X"0F",X"00",X"0F",X"00",X"00",X"0F",X"0B",X"0F",X"0B",X"00",X"0F",X"0F",X"0B",X"00",X"00",X"0F",
		X"0B",X"00",X"0F",X"0F",X"0B",X"0F",X"0B",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0F",X"0F",X"0A",X"08",X"00",X"00",X"00",X"00",X"0F",X"0A",X"08",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0A",X"08",X"0F",
		X"0A",X"00",X"00",X"0F",X"0F",X"0F",X"0A",X"00",X"00",X"00",X"00",X"0F",X"0B",X"07",X"00",X"00",
		X"05",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",X"00",X"00",X"00",X"0E",X"08",X"0F",X"0F",X"00",
		X"07",X"00",X"00",X"0F",X"00",X"0F",X"0C",X"09",X"08",X"00",X"00",X"0F",X"09",X"0F",X"0F",X"09",
		X"08",X"00",X"00",X"0F",X"09",X"0F",X"0C",X"0A",X"08",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"0A",X"08",X"06",X"06",X"00",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"05",X"08",X"00",X"08",X"05",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"05",X"08",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",
		X"00",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",X"08",X"00",X"00",X"0F",X"05",X"02",X"08",X"06",
		X"0F",X"00",X"0F",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0A",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0B",X"09",X"08",X"00",
		X"00",X"00",X"04",X"07",X"05",X"00",X"00",X"0B",X"08",X"00",X"03",X"07",X"05",X"00",X"00",X"0B",
		X"08",X"00",X"02",X"07",X"05",X"00",X"00",X"0B",X"08",X"00",X"01",X"07",X"05",X"00",X"00",X"0B",
		X"08",X"00",X"0F",X"07",X"05",X"00",X"00",X"0B",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"09",X"06",X"00",X"00",
		X"00",X"00",X"05",X"07",X"05",X"00",X"00",X"0B",X"08",X"00",X"0F",X"0F",X"0A",X"08",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"00",X"0F",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"00",X"0B",X"00",X"0B",X"0B",X"00",X"00",X"00",X"00",X"07",X"00",X"07",
		X"07",X"00",X"0F",X"00",X"00",X"04",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"07",X"06",X"05",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"04",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",
		X"09",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",X"0F",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",
		X"0F",X"00",X"0F",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",
		X"0F",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0C",X"0A",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"0A",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"0F",X"0F",X"0F",X"0B",X"07",
		X"00",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0E",X"00",X"00",X"00",X"0E",X"00",X"0F",X"00",X"00",
		X"0F",X"00",X"00",X"0F",X"0F",X"00",X"0C",X"09",X"08",X"00",X"00",X"0F",X"00",X"0F",X"0A",X"09",
		X"0F",X"00",X"00",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"0F",X"0B",X"0A",X"09",X"08",X"07",X"06",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"0C",X"07",X"00",X"0F",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"08",X"07",X"00",X"05",X"02",X"0F",X"00",X"00",X"0F",X"00",X"0F",
		X"0F",X"02",X"00",X"00",X"0F",X"00",X"08",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",X"00",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",
		X"0C",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",X"0F",X"00",X"00",X"0F",X"00",X"00",X"08",X"06",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0A",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0B",X"09",X"08",X"00",
		X"00",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",X"08",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",
		X"08",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",X"08",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",
		X"08",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"02",X"00",X"0F",X"09",X"06",X"00",X"00",
		X"00",X"02",X"00",X"0B",X"0A",X"08",X"00",X"0B",X"08",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"06",X"00",X"11",X"00",X"80",X"78",X"2F",
		X"3C",X"F5",X"21",X"09",X"1A",X"CD",X"50",X"20",X"4E",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"CB",
		X"21",X"F1",X"F5",X"21",X"09",X"1C",X"CD",X"50",X"20",X"7E",X"B1",X"12",X"13",X"F1",X"21",X"09",
		X"1E",X"CD",X"50",X"20",X"7E",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"12",X"13",X"10",
		X"CD",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"06",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"12",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"16",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"7B",X"C4",X"CB",
		X"DF",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"C9",X"3A",X"7B",X"C4",X"CB",X"9F",X"32",X"7B",X"C4",
		X"32",X"08",X"D0",X"C9",X"81",X"4F",X"D0",X"04",X"3F",X"C9",X"83",X"5F",X"D0",X"14",X"3F",X"C9",
		X"85",X"6F",X"D0",X"24",X"3F",X"C9",X"85",X"6F",X"30",X"01",X"24",X"5E",X"23",X"56",X"C9",X"7B",
		X"CD",X"77",X"20",X"08",X"E5",X"7A",X"CD",X"79",X"20",X"57",X"08",X"84",X"65",X"6B",X"5F",X"30",
		X"01",X"14",X"C1",X"09",X"D0",X"13",X"C9",X"1E",X"00",X"63",X"6B",X"87",X"30",X"02",X"09",X"8B",
		X"29",X"8F",X"30",X"02",X"09",X"8B",X"29",X"8F",X"30",X"02",X"09",X"8B",X"29",X"8F",X"30",X"02",
		X"09",X"8B",X"29",X"8F",X"30",X"02",X"09",X"8B",X"29",X"8F",X"30",X"02",X"09",X"8B",X"29",X"8F",
		X"30",X"02",X"09",X"8B",X"29",X"8F",X"D0",X"09",X"8B",X"C9",X"2E",X"00",X"67",X"48",X"06",X"00",
		X"3E",X"08",X"29",X"30",X"01",X"09",X"3D",X"20",X"F9",X"C9",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"F5",X"7C",X"E6",X"03",X"67",X"F1",
		X"C9",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"F5",X"7C",X"E6",
		X"07",X"67",X"F1",X"C9",X"C5",X"7A",X"2F",X"3C",X"E6",X"F8",X"06",X"08",X"CD",X"AA",X"20",X"7B",
		X"E6",X"F8",X"CB",X"3F",X"CB",X"3F",X"CD",X"50",X"20",X"11",X"00",X"E0",X"19",X"5E",X"23",X"56",
		X"2B",X"C1",X"C9",X"F5",X"7D",X"D6",X"41",X"6F",X"30",X"01",X"25",X"F1",X"C9",X"F5",X"7B",X"D6",
		X"41",X"5F",X"30",X"01",X"15",X"F1",X"C9",X"E5",X"D5",X"C5",X"21",X"00",X"E0",X"11",X"02",X"E0",
		X"01",X"FE",X"07",X"36",X"00",X"23",X"36",X"20",X"2B",X"ED",X"B0",X"C1",X"D1",X"E1",X"C9",X"21",
		X"04",X"E0",X"06",X"20",X"C5",X"E5",X"D1",X"13",X"13",X"01",X"3A",X"00",X"36",X"00",X"23",X"36",
		X"20",X"2B",X"E5",X"ED",X"B0",X"E1",X"11",X"40",X"00",X"19",X"C1",X"10",X"E7",X"C9",X"21",X"F0",
		X"08",X"CD",X"D1",X"20",X"7C",X"32",X"CB",X"C4",X"4D",X"21",X"86",X"E0",X"CD",X"6C",X"21",X"21",
		X"46",X"E7",X"CD",X"6C",X"21",X"21",X"44",X"E7",X"CD",X"80",X"21",X"C9",X"11",X"96",X"21",X"06",
		X"1D",X"3A",X"CB",X"C4",X"F6",X"48",X"77",X"23",X"1A",X"81",X"77",X"23",X"13",X"10",X"F2",X"C9",
		X"11",X"B4",X"21",X"06",X"1C",X"3A",X"CB",X"C4",X"F6",X"48",X"77",X"23",X"1A",X"81",X"13",X"77",
		X"CD",X"03",X"21",X"10",X"F0",X"C9",X"04",X"03",X"02",X"01",X"00",X"04",X"03",X"02",X"01",X"00",
		X"04",X"03",X"02",X"01",X"00",X"04",X"03",X"02",X"01",X"00",X"04",X"03",X"02",X"01",X"00",X"04",
		X"03",X"02",X"01",X"00",X"05",X"0A",X"0A",X"0A",X"0A",X"06",X"07",X"08",X"09",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"06",X"07",X"08",X"09",X"0A",X"0A",X"0A",X"0A",X"0B",
		X"E5",X"D5",X"C5",X"21",X"00",X"E8",X"11",X"01",X"E8",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",
		X"21",X"7D",X"C4",X"11",X"7E",X"C4",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"C1",X"D1",X"E1",
		X"C9",X"C5",X"F5",X"F5",X"1A",X"47",X"0E",X"FF",X"F1",X"07",X"07",X"07",X"13",X"EB",X"12",X"13",
		X"ED",X"A0",X"1B",X"CD",X"0D",X"21",X"10",X"F6",X"F1",X"C1",X"C9",X"C5",X"07",X"07",X"07",X"4F",
		X"1A",X"47",X"71",X"23",X"CD",X"03",X"21",X"10",X"F9",X"79",X"C1",X"C9",X"C5",X"1A",X"47",X"AF",
		X"77",X"23",X"36",X"20",X"CD",X"03",X"21",X"10",X"F7",X"C1",X"C9",X"F5",X"0A",X"03",X"32",X"C9",
		X"C4",X"DD",X"21",X"C9",X"C4",X"F1",X"07",X"07",X"07",X"F5",X"E5",X"F5",X"0A",X"03",X"CD",X"50",
		X"20",X"EB",X"F1",X"B2",X"77",X"23",X"73",X"CD",X"03",X"21",X"EB",X"E6",X"0F",X"E1",X"DD",X"35",
		X"00",X"20",X"E7",X"F1",X"C9",X"EB",X"C5",X"E5",X"CD",X"65",X"22",X"E1",X"01",X"40",X"00",X"09",
		X"C1",X"0D",X"20",X"F2",X"C9",X"F5",X"B2",X"77",X"F1",X"23",X"73",X"13",X"23",X"10",X"F6",X"C9",
		X"3A",X"72",X"ED",X"FE",X"20",X"20",X"0E",X"3E",X"08",X"32",X"CA",X"C4",X"21",X"D0",X"37",X"CD",
		X"D1",X"20",X"23",X"18",X"1A",X"3E",X"F8",X"32",X"CA",X"C4",X"21",X"00",X"0C",X"CD",X"D1",X"20",
		X"3A",X"72",X"ED",X"E6",X"03",X"11",X"C6",X"22",X"CD",X"4A",X"20",X"1A",X"CD",X"50",X"20",X"EB",
		X"3A",X"71",X"ED",X"3D",X"C8",X"FE",X"05",X"38",X"02",X"3E",X"05",X"47",X"21",X"3E",X"E7",X"D5",
		X"CD",X"BB",X"22",X"1B",X"CD",X"BB",X"22",X"D1",X"10",X"F5",X"C9",X"3A",X"CA",X"C4",X"82",X"77",
		X"23",X"73",X"CD",X"03",X"21",X"C9",X"05",X"03",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"FF",X"0E",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"0E",X"FF",X"00",X"00",X"FF",
		X"0A",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"0A",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"02",X"02",X"02",X"1E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"06",X"06",X"06",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1A",X"0A",X"0A",X"0A",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"0E",X"0E",X"0E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"12",X"12",
		X"12",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"16",X"16",X"16",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A8",X"FD",X"21",X"CC",X"C4",X"FD",X"34",X"00",X"CD",X"4E",X"24",X"CD",
		X"85",X"27",X"CD",X"F5",X"24",X"CD",X"9F",X"25",X"CD",X"CC",X"23",X"C9",X"3A",X"CE",X"C4",X"A7",
		X"C8",X"21",X"CD",X"C4",X"34",X"CB",X"46",X"C8",X"7E",X"F5",X"FE",X"0D",X"20",X"03",X"3E",X"07",
		X"77",X"F1",X"CB",X"3F",X"5F",X"CB",X"27",X"CB",X"27",X"83",X"83",X"5F",X"16",X"00",X"21",X"24",
		X"24",X"19",X"7E",X"32",X"CF",X"C4",X"23",X"EB",X"21",X"F0",X"08",X"CD",X"D1",X"20",X"01",X"B6",
		X"E0",X"3E",X"05",X"F5",X"E5",X"1A",X"FE",X"FF",X"20",X"06",X"3E",X"20",X"26",X"00",X"18",X"01",
		X"85",X"03",X"02",X"0B",X"3A",X"CF",X"C4",X"CE",X"00",X"84",X"02",X"03",X"03",X"13",X"E1",X"F1",
		X"3D",X"20",X"E0",X"C9",X"50",X"10",X"0F",X"0E",X"0D",X"0C",X"50",X"15",X"14",X"13",X"12",X"11",
		X"50",X"19",X"18",X"FF",X"17",X"16",X"60",X"1D",X"1C",X"FF",X"1B",X"1A",X"60",X"1F",X"22",X"21",
		X"20",X"1E",X"60",X"1F",X"25",X"24",X"23",X"1E",X"60",X"1F",X"2B",X"2A",X"29",X"1E",X"3A",X"D0",
		X"C4",X"A7",X"C8",X"CB",X"67",X"28",X"12",X"CB",X"47",X"28",X"38",X"3A",X"D1",X"C4",X"47",X"3A",
		X"32",X"C4",X"B8",X"C8",X"32",X"D1",X"C4",X"18",X"0F",X"CB",X"E7",X"32",X"D0",X"C4",X"21",X"FE",
		X"E2",X"11",X"A1",X"24",X"AF",X"CD",X"F1",X"21",X"3A",X"32",X"C4",X"DD",X"21",X"3E",X"E1",X"FE",
		X"0A",X"DD",X"36",X"01",X"20",X"38",X"06",X"DD",X"36",X"01",X"31",X"D6",X"0A",X"C6",X"30",X"DD",
		X"77",X"C1",X"C9",X"11",X"A1",X"24",X"21",X"FE",X"E2",X"CD",X"1C",X"22",X"AF",X"32",X"D0",X"C4",
		X"C9",X"09",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"20",X"20",X"11",X"D3",X"24",X"18",X"03",
		X"11",X"E4",X"24",X"31",X"FE",X"C7",X"21",X"20",X"E7",X"AF",X"CD",X"F1",X"21",X"01",X"00",X"00",
		X"16",X"03",X"32",X"10",X"D0",X"32",X"10",X"D0",X"0B",X"78",X"B1",X"20",X"F5",X"15",X"20",X"F2",
		X"C3",X"00",X"00",X"10",X"53",X"54",X"41",X"43",X"4B",X"20",X"4F",X"56",X"45",X"52",X"46",X"4C",
		X"4F",X"57",X"21",X"21",X"10",X"50",X"43",X"20",X"52",X"41",X"4E",X"47",X"45",X"20",X"45",X"52",
		X"52",X"4F",X"52",X"21",X"21",X"DD",X"21",X"D2",X"C4",X"DD",X"7E",X"00",X"A7",X"C8",X"CB",X"47",
		X"20",X"14",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"11",X"7D",X"25",X"21",
		X"20",X"E7",X"CD",X"1C",X"22",X"C9",X"CB",X"67",X"20",X"0D",X"CB",X"E7",X"DD",X"77",X"00",X"FD",
		X"7E",X"00",X"C6",X"05",X"DD",X"77",X"01",X"DD",X"7E",X"01",X"FD",X"BE",X"00",X"C0",X"3A",X"32",
		X"C4",X"A7",X"C8",X"3D",X"21",X"63",X"25",X"28",X"03",X"21",X"7D",X"25",X"DD",X"7E",X"02",X"DD",
		X"34",X"02",X"11",X"97",X"25",X"CD",X"4A",X"20",X"1A",X"FE",X"FF",X"20",X"06",X"AF",X"DD",X"77",
		X"02",X"18",X"E9",X"11",X"20",X"E7",X"EB",X"CD",X"F1",X"21",X"FD",X"7E",X"00",X"C6",X"05",X"DD",
		X"77",X"01",X"C9",X"19",X"50",X"55",X"53",X"48",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"19",X"50",X"55",
		X"53",X"48",X"20",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"FF",X"3A",
		X"D5",X"C4",X"A7",X"C8",X"CB",X"47",X"CA",X"A2",X"26",X"CB",X"67",X"CC",X"B0",X"25",X"18",X"57",
		X"CB",X"E7",X"32",X"D5",X"C4",X"21",X"80",X"E6",X"11",X"F2",X"26",X"3E",X"01",X"CD",X"F1",X"21",
		X"AF",X"21",X"42",X"E7",X"11",X"EA",X"26",X"CD",X"F1",X"21",X"CD",X"2C",X"26",X"21",X"00",X"E5",
		X"11",X"FA",X"26",X"3E",X"01",X"CD",X"F1",X"21",X"21",X"C2",X"E4",X"11",X"E2",X"26",X"AF",X"CD",
		X"F1",X"21",X"CD",X"40",X"26",X"3A",X"6F",X"ED",X"CB",X"47",X"28",X"1B",X"21",X"C0",X"E1",X"11",
		X"F6",X"26",X"3E",X"01",X"CD",X"F1",X"21",X"21",X"82",X"E2",X"11",X"EA",X"26",X"AF",X"CD",X"F1",
		X"21",X"CD",X"36",X"26",X"32",X"D6",X"C4",X"3A",X"6F",X"ED",X"CB",X"57",X"28",X"1D",X"CD",X"8E",
		X"26",X"CB",X"47",X"28",X"08",X"CD",X"2C",X"26",X"CD",X"36",X"26",X"18",X"08",X"CB",X"4F",X"CC",
		X"2C",X"26",X"C4",X"36",X"26",X"CD",X"4A",X"27",X"CD",X"40",X"26",X"C9",X"21",X"42",X"E7",X"11",
		X"D7",X"C4",X"CD",X"4A",X"26",X"C9",X"21",X"82",X"E2",X"11",X"DB",X"C4",X"CD",X"4A",X"26",X"C9",
		X"21",X"C2",X"E4",X"11",X"DF",X"C4",X"CD",X"4A",X"26",X"C9",X"F5",X"06",X"03",X"1A",X"4F",X"07",
		X"07",X"07",X"07",X"E6",X"0F",X"CD",X"6F",X"26",X"78",X"FE",X"01",X"20",X"03",X"32",X"E3",X"C4",
		X"79",X"E6",X"0F",X"CD",X"6F",X"26",X"13",X"10",X"E4",X"AF",X"32",X"E3",X"C4",X"F1",X"C9",X"23",
		X"A7",X"F5",X"20",X"0B",X"3A",X"E3",X"C4",X"A7",X"20",X"05",X"36",X"20",X"F1",X"18",X"07",X"F1",
		X"C6",X"30",X"77",X"32",X"E3",X"C4",X"2B",X"36",X"00",X"23",X"CD",X"03",X"21",X"C9",X"F5",X"3A",
		X"D6",X"C4",X"3C",X"32",X"D6",X"C4",X"FE",X"19",X"CC",X"BC",X"26",X"FE",X"32",X"CC",X"BC",X"26",
		X"F1",X"C9",X"AF",X"32",X"D5",X"C4",X"32",X"D6",X"C4",X"21",X"80",X"E6",X"11",X"05",X"27",X"CD",
		X"1C",X"22",X"21",X"42",X"E7",X"11",X"05",X"27",X"CD",X"1C",X"22",X"C9",X"F5",X"3A",X"6F",X"ED",
		X"21",X"80",X"E6",X"11",X"F2",X"26",X"CB",X"4F",X"28",X"06",X"11",X"F6",X"26",X"21",X"C0",X"E1",
		X"F1",X"FE",X"32",X"20",X"09",X"3E",X"01",X"CD",X"F1",X"21",X"32",X"D6",X"C4",X"C9",X"CD",X"1C",
		X"22",X"C9",X"07",X"20",X"20",X"20",X"20",X"20",X"30",X"30",X"07",X"20",X"20",X"20",X"20",X"20",
		X"30",X"30",X"03",X"31",X"55",X"50",X"03",X"32",X"55",X"50",X"0A",X"48",X"49",X"47",X"48",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"1A",X"21",X"12",X"27",X"11",X"DF",X"C4",X"01",X"03",X"00",X"ED",
		X"B0",X"C9",X"00",X"50",X"00",X"21",X"D7",X"C4",X"11",X"D8",X"C4",X"01",X"07",X"00",X"36",X"00",
		X"ED",X"B0",X"C9",X"F5",X"3A",X"66",X"EF",X"A7",X"20",X"1E",X"E5",X"3A",X"6F",X"ED",X"21",X"D9",
		X"C4",X"CB",X"4F",X"28",X"03",X"21",X"DD",X"C4",X"7B",X"86",X"27",X"77",X"7A",X"2B",X"8E",X"27",
		X"77",X"3E",X"00",X"2B",X"8E",X"27",X"77",X"E1",X"F1",X"C9",X"F5",X"D5",X"E5",X"3A",X"6F",X"ED",
		X"11",X"DF",X"C4",X"21",X"D7",X"C4",X"CB",X"4F",X"28",X"03",X"21",X"DB",X"C4",X"1A",X"BE",X"28",
		X"04",X"30",X"1E",X"18",X"12",X"23",X"13",X"1A",X"BE",X"28",X"04",X"30",X"14",X"18",X"0C",X"23",
		X"13",X"1A",X"BE",X"30",X"0C",X"18",X"08",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",
		X"12",X"E1",X"D1",X"F1",X"C9",X"3A",X"6F",X"ED",X"11",X"6C",X"EF",X"01",X"68",X"EF",X"21",X"D7",
		X"C4",X"CB",X"4F",X"28",X"09",X"21",X"DB",X"C4",X"11",X"6E",X"EF",X"01",X"69",X"EF",X"1A",X"BE",
		X"38",X"08",X"C0",X"23",X"13",X"1A",X"BE",X"38",X"02",X"C0",X"13",X"0A",X"CB",X"47",X"20",X"25",
		X"3A",X"71",X"ED",X"3C",X"32",X"71",X"ED",X"3E",X"10",X"CD",X"AE",X"67",X"E5",X"3A",X"6F",X"ED",
		X"21",X"6A",X"EF",X"CB",X"4F",X"28",X"03",X"21",X"6B",X"EF",X"34",X"E1",X"C5",X"D5",X"E5",X"CD",
		X"70",X"22",X"E1",X"D1",X"C1",X"3A",X"C1",X"C4",X"CB",X"67",X"20",X"04",X"0A",X"CB",X"C7",X"02",
		X"E5",X"3A",X"6F",X"ED",X"11",X"6C",X"EF",X"21",X"6A",X"EF",X"CB",X"4F",X"28",X"06",X"11",X"6E",
		X"EF",X"21",X"6B",X"EF",X"7E",X"FE",X"01",X"20",X"04",X"3E",X"40",X"18",X"02",X"3E",X"60",X"E1",
		X"EB",X"23",X"86",X"27",X"77",X"2B",X"3E",X"00",X"8E",X"27",X"77",X"C3",X"85",X"27",X"21",X"A0",
		X"1C",X"CD",X"BA",X"20",X"11",X"0E",X"00",X"19",X"01",X"B0",X"60",X"1E",X"03",X"16",X"00",X"CD",
		X"64",X"29",X"AF",X"32",X"E4",X"C4",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"3A",X"72",X"ED",X"3C",
		X"06",X"FF",X"D6",X"0A",X"04",X"30",X"FB",X"C6",X"0A",X"4F",X"C5",X"06",X"00",X"09",X"01",X"B0",
		X"90",X"3E",X"03",X"1E",X"00",X"CD",X"B9",X"BD",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"C1",X"48",
		X"79",X"FE",X"00",X"C8",X"06",X"00",X"09",X"01",X"B0",X"88",X"3E",X"04",X"1E",X"00",X"CD",X"B9",
		X"BD",X"C9",X"3A",X"6F",X"ED",X"CB",X"47",X"28",X"13",X"01",X"C0",X"48",X"CD",X"83",X"28",X"01",
		X"C0",X"78",X"CD",X"97",X"28",X"01",X"C0",X"90",X"CD",X"B5",X"28",X"C9",X"01",X"C0",X"6C",X"CD",
		X"B5",X"28",X"C9",X"C5",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"11",X"11",X"00",X"19",X"1E",X"03",
		X"16",X"05",X"C1",X"CD",X"64",X"29",X"C9",X"C5",X"3A",X"6F",X"ED",X"1E",X"01",X"CB",X"4F",X"28",
		X"02",X"1E",X"02",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"16",X"00",X"19",X"3E",X"08",X"1E",X"00",
		X"C1",X"CD",X"B9",X"BD",X"C9",X"C5",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"11",X"14",X"00",X"19",
		X"1E",X"03",X"16",X"09",X"C1",X"CD",X"64",X"29",X"C9",X"01",X"B0",X"38",X"CD",X"83",X"28",X"01",
		X"B0",X"68",X"CD",X"97",X"28",X"01",X"B0",X"80",X"CD",X"E2",X"28",X"01",X"B0",X"A8",X"CD",X"F6",
		X"28",X"C9",X"C5",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"11",X"0A",X"00",X"19",X"1E",X"02",X"16",
		X"0C",X"C1",X"CD",X"64",X"29",X"C9",X"C5",X"21",X"A0",X"1C",X"CD",X"BA",X"20",X"11",X"0C",X"00",
		X"19",X"1E",X"02",X"16",X"0E",X"C1",X"CD",X"64",X"29",X"C9",X"3A",X"6F",X"ED",X"CB",X"47",X"20",
		X"0D",X"01",X"B0",X"5E",X"CD",X"E2",X"28",X"01",X"B0",X"86",X"CD",X"F6",X"28",X"C9",X"01",X"70",
		X"5E",X"CD",X"E2",X"28",X"01",X"70",X"86",X"CD",X"F6",X"28",X"C9",X"21",X"54",X"29",X"3A",X"72",
		X"ED",X"E6",X"03",X"87",X"CD",X"56",X"20",X"3E",X"07",X"CD",X"50",X"20",X"7E",X"4F",X"EB",X"CD",
		X"D1",X"20",X"EB",X"21",X"2C",X"E5",X"06",X"0A",X"79",X"B2",X"77",X"23",X"73",X"CD",X"03",X"21",
		X"13",X"10",X"F5",X"C9",X"E0",X"37",X"30",X"38",X"80",X"38",X"D0",X"38",X"E0",X"00",X"E8",X"00",
		X"E8",X"00",X"F0",X"00",X"D5",X"7A",X"1E",X"00",X"D5",X"E5",X"C5",X"CD",X"B9",X"BD",X"C1",X"E1",
		X"D1",X"23",X"3E",X"10",X"80",X"47",X"D1",X"14",X"1D",X"20",X"E9",X"C9",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"16",X"0A",X"16",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"16",X"0A",X"02",X"0A",
		X"16",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"16",X"0A",X"02",X"0A",X"02",X"0A",X"16",X"00",
		X"00",X"00",X"FF",X"00",X"16",X"0A",X"02",X"0A",X"03",X"0A",X"02",X"0A",X"16",X"00",X"00",X"FF",
		X"00",X"00",X"16",X"0A",X"02",X"0A",X"02",X"0A",X"16",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"16",X"0A",X"02",X"0A",X"16",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"16",X"0A",
		X"16",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"CD",X"BF",X"95",X"CD",X"D0",X"21",X"CD",X"57",X"2D",
		X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",
		X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"01",X"00",X"08",X"0B",X"78",
		X"B1",X"20",X"FB",X"3A",X"0C",X"D0",X"CB",X"47",X"32",X"10",X"D0",X"20",X"D3",X"31",X"FE",X"C7",
		X"3E",X"80",X"32",X"08",X"D0",X"32",X"7B",X"C4",X"CD",X"17",X"21",X"3E",X"0F",X"32",X"00",X"D0",
		X"3A",X"01",X"D0",X"32",X"C1",X"C4",X"CD",X"BF",X"95",X"CD",X"2C",X"20",X"21",X"02",X"E5",X"11",
		X"50",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"8C",X"E3",X"11",X"5A",X"2E",X"AF",X"CD",X"F1",X"21",
		X"21",X"8C",X"E6",X"11",X"5F",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"10",X"E7",X"11",X"67",X"2E",
		X"AF",X"CD",X"F1",X"21",X"21",X"90",X"E3",X"11",X"71",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"88",
		X"E6",X"11",X"7B",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"88",X"E3",X"11",X"81",X"2E",X"AF",X"CD",
		X"F1",X"21",X"21",X"14",X"E7",X"11",X"87",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"94",X"E3",X"11",
		X"99",X"2E",X"AF",X"CD",X"F1",X"21",X"21",X"A6",X"E6",X"11",X"7C",X"2F",X"AF",X"CD",X"F1",X"21",
		X"21",X"24",X"E5",X"11",X"04",X"30",X"AF",X"CD",X"F1",X"21",X"21",X"E6",X"E2",X"11",X"F9",X"2F",
		X"AF",X"CD",X"F1",X"21",X"21",X"AC",X"E6",X"11",X"F0",X"2F",X"AF",X"CD",X"F1",X"21",X"21",X"B0",
		X"E6",X"11",X"D3",X"2F",X"AF",X"CD",X"F1",X"21",X"21",X"B4",X"E6",X"11",X"DC",X"2F",X"AF",X"CD",
		X"F1",X"21",X"21",X"1C",X"E7",X"11",X"E5",X"2F",X"AF",X"CD",X"F1",X"21",X"CD",X"DB",X"67",X"3A",
		X"7B",X"C4",X"CB",X"97",X"32",X"08",X"D0",X"3A",X"7C",X"C4",X"32",X"F5",X"C4",X"AF",X"32",X"F6",
		X"C4",X"3E",X"EF",X"CD",X"AE",X"67",X"CD",X"92",X"67",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",
		X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"3E",
		X"16",X"86",X"E1",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"7C",X"C4",X"32",X"18",X"D0",
		X"CB",X"76",X"28",X"FC",X"CB",X"7E",X"20",X"FC",X"11",X"7C",X"C4",X"E5",X"D5",X"21",X"7D",X"C4",
		X"11",X"00",X"E8",X"01",X"40",X"00",X"ED",X"B0",X"D1",X"E1",X"3A",X"18",X"D0",X"12",X"CB",X"7E",
		X"20",X"FC",X"D5",X"CD",X"92",X"67",X"E1",X"3A",X"18",X"D0",X"86",X"77",X"CD",X"DD",X"2B",X"32",
		X"10",X"D0",X"01",X"C0",X"0B",X"0B",X"78",X"B1",X"20",X"FB",X"C3",X"79",X"2B",X"3A",X"0C",X"D0",
		X"CB",X"47",X"11",X"77",X"2F",X"20",X"03",X"11",X"72",X"2F",X"21",X"D0",X"E4",X"AF",X"CD",X"F1",
		X"21",X"3A",X"0C",X"D0",X"CB",X"4F",X"11",X"77",X"2F",X"20",X"03",X"11",X"72",X"2F",X"21",X"50",
		X"E1",X"AF",X"CD",X"F1",X"21",X"3A",X"0C",X"D0",X"CB",X"57",X"11",X"77",X"2F",X"20",X"03",X"11",
		X"72",X"2F",X"21",X"CC",X"E4",X"AF",X"CD",X"F1",X"21",X"3A",X"0C",X"D0",X"CB",X"5F",X"11",X"77",
		X"2F",X"20",X"03",X"11",X"72",X"2F",X"21",X"4C",X"E2",X"AF",X"CD",X"F1",X"21",X"3A",X"0C",X"D0",
		X"CB",X"67",X"11",X"77",X"2F",X"28",X"03",X"11",X"72",X"2F",X"21",X"48",X"E5",X"AF",X"CD",X"F1",
		X"21",X"3A",X"0C",X"D0",X"CB",X"6F",X"11",X"77",X"2F",X"28",X"03",X"11",X"72",X"2F",X"21",X"48",
		X"E2",X"AF",X"CD",X"F1",X"21",X"3A",X"10",X"D0",X"CB",X"47",X"11",X"77",X"2F",X"20",X"03",X"11",
		X"72",X"2F",X"21",X"D4",X"E4",X"AF",X"CD",X"F1",X"21",X"3A",X"10",X"D0",X"CB",X"57",X"11",X"77",
		X"2F",X"20",X"03",X"11",X"72",X"2F",X"21",X"54",X"E1",X"AF",X"CD",X"F1",X"21",X"11",X"8F",X"2E",
		X"3A",X"0C",X"D0",X"CB",X"4F",X"20",X"03",X"11",X"A1",X"2E",X"21",X"18",X"E7",X"AF",X"CD",X"F1",
		X"21",X"3A",X"0C",X"D0",X"CB",X"4F",X"3A",X"7B",X"C4",X"CB",X"97",X"20",X"02",X"CB",X"D7",X"32",
		X"08",X"D0",X"3A",X"7C",X"C4",X"21",X"E5",X"C4",X"CD",X"2A",X"2D",X"21",X"D8",X"E4",X"11",X"E5",
		X"C4",X"AF",X"CD",X"F1",X"21",X"3A",X"0C",X"D0",X"CB",X"4F",X"3A",X"7B",X"C4",X"CB",X"97",X"20",
		X"02",X"CB",X"D7",X"32",X"08",X"D0",X"3A",X"F5",X"C4",X"47",X"3A",X"7C",X"C4",X"90",X"21",X"0C",
		X"D0",X"CB",X"46",X"20",X"11",X"21",X"F6",X"C4",X"CB",X"46",X"20",X"0F",X"CD",X"AE",X"67",X"21",
		X"F6",X"C4",X"CB",X"C6",X"18",X"05",X"21",X"F6",X"C4",X"CB",X"86",X"21",X"E5",X"C4",X"CD",X"2A",
		X"2D",X"21",X"9C",X"E4",X"11",X"E5",X"C4",X"AF",X"CD",X"F1",X"21",X"3E",X"0F",X"32",X"00",X"D0",
		X"3A",X"01",X"D0",X"21",X"E5",X"C4",X"36",X"08",X"23",X"06",X"08",X"36",X"4C",X"CB",X"47",X"28",
		X"02",X"36",X"48",X"23",X"0F",X"10",X"F4",X"11",X"E5",X"C4",X"21",X"26",X"E5",X"AF",X"CD",X"F1",
		X"21",X"C9",X"64",X"2F",X"56",X"2F",X"48",X"2F",X"3A",X"2F",X"36",X"04",X"23",X"36",X"3A",X"23",
		X"36",X"20",X"23",X"F5",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"0A",X"30",X"04",
		X"C6",X"30",X"18",X"02",X"C6",X"37",X"77",X"23",X"F1",X"E6",X"0F",X"FE",X"0A",X"30",X"04",X"C6",
		X"30",X"18",X"02",X"C6",X"37",X"77",X"C9",X"21",X"48",X"2E",X"11",X"00",X"E0",X"01",X"04",X"00",
		X"ED",X"B0",X"21",X"00",X"E0",X"01",X"3C",X"00",X"ED",X"B0",X"21",X"4C",X"2E",X"11",X"40",X"E0",
		X"01",X"04",X"00",X"ED",X"B0",X"21",X"40",X"E0",X"01",X"3C",X"00",X"ED",X"B0",X"21",X"00",X"E0",
		X"11",X"80",X"E0",X"01",X"80",X"07",X"ED",X"B0",X"21",X"10",X"E2",X"3E",X"18",X"16",X"66",X"CD",
		X"B1",X"2D",X"21",X"10",X"E3",X"3E",X"18",X"16",X"65",X"CD",X"B1",X"2D",X"21",X"10",X"E4",X"3E",
		X"18",X"16",X"64",X"CD",X"B1",X"2D",X"21",X"10",X"E5",X"3E",X"18",X"16",X"63",X"CD",X"B1",X"2D",
		X"C9",X"1E",X"04",X"0E",X"04",X"E5",X"D5",X"F5",X"06",X"04",X"77",X"23",X"72",X"23",X"10",X"FA",
		X"D6",X"08",X"0D",X"20",X"F3",X"F1",X"D1",X"E1",X"F5",X"3E",X"40",X"CD",X"50",X"20",X"F1",X"1D",
		X"20",X"E1",X"C9",X"D9",X"21",X"00",X"E0",X"01",X"00",X"08",X"AF",X"77",X"BE",X"20",X"39",X"3D",
		X"77",X"BE",X"20",X"34",X"23",X"0B",X"78",X"B1",X"20",X"F0",X"21",X"00",X"E8",X"01",X"40",X"00",
		X"AF",X"77",X"BE",X"20",X"23",X"3D",X"77",X"BE",X"20",X"1E",X"23",X"0B",X"78",X"B1",X"20",X"F0",
		X"21",X"00",X"C0",X"01",X"00",X"08",X"AF",X"77",X"BE",X"20",X"0D",X"3D",X"77",X"BE",X"20",X"08",
		X"23",X"0B",X"78",X"B1",X"20",X"F0",X"D9",X"E9",X"F3",X"31",X"FF",X"C7",X"D5",X"CD",X"17",X"21",
		X"CD",X"D0",X"21",X"E1",X"7C",X"FE",X"E8",X"28",X"0B",X"E6",X"F0",X"FE",X"E0",X"28",X"0A",X"11",
		X"BD",X"2F",X"18",X"08",X"11",X"AC",X"2F",X"18",X"03",X"11",X"9B",X"2F",X"21",X"20",X"E6",X"AF",
		X"CD",X"F1",X"21",X"32",X"10",X"D0",X"18",X"FB",X"00",X"60",X"00",X"61",X"00",X"5E",X"00",X"62",
		X"09",X"54",X"45",X"53",X"54",X"20",X"4D",X"4F",X"44",X"45",X"04",X"54",X"49",X"4C",X"54",X"07",
		X"53",X"45",X"52",X"56",X"49",X"43",X"45",X"09",X"31",X"50",X"20",X"53",X"45",X"4C",X"45",X"43",
		X"54",X"09",X"32",X"50",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"05",X"43",X"4F",X"49",X"4E",
		X"41",X"05",X"43",X"4F",X"49",X"4E",X"42",X"07",X"31",X"50",X"20",X"46",X"49",X"52",X"45",X"09",
		X"31",X"50",X"20",X"50",X"41",X"44",X"44",X"4C",X"45",X"07",X"32",X"50",X"20",X"46",X"49",X"52",
		X"45",X"09",X"32",X"50",X"20",X"50",X"41",X"44",X"44",X"4C",X"45",X"0A",X"49",X"4E",X"54",X"45",
		X"52",X"52",X"55",X"50",X"54",X"20",X"0A",X"47",X"41",X"4D",X"45",X"20",X"53",X"54",X"59",X"4C",
		X"45",X"06",X"53",X"43",X"52",X"45",X"45",X"4E",X"06",X"45",X"58",X"54",X"45",X"4E",X"44",X"06",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"04",X"43",X"4F",X"49",X"4E",X"0A",X"44",X"49",X"46",X"46",
		X"49",X"43",X"55",X"4C",X"54",X"59",X"09",X"54",X"45",X"53",X"54",X"20",X"4D",X"4F",X"44",X"45",
		X"07",X"3A",X"20",X"55",X"50",X"20",X"20",X"20",X"07",X"3A",X"20",X"54",X"41",X"42",X"4C",X"45",
		X"08",X"3A",X"20",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"08",X"3A",X"20",X"49",X"4E",X"56",X"45",
		X"52",X"54",X"0F",X"3A",X"20",X"4F",X"4E",X"4C",X"59",X"20",X"32",X"30",X"30",X"30",X"30",X"20",
		X"20",X"20",X"0F",X"3A",X"20",X"32",X"30",X"30",X"30",X"30",X"20",X"45",X"20",X"36",X"30",X"30",
		X"30",X"30",X"03",X"3A",X"20",X"33",X"03",X"3A",X"20",X"35",X"0D",X"3A",X"20",X"31",X"43",X"4F",
		X"49",X"4E",X"20",X"31",X"50",X"4C",X"41",X"59",X"0D",X"3A",X"20",X"31",X"43",X"4F",X"49",X"4E",
		X"20",X"32",X"50",X"4C",X"41",X"59",X"0D",X"3A",X"20",X"32",X"43",X"4F",X"49",X"4E",X"20",X"31",
		X"50",X"4C",X"41",X"59",X"0D",X"3A",X"20",X"32",X"43",X"4F",X"49",X"4E",X"20",X"33",X"50",X"4C",
		X"41",X"59",X"04",X"3A",X"4F",X"4E",X"20",X"04",X"3A",X"4F",X"46",X"46",X"06",X"44",X"49",X"50",
		X"53",X"57",X"3A",X"0B",X"3A",X"20",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",X"54",X"0B",
		X"3A",X"20",X"45",X"41",X"53",X"59",X"20",X"20",X"20",X"20",X"20",X"10",X"53",X"43",X"52",X"45",
		X"45",X"4E",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"10",X"4F",X"42",X"4A",
		X"45",X"43",X"54",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"0E",X"57",X"4F",
		X"52",X"4B",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"06",X"42",X"41",X"44",
		X"20",X"48",X"57",X"08",X"52",X"41",X"4D",X"20",X"20",X"20",X"4F",X"4B",X"08",X"52",X"4F",X"4D",
		X"20",X"20",X"20",X"4F",X"4B",X"0A",X"53",X"4F",X"55",X"4E",X"44",X"20",X"43",X"4F",X"44",X"45",
		X"08",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4F",X"4B",X"0A",X"4C",X"3A",X"4F",X"4E",X"20",X"48",
		X"3A",X"4F",X"46",X"46",X"08",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"03",X"03",X"00",X"03",X"00",
		X"03",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"00",
		X"03",X"00",X"03",X"00",X"03",X"03",X"03",X"00",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"D0",X"21",X"CD",X"17",X"21",X"21",X"98",X"E6",
		X"11",X"A9",X"5C",X"AF",X"CD",X"C3",X"32",X"E7",X"CD",X"12",X"33",X"3E",X"01",X"32",X"D5",X"C4",
		X"01",X"E0",X"01",X"26",X"D0",X"2E",X"0C",X"E7",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",
		X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"CD",
		X"90",X"32",X"C2",X"36",X"32",X"0B",X"78",X"B1",X"20",X"DD",X"CD",X"D0",X"21",X"CD",X"17",X"21",
		X"3A",X"7B",X"C4",X"CB",X"F7",X"CB",X"EF",X"32",X"7B",X"C4",X"CD",X"D9",X"A5",X"E7",X"CD",X"35",
		X"A6",X"CD",X"95",X"32",X"3E",X"01",X"32",X"D5",X"C4",X"32",X"D0",X"C4",X"3E",X"07",X"F7",X"AF",
		X"32",X"00",X"EC",X"E7",X"CD",X"B0",X"A7",X"CD",X"74",X"A7",X"CD",X"90",X"32",X"C2",X"36",X"32",
		X"3A",X"B3",X"EF",X"FE",X"1E",X"20",X"EC",X"3E",X"00",X"32",X"D5",X"C4",X"E7",X"CD",X"17",X"21",
		X"3E",X"07",X"CF",X"21",X"18",X"31",X"11",X"45",X"34",X"01",X"17",X"00",X"1A",X"ED",X"A1",X"20",
		X"07",X"13",X"78",X"B1",X"20",X"F6",X"18",X"0D",X"21",X"00",X"E0",X"11",X"00",X"C0",X"01",X"FF",
		X"0F",X"ED",X"B0",X"18",X"0C",X"E7",X"3A",X"7B",X"C4",X"CB",X"B7",X"CB",X"AF",X"32",X"7B",X"C4",
		X"E7",X"ED",X"5F",X"E6",X"1F",X"32",X"72",X"ED",X"21",X"8B",X"ED",X"22",X"88",X"ED",X"AF",X"32",
		X"6F",X"ED",X"32",X"CE",X"C4",X"32",X"62",X"EF",X"3A",X"C1",X"C4",X"E6",X"20",X"07",X"07",X"07",
		X"21",X"28",X"9A",X"CD",X"50",X"20",X"7E",X"32",X"71",X"ED",X"CD",X"5B",X"96",X"3E",X"04",X"F7",
		X"01",X"B8",X"0B",X"E7",X"CD",X"90",X"32",X"20",X"4D",X"0B",X"78",X"B1",X"20",X"F5",X"3E",X"04",
		X"CF",X"3E",X"03",X"CF",X"3E",X"06",X"CF",X"AF",X"32",X"CE",X"C4",X"32",X"C4",X"C4",X"CD",X"17",
		X"21",X"CD",X"D0",X"21",X"E7",X"CD",X"F8",X"9E",X"01",X"E0",X"01",X"26",X"D0",X"2E",X"0C",X"CB",
		X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",
		X"20",X"7E",X"E1",X"32",X"18",X"D0",X"E7",X"CD",X"90",X"32",X"C2",X"36",X"32",X"0B",X"79",X"B0",
		X"20",X"DD",X"E7",X"C3",X"F7",X"30",X"3E",X"04",X"CF",X"3E",X"03",X"CF",X"3E",X"06",X"CF",X"3E",
		X"07",X"CF",X"AF",X"32",X"CE",X"C4",X"32",X"C4",X"C4",X"E7",X"CD",X"A8",X"32",X"CD",X"17",X"21",
		X"CD",X"D0",X"21",X"3A",X"7B",X"C4",X"CB",X"B7",X"CB",X"AF",X"32",X"7B",X"C4",X"3E",X"01",X"32",
		X"D0",X"C4",X"32",X"D5",X"C4",X"CD",X"C3",X"32",X"E7",X"CD",X"12",X"33",X"21",X"0F",X"32",X"11",
		X"45",X"34",X"01",X"17",X"00",X"1A",X"ED",X"A1",X"20",X"07",X"13",X"78",X"B1",X"20",X"F6",X"18",
		X"09",X"ED",X"5F",X"32",X"18",X"D0",X"3E",X"ED",X"ED",X"47",X"3E",X"00",X"D7",X"AF",X"DF",X"E7",
		X"3A",X"32",X"C4",X"A7",X"C9",X"3A",X"F7",X"C4",X"3D",X"32",X"F7",X"C4",X"11",X"B7",X"32",X"21",
		X"18",X"E5",X"AF",X"CD",X"F1",X"21",X"18",X"0B",X"11",X"B7",X"32",X"21",X"18",X"E5",X"CD",X"1C",
		X"22",X"3E",X"10",X"32",X"F7",X"C4",X"C9",X"0B",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"43",
		X"4F",X"49",X"4E",X"AF",X"32",X"FA",X"C4",X"21",X"00",X"90",X"01",X"00",X"10",X"3A",X"FA",X"C4",
		X"86",X"32",X"FA",X"C4",X"23",X"0B",X"78",X"B1",X"20",X"F3",X"3A",X"FA",X"C4",X"21",X"73",X"A5",
		X"BE",X"28",X"0C",X"3E",X"EA",X"ED",X"47",X"E7",X"3E",X"ED",X"ED",X"47",X"ED",X"46",X"E7",X"21",
		X"80",X"03",X"CD",X"D1",X"20",X"EB",X"21",X"CC",X"E0",X"0E",X"19",X"06",X"06",X"E5",X"3E",X"B0",
		X"B2",X"77",X"23",X"73",X"23",X"13",X"10",X"F6",X"E1",X"3E",X"40",X"CD",X"50",X"20",X"0D",X"20",
		X"EA",X"C9",X"3A",X"FF",X"BF",X"FE",X"76",X"28",X"48",X"FE",X"92",X"28",X"24",X"FE",X"33",X"28",
		X"0A",X"3E",X"ED",X"ED",X"47",X"ED",X"5E",X"E7",X"C3",X"45",X"23",X"11",X"2D",X"34",X"21",X"F2",
		X"E6",X"AF",X"CD",X"F1",X"21",X"11",X"D6",X"33",X"21",X"76",X"E6",X"AF",X"CD",X"F1",X"21",X"18",
		X"34",X"11",X"EA",X"33",X"21",X"32",X"E7",X"AF",X"CD",X"F1",X"21",X"11",X"05",X"34",X"21",X"B6",
		X"E6",X"AF",X"CD",X"F1",X"21",X"11",X"19",X"34",X"21",X"BA",X"E6",X"AF",X"CD",X"F1",X"21",X"18",
		X"14",X"11",X"BD",X"33",X"21",X"F2",X"E6",X"AF",X"CD",X"F1",X"21",X"11",X"D6",X"33",X"21",X"76",
		X"E6",X"AF",X"CD",X"F1",X"21",X"21",X"30",X"08",X"CD",X"D1",X"20",X"01",X"A3",X"33",X"3E",X"FF",
		X"32",X"F8",X"C4",X"3A",X"F8",X"C4",X"3C",X"32",X"F8",X"C4",X"FE",X"02",X"C8",X"E5",X"21",X"9F",
		X"33",X"CB",X"27",X"CD",X"56",X"20",X"E1",X"3A",X"F9",X"C4",X"CD",X"2B",X"22",X"18",X"E4",X"6C",
		X"E5",X"6E",X"E5",X"0C",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",
		X"0C",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"40",X"20",
		X"54",X"41",X"49",X"54",X"4F",X"20",X"43",X"4F",X"52",X"50",X"4F",X"52",X"41",X"54",X"49",X"4F",
		X"4E",X"20",X"31",X"39",X"38",X"36",X"13",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",
		X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"1A",X"40",X"20",X"31",X"39",X"38",
		X"36",X"20",X"54",X"41",X"49",X"54",X"4F",X"20",X"41",X"4D",X"45",X"52",X"49",X"43",X"41",X"20",
		X"43",X"4F",X"52",X"50",X"2E",X"13",X"4C",X"49",X"43",X"45",X"4E",X"53",X"45",X"44",X"20",X"54",
		X"4F",X"20",X"52",X"4F",X"4D",X"53",X"54",X"41",X"52",X"13",X"20",X"20",X"20",X"20",X"20",X"46",
		X"4F",X"52",X"20",X"55",X"2E",X"53",X"2E",X"41",X"20",X"20",X"20",X"20",X"20",X"17",X"40",X"20",
		X"31",X"39",X"38",X"36",X"20",X"54",X"41",X"49",X"54",X"4F",X"20",X"43",X"4F",X"52",X"50",X"20",
		X"4A",X"41",X"50",X"41",X"4E",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",
		X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"1A",X"00",X"00",X"FF",X"02",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"0E",X"00",X"FF",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",
		X"00",X"06",X"FF",X"00",X"00",X"FF",X"00",X"16",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"12",X"FF",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"0A",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"1E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B2",X"18",X"C7",X"00",X"1B",X"C6",X"00",X"1B",X"C7",X"00",
		X"10",X"15",X"02",X"B6",X"00",X"14",X"02",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",X"00",
		X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"AE",X"FF",X"BF",X"04",X"CB",X"00",X"1A",X"24",X"02",
		X"3C",X"10",X"B7",X"00",X"17",X"02",X"16",X"17",X"C7",X"00",X"19",X"01",X"02",X"FD",X"2F",X"FB",
		X"15",X"02",X"B6",X"00",X"14",X"02",X"4D",X"27",X"0A",X"C7",X"00",X"17",X"CB",X"00",X"10",X"97",
		X"C7",X"00",X"16",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",X"00",
		X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"27",X"0A",X"C7",X"00",X"17",X"CB",X"00",X"10",X"97",
		X"C7",X"00",X"16",X"01",X"02",X"FD",X"2F",X"17",X"C7",X"00",X"19",X"01",X"02",X"FD",X"2F",X"FB",
		X"15",X"02",X"B6",X"00",X"14",X"02",X"4D",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",X"00",
		X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",X"00",
		X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"27",X"0A",X"C7",X"00",X"17",X"CB",X"00",X"10",X"97",
		X"C7",X"00",X"16",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",X"00",
		X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"A6",X"FF",X"B7",X"02",X"A6",X"FC",X"B7",X"06",X"A6",
		X"00",X"B7",X"05",X"AE",X"80",X"3F",X"10",X"CB",X"00",X"10",X"C7",X"00",X"10",X"5C",X"26",X"F6",
		X"A6",X"FF",X"B7",X"E7",X"AF",X"32",X"65",X"C5",X"21",X"00",X"10",X"01",X"00",X"10",X"3A",X"65",
		X"C5",X"86",X"32",X"65",X"C5",X"23",X"0B",X"78",X"B1",X"20",X"F3",X"3A",X"65",X"C5",X"21",X"B4",
		X"23",X"BE",X"28",X"06",X"32",X"64",X"C5",X"32",X"33",X"C4",X"E7",X"3A",X"72",X"ED",X"FE",X"20",
		X"CA",X"09",X"88",X"3A",X"64",X"EF",X"A7",X"28",X"F1",X"3A",X"49",X"C5",X"CB",X"67",X"20",X"06",
		X"3C",X"32",X"49",X"C5",X"18",X"E4",X"CD",X"B4",X"3D",X"3A",X"64",X"EF",X"32",X"5C",X"C5",X"32",
		X"65",X"EF",X"AF",X"32",X"5E",X"C5",X"32",X"5D",X"C5",X"3A",X"64",X"EF",X"47",X"3E",X"03",X"90",
		X"A7",X"47",X"28",X"0F",X"DD",X"21",X"07",X"C5",X"DD",X"CB",X"0B",X"C6",X"11",X"14",X"00",X"DD",
		X"19",X"10",X"F5",X"3A",X"FD",X"C4",X"21",X"9D",X"36",X"CD",X"A8",X"3D",X"E9",X"A5",X"36",X"D0",
		X"37",X"FB",X"38",X"90",X"3A",X"E7",X"CD",X"3C",X"3C",X"DD",X"21",X"07",X"C5",X"21",X"FE",X"C4",
		X"22",X"FB",X"C4",X"21",X"85",X"4B",X"22",X"44",X"C5",X"21",X"00",X"17",X"22",X"46",X"C5",X"AF",
		X"32",X"5F",X"C5",X"3A",X"5E",X"C5",X"A7",X"28",X"15",X"DD",X"CB",X"0B",X"46",X"28",X"0F",X"3D",
		X"32",X"5E",X"C5",X"3A",X"65",X"EF",X"3C",X"32",X"65",X"EF",X"DD",X"CB",X"0B",X"86",X"DD",X"7E",
		X"0D",X"E6",X"22",X"C4",X"44",X"40",X"DD",X"CB",X"0B",X"46",X"C2",X"B2",X"37",X"DD",X"CB",X"0B",
		X"5E",X"20",X"06",X"DD",X"CB",X"0B",X"7E",X"20",X"06",X"CD",X"AE",X"3E",X"C3",X"B2",X"37",X"CD",
		X"7A",X"3C",X"D2",X"B2",X"37",X"CD",X"3B",X"3D",X"FD",X"7E",X"00",X"FE",X"28",X"30",X"0E",X"DD",
		X"36",X"11",X"00",X"DD",X"36",X"13",X"00",X"CD",X"53",X"3D",X"C3",X"8F",X"37",X"DD",X"CB",X"11",
		X"5E",X"20",X"55",X"DD",X"CB",X"11",X"FE",X"CD",X"07",X"47",X"CD",X"D4",X"4A",X"DA",X"8F",X"37",
		X"DD",X"36",X"11",X"00",X"DD",X"CB",X"11",X"DE",X"DD",X"34",X"02",X"3E",X"10",X"DD",X"BE",X"02",
		X"20",X"04",X"DD",X"36",X"02",X"0F",X"FD",X"7E",X"01",X"FE",X"78",X"38",X"04",X"DD",X"CB",X"11",
		X"D6",X"DD",X"CB",X"11",X"56",X"28",X"05",X"21",X"DB",X"4C",X"18",X"03",X"21",X"0D",X"4D",X"7E",
		X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"12",X"DD",X"36",X"13",X"00",X"21",X"0D",X"4D",X"22",
		X"60",X"C5",X"21",X"DB",X"4C",X"22",X"62",X"C5",X"CD",X"0C",X"4B",X"CD",X"BB",X"3B",X"30",X"0F",
		X"21",X"0D",X"4D",X"22",X"60",X"C5",X"21",X"DB",X"4C",X"22",X"62",X"C5",X"CD",X"F5",X"3B",X"FD",
		X"E5",X"E1",X"CD",X"4A",X"11",X"E5",X"FD",X"E1",X"CD",X"DE",X"42",X"FD",X"7E",X"00",X"FE",X"F8",
		X"30",X"08",X"2A",X"FB",X"C4",X"CD",X"29",X"3E",X"18",X"05",X"CD",X"F6",X"3C",X"18",X"03",X"CD",
		X"41",X"3E",X"11",X"03",X"00",X"2A",X"FB",X"C4",X"19",X"22",X"FB",X"C4",X"11",X"14",X"00",X"DD",
		X"19",X"3A",X"5F",X"C5",X"3C",X"32",X"5F",X"C5",X"FE",X"03",X"CA",X"A5",X"36",X"C3",X"C3",X"36",
		X"E7",X"CD",X"3C",X"3C",X"DD",X"21",X"07",X"C5",X"21",X"FE",X"C4",X"22",X"FB",X"C4",X"21",X"A7",
		X"4B",X"22",X"44",X"C5",X"21",X"A0",X"15",X"22",X"46",X"C5",X"AF",X"32",X"5F",X"C5",X"3A",X"5E",
		X"C5",X"A7",X"28",X"15",X"DD",X"CB",X"0B",X"46",X"28",X"0F",X"3D",X"32",X"5E",X"C5",X"3A",X"65",
		X"EF",X"3C",X"32",X"65",X"EF",X"DD",X"CB",X"0B",X"86",X"DD",X"7E",X"0D",X"E6",X"22",X"C4",X"44",
		X"40",X"DD",X"CB",X"0B",X"46",X"C2",X"DD",X"38",X"DD",X"CB",X"0B",X"5E",X"20",X"06",X"DD",X"CB",
		X"0B",X"7E",X"20",X"06",X"CD",X"AE",X"3E",X"C3",X"DD",X"38",X"CD",X"7A",X"3C",X"D2",X"DD",X"38",
		X"CD",X"3B",X"3D",X"FD",X"7E",X"00",X"FE",X"28",X"30",X"0E",X"DD",X"36",X"11",X"00",X"DD",X"36",
		X"13",X"00",X"CD",X"53",X"3D",X"C3",X"BA",X"38",X"DD",X"CB",X"11",X"5E",X"20",X"55",X"DD",X"CB",
		X"11",X"FE",X"CD",X"07",X"47",X"CD",X"D4",X"4A",X"DA",X"BA",X"38",X"DD",X"36",X"11",X"00",X"DD",
		X"CB",X"11",X"DE",X"DD",X"35",X"02",X"3E",X"00",X"DD",X"BE",X"02",X"20",X"04",X"DD",X"36",X"02",
		X"01",X"FD",X"7E",X"01",X"FE",X"78",X"38",X"04",X"DD",X"CB",X"11",X"D6",X"DD",X"CB",X"11",X"56",
		X"28",X"05",X"21",X"7B",X"4D",X"18",X"03",X"21",X"5B",X"4D",X"7E",X"DD",X"77",X"03",X"23",X"7E",
		X"DD",X"77",X"12",X"DD",X"36",X"13",X"00",X"21",X"5B",X"4D",X"22",X"60",X"C5",X"21",X"7B",X"4D",
		X"22",X"62",X"C5",X"CD",X"0C",X"4B",X"CD",X"BB",X"3B",X"30",X"0F",X"21",X"5B",X"4D",X"22",X"60",
		X"C5",X"21",X"7B",X"4D",X"22",X"62",X"C5",X"CD",X"F5",X"3B",X"FD",X"E5",X"E1",X"CD",X"4A",X"11",
		X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",X"F8",X"30",X"0B",X"CD",X"DE",X"42",X"2A",X"FB",X"C4",
		X"CD",X"29",X"3E",X"18",X"05",X"CD",X"F6",X"3C",X"18",X"03",X"CD",X"41",X"3E",X"11",X"03",X"00",
		X"2A",X"FB",X"C4",X"19",X"22",X"FB",X"C4",X"11",X"14",X"00",X"DD",X"19",X"3A",X"5F",X"C5",X"3C",
		X"32",X"5F",X"C5",X"FE",X"03",X"CA",X"D0",X"37",X"C3",X"EE",X"37",X"E7",X"CD",X"3C",X"3C",X"DD",
		X"21",X"07",X"C5",X"21",X"FE",X"C4",X"22",X"FB",X"C4",X"21",X"D9",X"4B",X"22",X"44",X"C5",X"21",
		X"A0",X"12",X"22",X"46",X"C5",X"21",X"77",X"4B",X"22",X"4A",X"C5",X"3E",X"08",X"32",X"4C",X"C5",
		X"AF",X"32",X"5F",X"C5",X"3A",X"5E",X"C5",X"A7",X"28",X"15",X"DD",X"CB",X"0B",X"46",X"28",X"0F",
		X"3D",X"32",X"5E",X"C5",X"3A",X"65",X"EF",X"3C",X"32",X"65",X"EF",X"DD",X"CB",X"0B",X"86",X"DD",
		X"7E",X"0D",X"E6",X"22",X"C4",X"44",X"40",X"DD",X"CB",X"0B",X"46",X"C2",X"72",X"3A",X"DD",X"CB",
		X"0B",X"5E",X"20",X"06",X"DD",X"CB",X"0B",X"7E",X"20",X"06",X"CD",X"AE",X"3E",X"C3",X"72",X"3A",
		X"CD",X"7A",X"3C",X"D2",X"72",X"3A",X"DD",X"CB",X"0B",X"56",X"20",X"34",X"2A",X"FB",X"C4",X"CB",
		X"66",X"28",X"61",X"D5",X"11",X"50",X"00",X"CD",X"23",X"27",X"D1",X"3E",X"8E",X"A6",X"77",X"DD",
		X"CB",X"0B",X"D6",X"21",X"77",X"4B",X"7E",X"DD",X"77",X"0E",X"23",X"DD",X"77",X"0F",X"3E",X"08",
		X"DD",X"77",X"0C",X"DD",X"36",X"10",X"00",X"2A",X"46",X"C5",X"CD",X"73",X"3E",X"C3",X"72",X"3A",
		X"DD",X"35",X"0E",X"C2",X"72",X"3A",X"DD",X"34",X"10",X"DD",X"7E",X"10",X"CB",X"27",X"21",X"77",
		X"4B",X"16",X"00",X"5F",X"19",X"7E",X"FE",X"FF",X"28",X"14",X"DD",X"77",X"0E",X"23",X"7E",X"DD",
		X"77",X"0F",X"DD",X"34",X"0C",X"2A",X"46",X"C5",X"CD",X"73",X"3E",X"C3",X"72",X"3A",X"CD",X"F6",
		X"3C",X"C3",X"72",X"3A",X"CD",X"3B",X"3D",X"FD",X"7E",X"00",X"FE",X"28",X"30",X"0E",X"DD",X"36",
		X"11",X"00",X"DD",X"36",X"13",X"00",X"CD",X"53",X"3D",X"C3",X"4F",X"3A",X"DD",X"CB",X"11",X"5E",
		X"20",X"46",X"DD",X"CB",X"11",X"FE",X"CD",X"07",X"47",X"CD",X"D4",X"4A",X"38",X"51",X"DD",X"36",
		X"11",X"00",X"DD",X"CB",X"11",X"DE",X"FD",X"7E",X"01",X"FE",X"78",X"38",X"04",X"DD",X"CB",X"11",
		X"D6",X"DD",X"CB",X"11",X"56",X"28",X"05",X"21",X"AB",X"4D",X"18",X"03",X"21",X"9B",X"4D",X"7E",
		X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"12",X"DD",X"36",X"13",X"00",X"21",X"9B",X"4D",X"22",
		X"60",X"C5",X"21",X"AB",X"4D",X"22",X"62",X"C5",X"CD",X"0C",X"4B",X"CD",X"BB",X"3B",X"30",X"0F",
		X"21",X"9B",X"4D",X"22",X"60",X"C5",X"21",X"AB",X"4D",X"22",X"62",X"C5",X"CD",X"F5",X"3B",X"FD",
		X"E5",X"E1",X"CD",X"4A",X"11",X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",X"F8",X"30",X"0B",X"CD",
		X"DE",X"42",X"2A",X"FB",X"C4",X"CD",X"29",X"3E",X"18",X"05",X"CD",X"F6",X"3C",X"18",X"03",X"CD",
		X"41",X"3E",X"11",X"03",X"00",X"2A",X"FB",X"C4",X"19",X"22",X"FB",X"C4",X"11",X"14",X"00",X"DD",
		X"19",X"3A",X"5F",X"C5",X"3C",X"32",X"5F",X"C5",X"FE",X"03",X"CA",X"FB",X"38",X"C3",X"24",X"39",
		X"E7",X"CD",X"3C",X"3C",X"DD",X"21",X"07",X"C5",X"21",X"FE",X"C4",X"22",X"FB",X"C4",X"21",X"3B",
		X"4C",X"22",X"44",X"C5",X"21",X"60",X"14",X"22",X"46",X"C5",X"AF",X"32",X"5F",X"C5",X"3A",X"5E",
		X"C5",X"A7",X"28",X"15",X"DD",X"CB",X"0B",X"46",X"28",X"0F",X"3D",X"32",X"5E",X"C5",X"3A",X"65",
		X"EF",X"3C",X"32",X"65",X"EF",X"DD",X"CB",X"0B",X"86",X"DD",X"7E",X"0D",X"E6",X"22",X"C4",X"44",
		X"40",X"DD",X"CB",X"0B",X"46",X"C2",X"9D",X"3B",X"DD",X"CB",X"0B",X"5E",X"20",X"06",X"DD",X"CB",
		X"0B",X"7E",X"20",X"06",X"CD",X"AE",X"3E",X"C3",X"9D",X"3B",X"CD",X"7A",X"3C",X"D2",X"9D",X"3B",
		X"CD",X"3B",X"3D",X"FD",X"7E",X"00",X"FE",X"28",X"30",X"0E",X"DD",X"36",X"11",X"00",X"DD",X"36",
		X"13",X"00",X"CD",X"53",X"3D",X"C3",X"7A",X"3B",X"DD",X"CB",X"11",X"5E",X"20",X"55",X"DD",X"CB",
		X"11",X"FE",X"CD",X"07",X"47",X"CD",X"D4",X"4A",X"DA",X"7A",X"3B",X"DD",X"36",X"11",X"00",X"DD",
		X"CB",X"11",X"DE",X"DD",X"34",X"02",X"3E",X"0F",X"DD",X"BE",X"02",X"20",X"04",X"DD",X"36",X"02",
		X"0F",X"FD",X"7E",X"01",X"FE",X"78",X"38",X"04",X"DD",X"CB",X"11",X"D6",X"DD",X"CB",X"11",X"56",
		X"28",X"05",X"21",X"DD",X"4D",X"18",X"03",X"21",X"BB",X"4D",X"7E",X"DD",X"77",X"03",X"23",X"7E",
		X"DD",X"77",X"12",X"DD",X"36",X"13",X"00",X"21",X"BB",X"4D",X"22",X"60",X"C5",X"21",X"DD",X"4D",
		X"22",X"62",X"C5",X"CD",X"0C",X"4B",X"CD",X"BB",X"3B",X"30",X"0F",X"21",X"BB",X"4D",X"22",X"60",
		X"C5",X"21",X"DD",X"4D",X"22",X"62",X"C5",X"CD",X"F5",X"3B",X"FD",X"E5",X"E1",X"CD",X"4A",X"11",
		X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",X"F8",X"30",X"0B",X"CD",X"DE",X"42",X"2A",X"FB",X"C4",
		X"CD",X"29",X"3E",X"18",X"05",X"CD",X"F6",X"3C",X"18",X"03",X"CD",X"41",X"3E",X"11",X"03",X"00",
		X"2A",X"FB",X"C4",X"19",X"22",X"FB",X"C4",X"11",X"14",X"00",X"DD",X"19",X"3A",X"5F",X"C5",X"3C",
		X"32",X"5F",X"C5",X"FE",X"03",X"CA",X"90",X"3A",X"C3",X"AE",X"3A",X"DD",X"CB",X"11",X"46",X"20",
		X"23",X"FD",X"7E",X"04",X"FE",X"B8",X"D8",X"DD",X"CB",X"11",X"C6",X"DD",X"36",X"13",X"00",X"21",
		X"4D",X"4D",X"DD",X"CB",X"11",X"56",X"28",X"03",X"21",X"3F",X"4D",X"7E",X"DD",X"77",X"03",X"23",
		X"7E",X"DD",X"77",X"12",X"21",X"4D",X"4D",X"22",X"60",X"C5",X"21",X"3F",X"4D",X"22",X"62",X"C5",
		X"CD",X"F5",X"3B",X"A7",X"C9",X"DD",X"7E",X"12",X"DD",X"96",X"02",X"DD",X"77",X"12",X"D0",X"DD",
		X"34",X"13",X"DD",X"CB",X"11",X"56",X"28",X"05",X"2A",X"62",X"C5",X"18",X"03",X"2A",X"60",X"C5",
		X"DD",X"7E",X"13",X"CB",X"27",X"5F",X"16",X"00",X"19",X"3E",X"FF",X"BE",X"20",X"14",X"DD",X"CB",
		X"11",X"56",X"28",X"05",X"2A",X"62",X"C5",X"18",X"03",X"2A",X"60",X"C5",X"DD",X"36",X"13",X"00",
		X"18",X"00",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"77",X"12",X"C9",X"3A",X"64",X"EF",X"F5",
		X"3A",X"5C",X"C5",X"47",X"F1",X"F5",X"B8",X"28",X"18",X"30",X"19",X"C1",X"3A",X"5C",X"C5",X"32",
		X"65",X"EF",X"90",X"32",X"5D",X"C5",X"3A",X"64",X"EF",X"32",X"5C",X"C5",X"AF",X"32",X"5E",X"C5",
		X"C9",X"F1",X"AF",X"C9",X"3A",X"5C",X"C5",X"32",X"65",X"EF",X"F1",X"90",X"32",X"5E",X"C5",X"3A",
		X"64",X"EF",X"32",X"5C",X"C5",X"AF",X"32",X"5D",X"C5",X"C9",X"DD",X"CB",X"0B",X"76",X"20",X"46",
		X"2A",X"FB",X"C4",X"CB",X"46",X"28",X"08",X"CB",X"6E",X"20",X"09",X"CB",X"76",X"20",X"05",X"AF",
		X"37",X"C9",X"AF",X"C9",X"D5",X"11",X"10",X"00",X"CD",X"23",X"27",X"3E",X"14",X"CD",X"AE",X"67",
		X"D1",X"3E",X"8E",X"A6",X"77",X"DD",X"CB",X"0B",X"F6",X"21",X"8D",X"4C",X"7E",X"DD",X"77",X"0E",
		X"23",X"7E",X"DD",X"77",X"0F",X"23",X"7E",X"DD",X"77",X"0C",X"DD",X"36",X"10",X"00",X"21",X"E0",
		X"1B",X"CD",X"73",X"3E",X"AF",X"C9",X"DD",X"35",X"0E",X"20",X"C7",X"DD",X"34",X"10",X"DD",X"7E",
		X"10",X"CB",X"27",X"CB",X"27",X"21",X"8D",X"4C",X"16",X"00",X"5F",X"19",X"7E",X"FE",X"FF",X"28",
		X"15",X"DD",X"77",X"0E",X"23",X"7E",X"DD",X"77",X"0F",X"23",X"7E",X"DD",X"77",X"0C",X"21",X"E0",
		X"1B",X"CD",X"73",X"3E",X"AF",X"C9",X"CD",X"3B",X"3D",X"FD",X"E5",X"E1",X"06",X"08",X"36",X"00",
		X"23",X"10",X"FB",X"3E",X"30",X"DD",X"A6",X"0B",X"DD",X"77",X"0B",X"DD",X"36",X"11",X"00",X"DD",
		X"7E",X"0D",X"E6",X"22",X"DD",X"77",X"0D",X"2A",X"FB",X"C4",X"3E",X"8E",X"A6",X"77",X"23",X"36",
		X"00",X"23",X"36",X"00",X"3A",X"5D",X"C5",X"A7",X"28",X"0F",X"3D",X"32",X"5D",X"C5",X"3A",X"65",
		X"EF",X"3D",X"32",X"65",X"EF",X"DD",X"CB",X"0B",X"C6",X"AF",X"C9",X"DD",X"7E",X"0B",X"E6",X"30",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3D",X"21",X"71",X"4B",X"CD",X"A8",X"3D",X"E5",
		X"FD",X"E1",X"C9",X"FD",X"7E",X"01",X"FE",X"D9",X"38",X"13",X"ED",X"5F",X"E6",X"1F",X"CB",X"E7",
		X"DD",X"77",X"03",X"FD",X"36",X"01",X"D8",X"FD",X"36",X"05",X"D8",X"18",X"15",X"FE",X"17",X"30",
		X"11",X"ED",X"5F",X"E6",X"1F",X"CB",X"A7",X"DD",X"77",X"03",X"FD",X"36",X"01",X"18",X"FD",X"36",
		X"05",X"18",X"FD",X"7E",X"04",X"FE",X"19",X"D0",X"DD",X"7E",X"03",X"A7",X"20",X"04",X"ED",X"5F",
		X"E6",X"1F",X"CB",X"67",X"20",X"04",X"CB",X"DF",X"18",X"02",X"CB",X"9F",X"DD",X"77",X"03",X"FD",
		X"36",X"04",X"18",X"FD",X"36",X"00",X"20",X"C9",X"D5",X"07",X"16",X"00",X"5F",X"19",X"5E",X"23",
		X"56",X"EB",X"D1",X"C9",X"21",X"89",X"C4",X"11",X"8A",X"C4",X"01",X"17",X"00",X"36",X"00",X"ED",
		X"B0",X"21",X"07",X"C5",X"11",X"08",X"C5",X"01",X"3C",X"00",X"36",X"00",X"ED",X"B0",X"21",X"54",
		X"C5",X"11",X"55",X"C5",X"01",X"07",X"00",X"36",X"00",X"ED",X"B0",X"3E",X"00",X"32",X"67",X"C5",
		X"32",X"49",X"C5",X"3A",X"72",X"ED",X"E6",X"03",X"32",X"FD",X"C4",X"FE",X"03",X"20",X"02",X"C6",
		X"02",X"4F",X"3E",X"00",X"32",X"43",X"C5",X"79",X"FD",X"21",X"FE",X"C4",X"DD",X"21",X"07",X"C5",
		X"06",X"03",X"FD",X"77",X"00",X"F5",X"FD",X"77",X"01",X"FD",X"77",X"02",X"32",X"49",X"C5",X"3A",
		X"43",X"C5",X"0E",X"10",X"81",X"DD",X"77",X"0B",X"32",X"43",X"C5",X"F1",X"11",X"14",X"00",X"DD",
		X"19",X"11",X"03",X"00",X"FD",X"19",X"10",X"DA",X"C9",X"F5",X"DD",X"E5",X"E5",X"DD",X"E1",X"FD",
		X"7E",X"01",X"D6",X"08",X"DD",X"77",X"01",X"FD",X"7E",X"04",X"DD",X"77",X"02",X"DD",X"E1",X"F1",
		X"C9",X"DD",X"35",X"0E",X"C0",X"DD",X"34",X"10",X"DD",X"7E",X"10",X"2A",X"44",X"C5",X"CB",X"27",
		X"CB",X"27",X"16",X"00",X"5F",X"19",X"3E",X"FF",X"BE",X"20",X"07",X"2A",X"44",X"C5",X"DD",X"36",
		X"10",X"00",X"7E",X"DD",X"77",X"0E",X"23",X"7E",X"DD",X"77",X"0F",X"23",X"7E",X"DD",X"77",X"0C",
		X"2A",X"46",X"C5",X"FD",X"E5",X"D5",X"E5",X"CD",X"3B",X"3D",X"E1",X"CD",X"BA",X"20",X"DD",X"7E",
		X"0C",X"CB",X"27",X"16",X"00",X"5F",X"19",X"7D",X"FD",X"77",X"07",X"DD",X"7E",X"0F",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"84",X"FD",X"77",X"06",X"23",X"7D",X"FD",X"77",X"03",X"DD",X"7E",X"0F",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"84",X"FD",X"77",X"02",X"D1",X"FD",X"E1",X"C9",X"FD",X"21",
		X"54",X"C5",X"DD",X"CB",X"0D",X"46",X"C2",X"E9",X"3E",X"DD",X"CB",X"0D",X"66",X"C2",X"71",X"3F",
		X"DD",X"CB",X"0B",X"5E",X"C2",X"DF",X"3F",X"3A",X"3B",X"C4",X"FE",X"78",X"DA",X"57",X"3F",X"3A",
		X"54",X"C5",X"E6",X"0F",X"C0",X"3A",X"54",X"C5",X"CB",X"C7",X"32",X"54",X"C5",X"DD",X"CB",X"0D",
		X"C6",X"FD",X"36",X"02",X"FF",X"FD",X"36",X"01",X"01",X"FD",X"35",X"01",X"C0",X"FD",X"34",X"02",
		X"FD",X"7E",X"02",X"21",X"AB",X"4C",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"19",X"3E",X"FF",
		X"BE",X"CA",X"1E",X"3F",X"7E",X"FD",X"77",X"01",X"23",X"7E",X"FD",X"77",X"06",X"23",X"7E",X"FD",
		X"77",X"05",X"DD",X"E5",X"DD",X"21",X"82",X"E2",X"CD",X"D3",X"40",X"DD",X"E1",X"C9",X"DD",X"CB",
		X"0D",X"86",X"DD",X"CB",X"0B",X"DE",X"DD",X"36",X"10",X"FF",X"DD",X"36",X"0E",X"01",X"CD",X"41",
		X"3E",X"CD",X"3B",X"3D",X"FD",X"36",X"00",X"18",X"FD",X"36",X"04",X"10",X"FD",X"36",X"01",X"B0",
		X"FD",X"36",X"05",X"B0",X"DD",X"36",X"03",X"10",X"DD",X"36",X"04",X"02",X"3E",X"01",X"DD",X"77",
		X"02",X"2A",X"FB",X"C4",X"CB",X"C6",X"C9",X"3A",X"54",X"C5",X"E6",X"F0",X"C0",X"3A",X"54",X"C5",
		X"CB",X"E7",X"32",X"54",X"C5",X"DD",X"CB",X"0D",X"E6",X"FD",X"36",X"04",X"FF",X"FD",X"36",X"03",
		X"01",X"FD",X"35",X"03",X"C0",X"FD",X"34",X"04",X"FD",X"7E",X"04",X"21",X"AB",X"4C",X"CB",X"27",
		X"CB",X"27",X"16",X"00",X"5F",X"19",X"3E",X"FF",X"BE",X"CA",X"A6",X"3F",X"7E",X"FD",X"77",X"03",
		X"23",X"7E",X"FD",X"77",X"06",X"23",X"7E",X"FD",X"77",X"05",X"DD",X"E5",X"DD",X"21",X"02",X"E6",
		X"CD",X"D3",X"40",X"DD",X"E1",X"C9",X"DD",X"CB",X"0D",X"A6",X"DD",X"CB",X"0B",X"DE",X"DD",X"36",
		X"10",X"FF",X"DD",X"36",X"0E",X"01",X"CD",X"41",X"3E",X"CD",X"3B",X"3D",X"FD",X"36",X"00",X"18",
		X"FD",X"36",X"04",X"10",X"FD",X"36",X"01",X"40",X"FD",X"36",X"05",X"40",X"DD",X"36",X"03",X"10",
		X"DD",X"36",X"04",X"02",X"3E",X"01",X"DD",X"77",X"02",X"2A",X"FB",X"C4",X"CB",X"C6",X"C9",X"CD",
		X"41",X"3E",X"CD",X"3B",X"3D",X"FD",X"E5",X"E1",X"CD",X"4A",X"11",X"E5",X"FD",X"E1",X"2A",X"FB",
		X"C4",X"CD",X"29",X"3E",X"3E",X"18",X"FD",X"BE",X"04",X"38",X"01",X"C9",X"ED",X"5F",X"E6",X"1F",
		X"DD",X"77",X"03",X"DD",X"CB",X"0B",X"9E",X"DD",X"CB",X"0B",X"FE",X"FD",X"7E",X"01",X"FE",X"78",
		X"38",X"19",X"3A",X"54",X"C5",X"CB",X"CF",X"32",X"54",X"C5",X"DD",X"CB",X"0D",X"CE",X"FD",X"21",
		X"54",X"C5",X"FD",X"36",X"02",X"FF",X"FD",X"36",X"01",X"01",X"C9",X"3A",X"54",X"C5",X"CB",X"EF",
		X"32",X"54",X"C5",X"DD",X"CB",X"0D",X"EE",X"FD",X"21",X"54",X"C5",X"FD",X"36",X"04",X"FF",X"FD",
		X"36",X"03",X"01",X"C9",X"FD",X"21",X"54",X"C5",X"DD",X"CB",X"0D",X"6E",X"C2",X"84",X"40",X"FD",
		X"35",X"01",X"C0",X"FD",X"34",X"02",X"FD",X"7E",X"02",X"21",X"C1",X"4C",X"CB",X"27",X"CB",X"27",
		X"16",X"00",X"5F",X"19",X"3E",X"FF",X"BE",X"CA",X"B9",X"40",X"7E",X"FD",X"77",X"01",X"23",X"7E",
		X"FD",X"77",X"06",X"23",X"7E",X"FD",X"77",X"05",X"DD",X"E5",X"DD",X"21",X"82",X"E2",X"CD",X"D3",
		X"40",X"DD",X"E1",X"C9",X"FD",X"35",X"03",X"C0",X"FD",X"34",X"04",X"FD",X"7E",X"04",X"21",X"C1",
		X"4C",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"19",X"3E",X"FF",X"BE",X"CA",X"C6",X"40",X"7E",
		X"FD",X"77",X"03",X"23",X"7E",X"FD",X"77",X"06",X"23",X"7E",X"FD",X"77",X"05",X"DD",X"E5",X"DD",
		X"21",X"02",X"E6",X"CD",X"D3",X"40",X"DD",X"E1",X"C9",X"3A",X"54",X"C5",X"E6",X"F0",X"32",X"54",
		X"C5",X"DD",X"36",X"0D",X"00",X"C9",X"3A",X"54",X"C5",X"E6",X"0F",X"32",X"54",X"C5",X"DD",X"36",
		X"0D",X"00",X"C9",X"E5",X"D5",X"C5",X"21",X"F0",X"08",X"CD",X"D1",X"20",X"FD",X"7E",X"05",X"16",
		X"00",X"5F",X"19",X"11",X"40",X"00",X"06",X"04",X"7D",X"DD",X"77",X"03",X"FD",X"7E",X"06",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"84",X"DD",X"77",X"02",X"23",X"E5",X"DD",X"E5",X"E1",X"ED",X"52",
		X"E5",X"DD",X"E1",X"E1",X"10",X"E2",X"C1",X"D1",X"E1",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",
		X"1D",X"1D",X"00",X"01",X"01",X"01",X"00",X"1D",X"1D",X"1D",X"00",X"00",X"19",X"19",X"19",X"00",
		X"05",X"05",X"05",X"00",X"19",X"19",X"19",X"00",X"00",X"15",X"15",X"15",X"00",X"09",X"0A",X"09",
		X"00",X"15",X"15",X"15",X"00",X"00",X"11",X"11",X"11",X"00",X"0D",X"0D",X"0D",X"00",X"11",X"11",
		X"11",X"00",X"00",X"0D",X"0E",X"0D",X"00",X"11",X"12",X"11",X"00",X"0D",X"0E",X"0D",X"00",X"00",
		X"09",X"09",X"09",X"00",X"15",X"15",X"15",X"00",X"09",X"09",X"09",X"00",X"00",X"05",X"05",X"05",
		X"00",X"19",X"19",X"19",X"00",X"05",X"05",X"05",X"00",X"00",X"01",X"02",X"01",X"00",X"1D",X"1D",
		X"1D",X"00",X"01",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"15",X"15",X"15",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"15",X"15",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"16",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"06",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"0A",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"12",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"3A",X"5F",
		X"C5",X"21",X"6B",X"4B",X"CD",X"A8",X"3D",X"E9",X"3A",X"18",X"C5",X"CB",X"5F",X"C0",X"3A",X"2C",
		X"C5",X"CB",X"5F",X"C0",X"3A",X"14",X"C5",X"E6",X"11",X"28",X"12",X"ED",X"5B",X"91",X"C4",X"CD",
		X"E7",X"44",X"30",X"76",X"3A",X"67",X"C5",X"CB",X"47",X"20",X"79",X"18",X"5D",X"3A",X"28",X"C5",
		X"E6",X"11",X"28",X"11",X"2A",X"89",X"C4",X"CD",X"FB",X"44",X"30",X"5E",X"3A",X"67",X"C5",X"CB",
		X"47",X"20",X"61",X"18",X"4D",X"2A",X"89",X"C4",X"ED",X"5B",X"91",X"C4",X"CD",X"CA",X"45",X"30",
		X"49",X"3A",X"67",X"C5",X"CB",X"47",X"20",X"4C",X"3A",X"12",X"C5",X"CB",X"5F",X"20",X"2B",X"3A",
		X"26",X"C5",X"CB",X"5F",X"20",X"2C",X"21",X"0A",X"C5",X"11",X"1E",X"C5",X"CD",X"F6",X"45",X"21",
		X"18",X"C5",X"11",X"2C",X"C5",X"FD",X"E5",X"FD",X"21",X"1B",X"C5",X"CD",X"0F",X"45",X"FD",X"E1",
		X"3A",X"67",X"C5",X"CB",X"C7",X"32",X"67",X"C5",X"18",X"2C",X"11",X"1E",X"C5",X"CD",X"40",X"46",
		X"18",X"DD",X"21",X"0A",X"C5",X"CD",X"7C",X"46",X"18",X"D5",X"3A",X"67",X"C5",X"CB",X"87",X"32",
		X"67",X"C5",X"18",X"12",X"3A",X"0A",X"C5",X"47",X"3A",X"1E",X"C5",X"90",X"30",X"02",X"2F",X"3C",
		X"FE",X"03",X"30",X"02",X"18",X"B0",X"3A",X"40",X"C5",X"CB",X"5F",X"C0",X"3A",X"14",X"C5",X"E6",
		X"11",X"28",X"12",X"ED",X"5B",X"99",X"C4",X"CD",X"E7",X"44",X"30",X"75",X"3A",X"67",X"C5",X"CB",
		X"4F",X"20",X"77",X"18",X"5C",X"3A",X"3C",X"C5",X"E6",X"11",X"28",X"11",X"2A",X"89",X"C4",X"CD",
		X"FB",X"44",X"30",X"5D",X"3A",X"67",X"C5",X"CB",X"4F",X"20",X"5F",X"18",X"4C",X"2A",X"89",X"C4",
		X"ED",X"5B",X"99",X"C4",X"CD",X"CA",X"45",X"30",X"48",X"3A",X"67",X"C5",X"CB",X"4F",X"20",X"4A",
		X"3A",X"12",X"C5",X"CB",X"5F",X"20",X"2A",X"3A",X"3A",X"C5",X"CB",X"5F",X"20",X"2B",X"21",X"0A",
		X"C5",X"11",X"32",X"C5",X"CD",X"F6",X"45",X"21",X"18",X"C5",X"11",X"40",X"C5",X"FD",X"E5",X"FD",
		X"21",X"2F",X"C5",X"CD",X"0F",X"45",X"FD",X"E1",X"3A",X"67",X"C5",X"CB",X"CF",X"32",X"67",X"C5",
		X"C9",X"11",X"32",X"C5",X"CD",X"40",X"46",X"18",X"DE",X"21",X"0A",X"C5",X"CD",X"7C",X"46",X"18",
		X"D6",X"3A",X"67",X"C5",X"CB",X"8F",X"32",X"67",X"C5",X"C9",X"3A",X"0A",X"C5",X"47",X"3A",X"32",
		X"C5",X"90",X"30",X"02",X"2F",X"3C",X"FE",X"03",X"D0",X"18",X"B3",X"3A",X"2C",X"C5",X"CB",X"5F",
		X"C0",X"3A",X"40",X"C5",X"CB",X"5F",X"C0",X"3A",X"28",X"C5",X"E6",X"11",X"28",X"12",X"ED",X"5B",
		X"99",X"C4",X"CD",X"E7",X"44",X"30",X"75",X"3A",X"67",X"C5",X"CB",X"57",X"20",X"77",X"18",X"5C",
		X"3A",X"3C",X"C5",X"E6",X"11",X"28",X"11",X"2A",X"91",X"C4",X"CD",X"FB",X"44",X"30",X"5D",X"3A",
		X"67",X"C5",X"CB",X"57",X"20",X"5F",X"18",X"4C",X"2A",X"91",X"C4",X"ED",X"5B",X"99",X"C4",X"CD",
		X"CA",X"45",X"30",X"48",X"3A",X"67",X"C5",X"CB",X"57",X"20",X"4A",X"3A",X"26",X"C5",X"CB",X"5F",
		X"20",X"2A",X"3A",X"3A",X"C5",X"CB",X"5F",X"20",X"2B",X"21",X"1E",X"C5",X"11",X"32",X"C5",X"CD",
		X"F6",X"45",X"21",X"2C",X"C5",X"11",X"40",X"C5",X"FD",X"E5",X"FD",X"21",X"2F",X"C5",X"CD",X"0F",
		X"45",X"FD",X"E1",X"3A",X"67",X"C5",X"CB",X"D7",X"32",X"67",X"C5",X"C9",X"11",X"32",X"C5",X"CD",
		X"40",X"46",X"18",X"DE",X"21",X"1E",X"C5",X"CD",X"7C",X"46",X"18",X"D6",X"3A",X"67",X"C5",X"CB",
		X"97",X"32",X"67",X"C5",X"C9",X"3A",X"1E",X"C5",X"47",X"3A",X"32",X"C5",X"90",X"30",X"02",X"2F",
		X"3C",X"FE",X"03",X"D0",X"18",X"B3",X"C9",X"CB",X"47",X"20",X"08",X"26",X"40",X"2E",X"18",X"CD",
		X"CA",X"45",X"C9",X"26",X"B0",X"2E",X"18",X"CD",X"CA",X"45",X"C9",X"CB",X"47",X"20",X"08",X"16",
		X"40",X"1E",X"18",X"CD",X"CA",X"45",X"C9",X"16",X"B0",X"1E",X"18",X"CD",X"CA",X"45",X"C9",X"7E",
		X"CB",X"5F",X"C2",X"8A",X"45",X"CB",X"7F",X"CA",X"6B",X"45",X"E6",X"CC",X"F5",X"3A",X"66",X"C5",
		X"CB",X"47",X"20",X"10",X"F1",X"CB",X"EF",X"77",X"1A",X"CB",X"7F",X"28",X"17",X"E6",X"CC",X"CB",
		X"E7",X"12",X"18",X"10",X"F1",X"CB",X"E7",X"77",X"1A",X"CB",X"7F",X"28",X"07",X"E6",X"CC",X"CB",
		X"EF",X"12",X"18",X"00",X"3A",X"66",X"C5",X"CB",X"4F",X"20",X"10",X"7E",X"CB",X"77",X"20",X"03",
		X"CB",X"F7",X"77",X"1A",X"CB",X"77",X"C8",X"CB",X"B7",X"12",X"C9",X"7E",X"CB",X"77",X"28",X"03",
		X"CB",X"B7",X"77",X"1A",X"CB",X"77",X"C0",X"CB",X"F7",X"12",X"C9",X"1A",X"CB",X"5F",X"C2",X"AD",
		X"45",X"CB",X"7F",X"C8",X"E6",X"CC",X"F5",X"3A",X"66",X"C5",X"CB",X"47",X"20",X"06",X"F1",X"CB",
		X"E7",X"12",X"18",X"C0",X"F1",X"CB",X"EF",X"12",X"18",X"BA",X"C3",X"6B",X"45",X"CB",X"57",X"28",
		X"0E",X"CB",X"97",X"77",X"DD",X"36",X"13",X"00",X"DD",X"36",X"12",X"00",X"C3",X"6B",X"45",X"CB",
		X"D7",X"77",X"DD",X"36",X"13",X"00",X"DD",X"36",X"12",X"00",X"C3",X"6B",X"45",X"C9",X"CB",X"57",
		X"28",X"0C",X"CB",X"97",X"12",X"FD",X"36",X"13",X"00",X"FD",X"36",X"12",X"00",X"C9",X"CB",X"D7",
		X"12",X"FD",X"36",X"13",X"00",X"FD",X"36",X"12",X"00",X"C9",X"AF",X"32",X"66",X"C5",X"44",X"4D",
		X"7A",X"90",X"30",X"0C",X"2F",X"3C",X"F5",X"3A",X"66",X"C5",X"CB",X"C7",X"32",X"66",X"C5",X"F1",
		X"FE",X"0F",X"D0",X"7B",X"91",X"30",X"0C",X"2F",X"3C",X"F5",X"3A",X"66",X"C5",X"CB",X"CF",X"32",
		X"66",X"C5",X"F1",X"FE",X"0F",X"C9",X"E5",X"3A",X"66",X"C5",X"21",X"BF",X"46",X"CD",X"A8",X"3D",
		X"E9",X"E1",X"7E",X"A7",X"28",X"3A",X"FE",X"18",X"38",X"2B",X"18",X"34",X"E1",X"7E",X"A7",X"28",
		X"2F",X"FE",X"09",X"30",X"20",X"18",X"29",X"E1",X"7E",X"D6",X"10",X"38",X"18",X"A7",X"28",X"20",
		X"FE",X"09",X"30",X"11",X"18",X"1A",X"E1",X"7E",X"D6",X"08",X"38",X"09",X"A7",X"28",X"11",X"FE",
		X"09",X"30",X"02",X"18",X"0B",X"7E",X"E5",X"21",X"4B",X"4B",X"CD",X"50",X"20",X"7E",X"E1",X"77",
		X"3A",X"66",X"C5",X"21",X"CF",X"46",X"CD",X"A8",X"3D",X"E9",X"1A",X"A7",X"C8",X"FE",X"18",X"38",
		X"21",X"C9",X"1A",X"A7",X"C8",X"FE",X"09",X"30",X"19",X"C9",X"1A",X"D6",X"10",X"38",X"13",X"A7",
		X"C8",X"FE",X"09",X"30",X"0D",X"C9",X"1A",X"D6",X"08",X"38",X"07",X"A7",X"C8",X"FE",X"09",X"30",
		X"01",X"C9",X"1A",X"21",X"4B",X"4B",X"CD",X"50",X"20",X"7E",X"12",X"C9",X"E5",X"3A",X"66",X"C5",
		X"21",X"C7",X"46",X"CD",X"A8",X"3D",X"E9",X"E1",X"7E",X"A7",X"C8",X"FE",X"18",X"38",X"24",X"C9",
		X"E1",X"7E",X"A7",X"C8",X"FE",X"09",X"30",X"1B",X"C9",X"E1",X"7E",X"D6",X"10",X"38",X"14",X"A7",
		X"C8",X"FE",X"09",X"30",X"0E",X"C9",X"E1",X"7E",X"D6",X"08",X"38",X"07",X"A7",X"C8",X"FE",X"09",
		X"30",X"01",X"C9",X"7E",X"E5",X"21",X"4B",X"4B",X"CD",X"50",X"20",X"7E",X"E1",X"77",X"C9",X"01",
		X"46",X"0C",X"46",X"17",X"46",X"26",X"46",X"87",X"46",X"90",X"46",X"99",X"46",X"A6",X"46",X"66",
		X"46",X"5A",X"46",X"52",X"46",X"4A",X"46",X"7C",X"D6",X"18",X"38",X"29",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"FE",X"0D",X"30",X"1D",X"67",X"7D",X"D6",X"18",X"D8",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"6F",X"3E",X"11",X"95",X"D8",X"7D",X"A7",X"28",X"06",X"AF",X"C6",X"0D",X"2D",
		X"20",X"FB",X"84",X"A7",X"C9",X"37",X"C9",X"DD",X"7E",X"03",X"E6",X"07",X"28",X"0B",X"DD",X"7E",
		X"03",X"CB",X"67",X"C2",X"47",X"48",X"C3",X"AE",X"47",X"DD",X"7E",X"03",X"E6",X"1C",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"21",X"43",X"4B",X"CD",X"A8",X"3D",X"E9",X"DD",X"CB",X"11",X"4E",X"20",
		X"2F",X"DD",X"CB",X"11",X"46",X"20",X"3A",X"CD",X"3B",X"49",X"D0",X"DD",X"CB",X"11",X"6E",X"20",
		X"04",X"CD",X"87",X"49",X"D0",X"DD",X"CB",X"11",X"66",X"20",X"04",X"CD",X"1F",X"4A",X"D0",X"DD",
		X"CB",X"11",X"B6",X"DD",X"CB",X"11",X"A6",X"DD",X"CB",X"11",X"AE",X"DD",X"36",X"03",X"10",X"C9",
		X"CD",X"70",X"4A",X"38",X"D2",X"DD",X"CB",X"11",X"6E",X"20",X"CC",X"CD",X"87",X"49",X"38",X"C7",
		X"C9",X"CD",X"A4",X"4A",X"38",X"C1",X"DD",X"CB",X"11",X"66",X"20",X"BB",X"CD",X"1F",X"4A",X"38",
		X"B6",X"C9",X"CD",X"D3",X"49",X"D0",X"DD",X"CB",X"11",X"6E",X"20",X"04",X"CD",X"87",X"49",X"D0",
		X"DD",X"CB",X"11",X"66",X"20",X"04",X"CD",X"1F",X"4A",X"D0",X"CD",X"E0",X"48",X"DD",X"CB",X"11",
		X"AE",X"DD",X"CB",X"11",X"A6",X"DD",X"CB",X"11",X"F6",X"DD",X"36",X"03",X"00",X"C9",X"DD",X"CB",
		X"11",X"76",X"20",X"2C",X"CD",X"D3",X"49",X"D0",X"DD",X"CB",X"11",X"6E",X"20",X"04",X"CD",X"87",
		X"49",X"D0",X"DD",X"CB",X"11",X"66",X"20",X"04",X"CD",X"1F",X"4A",X"D0",X"CD",X"E0",X"48",X"DD",
		X"CB",X"11",X"AE",X"DD",X"CB",X"11",X"A6",X"DD",X"CB",X"11",X"F6",X"DD",X"36",X"03",X"00",X"C9",
		X"DD",X"CB",X"11",X"4E",X"20",X"2F",X"DD",X"CB",X"11",X"46",X"20",X"42",X"CD",X"3B",X"49",X"D0",
		X"DD",X"CB",X"11",X"6E",X"20",X"04",X"CD",X"87",X"49",X"D0",X"DD",X"CB",X"11",X"66",X"20",X"04",
		X"CD",X"1F",X"4A",X"D0",X"DD",X"CB",X"11",X"B6",X"DD",X"CB",X"11",X"A6",X"DD",X"CB",X"11",X"AE",
		X"DD",X"36",X"03",X"10",X"C9",X"DD",X"CB",X"11",X"6E",X"20",X"D1",X"CD",X"87",X"49",X"38",X"CC",
		X"FD",X"7E",X"01",X"DD",X"46",X"13",X"B8",X"C0",X"DD",X"CB",X"11",X"8E",X"18",X"D6",X"DD",X"CB",
		X"11",X"66",X"20",X"B8",X"CD",X"1F",X"4A",X"38",X"B3",X"FD",X"7E",X"01",X"DD",X"46",X"13",X"B8",
		X"C0",X"DD",X"CB",X"11",X"86",X"18",X"BD",X"DD",X"CB",X"11",X"76",X"20",X"2C",X"CD",X"D3",X"49",
		X"D0",X"DD",X"CB",X"11",X"66",X"20",X"04",X"CD",X"1F",X"4A",X"D0",X"DD",X"CB",X"11",X"6E",X"20",
		X"04",X"CD",X"87",X"49",X"D0",X"CD",X"E0",X"48",X"DD",X"CB",X"11",X"AE",X"DD",X"CB",X"11",X"A6",
		X"DD",X"CB",X"11",X"F6",X"DD",X"36",X"03",X"00",X"C9",X"DD",X"CB",X"11",X"4E",X"20",X"2F",X"DD",
		X"CB",X"11",X"46",X"20",X"42",X"CD",X"3B",X"49",X"D0",X"DD",X"CB",X"11",X"66",X"20",X"04",X"CD",
		X"1F",X"4A",X"D0",X"DD",X"CB",X"11",X"6E",X"20",X"04",X"CD",X"87",X"49",X"D0",X"DD",X"CB",X"11",
		X"B6",X"DD",X"CB",X"11",X"A6",X"DD",X"CB",X"11",X"AE",X"DD",X"36",X"03",X"10",X"C9",X"DD",X"CB",
		X"11",X"6E",X"20",X"D1",X"CD",X"87",X"49",X"38",X"CC",X"FD",X"7E",X"01",X"DD",X"46",X"13",X"B8",
		X"C0",X"DD",X"CB",X"13",X"8E",X"18",X"D6",X"DD",X"CB",X"11",X"66",X"20",X"B8",X"CD",X"1F",X"4A",
		X"38",X"B3",X"FD",X"7E",X"01",X"DD",X"46",X"13",X"B8",X"C0",X"DD",X"CB",X"11",X"86",X"18",X"BD",
		X"FD",X"7E",X"00",X"C6",X"08",X"6F",X"26",X"18",X"16",X"18",X"CD",X"D7",X"46",X"4F",X"06",X"0D",
		X"2A",X"88",X"ED",X"79",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"28",X"0B",X"0C",X"F5",X"3E",X"10",
		X"82",X"57",X"F1",X"10",X"EB",X"18",X"2B",X"FD",X"6E",X"00",X"FD",X"7E",X"01",X"C6",X"10",X"67",
		X"CD",X"D7",X"46",X"47",X"79",X"D6",X"0D",X"B8",X"38",X"0C",X"DD",X"CB",X"11",X"CE",X"DD",X"CB",
		X"11",X"86",X"DD",X"72",X"13",X"C9",X"DD",X"CB",X"11",X"C6",X"DD",X"CB",X"11",X"8E",X"DD",X"72",
		X"13",X"C9",X"3E",X"FC",X"DD",X"A6",X"11",X"DD",X"77",X"11",X"C9",X"FD",X"7E",X"00",X"D6",X"08",
		X"6F",X"FD",X"7E",X"01",X"C6",X"0F",X"67",X"CD",X"D7",X"46",X"DA",X"D2",X"4A",X"2A",X"88",X"ED",
		X"CD",X"50",X"20",X"7E",X"E6",X"03",X"C2",X"D2",X"4A",X"FD",X"7E",X"00",X"D6",X"08",X"6F",X"FD",
		X"7E",X"01",X"D6",X"0F",X"C6",X"10",X"67",X"CD",X"D7",X"46",X"DA",X"D2",X"4A",X"2A",X"88",X"ED",
		X"CD",X"50",X"20",X"7E",X"E6",X"03",X"C2",X"D2",X"4A",X"DD",X"36",X"03",X"00",X"DD",X"CB",X"11",
		X"AE",X"DD",X"CB",X"11",X"A6",X"A7",X"C9",X"FD",X"7E",X"00",X"C6",X"07",X"6F",X"FD",X"7E",X"01",
		X"3D",X"FE",X"D7",X"D2",X"CD",X"49",X"C6",X"10",X"67",X"CD",X"D7",X"46",X"DA",X"CD",X"49",X"2A",
		X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"C2",X"CD",X"49",X"FD",X"7E",X"00",X"D6",X"07",
		X"6F",X"FD",X"7E",X"01",X"3D",X"C6",X"10",X"67",X"CD",X"D7",X"46",X"2A",X"88",X"ED",X"CD",X"50",
		X"20",X"7E",X"E6",X"03",X"C2",X"CD",X"49",X"DD",X"36",X"03",X"08",X"A7",X"C9",X"DD",X"CB",X"11",
		X"EE",X"37",X"C9",X"FD",X"7E",X"00",X"C6",X"08",X"6F",X"FD",X"7E",X"01",X"C6",X"0F",X"67",X"CD",
		X"D7",X"46",X"DA",X"D2",X"4A",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"C2",X"D2",
		X"4A",X"FD",X"7E",X"00",X"C6",X"08",X"6F",X"FD",X"7E",X"01",X"D6",X"0F",X"C6",X"10",X"67",X"CD",
		X"D7",X"46",X"DA",X"D2",X"4A",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"C2",X"D2",
		X"4A",X"DD",X"36",X"03",X"10",X"DD",X"CB",X"11",X"AE",X"DD",X"CB",X"11",X"A6",X"A7",X"C9",X"FD",
		X"7E",X"00",X"C6",X"07",X"6F",X"FD",X"7E",X"01",X"D6",X"0F",X"FE",X"09",X"DA",X"6A",X"4A",X"C6",
		X"10",X"67",X"CD",X"D7",X"46",X"DA",X"6A",X"4A",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",
		X"03",X"C2",X"6A",X"4A",X"FD",X"7E",X"00",X"D6",X"07",X"6F",X"FD",X"7E",X"01",X"D6",X"0F",X"C6",
		X"10",X"67",X"CD",X"D7",X"46",X"DA",X"6A",X"4A",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",
		X"03",X"C2",X"6A",X"4A",X"DD",X"36",X"03",X"18",X"A7",X"C9",X"DD",X"CB",X"11",X"E6",X"37",X"C9",
		X"FD",X"7E",X"01",X"C6",X"10",X"67",X"FD",X"6E",X"00",X"CD",X"D7",X"46",X"38",X"54",X"2A",X"88",
		X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"20",X"49",X"FD",X"7E",X"01",X"C6",X"10",X"67",X"FD",
		X"6E",X"04",X"CD",X"D7",X"46",X"38",X"3B",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",
		X"20",X"30",X"A7",X"C9",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"CD",X"D7",X"46",X"38",X"23",X"2A",
		X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"20",X"18",X"FD",X"66",X"01",X"FD",X"6E",X"04",
		X"CD",X"D7",X"46",X"38",X"0D",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"20",X"02",
		X"A7",X"C9",X"37",X"C9",X"DD",X"CB",X"11",X"76",X"20",X"F8",X"FD",X"7E",X"00",X"FE",X"70",X"38",
		X"F1",X"C6",X"08",X"6F",X"26",X"18",X"CD",X"D7",X"46",X"38",X"1C",X"0E",X"00",X"06",X"0D",X"2A",
		X"88",X"ED",X"F5",X"CD",X"50",X"20",X"7E",X"E6",X"03",X"28",X"06",X"0C",X"3E",X"01",X"B9",X"28",
		X"08",X"F1",X"3C",X"10",X"EA",X"A7",X"C9",X"A7",X"C9",X"F1",X"37",X"C9",X"FD",X"7E",X"01",X"FE",
		X"D9",X"38",X"18",X"DD",X"7E",X"03",X"DD",X"36",X"12",X"00",X"DD",X"36",X"13",X"00",X"DD",X"CB",
		X"11",X"D6",X"FD",X"36",X"01",X"D8",X"FD",X"36",X"05",X"D8",X"C9",X"FE",X"17",X"D0",X"DD",X"36",
		X"12",X"00",X"DD",X"36",X"13",X"00",X"DD",X"CB",X"11",X"96",X"FD",X"36",X"01",X"18",X"FD",X"36",
		X"05",X"18",X"C9",X"2B",X"47",X"AE",X"47",X"82",X"47",X"47",X"48",X"10",X"11",X"12",X"13",X"14",
		X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",X"1D",X"1E",X"1F",X"00",X"01",X"02",X"03",X"04",
		X"05",X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"E8",X"42",X"3B",X"44",X"E6",
		X"44",X"89",X"C4",X"91",X"C4",X"99",X"C4",X"03",X"0D",X"04",X"0D",X"05",X"0D",X"08",X"0D",X"08",
		X"0D",X"08",X"0D",X"FF",X"FF",X"07",X"12",X"00",X"00",X"07",X"12",X"01",X"00",X"07",X"12",X"02",
		X"00",X"07",X"12",X"03",X"00",X"07",X"12",X"04",X"00",X"07",X"12",X"05",X"00",X"07",X"12",X"06",
		X"00",X"07",X"12",X"07",X"00",X"FF",X"FF",X"0A",X"11",X"00",X"00",X"0A",X"11",X"01",X"00",X"0A",
		X"11",X"02",X"00",X"0A",X"11",X"03",X"00",X"0A",X"11",X"04",X"00",X"0A",X"11",X"05",X"00",X"0A",
		X"11",X"06",X"00",X"0A",X"11",X"07",X"00",X"0A",X"11",X"08",X"00",X"0A",X"11",X"09",X"00",X"0A",
		X"11",X"0A",X"00",X"0A",X"11",X"05",X"00",X"FF",X"FF",X"05",X"0D",X"00",X"00",X"05",X"0D",X"01",
		X"00",X"05",X"0D",X"02",X"00",X"05",X"0D",X"03",X"00",X"05",X"0D",X"04",X"00",X"05",X"0D",X"05",
		X"00",X"05",X"0D",X"06",X"00",X"05",X"0D",X"07",X"00",X"05",X"0E",X"00",X"00",X"05",X"0E",X"01",
		X"00",X"05",X"0E",X"02",X"00",X"05",X"0E",X"03",X"00",X"05",X"0E",X"04",X"00",X"05",X"0E",X"05",
		X"00",X"05",X"0E",X"06",X"00",X"05",X"0E",X"07",X"00",X"05",X"0F",X"00",X"00",X"05",X"0F",X"01",
		X"00",X"05",X"0F",X"02",X"00",X"05",X"0F",X"03",X"00",X"05",X"0F",X"04",X"00",X"05",X"0F",X"05",
		X"00",X"05",X"0F",X"06",X"00",X"05",X"0F",X"07",X"00",X"FF",X"FF",X"0A",X"10",X"00",X"00",X"0A",
		X"10",X"01",X"00",X"0A",X"10",X"02",X"00",X"0A",X"10",X"03",X"00",X"0A",X"10",X"04",X"00",X"0A",
		X"10",X"05",X"00",X"0A",X"10",X"00",X"00",X"0A",X"10",X"01",X"00",X"0A",X"10",X"02",X"00",X"0A",
		X"10",X"03",X"00",X"0A",X"10",X"04",X"00",X"0A",X"10",X"05",X"00",X"05",X"10",X"06",X"00",X"05",
		X"10",X"07",X"00",X"05",X"10",X"08",X"00",X"0A",X"10",X"09",X"00",X"05",X"10",X"08",X"00",X"05",
		X"10",X"07",X"00",X"05",X"10",X"06",X"00",X"0A",X"10",X"05",X"00",X"FF",X"FF",X"05",X"13",X"00",
		X"00",X"05",X"13",X"01",X"00",X"05",X"13",X"02",X"00",X"05",X"13",X"03",X"00",X"05",X"13",X"00",
		X"00",X"05",X"13",X"04",X"00",X"05",X"13",X"05",X"00",X"FF",X"FF",X"04",X"09",X"2C",X"00",X"04",
		X"09",X"30",X"00",X"04",X"09",X"34",X"00",X"04",X"09",X"38",X"00",X"04",X"09",X"3C",X"00",X"FF",
		X"FF",X"04",X"09",X"3C",X"00",X"04",X"09",X"38",X"00",X"04",X"09",X"34",X"00",X"04",X"09",X"30",
		X"00",X"04",X"09",X"2C",X"00",X"04",X"09",X"06",X"00",X"FF",X"FF",X"15",X"30",X"16",X"10",X"17",
		X"20",X"18",X"38",X"19",X"08",X"1B",X"08",X"1C",X"08",X"1E",X"08",X"1F",X"08",X"00",X"08",X"04",
		X"08",X"06",X"08",X"07",X"08",X"08",X"2D",X"09",X"08",X"0A",X"08",X"0B",X"08",X"0C",X"08",X"0D",
		X"28",X"0E",X"08",X"0F",X"08",X"10",X"08",X"12",X"04",X"14",X"04",X"FF",X"FF",X"0B",X"30",X"0A",
		X"10",X"09",X"20",X"08",X"38",X"07",X"08",X"05",X"08",X"04",X"08",X"02",X"08",X"01",X"08",X"00",
		X"08",X"1C",X"08",X"1A",X"08",X"19",X"08",X"18",X"2D",X"17",X"08",X"16",X"08",X"15",X"08",X"14",
		X"08",X"13",X"28",X"12",X"08",X"11",X"08",X"10",X"08",X"0E",X"04",X"0C",X"04",X"FF",X"FF",X"18",
		X"08",X"17",X"10",X"15",X"0A",X"14",X"0B",X"13",X"0C",X"12",X"0D",X"11",X"1D",X"08",X"08",X"09",
		X"10",X"0B",X"0A",X"0C",X"0B",X"0D",X"0C",X"0E",X"0D",X"0F",X"1D",X"0E",X"28",X"0D",X"26",X"0A",
		X"15",X"09",X"18",X"08",X"1F",X"04",X"1A",X"01",X"0E",X"1C",X"0E",X"19",X"10",X"17",X"1A",X"16",
		X"28",X"14",X"13",X"12",X"15",X"10",X"0E",X"0D",X"1C",X"FF",X"FF",X"12",X"28",X"13",X"26",X"16",
		X"15",X"17",X"18",X"18",X"1F",X"1C",X"1A",X"1F",X"0E",X"04",X"0E",X"07",X"10",X"09",X"1A",X"0A",
		X"28",X"0C",X"13",X"0E",X"15",X"10",X"0E",X"13",X"1C",X"FF",X"FF",X"0A",X"11",X"0E",X"34",X"0B",
		X"11",X"08",X"11",X"05",X"11",X"02",X"34",X"06",X"11",X"FF",X"FF",X"16",X"11",X"12",X"34",X"15",
		X"11",X"18",X"11",X"1B",X"11",X"1E",X"34",X"1A",X"11",X"FF",X"FF",X"0F",X"24",X"0D",X"39",X"0A",
		X"1C",X"09",X"24",X"08",X"30",X"06",X"24",X"04",X"1C",X"01",X"10",X"1D",X"13",X"1A",X"18",X"19",
		X"26",X"18",X"21",X"16",X"28",X"15",X"26",X"13",X"15",X"11",X"26",X"FF",X"FF",X"11",X"24",X"13",
		X"39",X"16",X"1C",X"17",X"24",X"18",X"30",X"1A",X"24",X"1C",X"1C",X"1F",X"10",X"03",X"13",X"06",
		X"18",X"07",X"26",X"08",X"21",X"0A",X"28",X"0B",X"26",X"0D",X"15",X"0F",X"26",X"FF",X"FF",X"73",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"01",
		X"FF",X"09",X"09",X"09",X"0A",X"09",X"09",X"09",X"FF",X"01",X"09",X"09",X"01",X"1D",X"FF",X"09",
		X"0A",X"0A",X"0A",X"09",X"FF",X"0D",X"01",X"09",X"09",X"01",X"1D",X"1D",X"FF",X"09",X"0A",X"09",
		X"FF",X"0D",X"0D",X"01",X"09",X"09",X"01",X"1D",X"1D",X"1D",X"FF",X"02",X"FF",X"0D",X"0D",X"0D",
		X"01",X"09",X"09",X"01",X"1D",X"1D",X"1D",X"1D",X"01",X"0D",X"0D",X"0D",X"0D",X"01",X"09",X"09",
		X"01",X"1E",X"1D",X"1D",X"1D",X"01",X"0D",X"0D",X"0D",X"0E",X"01",X"09",X"09",X"01",X"1E",X"1D",
		X"1D",X"1D",X"01",X"0D",X"0D",X"0D",X"0E",X"01",X"09",X"09",X"03",X"1E",X"1D",X"1D",X"1D",X"02",
		X"0D",X"0D",X"0D",X"0E",X"03",X"09",X"0A",X"0A",X"03",X"1E",X"1D",X"1D",X"02",X"0D",X"0D",X"0E",
		X"03",X"0A",X"0A",X"09",X"09",X"09",X"03",X"1D",X"1D",X"02",X"0D",X"0D",X"03",X"09",X"09",X"09",
		X"09",X"09",X"09",X"09",X"03",X"1D",X"02",X"0D",X"03",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"09",X"09",X"03",X"02",X"03",X"09",X"09",X"09",X"09",X"09",X"E7",X"AF",X"32",X"69",X"C5",X"21",
		X"00",X"00",X"01",X"00",X"10",X"3A",X"69",X"C5",X"86",X"32",X"69",X"C5",X"23",X"0B",X"78",X"B1",
		X"20",X"F3",X"3A",X"69",X"C5",X"21",X"D3",X"14",X"BE",X"28",X"26",X"32",X"84",X"ED",X"2F",X"32",
		X"80",X"ED",X"28",X"1D",X"3E",X"E9",X"ED",X"47",X"E7",X"3E",X"EA",X"ED",X"47",X"E7",X"3E",X"EB",
		X"ED",X"47",X"E7",X"3E",X"EC",X"ED",X"47",X"E7",X"3E",X"ED",X"ED",X"47",X"E7",X"3E",X"EE",X"ED",
		X"47",X"E7",X"21",X"6E",X"C5",X"11",X"6F",X"C5",X"01",X"E9",X"00",X"36",X"00",X"ED",X"B0",X"E7",
		X"DD",X"21",X"6A",X"C5",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"03",X"00",X"CD",X"D0",X"4F",X"AF",X"06",X"7B",X"F5",X"4F",X"21",X"6E",X"C5",X"CD",
		X"50",X"20",X"7E",X"A7",X"C4",X"88",X"4F",X"F1",X"3C",X"10",X"EF",X"F5",X"E7",X"F1",X"06",X"6F",
		X"F5",X"4F",X"21",X"6E",X"C5",X"CD",X"50",X"20",X"7E",X"A7",X"C4",X"88",X"4F",X"F1",X"3C",X"10",
		X"EF",X"F5",X"3E",X"03",X"DF",X"F1",X"18",X"CF",X"E5",X"F5",X"2A",X"88",X"ED",X"79",X"CD",X"50",
		X"20",X"7E",X"A7",X"20",X"05",X"F1",X"E1",X"36",X"00",X"C9",X"F1",X"FE",X"05",X"28",X"12",X"79",
		X"C5",X"CD",X"CA",X"5A",X"C1",X"23",X"34",X"34",X"CD",X"03",X"21",X"23",X"34",X"34",X"E1",X"34",
		X"C9",X"21",X"F0",X"0A",X"CD",X"D1",X"20",X"3E",X"10",X"85",X"F5",X"79",X"C5",X"CD",X"CA",X"5A",
		X"C1",X"23",X"F1",X"F5",X"77",X"CD",X"03",X"21",X"23",X"F1",X"3C",X"77",X"E1",X"36",X"00",X"C9",
		X"E7",X"DD",X"34",X"00",X"DD",X"7E",X"00",X"FE",X"03",X"20",X"F5",X"AF",X"DD",X"77",X"00",X"DD",
		X"77",X"03",X"06",X"E9",X"DD",X"7E",X"03",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"7E",X"E6",X"03",
		X"FE",X"03",X"20",X"39",X"DD",X"7E",X"02",X"FE",X"05",X"28",X"13",X"DD",X"7E",X"03",X"C5",X"CD",
		X"CA",X"5A",X"C1",X"23",X"34",X"34",X"CD",X"03",X"21",X"23",X"34",X"34",X"18",X"1F",X"21",X"F0",
		X"0A",X"CD",X"D1",X"20",X"3E",X"10",X"85",X"F5",X"DD",X"7E",X"03",X"C5",X"CD",X"CA",X"5A",X"C1",
		X"23",X"F1",X"F5",X"77",X"CD",X"03",X"21",X"23",X"F1",X"3C",X"77",X"18",X"00",X"DD",X"34",X"03",
		X"10",X"B2",X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"06",X"C2",X"D0",X"4F",X"DD",X"36",X"02",
		X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"00",X"00",X"FF",X"00",X"00",X"02",X"02",X"00",X"00",X"02",X"02",X"00",
		X"00",X"06",X"06",X"00",X"06",X"06",X"00",X"00",X"02",X"02",X"00",X"00",X"06",X"06",X"00",X"00",
		X"FF",X"00",X"00",X"06",X"06",X"00",X"00",X"06",X"06",X"00",X"00",X"1E",X"1E",X"00",X"1E",X"1E",
		X"00",X"00",X"06",X"06",X"00",X"00",X"1E",X"1E",X"00",X"00",X"FF",X"00",X"00",X"1E",X"1E",X"00",
		X"00",X"1E",X"1E",X"00",X"00",X"0E",X"0E",X"00",X"0E",X"0E",X"00",X"00",X"1E",X"1E",X"00",X"00",
		X"0E",X"0E",X"00",X"00",X"FF",X"00",X"00",X"0E",X"0E",X"00",X"00",X"0E",X"0E",X"00",X"00",X"12",
		X"12",X"00",X"12",X"12",X"00",X"00",X"0E",X"0E",X"00",X"00",X"12",X"12",X"00",X"00",X"FF",X"00",
		X"00",X"12",X"12",X"00",X"00",X"12",X"12",X"00",X"00",X"16",X"16",X"00",X"16",X"16",X"00",X"00",
		X"12",X"12",X"00",X"00",X"16",X"16",X"00",X"00",X"00",X"00",X"00",X"16",X"16",X"00",X"00",X"16",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"16",X"CD",X"40",X"51",X"3A",
		X"58",X"C6",X"CB",X"7F",X"C2",X"29",X"53",X"47",X"3A",X"59",X"C6",X"B8",X"C2",X"7F",X"52",X"C9",
		X"3A",X"59",X"C6",X"FE",X"01",X"C0",X"21",X"65",X"C6",X"FD",X"21",X"B9",X"C4",X"CD",X"5B",X"51",
		X"21",X"67",X"C6",X"FD",X"21",X"85",X"C4",X"CD",X"5B",X"51",X"C9",X"CB",X"76",X"C2",X"5D",X"52",
		X"CB",X"7E",X"20",X"62",X"3A",X"65",X"C4",X"FE",X"01",X"C0",X"3A",X"6F",X"ED",X"CB",X"4F",X"28",
		X"1A",X"3A",X"FF",X"BF",X"FE",X"76",X"20",X"13",X"3A",X"C1",X"C4",X"CB",X"7F",X"28",X"0C",X"3A",
		X"C0",X"C4",X"CB",X"57",X"C0",X"CB",X"D7",X"CB",X"87",X"18",X"10",X"3A",X"66",X"EF",X"A7",X"20",
		X"06",X"3A",X"C0",X"C4",X"CB",X"47",X"C0",X"CB",X"C7",X"CB",X"97",X"32",X"C0",X"C4",X"CB",X"FE",
		X"23",X"36",X"E8",X"3A",X"3A",X"C4",X"D6",X"08",X"FD",X"77",X"01",X"FD",X"36",X"00",X"E3",X"21",
		X"B0",X"1B",X"CD",X"BA",X"20",X"3E",X"C8",X"23",X"23",X"B4",X"FD",X"77",X"02",X"FD",X"75",X"03",
		X"3E",X"06",X"CD",X"AE",X"67",X"C9",X"FD",X"35",X"00",X"FD",X"35",X"00",X"FD",X"35",X"00",X"FD",
		X"35",X"00",X"FD",X"35",X"00",X"FD",X"7E",X"00",X"FE",X"18",X"30",X"06",X"CB",X"F6",X"23",X"36",
		X"00",X"C9",X"11",X"FE",X"C4",X"CD",X"2E",X"52",X"11",X"01",X"C5",X"CD",X"2E",X"52",X"11",X"04",
		X"C5",X"CD",X"2E",X"52",X"E5",X"AF",X"32",X"69",X"C6",X"FD",X"66",X"01",X"FD",X"6E",X"00",X"CD",
		X"D7",X"46",X"CD",X"54",X"58",X"38",X"05",X"3E",X"FF",X"32",X"69",X"C6",X"FD",X"7E",X"01",X"FD",
		X"6E",X"00",X"C6",X"0C",X"67",X"CD",X"D7",X"46",X"CD",X"54",X"58",X"38",X"05",X"3E",X"FF",X"32",
		X"69",X"C6",X"E1",X"3A",X"69",X"C6",X"A7",X"C8",X"CB",X"F6",X"23",X"36",X"00",X"C9",X"1A",X"CB",
		X"47",X"C8",X"13",X"1A",X"D6",X"06",X"FD",X"BE",X"01",X"D0",X"C6",X"18",X"FD",X"BE",X"01",X"D8",
		X"13",X"1A",X"D6",X"03",X"FD",X"BE",X"00",X"D0",X"C6",X"10",X"FD",X"BE",X"00",X"D8",X"1B",X"1B",
		X"1A",X"CB",X"E7",X"CB",X"EF",X"12",X"CB",X"F6",X"23",X"36",X"00",X"2B",X"C9",X"23",X"34",X"7E",
		X"FE",X"01",X"20",X"04",X"FD",X"35",X"03",X"C9",X"FE",X"06",X"20",X"04",X"FD",X"35",X"03",X"C9",
		X"FE",X"0B",X"C0",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"2B",X"36",X"00",X"C9",X"3A",
		X"59",X"C6",X"FE",X"01",X"28",X"12",X"FE",X"02",X"28",X"0E",X"21",X"85",X"C4",X"22",X"5D",X"C6",
		X"21",X"A1",X"C4",X"22",X"5B",X"C6",X"18",X"0C",X"21",X"A9",X"C4",X"22",X"5D",X"C6",X"21",X"AD",
		X"C4",X"22",X"5B",X"C6",X"21",X"19",X"53",X"3A",X"58",X"C6",X"CB",X"FF",X"32",X"58",X"C6",X"3D",
		X"CB",X"27",X"CD",X"56",X"20",X"7B",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"32",X"60",X"C6",X"21",
		X"00",X"18",X"CD",X"BA",X"20",X"7A",X"CD",X"50",X"20",X"E5",X"3A",X"5A",X"C6",X"CD",X"CA",X"5A",
		X"C1",X"CB",X"22",X"CB",X"22",X"CB",X"22",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"3E",
		X"18",X"82",X"57",X"3E",X"18",X"83",X"5F",X"2A",X"5B",X"C6",X"72",X"23",X"73",X"23",X"3A",X"60",
		X"C6",X"B0",X"77",X"23",X"71",X"E5",X"21",X"63",X"C6",X"23",X"77",X"2B",X"71",X"E1",X"14",X"14",
		X"1C",X"1C",X"2A",X"5D",X"C6",X"72",X"23",X"73",X"23",X"3E",X"40",X"B0",X"77",X"23",X"71",X"3E",
		X"0A",X"32",X"61",X"C6",X"AF",X"32",X"62",X"C6",X"C9",X"13",X"10",X"13",X"18",X"14",X"08",X"14",
		X"00",X"15",X"28",X"15",X"20",X"0C",X"30",X"00",X"00",X"3A",X"61",X"C6",X"3D",X"32",X"61",X"C6",
		X"20",X"30",X"3A",X"62",X"C6",X"3C",X"32",X"62",X"C6",X"06",X"07",X"FE",X"05",X"20",X"02",X"06",
		X"0F",X"F5",X"78",X"32",X"61",X"C6",X"F1",X"FE",X"08",X"20",X"04",X"AF",X"32",X"62",X"C6",X"2A",
		X"5B",X"C6",X"23",X"23",X"EB",X"2A",X"63",X"C6",X"3A",X"62",X"C6",X"CD",X"50",X"20",X"EB",X"72",
		X"23",X"73",X"2A",X"5D",X"C6",X"34",X"2A",X"5B",X"C6",X"34",X"7E",X"FE",X"F8",X"D2",X"EB",X"53",
		X"7E",X"FE",X"E2",X"D8",X"FE",X"EC",X"D0",X"23",X"3A",X"3A",X"C4",X"C6",X"04",X"96",X"D8",X"3A",
		X"3B",X"C4",X"D6",X"04",X"96",X"D0",X"AF",X"32",X"48",X"C4",X"2A",X"5D",X"C6",X"CD",X"6B",X"54",
		X"2A",X"5B",X"C6",X"CD",X"6B",X"54",X"3A",X"59",X"C6",X"FE",X"01",X"20",X"2B",X"CD",X"E4",X"53",
		X"FD",X"21",X"B9",X"C4",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"00",
		X"FD",X"36",X"03",X"00",X"FD",X"21",X"85",X"C4",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"00",
		X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"3A",X"58",X"C6",X"CB",X"BF",X"32",X"58",X"C6",
		X"32",X"59",X"C6",X"3D",X"CB",X"27",X"21",X"74",X"54",X"CD",X"56",X"20",X"EB",X"11",X"00",X"01",
		X"CD",X"23",X"27",X"E9",X"21",X"65",X"C6",X"CD",X"6B",X"54",X"C9",X"AF",X"2A",X"5D",X"C6",X"CD",
		X"6B",X"54",X"2A",X"5B",X"C6",X"CD",X"6B",X"54",X"3A",X"59",X"C6",X"32",X"58",X"C6",X"C9",X"CD",
		X"E4",X"53",X"3E",X"00",X"32",X"69",X"C4",X"3E",X"01",X"32",X"63",X"C4",X"C9",X"3E",X"00",X"32",
		X"69",X"C4",X"3E",X"02",X"32",X"63",X"C4",X"C9",X"3E",X"00",X"32",X"69",X"C4",X"3E",X"03",X"32",
		X"63",X"C4",X"C9",X"3E",X"00",X"32",X"69",X"C4",X"32",X"63",X"C4",X"3A",X"62",X"C4",X"D6",X"02",
		X"D8",X"C8",X"32",X"62",X"C4",X"C9",X"3E",X"00",X"32",X"63",X"C4",X"3E",X"00",X"32",X"69",X"C4",
		X"3E",X"01",X"32",X"CE",X"C4",X"C9",X"3E",X"00",X"32",X"63",X"C4",X"3E",X"02",X"32",X"69",X"C4",
		X"C9",X"3E",X"10",X"CD",X"AE",X"67",X"3A",X"71",X"ED",X"3C",X"32",X"71",X"ED",X"CD",X"70",X"22",
		X"3E",X"00",X"32",X"63",X"C4",X"3E",X"00",X"32",X"69",X"C4",X"C9",X"AF",X"77",X"23",X"77",X"23",
		X"77",X"23",X"77",X"C9",X"FF",X"53",X"0D",X"54",X"18",X"54",X"23",X"54",X"36",X"54",X"46",X"54",
		X"51",X"54",X"AF",X"32",X"58",X"C6",X"32",X"59",X"C6",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"15",
		X"16",X"03",X"0E",X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"15",X"15",X"16",X"01",X"01",X"01",
		X"0D",X"0D",X"0E",X"00",X"00",X"00",X"00",X"15",X"16",X"01",X"01",X"02",X"01",X"01",X"0E",X"0D",
		X"00",X"00",X"00",X"15",X"16",X"15",X"01",X"01",X"01",X"01",X"02",X"0D",X"0D",X"0D",X"00",X"00",
		X"16",X"15",X"15",X"01",X"01",X"01",X"02",X"01",X"0D",X"0D",X"0D",X"00",X"00",X"15",X"15",X"15",
		X"01",X"01",X"02",X"01",X"01",X"0D",X"0D",X"0E",X"00",X"00",X"03",X"00",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"FE",X"FF",X"20",X"05",X"3E",X"01",X"32",X"73",X"C6",X"CB",X"27",
		X"CB",X"27",X"21",X"29",X"56",X"CD",X"50",X"20",X"5E",X"16",X"00",X"23",X"E5",X"21",X"30",X"0C",
		X"CD",X"D1",X"20",X"19",X"EB",X"E1",X"46",X"48",X"23",X"7E",X"32",X"71",X"C6",X"32",X"6B",X"C6",
		X"21",X"C6",X"E0",X"D5",X"CD",X"F6",X"55",X"D5",X"11",X"40",X"00",X"19",X"D1",X"3E",X"04",X"CD",
		X"4A",X"20",X"10",X"F0",X"41",X"E5",X"11",X"C6",X"E7",X"ED",X"52",X"E1",X"D1",X"38",X"E4",X"21",
		X"06",X"E7",X"06",X"1D",X"7E",X"E6",X"07",X"77",X"3A",X"6B",X"C6",X"D6",X"B8",X"B6",X"77",X"23",
		X"23",X"10",X"F1",X"3A",X"73",X"C6",X"A7",X"20",X"15",X"FD",X"21",X"83",X"ED",X"FD",X"36",X"00",
		X"00",X"06",X"EA",X"AF",X"F5",X"C5",X"CD",X"39",X"56",X"C1",X"F1",X"3C",X"10",X"F6",X"AF",X"32",
		X"71",X"C6",X"32",X"73",X"C6",X"C9",X"E5",X"D5",X"C5",X"06",X"1D",X"7B",X"C6",X"04",X"F5",X"3A",
		X"71",X"C6",X"D6",X"B8",X"30",X"02",X"C6",X"B8",X"B2",X"77",X"F1",X"23",X"73",X"23",X"1C",X"05",
		X"F5",X"3A",X"71",X"C6",X"B2",X"77",X"F1",X"23",X"73",X"23",X"1C",X"BB",X"20",X"05",X"F5",X"D6",
		X"04",X"5F",X"F1",X"10",X"EB",X"C1",X"D1",X"E1",X"C9",X"00",X"03",X"E0",X"00",X"0C",X"04",X"E8",
		X"00",X"1C",X"04",X"E8",X"00",X"2C",X"04",X"F0",X"00",X"F5",X"ED",X"5B",X"88",X"ED",X"CD",X"4A",
		X"20",X"1A",X"A7",X"28",X"65",X"FE",X"FF",X"28",X"03",X"FD",X"34",X"00",X"E6",X"03",X"28",X"5A",
		X"FE",X"03",X"20",X"0D",X"1A",X"11",X"BC",X"56",X"FE",X"FF",X"20",X"10",X"11",X"BE",X"56",X"18",
		X"0B",X"1A",X"CB",X"3F",X"E6",X"0E",X"11",X"AC",X"56",X"CD",X"4A",X"20",X"21",X"F0",X"0A",X"CD",
		X"D1",X"20",X"1A",X"85",X"6F",X"30",X"01",X"24",X"13",X"1A",X"B4",X"67",X"EB",X"F1",X"F5",X"D5",
		X"CD",X"CA",X"5A",X"D1",X"72",X"23",X"73",X"13",X"CD",X"03",X"21",X"72",X"23",X"73",X"23",X"7E",
		X"E6",X"07",X"57",X"3A",X"6B",X"C6",X"D6",X"B8",X"82",X"77",X"23",X"CD",X"03",X"21",X"7E",X"E6",
		X"07",X"57",X"3A",X"6B",X"C6",X"D6",X"B8",X"82",X"77",X"23",X"F1",X"C9",X"00",X"C0",X"02",X"C0",
		X"04",X"C0",X"06",X"C0",X"08",X"C0",X"0A",X"C0",X"0C",X"C8",X"0E",X"C8",X"10",X"C8",X"10",X"D8",
		X"1E",X"00",X"CD",X"DB",X"56",X"CD",X"00",X"57",X"7B",X"FE",X"03",X"CA",X"95",X"57",X"CB",X"43",
		X"C2",X"65",X"57",X"CB",X"4B",X"C2",X"3B",X"57",X"C3",X"3F",X"58",X"DD",X"7E",X"07",X"6F",X"E6",
		X"F8",X"4F",X"DD",X"7E",X"09",X"E6",X"F8",X"B9",X"28",X"12",X"CB",X"C3",X"DD",X"CB",X"00",X"46",
		X"28",X"06",X"79",X"C6",X"08",X"6F",X"18",X"04",X"79",X"D6",X"03",X"6F",X"DD",X"75",X"09",X"C9",
		X"DD",X"7E",X"08",X"67",X"E6",X"F8",X"28",X"2F",X"FE",X"F8",X"28",X"2B",X"47",X"DD",X"7E",X"0A",
		X"E6",X"F8",X"B8",X"28",X"22",X"E6",X"18",X"C5",X"F5",X"78",X"E6",X"18",X"47",X"F1",X"A8",X"C1",
		X"FE",X"18",X"28",X"13",X"60",X"CB",X"CB",X"DD",X"CB",X"00",X"4E",X"28",X"06",X"78",X"C6",X"08",
		X"67",X"18",X"04",X"78",X"D6",X"02",X"67",X"DD",X"74",X"0A",X"C9",X"D9",X"DD",X"6E",X"07",X"DD",
		X"66",X"08",X"CD",X"D7",X"46",X"CD",X"54",X"58",X"D9",X"DA",X"3F",X"58",X"FD",X"7E",X"00",X"DD",
		X"77",X"09",X"DD",X"7E",X"0A",X"FD",X"77",X"01",X"DD",X"7E",X"03",X"2F",X"3C",X"E6",X"1F",X"DD",
		X"77",X"03",X"C3",X"3A",X"58",X"D9",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"CD",X"D7",X"46",X"CD",
		X"54",X"58",X"D9",X"DA",X"3F",X"58",X"DD",X"7E",X"09",X"FD",X"77",X"00",X"FD",X"7E",X"01",X"DD",
		X"77",X"0A",X"DD",X"7E",X"03",X"F5",X"2F",X"3C",X"E6",X"0F",X"5F",X"F1",X"E6",X"10",X"B3",X"DD",
		X"77",X"03",X"C3",X"3A",X"58",X"D9",X"DD",X"6E",X"07",X"DD",X"66",X"08",X"CD",X"D7",X"46",X"D9",
		X"DA",X"3F",X"58",X"57",X"DD",X"7E",X"03",X"CB",X"3F",X"CB",X"3F",X"E6",X"06",X"21",X"4C",X"58",
		X"CD",X"50",X"20",X"1E",X"00",X"7E",X"82",X"FE",X"EA",X"3F",X"F5",X"38",X"0D",X"ED",X"4B",X"88",
		X"ED",X"CD",X"44",X"20",X"0A",X"A7",X"28",X"02",X"CB",X"CB",X"23",X"7E",X"82",X"FE",X"EA",X"3F",
		X"F5",X"38",X"0D",X"ED",X"4B",X"88",X"ED",X"CD",X"44",X"20",X"0A",X"A7",X"28",X"02",X"CB",X"C3",
		X"7B",X"A7",X"28",X"2E",X"FE",X"03",X"20",X"0C",X"D9",X"F1",X"CD",X"54",X"58",X"F1",X"CD",X"54",
		X"58",X"D9",X"18",X"2A",X"CB",X"43",X"28",X"0D",X"F1",X"D9",X"C1",X"CD",X"54",X"58",X"D9",X"DA",
		X"3F",X"58",X"C3",X"76",X"57",X"F1",X"F1",X"D9",X"CD",X"54",X"58",X"D9",X"DA",X"3F",X"58",X"C3",
		X"4C",X"57",X"F1",X"F1",X"7A",X"D9",X"A7",X"CD",X"54",X"58",X"D9",X"DA",X"3F",X"58",X"DD",X"7E",
		X"03",X"2F",X"E6",X"10",X"5F",X"DD",X"7E",X"03",X"E6",X"0F",X"B3",X"DD",X"77",X"03",X"DD",X"7E",
		X"09",X"FD",X"77",X"00",X"DD",X"7E",X"0A",X"FD",X"77",X"01",X"DD",X"CB",X"06",X"BE",X"C9",X"DD",
		X"7E",X"07",X"DD",X"77",X"09",X"DD",X"7E",X"08",X"DD",X"77",X"0A",X"C9",X"0D",X"FF",X"F3",X"FF",
		X"F3",X"01",X"0D",X"01",X"D8",X"DD",X"E5",X"F5",X"3A",X"C4",X"C4",X"32",X"74",X"C6",X"AF",X"32",
		X"C4",X"C4",X"21",X"0B",X"D0",X"23",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",
		X"7E",X"CD",X"50",X"20",X"3E",X"48",X"86",X"E1",X"CB",X"76",X"28",X"FC",X"32",X"18",X"D0",X"CB",
		X"76",X"28",X"FC",X"F1",X"F5",X"32",X"18",X"D0",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"D5",
		X"3A",X"6A",X"C6",X"5F",X"3A",X"6C",X"C6",X"57",X"CD",X"23",X"27",X"2A",X"71",X"C4",X"7E",X"6F",
		X"E5",X"3A",X"0C",X"D0",X"CB",X"7F",X"20",X"F9",X"3A",X"33",X"C4",X"5F",X"3A",X"34",X"C4",X"57",
		X"CD",X"23",X"27",X"2A",X"71",X"C4",X"7E",X"E1",X"67",X"D1",X"3A",X"74",X"C6",X"32",X"C4",X"C4",
		X"7E",X"A7",X"CA",X"E4",X"59",X"FE",X"FF",X"20",X"17",X"F1",X"F5",X"21",X"6E",X"C5",X"CD",X"50",
		X"20",X"7E",X"A7",X"C2",X"D8",X"59",X"36",X"01",X"3E",X"16",X"CD",X"AE",X"67",X"C3",X"D8",X"59",
		X"FE",X"E2",X"20",X"08",X"3E",X"01",X"32",X"CE",X"C4",X"C3",X"94",X"59",X"7E",X"E6",X"03",X"FE",
		X"03",X"20",X"23",X"5F",X"F1",X"F5",X"E5",X"21",X"6E",X"C5",X"CD",X"50",X"20",X"7E",X"A7",X"20",
		X"02",X"36",X"01",X"E1",X"7E",X"E6",X"FC",X"D6",X"04",X"DA",X"94",X"59",X"B3",X"77",X"3E",X"16",
		X"CD",X"AE",X"67",X"C3",X"D8",X"59",X"CB",X"4F",X"28",X"7A",X"3A",X"69",X"C4",X"FE",X"02",X"28",
		X"73",X"3A",X"58",X"C6",X"CB",X"7F",X"20",X"6C",X"E5",X"3A",X"6F",X"ED",X"21",X"D9",X"C4",X"CB",
		X"4F",X"28",X"03",X"21",X"DD",X"C4",X"3A",X"58",X"C6",X"47",X"3A",X"66",X"EF",X"A7",X"ED",X"5F",
		X"20",X"01",X"7E",X"E1",X"E6",X"07",X"28",X"4C",X"B8",X"20",X"02",X"3E",X"06",X"FE",X"05",X"28",
		X"04",X"FE",X"07",X"20",X"37",X"E5",X"3A",X"6F",X"ED",X"21",X"D9",X"C4",X"CB",X"4F",X"28",X"03",
		X"21",X"DD",X"C4",X"7E",X"E1",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E6",X"07",X"28",
		X"23",X"B8",X"20",X"04",X"3E",X"06",X"18",X"14",X"FE",X"07",X"20",X"10",X"3A",X"74",X"C4",X"FE",
		X"07",X"20",X"04",X"3E",X"02",X"18",X"05",X"3E",X"07",X"32",X"74",X"C4",X"32",X"58",X"C6",X"F1",
		X"32",X"5A",X"C6",X"F5",X"3E",X"04",X"CD",X"AE",X"67",X"7E",X"CD",X"3B",X"5A",X"AF",X"32",X"72",
		X"C6",X"77",X"F1",X"F5",X"CD",X"CA",X"5A",X"7B",X"A7",X"3E",X"01",X"20",X"03",X"32",X"72",X"C6",
		X"F1",X"F5",X"CD",X"EE",X"5A",X"E5",X"CD",X"40",X"5B",X"E1",X"DD",X"21",X"6D",X"C6",X"CD",X"E9",
		X"59",X"CD",X"03",X"21",X"CD",X"E9",X"59",X"23",X"CD",X"2C",X"5A",X"CD",X"03",X"21",X"CD",X"2C",
		X"5A",X"3A",X"83",X"ED",X"3D",X"32",X"83",X"ED",X"F1",X"DD",X"E1",X"3A",X"63",X"EF",X"3C",X"32",
		X"63",X"EF",X"A7",X"C9",X"F1",X"DD",X"E1",X"37",X"C9",X"CD",X"B7",X"5A",X"38",X"47",X"3A",X"72",
		X"C6",X"A7",X"20",X"04",X"CB",X"41",X"28",X"1D",X"EB",X"21",X"30",X"0C",X"CD",X"D1",X"20",X"DD",
		X"7E",X"00",X"CD",X"50",X"20",X"EB",X"3A",X"6B",X"C6",X"D6",X"B8",X"B2",X"77",X"23",X"73",X"AF",
		X"32",X"72",X"C6",X"18",X"21",X"EB",X"21",X"30",X"0C",X"CD",X"D1",X"20",X"DD",X"7E",X"00",X"CD",
		X"50",X"20",X"EB",X"3A",X"6B",X"C6",X"B2",X"77",X"23",X"73",X"18",X"0A",X"CD",X"B7",X"5A",X"38",
		X"04",X"CB",X"41",X"28",X"E0",X"23",X"DD",X"23",X"CB",X"39",X"C9",X"D9",X"F5",X"E6",X"03",X"FE",
		X"03",X"20",X"0D",X"F1",X"3A",X"72",X"ED",X"87",X"21",X"73",X"5A",X"CD",X"50",X"20",X"18",X"0B",
		X"F1",X"CB",X"3F",X"E6",X"0E",X"21",X"63",X"5A",X"CD",X"50",X"20",X"5E",X"23",X"56",X"CD",X"23",
		X"27",X"D9",X"C9",X"05",X"00",X"06",X"00",X"07",X"00",X"08",X"00",X"09",X"00",X"10",X"00",X"11",
		X"00",X"12",X"00",X"05",X"00",X"10",X"00",X"15",X"00",X"20",X"00",X"25",X"00",X"30",X"00",X"35",
		X"00",X"40",X"00",X"45",X"00",X"50",X"00",X"55",X"00",X"60",X"00",X"65",X"00",X"70",X"00",X"75",
		X"00",X"80",X"00",X"85",X"00",X"90",X"00",X"95",X"00",X"00",X"01",X"05",X"01",X"10",X"01",X"15",
		X"01",X"20",X"01",X"25",X"01",X"30",X"01",X"35",X"01",X"40",X"01",X"45",X"01",X"50",X"01",X"55",
		X"01",X"60",X"01",X"75",X"01",X"80",X"01",X"D5",X"EB",X"A7",X"21",X"40",X"E7",X"ED",X"52",X"38",
		X"06",X"21",X"C6",X"E0",X"ED",X"52",X"3F",X"EB",X"D1",X"C9",X"F5",X"C5",X"4F",X"01",X"FF",X"00",
		X"0C",X"D6",X"0D",X"30",X"FB",X"C6",X"0D",X"5F",X"51",X"CB",X"3F",X"CB",X"18",X"CB",X"21",X"69",
		X"48",X"47",X"7D",X"21",X"06",X"E7",X"CD",X"50",X"20",X"ED",X"42",X"C1",X"F1",X"C9",X"D5",X"01",
		X"00",X"04",X"ED",X"5B",X"88",X"ED",X"D6",X"0E",X"F5",X"CD",X"4A",X"20",X"F1",X"F5",X"CD",X"39",
		X"5B",X"CB",X"39",X"13",X"F1",X"F5",X"CD",X"39",X"5B",X"F1",X"CB",X"39",X"06",X"1B",X"80",X"FE",
		X"EA",X"30",X"03",X"3F",X"18",X"01",X"37",X"ED",X"5B",X"88",X"ED",X"F5",X"CD",X"4A",X"20",X"F1",
		X"F5",X"CD",X"39",X"5B",X"CB",X"39",X"13",X"F1",X"CD",X"39",X"5B",X"D1",X"7B",X"A7",X"20",X"02",
		X"CB",X"81",X"FE",X"0C",X"20",X"02",X"CB",X"99",X"C9",X"D8",X"1A",X"A7",X"C8",X"CB",X"D9",X"C9",
		X"C5",X"3A",X"72",X"ED",X"E6",X"03",X"01",X"04",X"04",X"20",X"03",X"01",X"03",X"04",X"CD",X"9C",
		X"5B",X"E5",X"28",X"04",X"0E",X"10",X"18",X"02",X"0E",X"0C",X"DD",X"21",X"6D",X"C6",X"CD",X"7D",
		X"5B",X"DD",X"23",X"DD",X"23",X"7B",X"E6",X"03",X"FE",X"03",X"7B",X"20",X"02",X"D6",X"04",X"D6",
		X"03",X"CB",X"7F",X"28",X"01",X"81",X"5F",X"CD",X"7D",X"5B",X"E1",X"C1",X"C9",X"D5",X"7B",X"D6",
		X"04",X"30",X"01",X"81",X"57",X"21",X"BB",X"5B",X"3A",X"72",X"ED",X"E6",X"03",X"CD",X"50",X"20",
		X"7E",X"83",X"DD",X"77",X"00",X"7E",X"82",X"DD",X"77",X"01",X"D1",X"C9",X"F5",X"7A",X"CD",X"B6",
		X"5B",X"57",X"3E",X"0C",X"93",X"CB",X"27",X"3C",X"41",X"CD",X"B6",X"5B",X"CB",X"27",X"CB",X"27",
		X"82",X"5F",X"16",X"00",X"F1",X"C9",X"90",X"30",X"FD",X"80",X"C9",X"00",X"0C",X"1C",X"2C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"FF",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"FF",X"00",X"05",
		X"05",X"00",X"FF",X"FF",X"1D",X"1D",X"1D",X"1D",X"1D",X"FF",X"FF",X"00",X"05",X"06",X"00",X"FF",
		X"00",X"FF",X"1D",X"1D",X"1D",X"FF",X"00",X"FF",X"00",X"06",X"06",X"00",X"FF",X"00",X"19",X"FF",
		X"1E",X"FF",X"09",X"00",X"FF",X"00",X"06",X"06",X"00",X"FF",X"00",X"1A",X"00",X"03",X"00",X"0A",
		X"00",X"FF",X"00",X"06",X"06",X"00",X"FF",X"00",X"1A",X"00",X"0E",X"00",X"0A",X"00",X"FF",X"00",
		X"06",X"06",X"00",X"FF",X"00",X"1A",X"00",X"0D",X"00",X"0A",X"00",X"FF",X"00",X"06",X"06",X"00",
		X"FF",X"00",X"1A",X"00",X"0E",X"00",X"0A",X"00",X"FF",X"00",X"06",X"06",X"00",X"FF",X"00",X"1A",
		X"00",X"0D",X"00",X"0A",X"00",X"FF",X"00",X"06",X"05",X"FF",X"FF",X"FF",X"19",X"00",X"0E",X"00",
		X"09",X"FF",X"FF",X"FF",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"46",X"52",X"49",X"2C",X"20",X"20",
		X"36",X"20",X"4A",X"55",X"4E",X"20",X"31",X"39",X"38",X"36",X"2C",X"20",X"31",X"35",X"3A",X"34",
		X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"0E",X"11",X"16",X"19",X"FF",X"19",X"16",X"11",X"0E",X"00",X"00",X"00",
		X"00",X"0E",X"11",X"16",X"19",X"FF",X"19",X"16",X"11",X"0E",X"00",X"00",X"00",X"00",X"0E",X"11",
		X"16",X"19",X"FF",X"19",X"16",X"11",X"0E",X"00",X"00",X"00",X"00",X"0E",X"11",X"16",X"19",X"1E",
		X"19",X"16",X"11",X"0E",X"00",X"00",X"00",X"00",X"0E",X"11",X"16",X"19",X"FF",X"19",X"16",X"11",
		X"0E",X"00",X"00",X"00",X"00",X"0E",X"11",X"16",X"19",X"FF",X"19",X"16",X"11",X"0E",X"00",X"00",
		X"00",X"00",X"0E",X"11",X"16",X"19",X"FF",X"19",X"16",X"11",X"0E",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"FF",X"06",X"FF",X"0A",X"FF",X"0E",X"FF",X"12",X"FF",X"16",X"FF",X"FF",X"1A",X"FF",X"03",
		X"FF",X"03",X"FF",X"03",X"FF",X"03",X"FF",X"1E",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"FF",X"00",X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1A",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"1A",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"1A",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"1A",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"1A",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"D0",X"11",X"94",X"E8",X"DD",X"21",X"80",X"E8",X"CD",
		X"14",X"5F",X"11",X"9F",X"E8",X"CD",X"3A",X"5F",X"DD",X"CB",X"00",X"4E",X"28",X"07",X"3E",X"01",
		X"32",X"94",X"E9",X"18",X"23",X"3A",X"94",X"E9",X"A7",X"28",X"0D",X"97",X"32",X"94",X"E9",X"3D",
		X"32",X"11",X"E9",X"3E",X"03",X"32",X"12",X"E9",X"11",X"14",X"E9",X"DD",X"21",X"00",X"E9",X"CD",
		X"14",X"5F",X"11",X"1F",X"E9",X"CD",X"3A",X"5F",X"DD",X"21",X"80",X"E8",X"21",X"80",X"E8",X"22",
		X"92",X"E9",X"CB",X"46",X"C4",X"67",X"5F",X"DD",X"CB",X"00",X"4E",X"28",X"09",X"DD",X"35",X"13",
		X"CC",X"3A",X"60",X"CD",X"7B",X"62",X"DD",X"21",X"00",X"E9",X"21",X"00",X"E9",X"22",X"92",X"E9",
		X"CB",X"46",X"C4",X"67",X"5F",X"DD",X"CB",X"00",X"4E",X"C8",X"DD",X"35",X"13",X"CC",X"3A",X"60",
		X"CD",X"7B",X"62",X"C9",X"DD",X"4E",X"11",X"97",X"DD",X"77",X"11",X"47",X"CD",X"4F",X"5F",X"CD",
		X"4F",X"5F",X"CD",X"4F",X"5F",X"79",X"A7",X"C8",X"18",X"02",X"04",X"13",X"1F",X"30",X"FB",X"4F",
		X"70",X"1A",X"23",X"77",X"2B",X"79",X"A7",X"20",X"F1",X"C9",X"DD",X"4E",X"12",X"DD",X"36",X"12",
		X"00",X"06",X"0B",X"CD",X"4F",X"5F",X"CB",X"39",X"D0",X"70",X"1A",X"23",X"77",X"2B",X"C9",X"CB",
		X"39",X"30",X"0F",X"70",X"1A",X"23",X"77",X"2B",X"04",X"13",X"70",X"1A",X"23",X"77",X"2B",X"04",
		X"13",X"C9",X"04",X"04",X"13",X"13",X"C9",X"36",X"02",X"23",X"5E",X"23",X"56",X"1A",X"23",X"23",
		X"77",X"13",X"1A",X"E6",X"0F",X"20",X"02",X"3E",X"10",X"23",X"23",X"77",X"13",X"1A",X"23",X"77",
		X"13",X"1A",X"23",X"77",X"13",X"DD",X"73",X"0D",X"DD",X"72",X"0E",X"CD",X"95",X"5F",X"2A",X"92",
		X"E9",X"CD",X"AC",X"5F",X"C9",X"1A",X"E6",X"F0",X"DD",X"77",X"05",X"1A",X"E6",X"0F",X"DD",X"77",
		X"0A",X"13",X"1A",X"DD",X"77",X"0B",X"13",X"1A",X"DD",X"77",X"0C",X"C9",X"11",X"10",X"00",X"19",
		X"97",X"77",X"23",X"36",X"FF",X"23",X"36",X"03",X"23",X"36",X"01",X"23",X"06",X"0E",X"77",X"23",
		X"10",X"FC",X"3E",X"3F",X"F6",X"00",X"DD",X"77",X"1B",X"11",X"0B",X"00",X"06",X"07",X"97",X"77",
		X"19",X"10",X"FC",X"C9",X"DD",X"7E",X"0A",X"A7",X"28",X"06",X"3D",X"28",X"18",X"DD",X"77",X"0A",
		X"DD",X"5E",X"0D",X"DD",X"56",X"0E",X"13",X"1A",X"DD",X"77",X"0B",X"13",X"1A",X"DD",X"77",X"0C",
		X"DD",X"36",X"13",X"01",X"C9",X"DD",X"35",X"07",X"28",X"17",X"DD",X"5E",X"0D",X"DD",X"56",X"0E",
		X"13",X"13",X"13",X"DD",X"73",X"0D",X"DD",X"72",X"0E",X"CD",X"95",X"5F",X"DD",X"36",X"13",X"01",
		X"C9",X"DD",X"35",X"06",X"20",X"09",X"CB",X"8E",X"CD",X"AC",X"5F",X"CD",X"9F",X"66",X"C9",X"DD",
		X"5E",X"01",X"DD",X"56",X"02",X"13",X"13",X"1A",X"DD",X"77",X"07",X"13",X"13",X"DD",X"73",X"0D",
		X"DD",X"72",X"0E",X"CD",X"95",X"5F",X"CD",X"AC",X"5F",X"C9",X"DD",X"4E",X"0B",X"DD",X"46",X"0C",
		X"0A",X"FE",X"F0",X"20",X"02",X"03",X"0A",X"A7",X"20",X"04",X"CD",X"D4",X"5F",X"C9",X"DD",X"77",
		X"13",X"CD",X"5B",X"60",X"DD",X"71",X"0B",X"DD",X"70",X"0C",X"C9",X"03",X"0A",X"E6",X"C0",X"C8",
		X"0A",X"E6",X"F0",X"D6",X"40",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"10",X"61",X"19",X"5E",
		X"23",X"56",X"EB",X"0A",X"E6",X"0F",X"E9",X"DD",X"77",X"15",X"03",X"0A",X"DD",X"77",X"14",X"11",
		X"01",X"00",X"C3",X"FF",X"60",X"DD",X"77",X"17",X"03",X"0A",X"DD",X"77",X"16",X"11",X"02",X"00",
		X"18",X"6D",X"DD",X"77",X"19",X"03",X"0A",X"DD",X"77",X"18",X"11",X"04",X"00",X"18",X"60",X"07",
		X"07",X"07",X"07",X"DD",X"77",X"1F",X"03",X"0A",X"DD",X"77",X"20",X"11",X"00",X"03",X"18",X"4F",
		X"DD",X"77",X"1C",X"11",X"20",X"00",X"7B",X"2F",X"DD",X"A6",X"10",X"DD",X"77",X"10",X"18",X"3F",
		X"DD",X"77",X"1D",X"11",X"40",X"00",X"7B",X"2F",X"DD",X"A6",X"10",X"DD",X"77",X"10",X"18",X"2F",
		X"DD",X"77",X"1E",X"11",X"80",X"00",X"7B",X"2F",X"DD",X"A6",X"10",X"DD",X"77",X"10",X"18",X"1F",
		X"11",X"00",X"00",X"18",X"1A",X"11",X"00",X"00",X"18",X"15",X"11",X"00",X"00",X"18",X"10",X"11",
		X"00",X"00",X"18",X"0B",X"CD",X"28",X"61",X"7A",X"B3",X"CA",X"5B",X"60",X"CB",X"7A",X"C0",X"DD",
		X"7E",X"11",X"B3",X"DD",X"77",X"11",X"DD",X"7E",X"12",X"B2",X"DD",X"77",X"12",X"C3",X"5B",X"60",
		X"77",X"60",X"85",X"60",X"92",X"60",X"9F",X"60",X"B0",X"60",X"C0",X"60",X"D0",X"60",X"E0",X"60",
		X"E5",X"60",X"EA",X"60",X"EF",X"60",X"F4",X"60",X"87",X"87",X"5F",X"16",X"00",X"21",X"DD",X"61",
		X"19",X"5E",X"23",X"56",X"D5",X"23",X"5E",X"23",X"56",X"03",X"0A",X"C9",X"0B",X"C9",X"E6",X"1F",
		X"DD",X"77",X"1A",X"C9",X"21",X"2F",X"6A",X"CD",X"2D",X"62",X"FD",X"CB",X"00",X"CE",X"11",X"00",
		X"00",X"C9",X"E6",X"07",X"F6",X"08",X"DD",X"77",X"21",X"0A",X"07",X"38",X"0F",X"07",X"38",X"06",
		X"DD",X"36",X"0F",X"00",X"18",X"13",X"DD",X"36",X"0F",X"01",X"18",X"0D",X"07",X"38",X"06",X"DD",
		X"36",X"0F",X"02",X"18",X"04",X"DD",X"36",X"0F",X"04",X"E6",X"E0",X"DD",X"77",X"10",X"07",X"30",
		X"0A",X"DD",X"36",X"1E",X"10",X"DD",X"36",X"64",X"00",X"CB",X"FB",X"07",X"30",X"0A",X"DD",X"36",
		X"1D",X"10",X"DD",X"36",X"59",X"00",X"CB",X"F3",X"07",X"30",X"0A",X"DD",X"36",X"1C",X"10",X"DD",
		X"36",X"4E",X"00",X"CB",X"EB",X"C9",X"21",X"47",X"6A",X"CD",X"2D",X"62",X"11",X"00",X"00",X"C9",
		X"E6",X"3F",X"F6",X"00",X"DD",X"77",X"1B",X"C9",X"21",X"2F",X"6A",X"CD",X"2D",X"62",X"11",X"00",
		X"00",X"C9",X"E6",X"F0",X"20",X"14",X"0A",X"E6",X"0F",X"5F",X"16",X"00",X"21",X"1D",X"62",X"19",
		X"7E",X"A7",X"28",X"06",X"2A",X"92",X"E9",X"5F",X"19",X"72",X"5A",X"C9",X"C9",X"3C",X"61",X"00",
		X"80",X"3E",X"61",X"08",X"00",X"44",X"61",X"43",X"00",X"52",X"61",X"00",X"02",X"A6",X"61",X"22",
		X"00",X"A6",X"61",X"2D",X"00",X"A6",X"61",X"38",X"00",X"B0",X"61",X"10",X"00",X"B8",X"61",X"4E",
		X"00",X"B8",X"61",X"59",X"00",X"B8",X"61",X"64",X"00",X"DC",X"61",X"00",X"00",X"DC",X"61",X"00",
		X"00",X"DC",X"61",X"00",X"00",X"DC",X"61",X"00",X"00",X"C2",X"61",X"00",X"00",X"00",X"00",X"43",
		X"00",X"22",X"2D",X"38",X"00",X"4E",X"59",X"64",X"00",X"00",X"00",X"00",X"00",X"FD",X"2A",X"92",
		X"E9",X"FD",X"19",X"16",X"C1",X"CB",X"7F",X"28",X"02",X"CB",X"EA",X"FD",X"72",X"00",X"E6",X"7F",
		X"FD",X"77",X"09",X"5F",X"03",X"0A",X"FD",X"77",X"01",X"FD",X"77",X"0A",X"CB",X"6A",X"28",X"01",
		X"97",X"FD",X"77",X"02",X"E5",X"16",X"00",X"62",X"6B",X"29",X"29",X"19",X"D1",X"19",X"7E",X"FD",
		X"77",X"03",X"23",X"7E",X"FD",X"77",X"07",X"23",X"7E",X"FD",X"77",X"08",X"23",X"5E",X"FD",X"73",
		X"04",X"23",X"56",X"FD",X"72",X"05",X"FD",X"36",X"06",X"00",X"C9",X"DD",X"7E",X"0F",X"DD",X"A6",
		X"11",X"28",X"04",X"DD",X"CB",X"12",X"CE",X"FD",X"2A",X"92",X"E9",X"11",X"22",X"00",X"FD",X"19",
		X"11",X"14",X"01",X"CD",X"E5",X"62",X"11",X"0B",X"00",X"FD",X"19",X"11",X"16",X"02",X"CD",X"E5",
		X"62",X"11",X"0B",X"00",X"FD",X"19",X"11",X"18",X"04",X"CD",X"E5",X"62",X"11",X"0B",X"00",X"FD",
		X"19",X"11",X"08",X"00",X"21",X"1A",X"00",X"CD",X"C1",X"63",X"11",X"0B",X"00",X"FD",X"19",X"11",
		X"20",X"00",X"21",X"1C",X"00",X"CD",X"C1",X"63",X"11",X"0B",X"00",X"FD",X"19",X"11",X"40",X"00",
		X"21",X"1D",X"00",X"CD",X"C1",X"63",X"11",X"0B",X"00",X"FD",X"19",X"11",X"80",X"00",X"21",X"1E",
		X"00",X"CD",X"C1",X"63",X"C9",X"D5",X"FD",X"E5",X"E1",X"CB",X"46",X"CB",X"86",X"C2",X"BF",X"63",
		X"DD",X"7E",X"11",X"A2",X"28",X"23",X"CB",X"76",X"CA",X"BF",X"63",X"FD",X"5E",X"09",X"FD",X"7E",
		X"0A",X"FD",X"77",X"01",X"CB",X"6E",X"28",X"01",X"97",X"FD",X"77",X"02",X"21",X"47",X"6A",X"CD",
		X"54",X"62",X"FD",X"CB",X"00",X"FE",X"C3",X"BF",X"63",X"CB",X"7E",X"CA",X"BF",X"63",X"CB",X"6E",
		X"28",X"14",X"FD",X"7E",X"0A",X"A7",X"28",X"0A",X"23",X"7E",X"23",X"86",X"77",X"38",X"0D",X"C3",
		X"BF",X"63",X"23",X"23",X"18",X"06",X"23",X"23",X"35",X"C2",X"BF",X"63",X"23",X"23",X"5E",X"23",
		X"56",X"23",X"7E",X"34",X"26",X"00",X"6F",X"19",X"4E",X"23",X"7E",X"A7",X"20",X"40",X"FD",X"7E",
		X"07",X"A7",X"28",X"32",X"FD",X"35",X"07",X"20",X"2D",X"FD",X"5E",X"08",X"CB",X"7B",X"20",X"20",
		X"FD",X"7E",X"0A",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"6E",X"28",X"01",X"97",X"FD",X"77",X"02",
		X"21",X"47",X"6A",X"CD",X"54",X"62",X"FD",X"36",X"06",X"01",X"EB",X"4E",X"23",X"7E",X"18",X"0E",
		X"FD",X"CB",X"00",X"BE",X"18",X"39",X"FD",X"36",X"06",X"01",X"EB",X"4E",X"23",X"7E",X"06",X"00",
		X"91",X"4F",X"F2",X"96",X"63",X"05",X"2A",X"92",X"E9",X"D1",X"7A",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"09",X"EB",X"72",X"2B",X"73",X"DD",X"B6",X"11",X"DD",X"77",X"11",X"FD",X"7E",X"03",
		X"FD",X"86",X"01",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"6E",X"C0",X"FD",X"77",X"02",X"C9",X"D1",
		X"C9",X"D5",X"E5",X"FD",X"E5",X"E1",X"CB",X"46",X"28",X"0E",X"CB",X"86",X"DD",X"7E",X"10",X"A3",
		X"CA",X"C6",X"64",X"36",X"00",X"C3",X"C6",X"64",X"DD",X"7E",X"11",X"A3",X"20",X"06",X"DD",X"7E",
		X"12",X"A2",X"28",X"27",X"CB",X"76",X"CA",X"C6",X"64",X"FD",X"5E",X"09",X"FD",X"7E",X"0A",X"FD",
		X"77",X"01",X"CB",X"6E",X"28",X"01",X"97",X"FD",X"77",X"02",X"21",X"2F",X"6A",X"CD",X"54",X"62",
		X"FD",X"CB",X"00",X"FE",X"FD",X"CB",X"00",X"9E",X"C3",X"C6",X"64",X"CB",X"7E",X"CA",X"C6",X"64",
		X"CB",X"6E",X"28",X"14",X"FD",X"7E",X"0A",X"A7",X"28",X"0A",X"23",X"7E",X"23",X"86",X"77",X"38",
		X"0D",X"C3",X"C6",X"64",X"23",X"23",X"18",X"06",X"23",X"23",X"35",X"C2",X"C6",X"64",X"23",X"23",
		X"5E",X"23",X"56",X"23",X"6E",X"26",X"00",X"19",X"CD",X"C9",X"64",X"30",X"44",X"FD",X"7E",X"07",
		X"A7",X"28",X"32",X"FD",X"35",X"07",X"20",X"2D",X"FD",X"5E",X"08",X"CB",X"7B",X"20",X"20",X"FD",
		X"7E",X"0A",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"6E",X"28",X"01",X"97",X"FD",X"77",X"02",X"21",
		X"2F",X"6A",X"CD",X"54",X"62",X"FD",X"CB",X"00",X"9E",X"EB",X"CD",X"C9",X"64",X"18",X"12",X"FD",
		X"CB",X"00",X"BE",X"18",X"51",X"FD",X"36",X"06",X"00",X"FD",X"CB",X"00",X"9E",X"EB",X"CD",X"C9",
		X"64",X"90",X"47",X"2A",X"92",X"E9",X"D1",X"19",X"7E",X"80",X"F2",X"90",X"64",X"97",X"18",X"14",
		X"FE",X"10",X"38",X"10",X"FD",X"CB",X"00",X"4E",X"28",X"08",X"FE",X"20",X"38",X"06",X"3E",X"1F",
		X"18",X"02",X"3E",X"0F",X"77",X"D1",X"DD",X"7E",X"11",X"B3",X"DD",X"77",X"11",X"DD",X"7E",X"12",
		X"B2",X"DD",X"77",X"12",X"FD",X"7E",X"03",X"FD",X"86",X"01",X"FD",X"77",X"01",X"FD",X"CB",X"00",
		X"6E",X"C0",X"FD",X"77",X"02",X"C9",X"E1",X"D1",X"C9",X"7E",X"FD",X"CB",X"00",X"5E",X"20",X"11",
		X"FD",X"CB",X"00",X"DE",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"47",X"7E",X"E6",X"0F",X"28",X"16",
		X"C9",X"FD",X"CB",X"00",X"9E",X"E6",X"0F",X"47",X"FD",X"34",X"06",X"23",X"7E",X"E6",X"F0",X"28",
		X"05",X"0F",X"0F",X"0F",X"0F",X"C9",X"37",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",
		X"FF",X"00",X"12",X"12",X"12",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"0E",
		X"0E",X"0E",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"16",X"16",X"16",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"02",X"02",X"02",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",
		X"00",X"FF",X"0A",X"0A",X"0A",X"0A",X"0A",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"8B",X"3A",X"80",X"E9",X"47",X"3A",X"81",X"E9",X"B8",X"C8",X"3C",X"E6",X"0F",X"32",
		X"81",X"E9",X"4F",X"06",X"00",X"21",X"82",X"E9",X"09",X"7E",X"FE",X"E0",X"30",X"07",X"FE",X"1E",
		X"D0",X"CD",X"0C",X"66",X"C9",X"FE",X"F0",X"D0",X"CD",X"8C",X"66",X"C9",X"6F",X"26",X"00",X"29",
		X"11",X"23",X"69",X"19",X"4E",X"23",X"46",X"57",X"0A",X"A7",X"C8",X"FE",X"08",X"38",X"04",X"CD",
		X"38",X"66",X"C9",X"5F",X"60",X"69",X"23",X"4E",X"23",X"46",X"0A",X"CB",X"7F",X"28",X"05",X"E5",
		X"CD",X"38",X"66",X"E1",X"1D",X"20",X"EF",X"C9",X"6F",X"3A",X"95",X"E9",X"A7",X"C0",X"7D",X"D5",
		X"E6",X"FE",X"FE",X"84",X"11",X"80",X"E8",X"28",X"22",X"FE",X"86",X"11",X"00",X"E9",X"28",X"1B",
		X"FE",X"F0",X"20",X"36",X"03",X"0A",X"FE",X"84",X"DD",X"21",X"80",X"E8",X"28",X"08",X"FE",X"86",
		X"DD",X"21",X"00",X"E9",X"20",X"24",X"CD",X"5B",X"60",X"18",X"1F",X"1A",X"CB",X"4F",X"28",X"0F",
		X"21",X"05",X"00",X"19",X"6E",X"03",X"0A",X"0B",X"E6",X"F0",X"67",X"7D",X"BC",X"38",X"0B",X"EB",
		X"36",X"01",X"23",X"71",X"23",X"70",X"23",X"D1",X"72",X"C9",X"D1",X"C9",X"FE",X"EE",X"D8",X"FE",
		X"EE",X"20",X"06",X"3E",X"FF",X"32",X"95",X"E9",X"C9",X"3E",X"00",X"32",X"95",X"E9",X"C9",X"DD",
		X"7E",X"08",X"CD",X"AE",X"67",X"38",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"1D",X"1D",X"1D",
		X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"11",X"FF",X"00",X"FF",X"12",X"11",X"12",X"FF",X"00",X"FF",X"12",X"11",
		X"11",X"11",X"FF",X"00",X"FF",X"12",X"12",X"12",X"FF",X"00",X"FF",X"12",X"11",X"11",X"11",X"FF",
		X"00",X"FF",X"12",X"12",X"12",X"FF",X"00",X"FF",X"12",X"11",X"11",X"11",X"FF",X"00",X"FF",X"12",
		X"11",X"12",X"FF",X"00",X"FF",X"12",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CD",X"95",X"5E",X"CD",X"E3",X"65",X"C9",X"C5",X"E5",X"47",X"18",X"09",X"78",X"CD",
		X"2D",X"E0",X"0E",X"20",X"CD",X"0C",X"E0",X"78",X"CD",X"AE",X"67",X"E1",X"C1",X"C9",X"FE",X"F0",
		X"30",X"27",X"E5",X"C5",X"47",X"3A",X"81",X"E9",X"4F",X"3A",X"80",X"E9",X"3C",X"E6",X"0F",X"B9",
		X"20",X"01",X"0C",X"6F",X"26",X"00",X"32",X"80",X"E9",X"79",X"E6",X"0F",X"32",X"81",X"E9",X"78",
		X"01",X"82",X"E9",X"09",X"77",X"A7",X"C1",X"E1",X"C9",X"37",X"C9",X"21",X"00",X"20",X"01",X"00",
		X"10",X"AF",X"32",X"95",X"E9",X"3A",X"95",X"E9",X"86",X"32",X"95",X"E9",X"23",X"0B",X"78",X"B1",
		X"20",X"F3",X"3A",X"95",X"E9",X"21",X"46",X"35",X"BE",X"28",X"1C",X"AF",X"32",X"95",X"E9",X"3A",
		X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"21",X"98",X"7E",X"CD",X"50",X"20",X"3E",X"33",X"86",X"32",
		X"18",X"D0",X"3E",X"EF",X"ED",X"47",X"C9",X"3E",X"FF",X"32",X"95",X"E9",X"3E",X"FF",X"32",X"91",
		X"E8",X"3E",X"03",X"32",X"92",X"E8",X"3E",X"3F",X"F6",X"00",X"32",X"9B",X"E8",X"32",X"1B",X"E9",
		X"3E",X"01",X"32",X"93",X"E8",X"32",X"13",X"E9",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",
		X"00",X"03",X"03",X"03",X"00",X"00",X"03",X"0E",X"03",X"00",X"03",X"0E",X"03",X"00",X"03",X"0E",
		X"03",X"00",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"00",
		X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"00",X"03",X"12",X"03",X"00",X"03",X"12",X"03",
		X"00",X"03",X"12",X"03",X"00",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"03",X"03",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"00",X"00",X"03",X"16",X"03",X"00",
		X"03",X"16",X"03",X"00",X"03",X"16",X"03",X"00",X"00",X"03",X"03",X"03",X"00",X"03",X"03",X"03",
		X"00",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"5F",X"69",X"64",X"69",X"6B",X"69",X"72",X"69",X"87",X"69",X"8E",X"69",X"95",
		X"69",X"9C",X"69",X"AA",X"69",X"B1",X"69",X"BF",X"69",X"C6",X"69",X"D4",X"69",X"DB",X"69",X"E2",
		X"69",X"E9",X"69",X"F0",X"69",X"F7",X"69",X"FE",X"69",X"05",X"6A",X"1A",X"6A",X"21",X"6A",X"A3",
		X"69",X"28",X"6A",X"79",X"69",X"80",X"69",X"B8",X"69",X"0C",X"6A",X"13",X"6A",X"CD",X"69",X"02",
		X"64",X"69",X"6B",X"69",X"84",X"01",X"01",X"FF",X"01",X"B1",X"6A",X"86",X"01",X"01",X"FF",X"01",
		X"B1",X"6A",X"84",X"81",X"01",X"FF",X"81",X"B8",X"6A",X"84",X"71",X"01",X"FF",X"71",X"1A",X"6C",
		X"84",X"81",X"01",X"FF",X"81",X"38",X"6C",X"84",X"81",X"01",X"FF",X"81",X"C5",X"6A",X"84",X"31",
		X"01",X"FF",X"31",X"D2",X"6A",X"84",X"71",X"01",X"FF",X"71",X"21",X"6B",X"84",X"91",X"01",X"FF",
		X"91",X"DB",X"6B",X"84",X"81",X"01",X"FF",X"81",X"A4",X"6B",X"84",X"61",X"01",X"FF",X"61",X"D2",
		X"6A",X"84",X"61",X"01",X"FF",X"61",X"0A",X"6C",X"84",X"51",X"01",X"FF",X"51",X"F2",X"6A",X"86",
		X"81",X"01",X"FF",X"81",X"8B",X"6C",X"84",X"01",X"01",X"1D",X"01",X"B1",X"6A",X"86",X"81",X"01",
		X"FF",X"81",X"79",X"6D",X"84",X"21",X"01",X"FF",X"21",X"08",X"6E",X"86",X"81",X"01",X"FF",X"81",
		X"ED",X"6E",X"86",X"71",X"01",X"FF",X"71",X"3E",X"6F",X"86",X"8F",X"01",X"FF",X"7F",X"95",X"6F",
		X"84",X"41",X"01",X"FF",X"41",X"D4",X"72",X"84",X"81",X"01",X"FF",X"81",X"B1",X"6B",X"84",X"81",
		X"01",X"FF",X"81",X"C5",X"6A",X"84",X"81",X"01",X"FF",X"81",X"46",X"6B",X"84",X"81",X"01",X"FF",
		X"81",X"3F",X"6C",X"84",X"81",X"01",X"FF",X"81",X"5F",X"6C",X"84",X"71",X"01",X"FF",X"71",X"6D",
		X"6B",X"86",X"91",X"01",X"FF",X"91",X"8C",X"6B",X"84",X"81",X"01",X"FF",X"81",X"08",X"73",X"00",
		X"00",X"FF",X"3E",X"6A",X"00",X"00",X"FF",X"43",X"6A",X"00",X"00",X"FF",X"45",X"6A",X"FA",X"C8",
		X"63",X"10",X"00",X"21",X"00",X"12",X"00",X"00",X"00",X"FF",X"83",X"6A",X"00",X"00",X"FF",X"87",
		X"6A",X"00",X"00",X"FF",X"8A",X"6A",X"00",X"00",X"FF",X"8D",X"6A",X"00",X"00",X"FF",X"90",X"6A",
		X"00",X"00",X"FF",X"98",X"6A",X"00",X"00",X"FF",X"9C",X"6A",X"00",X"00",X"FF",X"9F",X"6A",X"00",
		X"00",X"FF",X"A3",X"6A",X"00",X"00",X"FF",X"A7",X"6A",X"00",X"00",X"FF",X"AB",X"6A",X"00",X"00",
		X"FF",X"AE",X"6A",X"80",X"81",X"80",X"00",X"80",X"FF",X"00",X"80",X"B0",X"00",X"F0",X"E0",X"00",
		X"80",X"7C",X"85",X"7F",X"81",X"7F",X"80",X"00",X"F0",X"F1",X"F0",X"00",X"80",X"D0",X"00",X"F0",
		X"D0",X"F0",X"00",X"F0",X"90",X"F0",X"00",X"F0",X"B0",X"F0",X"00",X"80",X"B0",X"00",X"B0",X"80",
		X"00",X"01",X"80",X"90",X"A0",X"F7",X"FF",X"00",X"3F",X"40",X"60",X"8F",X"F4",X"08",X"02",X"F8",
		X"01",X"05",X"F7",X"FE",X"00",X"3F",X"40",X"40",X"8F",X"F4",X"09",X"02",X"F8",X"01",X"06",X"F7",
		X"FE",X"00",X"18",X"40",X"20",X"8E",X"50",X"24",X"F7",X"FC",X"9E",X"F4",X"01",X"01",X"F5",X"01",
		X"01",X"F8",X"01",X"18",X"F9",X"01",X"18",X"18",X"40",X"20",X"50",X"24",X"18",X"40",X"20",X"50",
		X"24",X"00",X"10",X"40",X"00",X"8F",X"50",X"10",X"F7",X"FC",X"9F",X"F4",X"01",X"01",X"F5",X"01",
		X"01",X"F8",X"01",X"0C",X"F9",X"01",X"0C",X"10",X"40",X"00",X"50",X"10",X"10",X"40",X"00",X"50",
		X"10",X"10",X"40",X"00",X"50",X"10",X"10",X"40",X"00",X"50",X"10",X"10",X"40",X"00",X"50",X"10",
		X"00",X"08",X"40",X"60",X"8E",X"50",X"50",X"F7",X"FC",X"9E",X"F4",X"02",X"01",X"F5",X"02",X"01",
		X"F8",X"01",X"07",X"F9",X"01",X"07",X"08",X"40",X"60",X"50",X"50",X"08",X"40",X"60",X"50",X"50",
		X"08",X"40",X"60",X"50",X"50",X"00",X"05",X"40",X"10",X"50",X"12",X"60",X"14",X"8E",X"9E",X"AE",
		X"F4",X"04",X"01",X"F5",X"04",X"01",X"F6",X"04",X"01",X"F8",X"01",X"06",X"F9",X"01",X"06",X"FA",
		X"01",X"06",X"F7",X"F8",X"F0",X"34",X"40",X"20",X"50",X"22",X"60",X"24",X"00",X"1C",X"41",X"80",
		X"51",X"84",X"8E",X"9E",X"F7",X"F8",X"F4",X"06",X"01",X"F5",X"06",X"01",X"60",X"85",X"F6",X"06",
		X"01",X"AE",X"F8",X"01",X"07",X"F9",X"01",X"07",X"FA",X"01",X"07",X"00",X"22",X"46",X"80",X"56",
		X"90",X"80",X"90",X"F7",X"FC",X"F8",X"02",X"02",X"F9",X"02",X"02",X"3F",X"F8",X"01",X"07",X"F9",
		X"01",X"07",X"20",X"00",X"3F",X"40",X"30",X"8F",X"F4",X"05",X"02",X"F8",X"01",X"04",X"F7",X"FE",
		X"00",X"08",X"40",X"60",X"8E",X"50",X"50",X"F7",X"FC",X"9E",X"F4",X"02",X"01",X"F5",X"02",X"01",
		X"F8",X"01",X"06",X"F9",X"01",X"06",X"09",X"40",X"60",X"50",X"50",X"08",X"40",X"60",X"50",X"50",
		X"08",X"40",X"60",X"50",X"50",X"08",X"40",X"60",X"50",X"50",X"00",X"08",X"40",X"00",X"8E",X"50",
		X"10",X"F7",X"FC",X"9E",X"F4",X"01",X"01",X"F5",X"01",X"01",X"F8",X"01",X"06",X"F9",X"01",X"06",
		X"09",X"40",X"00",X"50",X"10",X"08",X"40",X"00",X"50",X"10",X"08",X"40",X"00",X"50",X"10",X"08",
		X"40",X"00",X"50",X"10",X"08",X"40",X"00",X"50",X"10",X"00",X"18",X"47",X"40",X"8F",X"57",X"50",
		X"F7",X"FC",X"9F",X"F4",X"03",X"01",X"F5",X"03",X"01",X"00",X"3F",X"40",X"10",X"50",X"13",X"8E",
		X"9E",X"F7",X"FC",X"F4",X"0A",X"01",X"F5",X"0A",X"01",X"14",X"F8",X"01",X"04",X"F9",X"01",X"04",
		X"F4",X"0B",X"01",X"F5",X"0B",X"01",X"29",X"00",X"01",X"40",X"60",X"8E",X"F7",X"FE",X"00",X"3F",
		X"40",X"10",X"50",X"14",X"60",X"24",X"8E",X"9E",X"AE",X"F4",X"04",X"01",X"F5",X"04",X"01",X"F6",
		X"04",X"01",X"F8",X"01",X"05",X"F9",X"01",X"05",X"F7",X"F8",X"FA",X"01",X"05",X"3F",X"00",X"3F",
		X"40",X"10",X"50",X"14",X"60",X"24",X"80",X"90",X"A0",X"F4",X"04",X"01",X"F5",X"04",X"01",X"F6",
		X"04",X"01",X"F8",X"02",X"04",X"F9",X"02",X"04",X"FA",X"02",X"04",X"F7",X"F8",X"3F",X"3F",X"F8",
		X"01",X"17",X"F9",X"01",X"17",X"FA",X"01",X"17",X"F0",X"A0",X"00",X"0C",X"F7",X"F8",X"8E",X"9E",
		X"AE",X"F8",X"00",X"05",X"F9",X"00",X"05",X"FA",X"00",X"05",X"41",X"66",X"51",X"DE",X"62",X"CD",
		X"F4",X"00",X"08",X"F5",X"00",X"08",X"06",X"F7",X"FC",X"41",X"66",X"51",X"DE",X"8E",X"9E",X"12",
		X"F7",X"F8",X"8E",X"9E",X"AE",X"40",X"EF",X"51",X"66",X"63",X"BD",X"12",X"F7",X"FB",X"AE",X"62",
		X"CD",X"06",X"F7",X"F8",X"8E",X"9E",X"AE",X"40",X"FD",X"51",X"2D",X"63",X"BD",X"06",X"F7",X"FC",
		X"8E",X"9E",X"40",X"EF",X"51",X"1C",X"06",X"F3",X"39",X"8D",X"9D",X"40",X"D5",X"51",X"0C",X"12",
		X"F7",X"F8",X"40",X"EF",X"51",X"1C",X"62",X"CD",X"8E",X"9E",X"AE",X"F8",X"00",X"06",X"F9",X"00",
		X"06",X"FA",X"00",X"06",X"12",X"AE",X"63",X"BD",X"F8",X"00",X"05",X"F9",X"00",X"05",X"FA",X"00",
		X"05",X"09",X"AE",X"62",X"CD",X"09",X"AE",X"63",X"BD",X"09",X"AE",X"63",X"54",X"09",X"AE",X"62",
		X"F7",X"0C",X"8D",X"9D",X"AE",X"41",X"66",X"51",X"DE",X"62",X"CD",X"06",X"8E",X"9E",X"41",X"66",
		X"51",X"DE",X"12",X"8E",X"9E",X"AE",X"40",X"EF",X"51",X"66",X"63",X"BD",X"F8",X"00",X"06",X"F9",
		X"00",X"06",X"FA",X"00",X"06",X"12",X"AE",X"62",X"CD",X"AE",X"FA",X"00",X"05",X"04",X"8E",X"9E",
		X"AE",X"F8",X"00",X"05",X"F9",X"00",X"05",X"FA",X"00",X"05",X"40",X"D5",X"51",X"0C",X"63",X"BD",
		X"05",X"8E",X"9E",X"40",X"EF",X"51",X"1C",X"05",X"8E",X"9E",X"40",X"FD",X"51",X"2D",X"05",X"8E",
		X"9E",X"40",X"D5",X"51",X"0C",X"36",X"8E",X"9E",X"AE",X"40",X"EF",X"51",X"1C",X"62",X"CD",X"F8",
		X"00",X"08",X"F9",X"00",X"08",X"FA",X"00",X"08",X"00",X"0C",X"F7",X"F8",X"8E",X"9E",X"40",X"EF",
		X"50",X"EC",X"F8",X"00",X"04",X"F9",X"00",X"04",X"06",X"8E",X"9E",X"40",X"EF",X"50",X"EC",X"06",
		X"8F",X"9F",X"AE",X"40",X"C9",X"50",X"C7",X"64",X"B5",X"F8",X"00",X"07",X"F9",X"00",X"07",X"FA",
		X"00",X"04",X"06",X"AE",X"64",X"B5",X"06",X"AE",X"64",X"B5",X"12",X"AE",X"64",X"B5",X"09",X"8E",
		X"9E",X"AF",X"F8",X"00",X"08",X"F9",X"00",X"08",X"40",X"D5",X"50",X"D3",X"64",X"32",X"FA",X"00",
		X"06",X"09",X"8E",X"9E",X"40",X"EF",X"50",X"EC",X"09",X"8E",X"9E",X"AF",X"41",X"0C",X"51",X"0A",
		X"63",X"54",X"09",X"8E",X"9E",X"40",X"D5",X"50",X"D3",X"09",X"F7",X"F8",X"8F",X"9F",X"AF",X"F4",
		X"00",X"04",X"F9",X"00",X"04",X"F8",X"00",X"0F",X"F9",X"00",X"0F",X"FA",X"00",X"04",X"40",X"EF",
		X"50",X"EC",X"62",X"CD",X"09",X"AF",X"63",X"BD",X"09",X"AF",X"62",X"CD",X"09",X"AF",X"63",X"BD",
		X"24",X"AF",X"62",X"CD",X"FA",X"00",X"04",X"00",X"0A",X"F7",X"F8",X"F3",X"39",X"70",X"20",X"41",
		X"66",X"50",X"EF",X"65",X"99",X"0A",X"F3",X"39",X"50",X"FD",X"62",X"CD",X"0A",X"F3",X"39",X"51",
		X"2D",X"65",X"99",X"0A",X"F3",X"39",X"52",X"19",X"61",X"0C",X"0A",X"65",X"99",X"0A",X"F3",X"39",
		X"50",X"FD",X"62",X"CD",X"0A",X"F3",X"39",X"50",X"EF",X"65",X"99",X"0A",X"62",X"CD",X"0A",X"F3",
		X"39",X"50",X"FD",X"64",X"B5",X"0A",X"F3",X"39",X"62",X"5B",X"0A",X"64",X"B5",X"0A",X"F3",X"39",
		X"62",X"5B",X"0A",X"F3",X"39",X"64",X"B5",X"0A",X"62",X"5B",X"0A",X"F3",X"39",X"64",X"B5",X"0A",
		X"F3",X"39",X"62",X"5B",X"0A",X"05",X"F7",X"F8",X"8C",X"9C",X"AC",X"40",X"7F",X"50",X"7C",X"60",
		X"7A",X"05",X"41",X"2D",X"51",X"2B",X"61",X"2A",X"05",X"41",X"66",X"51",X"64",X"61",X"62",X"05",
		X"41",X"AA",X"51",X"A8",X"61",X"A6",X"05",X"41",X"FB",X"51",X"F9",X"61",X"F8",X"05",X"42",X"5B",
		X"52",X"59",X"62",X"58",X"05",X"42",X"CD",X"52",X"CA",X"62",X"C8",X"05",X"43",X"54",X"53",X"52",
		X"63",X"50",X"05",X"43",X"F6",X"53",X"F4",X"63",X"F2",X"05",X"43",X"54",X"53",X"52",X"63",X"50",
		X"05",X"42",X"CD",X"52",X"CB",X"62",X"CA",X"05",X"42",X"5B",X"52",X"59",X"62",X"57",X"05",X"41",
		X"FB",X"51",X"F9",X"61",X"F7",X"05",X"41",X"AA",X"51",X"A8",X"61",X"A6",X"05",X"41",X"66",X"51",
		X"64",X"61",X"62",X"05",X"41",X"2D",X"51",X"2B",X"61",X"29",X"05",X"F7",X"F8",X"F3",X"39",X"70",
		X"10",X"41",X"66",X"50",X"FD",X"63",X"F6",X"20",X"F3",X"39",X"70",X"10",X"00",X"08",X"F7",X"F8",
		X"8F",X"9F",X"AF",X"40",X"B3",X"F8",X"00",X"07",X"08",X"50",X"A9",X"F9",X"00",X"07",X"9F",X"08",
		X"60",X"97",X"FA",X"00",X"07",X"AF",X"08",X"40",X"86",X"F8",X"00",X"07",X"8F",X"08",X"50",X"7F",
		X"F9",X"00",X"07",X"9F",X"08",X"60",X"71",X"FA",X"00",X"07",X"AF",X"08",X"40",X"65",X"F8",X"00",
		X"07",X"8F",X"08",X"50",X"5F",X"F9",X"00",X"07",X"9F",X"08",X"60",X"5A",X"FA",X"00",X"07",X"AF",
		X"F0",X"20",X"40",X"55",X"8F",X"F0",X"48",X"57",X"EB",X"9F",X"67",X"E0",X"AF",X"00",X"08",X"F7",
		X"F8",X"8F",X"9F",X"AF",X"40",X"C9",X"F8",X"00",X"07",X"08",X"50",X"FD",X"F9",X"00",X"07",X"08",
		X"60",X"EF",X"FA",X"00",X"07",X"08",X"41",X"3F",X"F8",X"00",X"07",X"8F",X"08",X"51",X"0C",X"F9",
		X"00",X"07",X"9F",X"08",X"61",X"52",X"FA",X"00",X"07",X"AF",X"08",X"41",X"3F",X"F8",X"00",X"07",
		X"8F",X"08",X"51",X"92",X"F9",X"00",X"07",X"9F",X"08",X"61",X"DE",X"FA",X"00",X"03",X"AF",X"08",
		X"41",X"DD",X"F8",X"00",X"03",X"8F",X"08",X"51",X"DC",X"F9",X"00",X"05",X"9F",X"38",X"61",X"DE",
		X"FA",X"00",X"07",X"AF",X"00",X"08",X"F7",X"F8",X"F3",X"21",X"70",X"0A",X"8D",X"9D",X"40",X"EF",
		X"50",X"EC",X"63",X"BD",X"08",X"F3",X"21",X"63",X"BD",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",
		X"61",X"DE",X"08",X"F3",X"21",X"40",X"C9",X"50",X"C7",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",
		X"63",X"BD",X"8E",X"9E",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"EF",X"50",X"EC",
		X"61",X"DE",X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",
		X"64",X"32",X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"A0",X"50",X"9D",
		X"62",X"19",X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",
		X"64",X"32",X"8D",X"9D",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"19",X"08",X"F3",X"21",X"80",
		X"90",X"08",X"F3",X"21",X"40",X"EF",X"50",X"EC",X"64",X"B5",X"8D",X"9D",X"08",X"F3",X"21",X"08",
		X"F3",X"21",X"40",X"D5",X"50",X"D3",X"62",X"5B",X"08",X"F3",X"21",X"40",X"C9",X"50",X"C7",X"08",
		X"F3",X"21",X"40",X"D5",X"50",X"D3",X"64",X"B5",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",
		X"40",X"EF",X"50",X"EC",X"62",X"5B",X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",
		X"40",X"EF",X"50",X"EC",X"64",X"FD",X"8D",X"9D",X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"FD",
		X"50",X"FB",X"62",X"7E",X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"EF",X"50",X"EC",X"64",X"FD",
		X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",X"62",X"7E",X"08",X"F3",X"21",X"08",
		X"F7",X"F8",X"F3",X"21",X"70",X"0A",X"8D",X"9D",X"40",X"EF",X"50",X"EC",X"63",X"BD",X"08",X"F3",
		X"21",X"63",X"BD",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",X"61",X"DE",X"08",X"F3",X"21",X"40",
		X"C9",X"50",X"C7",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",X"63",X"BD",X"8E",X"9E",X"08",X"F3",
		X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"EF",X"50",X"EC",X"61",X"DE",X"8D",X"9D",X"08",X"F3",
		X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",X"64",X"32",X"8D",X"9D",X"08",X"F3",
		X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"A0",X"50",X"9D",X"62",X"19",X"8D",X"9D",X"08",X"F3",
		X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"D5",X"50",X"D3",X"64",X"32",X"8D",X"9D",X"08",X"F3",
		X"21",X"08",X"F3",X"21",X"62",X"19",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"C9",
		X"50",X"C7",X"64",X"B5",X"8D",X"9D",X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",
		X"62",X"5B",X"08",X"F3",X"21",X"40",X"A0",X"50",X"9E",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",
		X"64",X"B5",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"C9",X"50",X"C7",X"62",X"5B",
		X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",X"64",X"32",
		X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"86",X"50",X"84",X"62",X"19",
		X"8D",X"9D",X"08",X"F3",X"21",X"80",X"90",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",X"64",X"32",
		X"8D",X"9D",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"19",X"80",X"90",X"08",X"F3",X"21",X"08",
		X"F7",X"F8",X"F3",X"39",X"70",X"0B",X"40",X"6A",X"50",X"00",X"63",X"BD",X"F4",X"00",X"03",X"08",
		X"F3",X"39",X"08",X"F3",X"21",X"80",X"90",X"61",X"DE",X"08",X"F3",X"21",X"08",X"F3",X"39",X"40",
		X"6A",X"50",X"00",X"63",X"BD",X"08",X"F3",X"39",X"08",X"F3",X"21",X"80",X"90",X"61",X"DE",X"08",
		X"F3",X"21",X"08",X"F3",X"39",X"40",X"6A",X"50",X"00",X"64",X"32",X"08",X"F3",X"39",X"08",X"F3",
		X"21",X"80",X"90",X"62",X"19",X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"6A",X"50",X"00",X"64",
		X"32",X"8D",X"9D",X"FF",X"04",X"08",X"F3",X"21",X"40",X"78",X"50",X"76",X"08",X"F3",X"21",X"40",
		X"86",X"50",X"84",X"62",X"19",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",X"08",X"F3",X"21",X"40",
		X"A0",X"50",X"9D",X"64",X"B5",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"5B",X"08",X"F3",X"21",
		X"08",X"F3",X"21",X"64",X"B5",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"5B",X"08",X"F3",X"21",
		X"08",X"F3",X"21",X"64",X"FD",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"7E",X"08",X"F3",X"21",
		X"08",X"F3",X"21",X"64",X"FD",X"80",X"90",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"7E",X"08",
		X"F3",X"21",X"08",X"F3",X"39",X"70",X"0A",X"40",X"6A",X"50",X"00",X"63",X"BD",X"F4",X"00",X"03",
		X"08",X"F3",X"39",X"08",X"F3",X"21",X"80",X"90",X"61",X"DE",X"08",X"F3",X"21",X"08",X"F3",X"39",
		X"40",X"6A",X"50",X"00",X"63",X"BD",X"08",X"F3",X"39",X"08",X"F3",X"21",X"80",X"90",X"61",X"DE",
		X"08",X"F3",X"21",X"08",X"F3",X"39",X"40",X"6A",X"50",X"00",X"64",X"32",X"08",X"F3",X"39",X"08",
		X"F3",X"21",X"80",X"90",X"62",X"19",X"08",X"F3",X"21",X"08",X"F3",X"21",X"40",X"6A",X"50",X"00",
		X"64",X"32",X"8D",X"9D",X"FF",X"04",X"08",X"F3",X"21",X"40",X"78",X"50",X"76",X"08",X"F3",X"21",
		X"40",X"86",X"50",X"84",X"62",X"19",X"08",X"F3",X"21",X"40",X"B3",X"50",X"B0",X"08",X"F3",X"21",
		X"40",X"A0",X"50",X"9D",X"64",X"B5",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"5B",X"08",X"F3",
		X"21",X"08",X"F3",X"21",X"64",X"B5",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"5B",X"08",X"F3",
		X"21",X"08",X"F3",X"21",X"64",X"FD",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"7E",X"08",X"F3",
		X"21",X"08",X"F3",X"21",X"64",X"FD",X"80",X"90",X"08",X"F3",X"21",X"08",X"F3",X"21",X"62",X"7E",
		X"07",X"F3",X"21",X"00",X"07",X"F7",X"F8",X"8F",X"9F",X"AF",X"40",X"EF",X"F8",X"00",X"07",X"07",
		X"50",X"A9",X"F9",X"00",X"07",X"07",X"60",X"A0",X"FA",X"00",X"07",X"07",X"40",X"86",X"8F",X"F8",
		X"00",X"07",X"07",X"50",X"78",X"9F",X"F9",X"00",X"07",X"07",X"60",X"5F",X"FA",X"00",X"07",X"AF",
		X"0E",X"40",X"50",X"F8",X"00",X"07",X"8F",X"00",X"05",X"F7",X"F8",X"8D",X"9D",X"AD",X"F8",X"00",
		X"02",X"F9",X"00",X"02",X"FA",X"00",X"03",X"40",X"EF",X"50",X"77",X"05",X"8D",X"9D",X"40",X"EF",
		X"50",X"77",X"14",X"8D",X"9D",X"AD",X"40",X"EF",X"50",X"77",X"62",X"CD",X"F8",X"00",X"05",X"F9",
		X"00",X"05",X"FA",X"00",X"03",X"14",X"8D",X"9D",X"AD",X"40",X"B3",X"50",X"59",X"63",X"BD",X"14",
		X"8D",X"9D",X"AD",X"40",X"BE",X"50",X"5E",X"62",X"CD",X"14",X"8D",X"9D",X"AD",X"40",X"A0",X"50",
		X"4F",X"63",X"BD",X"14",X"8D",X"9D",X"AD",X"40",X"B3",X"50",X"59",X"62",X"CD",X"05",X"8D",X"9D",
		X"AD",X"F8",X"00",X"08",X"F9",X"00",X"02",X"FA",X"00",X"03",X"40",X"EF",X"50",X"47",X"63",X"BD",
		X"05",X"9D",X"50",X"47",X"0A",X"9D",X"50",X"47",X"05",X"9D",X"AD",X"50",X"43",X"62",X"CD",X"05",
		X"9D",X"50",X"43",X"0A",X"9D",X"50",X"43",X"05",X"9D",X"AD",X"50",X"47",X"63",X"BD",X"05",X"9D",
		X"50",X"47",X"05",X"8D",X"9D",X"F8",X"00",X"02",X"F9",X"00",X"02",X"FA",X"00",X"03",X"40",X"EF",
		X"50",X"47",X"05",X"8D",X"9D",X"40",X"EF",X"50",X"77",X"14",X"8D",X"9D",X"AD",X"F8",X"00",X"05",
		X"F9",X"00",X"05",X"FA",X"00",X"03",X"40",X"EF",X"50",X"77",X"62",X"CD",X"14",X"8D",X"9D",X"AD",
		X"40",X"B3",X"50",X"59",X"63",X"BD",X"14",X"8D",X"9D",X"AD",X"40",X"BE",X"50",X"5E",X"62",X"CD",
		X"14",X"8D",X"9D",X"AD",X"40",X"A0",X"50",X"4F",X"63",X"BD",X"0E",X"8D",X"9D",X"AD",X"40",X"B3",
		X"50",X"8E",X"62",X"CD",X"06",X"8D",X"9D",X"AD",X"40",X"BE",X"50",X"A0",X"63",X"BD",X"F0",X"30",
		X"8D",X"9D",X"AD",X"40",X"8F",X"50",X"B3",X"62",X"CD",X"F8",X"00",X"06",X"F9",X"00",X"06",X"FA",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"15",X"02",X"15",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"15",X"15",X"02",X"15",X"15",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"15",X"15",X"15",X"15",X"15",X"15",X"00",X"00",X"00",X"00",X"00",X"15",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"15",X"00",X"00",X"00",X"00",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",
		X"15",X"00",X"00",X"00",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"00",
		X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"12",X"12",X"11",X"12",X"11",X"12",X"11",X"11",X"11",X"12",X"11",X"11",X"0D",X"0E",
		X"0E",X"0D",X"0E",X"0E",X"0D",X"0E",X"0D",X"0D",X"0E",X"0D",X"0D",X"15",X"16",X"16",X"15",X"16",
		X"15",X"16",X"15",X"15",X"15",X"16",X"15",X"15",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"FF",X"15",X"15",
		X"15",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"00",X"00",X"00",X"FF",X"15",X"15",X"15",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"0D",X"0D",
		X"0D",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"0D",X"0D",X"0D",X"FF",X"00",
		X"00",X"00",X"FF",X"FF",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"03",X"03",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"52",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",
		X"03",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"0A",X"0A",X"0A",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"16",X"16",X"16",X"16",X"16",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"1A",X"1A",X"1A",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"E7",X"DD",X"79",X"06",X"E7",X"09",X"7A",X"06",X"E7",X"67",X"7A",X"06",X"E7",
		X"A3",X"7A",X"06",X"E7",X"04",X"7B",X"06",X"E7",X"38",X"7B",X"88",X"E4",X"81",X"7B",X"50",X"E7",
		X"88",X"7B",X"AF",X"32",X"00",X"EC",X"32",X"04",X"EC",X"E7",X"26",X"D0",X"2E",X"0C",X"CB",X"76",
		X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",
		X"7E",X"E1",X"32",X"18",X"D0",X"3A",X"00",X"EC",X"A7",X"28",X"DE",X"F5",X"E6",X"C0",X"FE",X"40",
		X"CA",X"C4",X"77",X"F1",X"FE",X"87",X"20",X"08",X"3E",X"08",X"32",X"04",X"EC",X"3A",X"00",X"EC",
		X"CB",X"7F",X"0E",X"00",X"20",X"05",X"3D",X"28",X"02",X"0E",X"FF",X"3A",X"00",X"EC",X"21",X"C2",
		X"76",X"E6",X"0F",X"3D",X"CB",X"41",X"28",X"01",X"3D",X"CB",X"27",X"CB",X"27",X"CD",X"56",X"20",
		X"ED",X"53",X"02",X"EC",X"AF",X"23",X"CD",X"56",X"20",X"2A",X"02",X"EC",X"3E",X"02",X"32",X"01",
		X"EC",X"1A",X"47",X"13",X"1A",X"13",X"FE",X"40",X"20",X"10",X"2A",X"02",X"EC",X"23",X"23",X"23",
		X"23",X"22",X"02",X"EC",X"CB",X"41",X"20",X"41",X"18",X"1E",X"CB",X"41",X"28",X"0F",X"36",X"E3",
		X"23",X"36",X"38",X"CD",X"03",X"21",X"10",X"DC",X"0E",X"00",X"C3",X"2B",X"77",X"F5",X"3A",X"04",
		X"EC",X"77",X"23",X"F1",X"77",X"CD",X"03",X"21",X"3A",X"01",X"EC",X"DF",X"E5",X"26",X"D0",X"2E",
		X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",
		X"CD",X"50",X"20",X"7E",X"E1",X"E1",X"32",X"18",X"D0",X"10",X"A9",X"C3",X"E2",X"76",X"20",X"39",
		X"E0",X"3A",X"A0",X"3C",X"40",X"70",X"00",X"72",X"C0",X"73",X"80",X"75",X"40",X"77",X"00",X"79",
		X"C0",X"7A",X"80",X"7C",X"F1",X"AF",X"32",X"05",X"EC",X"3E",X"01",X"32",X"06",X"EC",X"CD",X"17",
		X"21",X"21",X"A0",X"E4",X"11",X"47",X"7C",X"AF",X"CD",X"B1",X"79",X"3E",X"3C",X"DF",X"CD",X"17",
		X"21",X"3E",X"FF",X"3A",X"7B",X"C4",X"CB",X"AF",X"CB",X"B7",X"32",X"7B",X"C4",X"21",X"0C",X"E4",
		X"AF",X"CD",X"98",X"79",X"21",X"E4",X"E3",X"11",X"4F",X"7C",X"AF",X"CD",X"B1",X"79",X"21",X"2E",
		X"E3",X"11",X"69",X"7C",X"AF",X"CD",X"B1",X"79",X"3E",X"96",X"DF",X"CD",X"17",X"21",X"3E",X"FF",
		X"21",X"24",X"E4",X"3E",X"01",X"CD",X"98",X"79",X"21",X"10",X"E6",X"11",X"72",X"7C",X"AF",X"CD",
		X"B1",X"79",X"21",X"5A",X"E4",X"11",X"97",X"7C",X"AF",X"CD",X"B1",X"79",X"3E",X"96",X"DF",X"CD",
		X"17",X"21",X"3E",X"FF",X"21",X"4C",X"E1",X"3E",X"02",X"CD",X"98",X"79",X"21",X"26",X"E7",X"11",
		X"A0",X"7C",X"AF",X"CD",X"B1",X"79",X"21",X"6C",X"E5",X"11",X"B5",X"7C",X"AF",X"CD",X"B1",X"79",
		X"3E",X"96",X"DF",X"CD",X"17",X"21",X"3E",X"FF",X"3A",X"7B",X"C4",X"CB",X"EF",X"32",X"7B",X"C4",
		X"21",X"64",X"E1",X"3E",X"03",X"CD",X"98",X"79",X"21",X"12",X"E7",X"11",X"BC",X"7C",X"AF",X"CD",
		X"B1",X"79",X"21",X"1A",X"E6",X"11",X"CD",X"7C",X"AF",X"CD",X"B1",X"79",X"3E",X"96",X"DF",X"CD",
		X"17",X"21",X"3E",X"FF",X"21",X"4C",X"E1",X"3E",X"04",X"CD",X"98",X"79",X"21",X"0C",X"E7",X"11",
		X"D7",X"7C",X"AF",X"CD",X"B1",X"79",X"21",X"D6",X"E6",X"11",X"E6",X"7C",X"AF",X"CD",X"B1",X"79",
		X"3E",X"32",X"DF",X"21",X"24",X"E4",X"3E",X"05",X"CD",X"98",X"79",X"21",X"A8",X"E2",X"11",X"EE",
		X"7C",X"AF",X"CD",X"B1",X"79",X"21",X"32",X"E3",X"11",X"FC",X"7C",X"AF",X"CD",X"B1",X"79",X"3E",
		X"64",X"DF",X"CD",X"17",X"21",X"3E",X"FF",X"21",X"0C",X"E4",X"3E",X"06",X"CD",X"98",X"79",X"21",
		X"8A",X"E2",X"11",X"07",X"7D",X"AF",X"CD",X"B1",X"79",X"21",X"56",X"E2",X"11",X"18",X"7D",X"AF",
		X"CD",X"B1",X"79",X"3E",X"32",X"DF",X"21",X"64",X"E1",X"3E",X"07",X"CD",X"98",X"79",X"21",X"28",
		X"E7",X"11",X"1F",X"7D",X"AF",X"CD",X"B1",X"79",X"21",X"32",X"E7",X"11",X"31",X"7D",X"AF",X"CD",
		X"B1",X"79",X"3E",X"64",X"DF",X"CD",X"17",X"21",X"3E",X"FF",X"21",X"4C",X"E1",X"3E",X"09",X"CD",
		X"98",X"79",X"21",X"0C",X"E7",X"11",X"57",X"7D",X"AF",X"CD",X"B1",X"79",X"21",X"16",X"E7",X"11",
		X"6B",X"7D",X"AF",X"CD",X"B1",X"79",X"3E",X"32",X"DF",X"21",X"24",X"E4",X"3E",X"08",X"CD",X"98",
		X"79",X"21",X"28",X"E3",X"11",X"3A",X"7D",X"AF",X"CD",X"B1",X"79",X"21",X"B2",X"E2",X"11",X"4F",
		X"7D",X"AF",X"CD",X"B1",X"79",X"3E",X"64",X"DF",X"CD",X"17",X"21",X"3E",X"FF",X"21",X"0C",X"E4",
		X"3E",X"0A",X"CD",X"98",X"79",X"21",X"A6",X"E4",X"11",X"77",X"7D",X"AF",X"CD",X"B1",X"79",X"21",
		X"6C",X"E3",X"11",X"88",X"7D",X"AF",X"CD",X"B1",X"79",X"3E",X"C8",X"DF",X"CD",X"17",X"21",X"3A",
		X"7B",X"C4",X"CB",X"AF",X"32",X"7B",X"C4",X"21",X"32",X"E5",X"11",X"90",X"7D",X"AF",X"CD",X"B1",
		X"79",X"21",X"F8",X"E5",X"11",X"9C",X"7D",X"AF",X"CD",X"B1",X"79",X"3E",X"FA",X"DF",X"CD",X"17",
		X"21",X"AF",X"32",X"00",X"EC",X"C3",X"E2",X"76",X"E5",X"E6",X"0F",X"CB",X"27",X"21",X"AE",X"77",
		X"CD",X"56",X"20",X"E1",X"01",X"07",X"08",X"EB",X"CD",X"D1",X"20",X"3E",X"B8",X"CD",X"55",X"22",
		X"C9",X"32",X"04",X"EC",X"1A",X"47",X"13",X"22",X"02",X"EC",X"1A",X"13",X"FE",X"40",X"20",X"0C",
		X"2A",X"02",X"EC",X"23",X"23",X"23",X"23",X"22",X"02",X"EC",X"18",X"0B",X"F5",X"3A",X"04",X"EC",
		X"77",X"23",X"F1",X"77",X"CD",X"03",X"21",X"3E",X"02",X"DF",X"10",X"DE",X"C9",X"2B",X"54",X"48",
		X"45",X"20",X"45",X"52",X"41",X"20",X"41",X"4E",X"44",X"20",X"54",X"49",X"4D",X"45",X"20",X"4F",
		X"46",X"20",X"40",X"54",X"48",X"49",X"53",X"20",X"53",X"54",X"4F",X"52",X"59",X"20",X"49",X"53",
		X"20",X"55",X"4E",X"4B",X"4E",X"4F",X"57",X"4E",X"2E",X"5D",X"41",X"46",X"54",X"45",X"52",X"20",
		X"54",X"48",X"45",X"20",X"4D",X"4F",X"54",X"48",X"45",X"52",X"53",X"48",X"49",X"50",X"20",X"40",
		X"22",X"41",X"52",X"4B",X"41",X"4E",X"4F",X"49",X"44",X"22",X"20",X"57",X"41",X"53",X"20",X"44",
		X"45",X"53",X"54",X"52",X"4F",X"59",X"45",X"44",X"2C",X"20",X"40",X"41",X"20",X"53",X"50",X"41",
		X"43",X"45",X"43",X"52",X"41",X"46",X"54",X"20",X"22",X"56",X"41",X"55",X"53",X"22",X"20",X"40",
		X"53",X"43",X"52",X"41",X"4D",X"42",X"4C",X"45",X"44",X"20",X"41",X"57",X"41",X"59",X"20",X"46",
		X"52",X"4F",X"4D",X"20",X"49",X"54",X"2E",X"3B",X"42",X"55",X"54",X"20",X"4F",X"4E",X"4C",X"59",
		X"20",X"54",X"4F",X"20",X"42",X"45",X"20",X"40",X"54",X"52",X"41",X"50",X"50",X"45",X"44",X"20",
		X"49",X"4E",X"20",X"53",X"50",X"41",X"43",X"45",X"20",X"57",X"41",X"52",X"50",X"45",X"44",X"20",
		X"40",X"42",X"59",X"20",X"53",X"4F",X"4D",X"45",X"4F",X"4E",X"45",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"60",X"44",X"49",X"4D",X"45",X"4E",X"53",X"49",X"4F",X"4E",X"2D",X"43",X"4F",
		X"4E",X"54",X"52",X"4F",X"4C",X"4C",X"49",X"4E",X"47",X"20",X"46",X"4F",X"52",X"54",X"20",X"40",
		X"22",X"44",X"4F",X"48",X"22",X"20",X"48",X"41",X"53",X"20",X"4E",X"4F",X"57",X"20",X"42",X"45",
		X"45",X"4E",X"20",X"40",X"44",X"45",X"4D",X"4F",X"4C",X"49",X"53",X"48",X"45",X"44",X"2C",X"20",
		X"41",X"4E",X"44",X"20",X"54",X"49",X"4D",X"45",X"20",X"40",X"53",X"54",X"41",X"52",X"54",X"45",
		X"44",X"20",X"46",X"4C",X"4F",X"57",X"49",X"4E",X"47",X"20",X"52",X"45",X"56",X"45",X"52",X"53",
		X"45",X"4C",X"59",X"2E",X"33",X"22",X"56",X"41",X"55",X"53",X"22",X"20",X"4D",X"41",X"4E",X"41",
		X"47",X"45",X"44",X"20",X"54",X"4F",X"20",X"45",X"53",X"43",X"41",X"50",X"45",X"20",X"40",X"46",
		X"52",X"4F",X"4D",X"20",X"54",X"48",X"45",X"20",X"44",X"49",X"53",X"54",X"4F",X"52",X"54",X"45",
		X"44",X"20",X"53",X"50",X"41",X"43",X"45",X"2E",X"48",X"42",X"55",X"54",X"20",X"54",X"48",X"45",
		X"20",X"52",X"45",X"41",X"4C",X"20",X"56",X"4F",X"59",X"41",X"47",X"45",X"20",X"4F",X"46",X"20",
		X"40",X"22",X"41",X"52",X"4B",X"41",X"4E",X"4F",X"49",X"44",X"22",X"20",X"49",X"4E",X"20",X"54",
		X"48",X"45",X"20",X"47",X"41",X"4C",X"41",X"58",X"59",X"20",X"40",X"48",X"41",X"53",X"20",X"4F",
		X"4E",X"4C",X"59",X"20",X"53",X"54",X"41",X"52",X"54",X"45",X"44",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"06",X"4E",X"4F",X"54",X"49",X"43",X"45",X"BE",X"54",X"48",X"49",X"53",X"20",X"47",X"41",
		X"4D",X"45",X"20",X"49",X"53",X"20",X"46",X"4F",X"52",X"20",X"55",X"53",X"45",X"20",X"49",X"4E",
		X"20",X"40",X"4A",X"41",X"50",X"41",X"4E",X"20",X"4F",X"4E",X"4C",X"59",X"2E",X"40",X"53",X"41",
		X"4C",X"45",X"53",X"2C",X"20",X"45",X"58",X"50",X"4F",X"52",X"54",X"2C",X"20",X"4F",X"52",X"20",
		X"4F",X"50",X"45",X"52",X"41",X"54",X"49",X"4F",X"4E",X"40",X"4F",X"55",X"54",X"53",X"49",X"44",
		X"45",X"20",X"54",X"48",X"49",X"53",X"20",X"54",X"45",X"52",X"52",X"49",X"54",X"4F",X"52",X"59",
		X"20",X"40",X"4D",X"41",X"59",X"20",X"56",X"49",X"4F",X"4C",X"41",X"54",X"45",X"20",X"49",X"4E",
		X"54",X"45",X"52",X"4E",X"41",X"54",X"49",X"4F",X"4E",X"41",X"4C",X"40",X"43",X"4F",X"50",X"59",
		X"52",X"49",X"47",X"48",X"54",X"20",X"41",X"4E",X"44",X"20",X"54",X"52",X"41",X"44",X"45",X"4D",
		X"41",X"52",X"4B",X"40",X"4C",X"41",X"57",X"53",X"20",X"41",X"4E",X"44",X"20",X"54",X"48",X"45",
		X"20",X"56",X"49",X"4F",X"4C",X"41",X"54",X"4F",X"52",X"20",X"40",X"53",X"55",X"42",X"4A",X"45",
		X"43",X"54",X"20",X"54",X"4F",X"20",X"53",X"45",X"56",X"45",X"52",X"45",X"20",X"50",X"45",X"4E",
		X"41",X"4C",X"54",X"49",X"45",X"53",X"2E",X"07",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"19",
		X"44",X"49",X"52",X"45",X"43",X"54",X"45",X"44",X"20",X"26",X"20",X"40",X"50",X"52",X"4F",X"47",
		X"52",X"41",X"4D",X"4D",X"45",X"44",X"20",X"42",X"59",X"08",X"59",X"2E",X"53",X"41",X"53",X"41",
		X"42",X"45",X"24",X"44",X"49",X"52",X"45",X"43",X"54",X"45",X"52",X"20",X"4F",X"46",X"20",X"48",
		X"41",X"52",X"44",X"57",X"41",X"52",X"45",X"20",X"26",X"40",X"43",X"4F",X"2D",X"50",X"52",X"4F",
		X"47",X"52",X"41",X"4D",X"4D",X"45",X"52",X"08",X"54",X"2E",X"53",X"41",X"4E",X"41",X"44",X"41",
		X"14",X"41",X"53",X"53",X"49",X"53",X"54",X"41",X"4E",X"54",X"20",X"50",X"52",X"4F",X"47",X"52",
		X"41",X"4D",X"4D",X"45",X"52",X"06",X"54",X"4F",X"52",X"55",X"2E",X"54",X"10",X"47",X"52",X"41",
		X"50",X"48",X"49",X"43",X"20",X"44",X"45",X"53",X"49",X"47",X"4E",X"45",X"52",X"09",X"4F",X"4E",
		X"49",X"4A",X"55",X"53",X"54",X"2E",X"48",X"0E",X"53",X"4F",X"55",X"4E",X"44",X"40",X"43",X"4F",
		X"4D",X"50",X"4F",X"53",X"45",X"52",X"07",X"48",X"2E",X"4F",X"47",X"55",X"52",X"41",X"0D",X"53",
		X"4F",X"55",X"4E",X"44",X"40",X"45",X"46",X"46",X"45",X"43",X"54",X"53",X"0A",X"54",X"2E",X"4B",
		X"49",X"4D",X"49",X"4A",X"49",X"4D",X"41",X"10",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"40",
		X"44",X"45",X"53",X"49",X"47",X"4E",X"45",X"52",X"06",X"41",X"2E",X"49",X"57",X"41",X"49",X"11",
		X"53",X"4F",X"46",X"54",X"57",X"41",X"52",X"45",X"40",X"41",X"4E",X"41",X"4C",X"59",X"5A",X"45",
		X"52",X"08",X"48",X"49",X"44",X"45",X"47",X"4F",X"4E",X"53",X"14",X"50",X"55",X"42",X"4C",X"49",
		X"43",X"49",X"54",X"59",X"40",X"53",X"55",X"50",X"45",X"52",X"56",X"49",X"53",X"4F",X"52",X"07",
		X"56",X"41",X"52",X"49",X"53",X"2E",X"49",X"13",X"4D",X"45",X"43",X"48",X"41",X"4E",X"49",X"43",
		X"41",X"4C",X"40",X"45",X"4E",X"47",X"49",X"4E",X"45",X"45",X"52",X"0B",X"48",X"2E",X"59",X"41",
		X"4D",X"41",X"47",X"55",X"43",X"48",X"49",X"10",X"47",X"41",X"4D",X"45",X"20",X"44",X"45",X"53",
		X"49",X"47",X"4E",X"45",X"44",X"20",X"42",X"59",X"07",X"41",X"4B",X"49",X"52",X"41",X"2E",X"46",
		X"0B",X"50",X"52",X"4F",X"44",X"55",X"43",X"45",X"44",X"20",X"42",X"59",X"11",X"54",X"41",X"49",
		X"54",X"4F",X"20",X"43",X"4F",X"52",X"50",X"4F",X"52",X"41",X"54",X"49",X"4F",X"4E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"1E",X"1D",X"1D",X"1D",X"1D",X"1D",
		X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1E",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"18",X"C7",X"00",X"1B",X"C6",X"00",X"1B",X"C7",
		X"00",X"10",X"15",X"02",X"B6",X"00",X"14",X"02",X"AE",X"FF",X"BF",X"04",X"CB",X"00",X"1A",X"24",
		X"02",X"3C",X"10",X"B7",X"00",X"17",X"02",X"16",X"02",X"03",X"02",X"FD",X"C6",X"00",X"10",X"B7",
		X"00",X"17",X"02",X"16",X"02",X"03",X"02",X"FD",X"80",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"02",
		X"B6",X"00",X"14",X"02",X"97",X"47",X"CB",X"00",X"17",X"C7",X"00",X"19",X"01",X"02",X"FD",X"2F",
		X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"4D",X"27",X"0A",X"C7",X"00",X"17",X"CB",X"00",X"10",
		X"97",X"C7",X"00",X"16",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"02",X"B6",X"00",X"14",X"02",X"C7",
		X"00",X"1A",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"A6",X"FF",X"B7",X"02",X"A6",X"FC",X"B7",X"06",
		X"A6",X"00",X"B7",X"05",X"AE",X"80",X"3F",X"10",X"F6",X"CB",X"00",X"10",X"C7",X"00",X"10",X"5C",
		X"26",X"F6",X"A6",X"FF",X"B7",X"04",X"C6",X"00",X"10",X"B7",X"00",X"17",X"02",X"16",X"02",X"03",
		X"02",X"FD",X"AE",X"13",X"7F",X"A6",X"C0",X"E7",X"01",X"3F",X"11",X"3F",X"12",X"3F",X"15",X"3F",
		X"16",X"3F",X"17",X"12",X"11",X"9A",X"02",X"11",X"FD",X"9B",X"A6",X"FF",X"B7",X"04",X"A6",X"55",
		X"B7",X"00",X"17",X"02",X"16",X"02",X"03",X"02",X"FD",X"4F",X"B7",X"00",X"17",X"02",X"16",X"02",
		X"03",X"02",X"FD",X"9A",X"21",X"FE",X"20",X"FC",X"01",X"02",X"FD",X"2F",X"FB",X"15",X"02",X"B6",
		X"00",X"14",X"02",X"97",X"A6",X"FF",X"B7",X"04",X"C6",X"00",X"16",X"CA",X"00",X"17",X"27",X"08",
		X"C6",X"00",X"18",X"C7",X"00",X"19",X"20",X"0A",X"02",X"03",X"02",X"FD",X"C6",X"00",X"10",X"A4",
		X"0F",X"97",X"D6",X"03",X"5D",X"B7",X"00",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",
		X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"15",X"15",X"15",X"15",X"15",X"15",X"FF",X"FF",X"FF",
		X"FF",X"19",X"FF",X"19",X"FF",X"FF",X"FF",X"FF",X"15",X"15",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"15",X"15",X"FF",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"FF",X"16",X"15",X"FF",X"19",X"1A",X"00",X"00",X"00",X"00",X"00",X"1A",X"19",X"FF",X"15");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
