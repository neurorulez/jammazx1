-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "E3FF7FFFFF80F000F3FFF3FF0850BD7F41FFFFFF3FFFCFFFFFFFFFFFFFFF3FFF";
    attribute INIT_01 of inst : label is "0F000A00FFFFFFFFFFFEFA00FFF0F87F004AD00CC800C000F400FFFFFFFFFFFF";
    attribute INIT_02 of inst : label is "C400C100FFFF0002FFE1E80F044A01CC0000001F0000D0002430010001E0A000";
    attribute INIT_03 of inst : label is "C000F500003A05F0FF63FFFEC000F500003A05F0FF00FF00FFFFFFF8FFFF0000";
    attribute INIT_04 of inst : label is "1CF07FFCBE003F99805F1FFFFC0AA0000080021F0000D0802430010000000000";
    attribute INIT_05 of inst : label is "01E0A000FFFFFFFFFFF3D52FFFFF7E163FEFC5FF3FFFFFFF000000003FA2FFFB";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "2F08F5473FFFCFFF3E07687FFEA42A002FFF8D400F000A002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A1FA002FF";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "F7F3FFFFF3FDFFFFCFCFFFFFFFCFFFFFFFFFFFFF01F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFE8F2FFFFFF75FFBEF02BAFB8BAAD1FFFF413FCCFFFFFF6CFCFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFF4ABFFD2FFFF2FFFF4FFFFFFC57FFFFCE11BFFFFDA8FFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFCFE1F7FFF5FFFFFFFFFFFFFA8AA15FFFFAAAAFFFFD552FFFF";
    attribute INIT_0F of inst : label is "FFFCFFF3FFFFFFFFFFFFFFFFFCFFFF3FFF3FFFCFFFF3FFF3FFFCFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "00000000FFFCFFFFFFFFFFFF3FFF3FFFF3FFCFFFFCFFF3FFFF3FFF3FFFF3FFCF";
    attribute INIT_11 of inst : label is "00000000C000C00000030003C000C0000003000300C0AA80030002AA00000000";
    attribute INIT_12 of inst : label is "FC00FF00C000F0000003000F0000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFCFFFFFFC0FFF003FF0FFF003F00FF";
    attribute INIT_14 of inst : label is "00FF1FFF0780F7000003000BFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF";
    attribute INIT_15 of inst : label is "1110FF80F400E0007FFFFFFF001F07FF00000001F508FFFFFCB8FDFD7FF84007";
    attribute INIT_16 of inst : label is "FFFFFFFF21BF0C7FFEB9FCC2FF1D09FFFFFFFFFF7CFF87FFFF4BFFF441DEFCFF";
    attribute INIT_17 of inst : label is "35000EFFFFFFFD6AFF9B5000FFFFFFFF0000000067FF2FFF00000000CC5BDD5F";
    attribute INIT_18 of inst : label is "C2177FFF00000000DBEE5555D0AFFFFDFFFD2F5BFFA5CDBFFF6FFA00002A0000";
    attribute INIT_19 of inst : label is "F000E0003F317F7700020000F00080006FFFFF6B000707FF5AFF2FF3FF5AFFFC";
    attribute INIT_1A of inst : label is "F000F00017FF57FF33337DFFFFFCFFFF0000000000000554F000F0000000FFFC";
    attribute INIT_1B of inst : label is "0F400FFF3C003C00F000F0000FE03C00FFFFEFFF000010000FFF0FFF0FFF0FFF";
    attribute INIT_1C of inst : label is "F3C0F0BDFFFFFFFFF000F5550000F000000000000000000403FC03FCFFFFFFFF";
    attribute INIT_1D of inst : label is "F0BF0342FFACC2D0A00B55FF1FFFFFFFE00F001FFFFF2F2FA050FFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "CCB8FFFFFFAF015F00FFFFFF0000FFFFFFFFBFE800FFFFFFFFFF0BFFFFFF8000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC2FFF0FFFFFFFFFFFA";
    attribute INIT_20 of inst : label is "002A00E000000000A0006C000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0B4BBF7FFC0000F08380F7F000FE0C0012D50415000000005784540400000000";
    attribute INIT_22 of inst : label is "034A3FFF0FF800308380FBF02FF00C000FC003F800FF2E00E4002FC0FF000000";
    attribute INIT_23 of inst : label is "003F003F003F01D7E000FC00FC0099807FB0006F003FBF340E3FEAD0F0001CA8";
    attribute INIT_24 of inst : label is "03F001AF007FFFB47FFCEA90F0001C001FF0006A003F0AB00EFFAAD0F0000FE0";
    attribute INIT_25 of inst : label is "01F001AF007F0A3403FFEA90F0003FE0000F03FF003F004EF4C0D000FC005990";
    attribute INIT_26 of inst : label is "04F0001B01FFFEB00C3FE024F0000C2603F20FFF007F0B76A000D630FC006600";
    attribute INIT_27 of inst : label is "1F70005B01FF00300EFFEA50F0003FE001F8003F003FAD39FF8BF014F8008400";
    attribute INIT_28 of inst : label is "02F9FDBF2FD1003081C0EFE0FFD01C00000B03FF00FF0007F700FED0FC006E64";
    attribute INIT_29 of inst : label is "00DC003F003F0000BB00FC00FC000800002B03FF007F0000FDE0FE40FC000098";
    attribute INIT_2A of inst : label is "000F03FF003F0000F200D000FC002D30090BBF7FFC0000F08380F7F000FC0C00";
    attribute INIT_2B of inst : label is "00DC003F003F0000CE000FD0FF000000034A3FFF07FE003081C0FFFC00BF0C00";
    attribute INIT_2C of inst : label is "03F00FFF007F2936B700D400FC00660001FF01AA003F0A3447FCAA40FC001E80";
    attribute INIT_2D of inst : label is "019F0BFF01FF0226FC00C000FC0059900BFC07AA003FFFB40DF0A900FC001C00";
    attribute INIT_2E of inst : label is "02CC0FF000FF00002FC0FF00FC0003600B40BF7FFC0000F00380F7F000FE0C00";
    attribute INIT_2F of inst : label is "000F03FF003F0000F200D000FC002D300D00BF7FFC0000F00380FBC0FD000C00";
    attribute INIT_30 of inst : label is "090BBF7FFC3F00F0A380FD0040000C000B4B3F7F0FC000F08380F7F02F400C00";
    attribute INIT_31 of inst : label is "00FC003F003F02660FC03F00FD0069B903F000FC003F2D790FC03F00FD00995A";
    attribute INIT_32 of inst : label is "BC0AFC3F01F400B082BCF3FC00000CA000FC003F003F02C4FC00FC00FC00EE20";
    attribute INIT_33 of inst : label is "00BF07D3000302B0FFC0FB40FFC01C001E40017F0000283000E0FE7F03F40C00";
    attribute INIT_34 of inst : label is "3EAFFC3F07D000F0EBF8F0FC1F400C00F66F003F00052BF2D15CFD005000FF80";
    attribute INIT_35 of inst : label is "000F03FF34400003DB00E8000240300001AF003F000017F0BF40FFF700007CBD";
    attribute INIT_36 of inst : label is "03FF003F01900D80E400E8000290280001AF003F000003F0BF40FF4100007CFC";
    attribute INIT_37 of inst : label is "002B03FF01A00000FD40FFC900C0009801AF007F000003F0BF40FF0000007CFC";
    attribute INIT_38 of inst : label is "002B03FF091F0000FDE0FE40F158009803EF3FFF1FDF0090BFE0FE7FF6507C00";
    attribute INIT_39 of inst : label is "00803A2A0000000800002A280000880003003A2A0000000000002A2800000000";
    attribute INIT_3A of inst : label is "03AF003F00003F30BFC0FF0000007CBD18003A2A0000008000002A2800000000";
    attribute INIT_3B of inst : label is "1FAF003F00002CB0BFC0FF00000078FC01FC00FE01C00330FC00FC000240CC00";
    attribute INIT_3C of inst : label is "03AF003F00003F30FBC0FF0000000CBD00FE00FE01C000CCF800FC0002400000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000EC00FE01800000FC00FC0002403300";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "53FF8FFFFFFAF800CFFFF3FFFC0B50B40BFFFFFF3FFFCFFFFFFFFFFFFFFFFFFF";
    attribute INIT_01 of inst : label is "00000500FFFFFFFF07FFFFF0FFFEFF810037188CE180C000F000FF40FFFFFFFF";
    attribute INIT_02 of inst : label is "E000C240FFFF00AFFFFEFF8700378CCC00000000000000000540018000141E00";
    attribute INIT_03 of inst : label is "D000C000A00C0030FF14FFF4D200C00002CC0030FFC0FF00FFFFFFFFFFFFA000";
    attribute INIT_04 of inst : label is "C11CF7FC07E03110F00101FF5E0FFC0010048220000000C00540018000000000";
    attribute INIT_05 of inst : label is "00141E00FFFFFFFFFFFFBFADFFFF07ABBFFF6A8F1555FFFF000000004FFBDA97";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "55D0FE853FFF0FFF1FF8A027E008FFF03CBF12BF000005001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF01F50FD7";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "5242FFF70000F7FF8123F7F7F808FFDFFFFFFFFF2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "FFFFFFF8E0037FD2FFD7471FFFFFFD1FFFFC5FDF2FFFFFFF4782CDFF0200DDFD";
    attribute INIT_0D of inst : label is "FFF5FFFFFFFF2BFFFD2FFFFD1555CBFFFFFF4FE7FFFFBEABFFFFBFFFFFFFFFFD";
    attribute INIT_0E of inst : label is "FFFFFFFF5555FFFFFFE1A1FFE17FFFFFFFFFFFFFFFFFFFFFFFFFFFFF2FFFFFFF";
    attribute INIT_0F of inst : label is "5554FFFC5555FFFFFFFFFFFF5455FCFFFF3FFFCFFFCFFFF3FFFCFFFCFFFFFFFF";
    attribute INIT_10 of inst : label is "000000005554FFFF5555FFFFCFFF3FFFF3FFCFFFFCFFFCFFFFCFFF3FFFF3FFCF";
    attribute INIT_11 of inst : label is "00000000C000C000000300034000C00000010003AAC000C003AA030000000000";
    attribute INIT_12 of inst : label is "FC00FF00C000F0000003000F0000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFCFFFFFFC0FFF003FF0FFF003F00FF";
    attribute INIT_14 of inst : label is "C03F07FF0060FD800000000FFFFFFFFF00000000FFFFFFFF00000000FFFFFFFF";
    attribute INIT_15 of inst : label is "2FFE5FC0AB00F0000FFFFFFF000A00FF000000002BFDFFFFFFFFFCDC1FFFF801";
    attribute INIT_16 of inst : label is "1FFFFFFFFFFF163FFFFFFCC355449B3FFFFFFFFFCCFFE9FFFE14FFC3BCC0D097";
    attribute INIT_17 of inst : label is "00003FF5FFFF6BFFFFFD0290FFFFFFFFAAAA00000FFF3BFF00000000FFFFCCF3";
    attribute INIT_18 of inst : label is "BFC1017F2AA80000BFFDA22043FDFD403FDB5AFFFFFFF9FFAAAAFE6202FF0000";
    attribute INIT_19 of inst : label is "F000F000FFFF2631002F0000F000F000FE51F6FF0000007FFFFFEF6F6AFCFFFF";
    attribute INIT_1A of inst : label is "FAAAF000FFFF53FFFFFF347FD7F0FFFFAAA80000AAAA0000F000F00000000000";
    attribute INIT_1B of inst : label is "2D000FF43C003C00FAAAF0000FFE1F00FFFFFFFFA00000000FFF0FFF0FFF0FFF";
    attribute INIT_1C of inst : label is "CB4BF0F0FFFFFFFFFAAAF000AAAA000000000000AAAA000003FC03FCFFFFFFFF";
    attribute INIT_1D of inst : label is "42FC2D08FFFF0B40F0BD001500FFFFFFF03F800F7FFFBFFFFE815FFCFFFFFFFF";
    attribute INIT_1E of inst : label is "ABFFDDDDFFFFE80F2BFF57FF0000555FFFFFFFFF00FF07FFFFFFBFFFFFFFFEAA";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFD0FFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "00D00015000000001C0050000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0FFFFF1FFC0002F0F8C0D3F8003F070041800000000000008241000000000000";
    attribute INIT_22 of inst : label is "0D3F3FC500FC00D0F1C04FF0FF40070007F001FF003F3B001F00BFC0FC00A000";
    attribute INIT_23 of inst : label is "003F003F003F00633800FC00FC0090000652002F001FF430017DE000D0000CFE";
    attribute INIT_24 of inst : label is "0C42002F001F17F0015CE000D000BFFC0610002F001F2FF0017CE000D0000FFE";
    attribute INIT_25 of inst : label is "0242002F001F3FF0015CE000D0001FFC00BF007F003F000BFE40F800FC00FB80";
    attribute INIT_26 of inst : label is "019200BF00FF7FF007FFF540D0000C7F0BFF07FF003FB630FEDCF840FC000000";
    attribute INIT_27 of inst : label is "00D200BF00FF3FF0047DF000D0001DFE00FF003F003F43B0F19DF000FC002800";
    attribute INIT_28 of inst : label is "2FEFFFFFFD00003002C0FFF000000700002F01FF003F0000F9E0E000FC00EB40";
    attribute INIT_29 of inst : label is "00EC003F003F0020FF00FC00FC00370000FF01FF003F0000E930E000FC002934";
    attribute INIT_2A of inst : label is "00BF007F003F0002FD00F800FC00DE403FFFFF1FFC0002D0F870D3F803FC0700";
    attribute INIT_2B of inst : label is "00EE003F003F00206B80BFC0FC00A8000D3F3FC5005500D0FBF854FF007F0700";
    attribute INIT_2C of inst : label is "0BFF07FF003F7BB0E300F800FC000000035F002F001F3FFE0174E000F4000FF8";
    attribute INIT_2D of inst : label is "00EF0FFF003F02A0F000E000FC00E9000C54002F001F1FF804D0E000F4000FF0";
    attribute INIT_2E of inst : label is "0BF403FE003F009C3F00FC00FC000B300FFFFF1FFC0002F0F8C0D3F8003F0700";
    attribute INIT_2F of inst : label is "00BF007F003F0002FD00F800FC00DE403FFFFF1FFC0302D0D8C0FFC0F4000700";
    attribute INIT_30 of inst : label is "3FFFFD1FFC1502D0FEC0F400000007002FFF3F9F01F802F0F8E0D3F074000700";
    attribute INIT_31 of inst : label is "00FC003F003F05CF0FC0BF00FC004ED003F800FE003F07B12FC03F00FC001ED0";
    attribute INIT_32 of inst : label is "FF7F1FA500000A40F5FC405000000D7C00FE003F003F00EFFC00FC00FC00CA40";
    attribute INIT_33 of inst : label is "0BFF000F00000FFB94F0FFC05500FF0007EF001F00003FD0FEFEF4BD00002E00";
    attribute INIT_34 of inst : label is "FD3F1F9F00000B42F0FFDBD00000078001BF003F0000BFDBFAB4FC000000FFE0";
    attribute INIT_35 of inst : label is "02FF0B5C056A0003D00001D02C2EBA00002F001F00000251FA98F50400005FF4";
    attribute INIT_36 of inst : label is "00FF02D102BA0660C00081802CB89100002F001F00000251FBF9D50000005FF0";
    attribute INIT_37 of inst : label is "00FF0DFF02AE0000402657D029A8293400EF001F00000251FB40D40000005FF0";
    attribute INIT_38 of inst : label is "00FF01FF016A0000E930E800295029340F6F3F3F01460301FBF8FEFD58000F00";
    attribute INIT_39 of inst : label is "09003FFF000000800000FFFC0000000009003FFF000000880000FFFC00008800";
    attribute INIT_3A of inst : label is "007F001F00000751FF00F40000005FF409003FFF000010000000FFFC00000000";
    attribute INIT_3B of inst : label is "007F001F0000FE51FF00F40000005FF000FC0B462E3A03F0FC000DC02C2EFC00";
    attribute INIT_3C of inst : label is "007F001F00000752FF00F4000000C5F400FC0B46003A00FDFC000DC02C2E8000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000FC09412E3A0098FC0025C02C2E3F00";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFE0000000FFFFFFFF0850BD7F41FFFFEAFFFFFFFFFFFFAAAAFFFFFFFF";
    attribute INIT_01 of inst : label is "0F000A00FFFFFFFF00000007FFFEFF800150B03FF800F0000000A800FFFFFFFF";
    attribute INIT_02 of inst : label is "D500F080FFFFFEAFFFFEFEF0055008FF0000001A0000D0002430010001E0A000";
    attribute INIT_03 of inst : label is "C000F500003A05F0FFD4FFFFC000F500003A05F0FFFFFFFFFFFFFFFFFFFFFEAA";
    attribute INIT_04 of inst : label is "FFFDFFFF01FE400017FFFFFF0000003F0080021A0000D0C02430010000000000";
    attribute INIT_05 of inst : label is "01E0A00044C455DDFAFFFFFFC3AFFFFFF0DFFFFFFFFFFFFF00030003C001FFFF";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "00140000FFFF3FFFFFF896000000D57F1000C02A0F000A002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00054000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "FFF3FFFFF3FFFFFFFFFFFFFFFFCFFFFFCF33D75D01F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFF5FFD7F0FFF7FD7FFFDF5FFFD7FFEBFFFFFFFCFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFEFFFFEBAF7FFFFFFFFFFFFFFBFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_11 of inst : label is "0000000F00000000000000000000000000000000FF3F557FFCFFFD550000FFFF";
    attribute INIT_12 of inst : label is "FF00FFC0F000FC00000F003F000000030000C000F000F000000F000F0000F000";
    attribute INIT_13 of inst : label is "FFBBFFF7FFFFFF7FFEFFFFFFFFFFFFFFFFFFFFFFFFF0FFFC0FFF3FFF00FF03FF";
    attribute INIT_14 of inst : label is "7FFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFF0000000000000000FFDFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFF00BC01600FFFFFFFF01E078000003001FFFF5FFFF3FFFFFFF0007BDFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFEFF01FFFFFEFF0C00FF07FFFFFFFFFF03FF7FFFFFF0FFFDBE000300";
    attribute INIT_17 of inst : label is "CAFFC000FFFF02BF0000F500FFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "DB8000000000FFFFDBFF000002FF0000FFFD3F5B00050DBFFF6FFFFFF500FFFF";
    attribute INIT_19 of inst : label is "00001FFFFFFFFFFF00BF000F00007FFF6FFFFF6B007FFFFF5000FFF0FF5AFFFC";
    attribute INIT_1A of inst : label is "00000000FFFFFFFFFFFFFFFFFFFCAAAA000F555F00003FFD0000000000001550";
    attribute INIT_1B of inst : label is "F400FFF4C000C00000000000FE00C000FFFFBFFF0000E000FFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "F3C0F0BDFFFFFFFF0000000000000000000F000F00003FF83FC03FC0FFFFFFFF";
    attribute INIT_1D of inst : label is "F0BF0342FFACC2D0A00B55FF1FFFFFFFE00F001FFFFF2F2FA050FFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "CCA8FFFFFFAF015F00FFAAAA0000FFFFFFFFBFE800FFFFFFFFFF0BFFFFFF8000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC2FFF0FFFFFFFFFFFA";
    attribute INIT_20 of inst : label is "002A00FF00000000A000BC000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0BFFB374CC0000FFFF80777000CEFC0012FF041500000000FF84540400000000";
    attribute INIT_22 of inst : label is "03FD34FF0E18003FFF80FC7024F0FC000DC0031800EF2E00FC002FC083000000";
    attribute INIT_23 of inst : label is "00330033003B01FFE0008C00CC00998067BF007F0034933FFE33FFD07000FCA8";
    attribute INIT_24 of inst : label is "03BF01FF006085BFEBCCFFD0F000FC001AFF007F003F0ABFFED3FFD0F000FFE0";
    attribute INIT_25 of inst : label is "01FF01FF00600A3FFFCFFFD0F000F4E0000E034B003F004FFFC0D000AC00F990";
    attribute INIT_26 of inst : label is "04FF001D01A2D6BFFC31FFF4F000FC2603720CF9006F0BF6A000D7F0BC006600";
    attribute INIT_27 of inst : label is "1A7F005D01A2003FFED3FF50F000F06001980033003EAFF9D98BB014B8008400";
    attribute INIT_28 of inst : label is "027FC9B42491003FFFC07FE0AFD0FC000009035500EC00073F00ABD03C00EE64";
    attribute INIT_29 of inst : label is "00FC0037003B0000BF00DC00EC00080000290355007C000069E0AB403C0000B8";
    attribute INIT_2A of inst : label is "000F034B003A0000BE00D000BC002FF00BFFB360CC0000FFFF80F73000CCFC00";
    attribute INIT_2B of inst : label is "00FC0037003F0000FE000D90EB00000003FD34FF0616003FFFC0CF8C00B3FC00";
    attribute INIT_2C of inst : label is "03700C7900622BF6BF00D400FC00660001C201FF00330A3FFFCCFF40FC00FE80";
    attribute INIT_2D of inst : label is "01FF0B6C01FA02276C00C000FC00F9900B0F07FF003385BFFF30FD00FC00FC00";
    attribute INIT_2E of inst : label is "02FC0E7000FF00002CC0DB00EC0003E00BFFB36FCC0000FFFF80E77000CEFC00";
    attribute INIT_2F of inst : label is "000D0373003A00003E00D000BC002FF00FFFB367CC0000FFFF80FAC0CD00FC00";
    attribute INIT_30 of inst : label is "0BFFB36FCC3300FFFF806D004000FC000BFF33740CC000FFFF8077702640FC00";
    attribute INIT_31 of inst : label is "00DC0033003F02660CC03300FD006BB9033000CC003F2FF90CC03300FD009BFA";
    attribute INIT_32 of inst : label is "B7FDCC3F01A400BFFFCCF34C0000FCA000CC0033003B02EEDC00CC00EC00EE20";
    attribute INIT_33 of inst : label is "00B40693000302BFE3C07F40AFC0FC001FFF017F0000283FFF60C67303A4FC00";
    attribute INIT_34 of inst : label is "35FFCC34079000FFFE1870CC1A40FC00E6F40032000529EFFFBCFD005000DF80";
    attribute INIT_35 of inst : label is "000D032E3FFF0003BF00E800FF40F00001FF00360000127FFE40FFF70000FC99";
    attribute INIT_36 of inst : label is "039F003A01FF0F807400E800FFD0280001FF00360000033FFE40FF410000FCCC";
    attribute INIT_37 of inst : label is "0029035501FF00006940557DFFC000B801FF00760000033FFE40FF000000FCCC";
    attribute INIT_38 of inst : label is "002903550BFE000069E0AB40BFF800B8037F36F61CDF00BFFC607E73F650FC00";
    attribute INIT_39 of inst : label is "00913BBB000000089100BBB80000880003993BBB000000001980BBB800000000";
    attribute INIT_3A of inst : label is "03FF00360000333FFEC0FF000000FC9919893BBB000008809800BBB800000000";
    attribute INIT_3B of inst : label is "1BFF0036000024BFFEC0FF000000F8CC018C00EE01FF03F0CC00EC00FF40FC00";
    attribute INIT_3C of inst : label is "03FF003F0000333FFFC0FF000000FC9900CF00EE01FF00FC9800EC00FF400000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000FC00FE01FF0000CC00EC00FF403F00";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFE000000FFFFFFFFFC0B50B40BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_01 of inst : label is "00000500FFFFFFFFE0000001FFFFFFF400001EBFA780F0000000D000FFFFFFFF";
    attribute INIT_02 of inst : label is "A000F2D0FFFFFFFFFFFFFFF80000BEFF00000000000000000540018000141E00";
    attribute INIT_03 of inst : label is "F000C000203F0030FFC2FFFFF000C00000FF0030FFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_04 of inst : label is "1FFFFFFFA0170680007FFFFFA0E0000F10048220000000000540018000000000";
    attribute INIT_05 of inst : label is "00141E00FFFFC4C4FFEFF5FFFFFFFF5F7FFFFFFFFFFFFFFF000300030000F57F";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "80020000FFFFBFFF7FFFFF8005400003C0004940000005001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAFC0020000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "FE80FFF70003F7FF9BA9F7F7F802FFDFFFFFCF342ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "FFFFFFF8E0037AD2EBFFFFFFFEBFC3FEAF0CEBEF2FFFD7FFDF12FDFFFF01FFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFFED75FFFFFF0FFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_11 of inst : label is "0000000F00000000000000000000000000000000553FFF3FFC55FCFF0000FFFF";
    attribute INIT_12 of inst : label is "FF00FFC0F000FC00000F003F000000030000C000F000F000000F000F0000F000";
    attribute INIT_13 of inst : label is "EFEFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFF0FFFC0FFF3FFF00FF03FF";
    attribute INIT_14 of inst : label is "1FFFFFFF2FFFFFFFFDFF2FFFFFFFFFFFFFFFFFFF0000000000000000FBFFFFFF";
    attribute INIT_15 of inst : label is "D001FFFCFFE00F007FFFFFFF00FF0F0000020007D400FFFFFFFF7FFFC000011F";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFF60FFFFFFFF2CAABF00FFFFFFFFFF03FF07FFFFABFFF4FF080460";
    attribute INIT_17 of inst : label is "FFFFC00AFFFFBFFF00000000FFFFFFFF000000007FFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "BFF0A00000000000BFFDF6FF0FFD000A3FDB5AFF000001FF0000FFFFC000FFF5";
    attribute INIT_19 of inst : label is "00000000FFFFFFFFABFF000F00000000FFFFF6FF000F07FF0000FF40FAFCFFFF";
    attribute INIT_1A of inst : label is "00000000FFFFFFFFFFFFFFFFD7F0FFFF0007000F00000000000000002AAA0000";
    attribute INIT_1B of inst : label is "D000FF40C000C00000000000FFE0E000FFFFFFFF00000000FFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "CB4BF0F05555FFFF0000000000000000000F000F000000003FC03FC0FFFFFFFF";
    attribute INIT_1D of inst : label is "42FC2D08FFFF0B40F0BD001500FFFFFFF03F800F7FFFBFFFFE815FFCFFFFFFFF";
    attribute INIT_1E of inst : label is "ABFFCCDCFFFFE80F2BFF57FF0000555FFFFFFFFF00FF07FFFFFFBFFFFFFFFEAA";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFD0FFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "00FF001500000000FC0050000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0CB4CB1FDC0002FF7FC0D3180033FF0041FF0000000000007F41000000000000";
    attribute INIT_22 of inst : label is "0FFF31C500EC00FFFFC04D30C340FF0007700187003F3F001F0090C0FC00A000";
    attribute INIT_23 of inst : label is "00330033003F007FF800CC00FC00900007FF0024001F643FFFED6000D000FCCE";
    attribute INIT_24 of inst : label is "0FFF0024001F163FFFEC6000D000D55C07FF002E001F26FFFFACE000D000FF9E";
    attribute INIT_25 of inst : label is "02FF0024001F387FFFEC6000D000FE1C00BD0061003F000B2F407800FC007F80";
    attribute INIT_26 of inst : label is "01FF009200EB62BFFFD3F540D000FC630B34073C003FBFF09EFC3840FC000000";
    attribute INIT_27 of inst : label is "00FF009200EB357FFFADF000D000FD8600CF0038003F537031FD7000FC002800";
    attribute INIT_28 of inst : label is "24BFCF4AC900003FFFC0D3F00000FF00002601E1003F0000FFE0E000FC00DF40";
    attribute INIT_29 of inst : label is "00FC0033003F0020DB00CC00FC003F0000EB01E1003F0000EBF0E000FC002BF4";
    attribute INIT_2A of inst : label is "00BD0061003F00026D00F800FC00FF4034B4CB1FDC0002FF7FF0D318032CFF00";
    attribute INIT_2B of inst : label is "00FE0033003F00207F80B2C0FC00A8000FFF31C5005500FFDE3854E7006BFF00";
    attribute INIT_2C of inst : label is "0B3D0707003F7FF05F009800FC00000003EB0026001F3857FFE4E000F400FF18";
    attribute INIT_2D of inst : label is "00FC0E70003F02A0B000E000FC00DD000FFF0026001F1E3FFFD0E000F400FD70";
    attribute INIT_2E of inst : label is "0B34039E003F00BC3300CC00FC000BF00CBFCB1FDC0002FFFFC0D3180033FF00";
    attribute INIT_2F of inst : label is "00B40071003F0002ED00F800FC00FF4034B7CB1FEC0302FFDFC0F6C0B400FF00";
    attribute INIT_30 of inst : label is "34B6C91CEC1502FFD3C0F4000000FF002CB4339F019802FF7FE0D3306400FF00";
    attribute INIT_31 of inst : label is "00CC0033003F05FF0CC0B300FC004FD0031800E6003F07F124C03300FC001FD0";
    attribute INIT_32 of inst : label is "CB7F19A500000AFFF5CC40500000FFCC00CE0033003F00FFCC00CC00FC00FF40";
    attribute INIT_33 of inst : label is "0B6B000D00000FBFFFF087C055005F00067E001F000031FFDF86E4990000FE00";
    attribute INIT_34 of inst : label is "C934199F00000BFF70E3D9900000FF8001FD003A00009BFFFFF4FC00000029E0";
    attribute INIT_35 of inst : label is "02DC0BFF057F0003D000FFD0FC267A000024001F000002FF7A98F5040000FF64";
    attribute INIT_36 of inst : label is "00E602FF023F07E0C000FF80FC98BD000024001F000002FF7BF9D5000000FF30";
    attribute INIT_37 of inst : label is "00EB0FEB022F0000402EFFD0FD882BF400E4001F000002FF7B40D4000000FF30";
    attribute INIT_38 of inst : label is "00EB01E1017F0000EBF0E800FD502BF40C64333F014603FF7B98FE6D5800FF00";
    attribute INIT_39 of inst : label is "09993AAA000000991980AAAC0000190009913AAA000000889180AAAC00008800";
    attribute INIT_3A of inst : label is "0074001F000006FF7F00F4000000FF6409913AAA000019988980AAAC00000000";
    attribute INIT_3B of inst : label is "0074001F0000CEFF7F00F4000000FF3000CC0BFF263F0330CC00FFC0FC26CC00";
    attribute INIT_3C of inst : label is "007F001F000006FFFF00F4000000FF6400CC0BFF003F00CFCC00FFC0FC268000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000CC0BFF263F00B8CC00FFC0FC263300";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
