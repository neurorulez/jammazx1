library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bubbles_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bubbles_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"34",X"07",X"1A",X"50",X"DE",X"0C",X"EC",X"C4",X"26",X"03",X"BD",X"01",X"C1",X"DD",X"0C",X"35",
		X"87",X"B6",X"BF",X"FF",X"8A",X"01",X"B7",X"C9",X"00",X"7E",X"01",X"E7",X"B6",X"BF",X"FF",X"B7",
		X"C9",X"00",X"10",X"DE",X"20",X"3B",X"1A",X"50",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",
		X"12",X"12",X"12",X"7E",X"0C",X"7F",X"34",X"10",X"8B",X"15",X"46",X"1F",X"01",X"B6",X"BF",X"FF",
		X"84",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"86",X"0F",X"24",X"02",X"86",X"F0",X"A4",X"84",
		X"A7",X"84",X"86",X"01",X"BA",X"BF",X"FF",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"90",X"BD",
		X"15",X"B9",X"84",X"01",X"8E",X"CD",X"00",X"30",X"8B",X"BD",X"15",X"BD",X"C4",X"F0",X"34",X"04",
		X"1A",X"50",X"E6",X"84",X"C4",X"0F",X"EA",X"E4",X"E7",X"84",X"E6",X"84",X"1C",X"EF",X"E8",X"E0",
		X"C4",X"F0",X"27",X"07",X"BD",X"00",X"AD",X"2F",X"FF",X"D0",X"8C",X"39",X"BD",X"15",X"BD",X"86",
		X"C8",X"BD",X"01",X"48",X"5A",X"26",X"F8",X"6E",X"9F",X"98",X"0A",X"0A",X"3F",X"0A",X"3F",X"0D",
		X"A5",X"34",X"56",X"B6",X"BF",X"FF",X"84",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"4F",X"A6",
		X"C0",X"49",X"89",X"00",X"49",X"89",X"00",X"49",X"89",X"00",X"49",X"89",X"00",X"A7",X"80",X"5A",
		X"26",X"EC",X"35",X"56",X"33",X"C9",X"01",X"00",X"30",X"89",X"FF",X"00",X"4A",X"26",X"D2",X"86",
		X"01",X"BA",X"BF",X"FF",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"39",X"86",X"03",X"BD",X"00",X"5C",
		X"CE",X"00",X"89",X"8E",X"D0",X"EE",X"4F",X"5F",X"35",X"20",X"34",X"56",X"6E",X"A4",X"80",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"7E",X"D3",X"C7",X"7E",X"D4",X"40",X"7E",X"D2",X"54",X"7E",X"D2",X"DC",X"7E",X"D6",X"54",X"7E",
		X"D4",X"9C",X"7E",X"D4",X"7C",X"7E",X"D4",X"4E",X"7E",X"D7",X"B6",X"7E",X"D7",X"B0",X"7E",X"D7",
		X"5C",X"7E",X"D7",X"81",X"7E",X"D7",X"92",X"7E",X"D7",X"90",X"7E",X"D7",X"9A",X"7E",X"D7",X"A8",
		X"7E",X"D7",X"A6",X"7E",X"D7",X"EF",X"7E",X"D9",X"B4",X"7E",X"D9",X"D8",X"7E",X"D9",X"D2",X"7E",
		X"D9",X"CC",X"7E",X"DA",X"3D",X"7E",X"DA",X"53",X"7E",X"DA",X"68",X"7E",X"DA",X"D2",X"7E",X"DB",
		X"ED",X"7E",X"DD",X"7D",X"34",X"02",X"A6",X"80",X"1E",X"12",X"BD",X"D7",X"9A",X"1E",X"12",X"5A",
		X"26",X"F4",X"35",X"82",X"8E",X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",
		X"36",X"8E",X"D2",X"96",X"10",X"8E",X"CC",X"00",X"C6",X"12",X"8D",X"D8",X"35",X"B6",X"34",X"36",
		X"8E",X"D2",X"A8",X"10",X"8E",X"CC",X"24",X"C6",X"34",X"8D",X"C9",X"BD",X"D3",X"9E",X"8E",X"CC",
		X"8E",X"BD",X"D7",X"9A",X"35",X"B6",X"25",X"03",X"01",X"03",X"01",X"04",X"01",X"01",X"00",X"00",
		X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"1A",
		X"1C",X"0F",X"1D",X"0F",X"18",X"1E",X"0F",X"0E",X"0A",X"0C",X"23",X"32",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",
		X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"2E",X"25",X"29",X"BD",X"D3",X"85",X"BD",
		X"D7",X"5C",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1B",X"84",X"0F",X"27",X"11",
		X"7F",X"CC",X"1B",X"BD",X"D3",X"85",X"BD",X"D7",X"5C",X"BD",X"D4",X"29",X"86",X"40",X"BD",X"F0",
		X"09",X"B6",X"CC",X"1D",X"84",X"0F",X"27",X"0D",X"7F",X"CC",X"1D",X"8D",X"78",X"BD",X"D2",X"0F",
		X"86",X"40",X"BD",X"F0",X"09",X"B6",X"CC",X"21",X"84",X"0F",X"27",X"24",X"7F",X"CC",X"21",X"8D",
		X"64",X"BD",X"D7",X"5C",X"86",X"0A",X"BD",X"7B",X"12",X"86",X"2B",X"BD",X"7B",X"12",X"BD",X"DC",
		X"77",X"B6",X"00",X"20",X"BD",X"F0",X"09",X"BD",X"D3",X"9E",X"8E",X"CC",X"8E",X"BD",X"D7",X"9A",
		X"B6",X"CC",X"23",X"84",X"0F",X"27",X"18",X"7F",X"CC",X"23",X"8D",X"39",X"BD",X"D7",X"5C",X"86",
		X"10",X"BD",X"7B",X"12",X"86",X"2B",X"BD",X"7B",X"12",X"BD",X"DA",X"7F",X"BD",X"D6",X"1B",X"B6",
		X"CC",X"1F",X"84",X"0F",X"27",X"0A",X"7F",X"CC",X"1F",X"8D",X"1A",X"8D",X"07",X"7E",X"F0",X"06",
		X"8D",X"02",X"20",X"53",X"B6",X"CC",X"19",X"84",X"0F",X"27",X"09",X"7C",X"CC",X"8C",X"7C",X"CC",
		X"8C",X"7F",X"CC",X"19",X"39",X"34",X"12",X"8D",X"08",X"8E",X"CC",X"8C",X"BD",X"D7",X"9A",X"35",
		X"92",X"34",X"34",X"8E",X"CC",X"00",X"10",X"8E",X"CC",X"24",X"8D",X"09",X"35",X"B4",X"8E",X"CC",
		X"24",X"10",X"8E",X"CC",X"8C",X"10",X"BF",X"BF",X"06",X"4F",X"E6",X"80",X"C4",X"0F",X"34",X"04",
		X"AB",X"E0",X"BC",X"BF",X"06",X"26",X"F3",X"8B",X"37",X"39",X"8D",X"D5",X"34",X"02",X"8E",X"CC",
		X"8C",X"BD",X"D7",X"81",X"A1",X"E0",X"39",X"8D",X"70",X"8D",X"EF",X"27",X"3D",X"86",X"39",X"B7",
		X"CB",X"FF",X"BD",X"D2",X"6F",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"A9",X"86",X"39",X"B7",X"CB",
		X"FF",X"BD",X"D7",X"5C",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"28",X"BD",X"D2",X"12",X"BD",X"D2",
		X"0C",X"8D",X"C7",X"27",X"1A",X"86",X"0B",X"BD",X"7B",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"B6",
		X"C8",X"0C",X"85",X"02",X"27",X"F4",X"6E",X"9F",X"EF",X"FE",X"BD",X"D2",X"0C",X"20",X"F7",X"86",
		X"0C",X"20",X"E4",X"8E",X"CD",X"02",X"C6",X"04",X"A6",X"80",X"84",X"0F",X"81",X"09",X"23",X"03",
		X"5A",X"27",X"06",X"8C",X"CD",X"3E",X"26",X"F0",X"39",X"86",X"0D",X"BD",X"7B",X"12",X"8E",X"CD",
		X"02",X"6F",X"80",X"8C",X"CD",X"3E",X"26",X"F9",X"39",X"8D",X"05",X"27",X"FB",X"7E",X"D2",X"7E",
		X"BD",X"D3",X"9E",X"34",X"02",X"8E",X"CC",X"8E",X"BD",X"D7",X"81",X"A1",X"E0",X"39",X"86",X"18",
		X"B7",X"BF",X"13",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"08",X"BD",X"F0",X"09",X"B6",X"C8",X"0C",
		X"85",X"08",X"27",X"17",X"7A",X"BF",X"13",X"26",X"EF",X"10",X"8E",X"CD",X"3E",X"8E",X"D4",X"D5",
		X"C6",X"17",X"BD",X"D2",X"06",X"BD",X"D6",X"1B",X"7F",X"C8",X"0E",X"39",X"10",X"8E",X"CD",X"74",
		X"C6",X"08",X"BD",X"D6",X"42",X"A8",X"26",X"84",X"0F",X"27",X"03",X"5A",X"27",X"0E",X"86",X"39",
		X"B7",X"CB",X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"E7",X"39",X"86",X"39",X"B7",X"CB",
		X"FF",X"8E",X"D4",X"D5",X"10",X"8E",X"CD",X"3E",X"C6",X"7D",X"BD",X"D2",X"06",X"8E",X"D5",X"52",
		X"10",X"8E",X"CE",X"38",X"C6",X"B6",X"BD",X"D2",X"06",X"BD",X"D6",X"1B",X"10",X"8E",X"CD",X"74",
		X"BD",X"D6",X"3A",X"86",X"39",X"B7",X"CB",X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"F0",
		X"86",X"0E",X"7E",X"7B",X"12",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"1D",X"0A",X"21",X"13",X"16",
		X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0A",X"0A",X"0A",X"21",X"13",X"16",X"00",X"10",X"91",X"02",
		X"17",X"1C",X"1D",X"00",X"04",X"84",X"93",X"14",X"14",X"15",X"00",X"04",X"71",X"13",X"1E",X"13",
		X"17",X"00",X"04",X"61",X"75",X"0B",X"18",X"11",X"00",X"04",X"52",X"22",X"0C",X"10",X"0E",X"00",
		X"04",X"42",X"10",X"15",X"10",X"16",X"00",X"04",X"32",X"17",X"15",X"0F",X"18",X"00",X"04",X"29",
		X"99",X"1C",X"19",X"18",X"00",X"04",X"10",X"11",X"1A",X"10",X"24",X"00",X"04",X"05",X"23",X"14",
		X"0F",X"18",X"00",X"03",X"99",X"09",X"0D",X"1C",X"0C",X"00",X"03",X"80",X"01",X"1A",X"20",X"0B",
		X"00",X"03",X"72",X"10",X"11",X"21",X"21",X"00",X"03",X"61",X"91",X"14",X"0B",X"18",X"00",X"03",
		X"51",X"01",X"14",X"19",X"0F",X"00",X"03",X"42",X"11",X"1E",X"13",X"17",X"00",X"03",X"35",X"67",
		X"0F",X"0A",X"0B",X"00",X"03",X"28",X"90",X"14",X"13",X"17",X"00",X"03",X"19",X"01",X"21",X"0F",
		X"1D",X"00",X"03",X"01",X"57",X"16",X"0F",X"19",X"00",X"02",X"92",X"30",X"0C",X"1F",X"24",X"00",
		X"02",X"87",X"77",X"14",X"14",X"15",X"00",X"02",X"79",X"87",X"1D",X"0B",X"15",X"00",X"02",X"69",
		X"59",X"0E",X"0F",X"0C",X"00",X"02",X"58",X"88",X"18",X"0A",X"10",X"00",X"02",X"46",X"75",X"14",
		X"14",X"15",X"00",X"02",X"33",X"10",X"1E",X"13",X"17",X"00",X"02",X"29",X"17",X"0B",X"18",X"11",
		X"00",X"02",X"25",X"52",X"0C",X"10",X"0E",X"00",X"02",X"05",X"22",X"1C",X"19",X"18",X"00",X"01",
		X"76",X"35",X"17",X"1C",X"1D",X"00",X"01",X"65",X"35",X"15",X"0B",X"23",X"00",X"01",X"55",X"05",
		X"14",X"11",X"16",X"00",X"01",X"43",X"15",X"1C",X"0B",X"17",X"00",X"01",X"31",X"09",X"12",X"0F",
		X"0D",X"00",X"01",X"20",X"10",X"15",X"20",X"0E",X"00",X"01",X"17",X"55",X"0F",X"14",X"1D",X"00",
		X"01",X"05",X"02",X"20",X"0B",X"22",X"00",X"00",X"94",X"05",X"0E",X"1C",X"14",X"00",X"00",X"83",
		X"11",X"14",X"0B",X"23",X"00",X"00",X"70",X"01",X"0A",X"0A",X"0A",X"00",X"00",X"40",X"00",X"34",
		X"34",X"8E",X"D6",X"08",X"C6",X"07",X"BD",X"D2",X"06",X"35",X"B4",X"34",X"02",X"8D",X"05",X"B7",
		X"CD",X"6C",X"35",X"82",X"34",X"10",X"8E",X"CD",X"3E",X"4F",X"AB",X"84",X"30",X"01",X"8C",X"CD",
		X"6C",X"27",X"F9",X"8C",X"CD",X"74",X"26",X"F2",X"35",X"90",X"34",X"02",X"8D",X"04",X"A7",X"26",
		X"35",X"82",X"34",X"24",X"C6",X"0E",X"4F",X"C1",X"08",X"27",X"02",X"AB",X"A4",X"31",X"21",X"5A",
		X"26",X"F5",X"35",X"A4",X"86",X"AA",X"B7",X"CF",X"FF",X"B1",X"CF",X"FF",X"27",X"03",X"7E",X"90",
		X"00",X"86",X"32",X"34",X"02",X"10",X"8E",X"CD",X"74",X"8D",X"D7",X"A8",X"26",X"84",X"0F",X"27",
		X"0F",X"BD",X"D7",X"31",X"7F",X"CD",X"00",X"7F",X"CD",X"01",X"6A",X"E4",X"27",X"12",X"20",X"E9",
		X"86",X"03",X"C6",X"04",X"8D",X"65",X"25",X"E9",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"D9",
		X"35",X"02",X"8E",X"D5",X"9F",X"10",X"8E",X"CF",X"A4",X"C6",X"2A",X"BD",X"D2",X"06",X"8D",X"84",
		X"B8",X"CD",X"6C",X"84",X"0F",X"27",X"02",X"8D",X"0F",X"10",X"8E",X"CD",X"3E",X"86",X"17",X"C6",
		X"04",X"8D",X"38",X"24",X"02",X"8D",X"01",X"39",X"8E",X"CD",X"3E",X"86",X"0A",X"BD",X"D7",X"9A",
		X"8C",X"CD",X"66",X"25",X"F8",X"8E",X"CD",X"74",X"10",X"8E",X"CD",X"3E",X"86",X"06",X"BD",X"D7",
		X"51",X"10",X"8E",X"CD",X"66",X"8D",X"7A",X"8E",X"CD",X"7A",X"10",X"8E",X"CD",X"6C",X"86",X"08",
		X"8D",X"6F",X"BD",X"D6",X"1B",X"10",X"8E",X"CD",X"74",X"20",X"46",X"34",X"16",X"C6",X"39",X"F7",
		X"CB",X"FF",X"1F",X"21",X"BD",X"D7",X"92",X"C1",X"0A",X"25",X"32",X"C1",X"24",X"22",X"2E",X"4A",
		X"26",X"F2",X"A6",X"61",X"BD",X"D7",X"92",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",X"D7",
		X"92",X"34",X"04",X"C4",X"0F",X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",X"22",
		X"0C",X"4A",X"26",X"EA",X"1C",X"FE",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"96",X"1A",X"01",X"20",
		X"F5",X"34",X"36",X"30",X"2E",X"8C",X"CF",X"A4",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",X"2E",
		X"30",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"EC",X"BD",X"D6",X"0F",X"BD",X"D6",X"3A",X"35",
		X"B6",X"34",X"36",X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"34",X"76",X"CC",X"00",
		X"00",X"1F",X"01",X"1F",X"02",X"CE",X"98",X"00",X"86",X"39",X"36",X"34",X"36",X"34",X"36",X"34",
		X"36",X"34",X"36",X"34",X"36",X"34",X"B7",X"CB",X"FF",X"11",X"83",X"A0",X"00",X"25",X"EB",X"35",
		X"F6",X"A6",X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",
		X"8D",X"EF",X"34",X"02",X"8D",X"EB",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",
		X"44",X"44",X"A7",X"81",X"35",X"82",X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",
		X"34",X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"0F",X"58",X"34",X"04",X"58",X"EB",X"E0",
		X"8E",X"CC",X"FC",X"3A",X"8D",X"CC",X"34",X"04",X"8D",X"C8",X"34",X"04",X"8D",X"C4",X"34",X"04",
		X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",X"89",X"00",
		X"19",X"30",X"1A",X"8D",X"B5",X"35",X"04",X"35",X"02",X"8D",X"BB",X"35",X"02",X"35",X"96",X"12",
		X"12",X"12",X"86",X"0F",X"BD",X"7B",X"12",X"7F",X"BF",X"06",X"8E",X"11",X"74",X"86",X"F1",X"C6",
		X"AA",X"10",X"8E",X"CD",X"3E",X"10",X"BC",X"BF",X"1B",X"26",X"04",X"C6",X"AA",X"20",X"08",X"10",
		X"BC",X"BF",X"1F",X"26",X"02",X"C6",X"AA",X"BD",X"7B",X"06",X"86",X"2B",X"BD",X"7B",X"00",X"30",
		X"89",X"03",X"00",X"86",X"15",X"B7",X"BF",X"0D",X"7A",X"BF",X"0D",X"27",X"1E",X"1E",X"12",X"BD",
		X"D2",X"21",X"81",X"0A",X"2E",X"0B",X"7D",X"BF",X"06",X"26",X"09",X"10",X"BF",X"BF",X"06",X"20",
		X"03",X"7F",X"BF",X"06",X"1E",X"12",X"BD",X"7B",X"00",X"20",X"DD",X"7D",X"BF",X"06",X"27",X"03",
		X"BE",X"BF",X"06",X"86",X"04",X"B7",X"BF",X"0D",X"10",X"8E",X"CD",X"6C",X"1E",X"12",X"BD",X"D2",
		X"21",X"1E",X"12",X"8A",X"F0",X"85",X"0F",X"26",X"02",X"8A",X"0F",X"BD",X"7B",X"06",X"7A",X"BF",
		X"0D",X"1E",X"12",X"BD",X"D2",X"21",X"1E",X"12",X"BD",X"7B",X"06",X"7A",X"BF",X"0D",X"26",X"F1",
		X"8E",X"13",X"80",X"C6",X"33",X"CE",X"7B",X"0F",X"FF",X"BF",X"10",X"CE",X"7B",X"09",X"86",X"0D",
		X"B7",X"BF",X"0D",X"86",X"02",X"B7",X"BF",X"13",X"86",X"07",X"B7",X"BF",X"12",X"86",X"0E",X"B7",
		X"BF",X"18",X"8D",X"55",X"8E",X"3D",X"80",X"86",X"0D",X"B7",X"BF",X"0D",X"86",X"15",X"B7",X"BF",
		X"13",X"8D",X"46",X"8E",X"67",X"80",X"86",X"0D",X"B7",X"BF",X"0D",X"86",X"28",X"B7",X"BF",X"13",
		X"8D",X"37",X"8E",X"13",X"41",X"10",X"8E",X"CF",X"A4",X"C6",X"11",X"CE",X"7B",X"06",X"FF",X"BF",
		X"10",X"CE",X"7B",X"00",X"86",X"03",X"B7",X"BF",X"0D",X"86",X"01",X"B7",X"BF",X"13",X"86",X"0A",
		X"B7",X"BF",X"12",X"86",X"15",X"B7",X"BF",X"18",X"8D",X"0F",X"8E",X"53",X"41",X"86",X"03",X"B7",
		X"BF",X"0D",X"86",X"04",X"B7",X"BF",X"13",X"20",X"00",X"BF",X"BF",X"0A",X"34",X"04",X"C6",X"03",
		X"F7",X"BF",X"1A",X"5C",X"F7",X"BF",X"17",X"E6",X"E4",X"10",X"BC",X"BF",X"1B",X"27",X"06",X"10",
		X"BC",X"BF",X"1D",X"26",X"02",X"C6",X"AA",X"10",X"BC",X"BF",X"1F",X"27",X"06",X"10",X"BC",X"BF",
		X"21",X"26",X"02",X"C6",X"77",X"B6",X"BF",X"13",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"AD",X"9F",
		X"BF",X"10",X"86",X"2B",X"AD",X"C4",X"86",X"0A",X"AD",X"C4",X"1E",X"12",X"BD",X"D2",X"21",X"1E",
		X"12",X"AD",X"C4",X"7A",X"BF",X"1A",X"26",X"F2",X"BF",X"BF",X"06",X"BE",X"BF",X"0A",X"1E",X"01",
		X"F6",X"BF",X"07",X"BB",X"BF",X"18",X"1E",X"01",X"7F",X"BF",X"0E",X"1E",X"12",X"BD",X"D2",X"21",
		X"1E",X"12",X"7D",X"BF",X"0E",X"26",X"1B",X"34",X"02",X"86",X"04",X"B1",X"BF",X"17",X"26",X"04",
		X"35",X"02",X"20",X"06",X"35",X"02",X"85",X"F0",X"26",X"08",X"8A",X"F0",X"85",X"0F",X"26",X"02",
		X"8A",X"0F",X"B7",X"BF",X"0E",X"73",X"BF",X"0E",X"AD",X"9F",X"BF",X"10",X"7A",X"BF",X"17",X"26",
		X"CA",X"BF",X"BF",X"06",X"BE",X"BF",X"0A",X"1E",X"01",X"F6",X"BF",X"07",X"FB",X"BF",X"12",X"1E",
		X"01",X"B6",X"BF",X"13",X"8B",X"01",X"19",X"B7",X"BF",X"13",X"7A",X"BF",X"0D",X"35",X"04",X"10",
		X"26",X"FF",X"49",X"39",X"34",X"12",X"BB",X"BF",X"23",X"19",X"24",X"02",X"86",X"99",X"B7",X"BF",
		X"23",X"8E",X"CD",X"00",X"BD",X"D7",X"9A",X"35",X"12",X"7E",X"00",X"18",X"34",X"16",X"C6",X"03",
		X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",X"C6",X"01",X"BD",X"D7",X"B0",X"58",
		X"8E",X"CC",X"06",X"3A",X"BD",X"D7",X"92",X"8D",X"6A",X"B6",X"BF",X"25",X"34",X"04",X"AB",X"E4",
		X"B7",X"BF",X"25",X"B6",X"BF",X"24",X"AB",X"E0",X"B7",X"BF",X"24",X"8E",X"CC",X"12",X"BD",X"D7",
		X"92",X"8D",X"50",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",X"96",X"8E",X"CC",X"0E",X"BD",X"D7",
		X"92",X"8D",X"40",X"8D",X"28",X"34",X"02",X"F7",X"BF",X"24",X"8E",X"CC",X"10",X"BD",X"D7",X"92",
		X"B6",X"BF",X"25",X"8D",X"2E",X"8D",X"16",X"4D",X"27",X"06",X"7F",X"BF",X"24",X"7F",X"BF",X"25",
		X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"D7",X"B6",X"BD",X"D9",X"B4",X"35",X"96",X"34",X"04",X"5D",
		X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",X"01",X"19",X"E0",X"E4",X"24",X"F9",
		X"EB",X"E0",X"39",X"34",X"02",X"4F",X"C1",X"10",X"25",X"06",X"8B",X"0A",X"C0",X"10",X"20",X"F6",
		X"34",X"04",X"AB",X"E0",X"1F",X"89",X"35",X"82",X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",
		X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"10",
		X"8E",X"B0",X"00",X"8E",X"CC",X"16",X"BD",X"D7",X"92",X"8D",X"C8",X"E7",X"A4",X"C6",X"14",X"86",
		X"0A",X"30",X"2F",X"A7",X"80",X"5A",X"26",X"FB",X"8E",X"DA",X"D2",X"AF",X"26",X"C6",X"02",X"E7",
		X"2E",X"8E",X"20",X"80",X"AF",X"28",X"C6",X"0A",X"E7",X"22",X"6F",X"21",X"86",X"25",X"A7",X"23",
		X"86",X"3C",X"A7",X"24",X"86",X"77",X"A7",X"25",X"AD",X"B8",X"06",X"25",X"05",X"BD",X"DB",X"E4",
		X"20",X"F6",X"C6",X"14",X"8E",X"CD",X"3E",X"31",X"2F",X"A6",X"A0",X"BD",X"D7",X"9A",X"5A",X"26",
		X"F8",X"39",X"4F",X"E6",X"21",X"27",X"11",X"34",X"04",X"CB",X"0E",X"E6",X"A5",X"58",X"BE",X"7B",
		X"18",X"AB",X"95",X"35",X"04",X"5A",X"26",X"EF",X"AE",X"28",X"30",X"8B",X"AF",X"2A",X"C6",X"0F",
		X"EB",X"21",X"A6",X"A5",X"BD",X"DB",X"9A",X"E6",X"24",X"F7",X"C8",X"07",X"F6",X"C8",X"04",X"C4",
		X"0F",X"26",X"08",X"E6",X"2E",X"27",X"78",X"6A",X"2E",X"20",X"74",X"8E",X"DB",X"13",X"AF",X"26",
		X"1C",X"FE",X"39",X"34",X"04",X"E6",X"24",X"F7",X"C8",X"07",X"F6",X"C8",X"04",X"C4",X"0F",X"E1",
		X"E4",X"35",X"04",X"26",X"5A",X"C5",X"02",X"27",X"0D",X"8D",X"67",X"A1",X"22",X"26",X"04",X"A6",
		X"23",X"20",X"12",X"4A",X"20",X"0F",X"C5",X"01",X"27",X"13",X"8D",X"56",X"A1",X"23",X"26",X"04",
		X"A6",X"22",X"20",X"01",X"4C",X"E6",X"2E",X"27",X"36",X"6A",X"2E",X"20",X"32",X"6D",X"2E",X"26",
		X"F8",X"C5",X"04",X"26",X"08",X"C6",X"02",X"E7",X"2E",X"81",X"25",X"26",X"12",X"C6",X"02",X"E7",
		X"2E",X"6D",X"21",X"27",X"1A",X"8D",X"2B",X"8D",X"2C",X"6C",X"A4",X"6A",X"21",X"20",X"12",X"8D",
		X"24",X"6C",X"21",X"6A",X"A4",X"26",X"08",X"1A",X"01",X"8E",X"DA",X"D2",X"AF",X"26",X"39",X"8D",
		X"04",X"1C",X"FE",X"20",X"F4",X"C6",X"0F",X"EB",X"21",X"A7",X"A5",X"E6",X"25",X"AE",X"2A",X"7E",
		X"7B",X"00",X"5F",X"20",X"F8",X"34",X"27",X"5F",X"20",X"04",X"34",X"27",X"E6",X"25",X"1A",X"F0",
		X"F7",X"CA",X"01",X"CC",X"DB",X"DC",X"FD",X"CA",X"02",X"AE",X"2A",X"30",X"08",X"CC",X"00",X"06",
		X"8D",X"19",X"CC",X"DB",X"DD",X"FD",X"CA",X"02",X"E6",X"A4",X"5A",X"2F",X"0C",X"4F",X"1F",X"02",
		X"CC",X"07",X"05",X"8D",X"06",X"31",X"3F",X"26",X"F7",X"35",X"A7",X"FD",X"CA",X"06",X"BF",X"CA",
		X"04",X"C6",X"1A",X"F7",X"CA",X"00",X"5F",X"88",X"04",X"30",X"8B",X"39",X"11",X"11",X"11",X"10",
		X"11",X"11",X"11",X"10",X"34",X"06",X"86",X"04",X"BD",X"F0",X"09",X"35",X"86",X"C6",X"11",X"F7",
		X"BF",X"1A",X"C6",X"4A",X"8D",X"04",X"C6",X"58",X"20",X"21",X"34",X"36",X"8E",X"CC",X"88",X"BD",
		X"D2",X"21",X"1F",X"02",X"8E",X"CC",X"24",X"F6",X"BF",X"1A",X"BD",X"D2",X"21",X"1E",X"12",X"BD",
		X"7B",X"00",X"1E",X"12",X"8C",X"CC",X"56",X"26",X"F1",X"35",X"B6",X"34",X"36",X"8E",X"CC",X"8A",
		X"BD",X"D2",X"21",X"1F",X"02",X"8E",X"CC",X"56",X"F6",X"BF",X"1A",X"BD",X"D2",X"21",X"1E",X"12",
		X"BD",X"7B",X"00",X"1E",X"12",X"8C",X"CC",X"88",X"26",X"F1",X"35",X"B6",X"10",X"8E",X"B0",X"00",
		X"AF",X"28",X"C6",X"02",X"E7",X"2E",X"CC",X"DA",X"D2",X"ED",X"26",X"C6",X"19",X"E7",X"A4",X"C6",
		X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",X"5A",X"26",X"FB",X"E7",X"21",X"E7",X"22",X"6F",X"2F",
		X"86",X"32",X"A7",X"23",X"86",X"3C",X"A7",X"24",X"86",X"77",X"A7",X"25",X"AD",X"B8",X"06",X"25",
		X"05",X"BD",X"DB",X"E4",X"20",X"F6",X"39",X"8E",X"25",X"60",X"8D",X"C0",X"C6",X"19",X"8E",X"CC",
		X"24",X"31",X"2F",X"A6",X"A0",X"BD",X"D7",X"9A",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"88",
		X"BD",X"D7",X"9A",X"C6",X"88",X"8D",X"34",X"86",X"34",X"C6",X"22",X"8E",X"48",X"6A",X"BD",X"7B",
		X"00",X"CE",X"DC",X"DB",X"8E",X"CC",X"88",X"BD",X"D7",X"92",X"BD",X"DD",X"3C",X"F7",X"BF",X"28",
		X"7F",X"BF",X"1A",X"C6",X"60",X"BD",X"DB",X"FA",X"B6",X"BF",X"28",X"8E",X"CC",X"88",X"BD",X"D7",
		X"9A",X"86",X"22",X"B7",X"BF",X"1A",X"BD",X"DB",X"FA",X"20",X"D9",X"86",X"51",X"8E",X"25",X"90",
		X"BD",X"7B",X"03",X"86",X"52",X"8E",X"25",X"A0",X"7E",X"7B",X"03",X"86",X"34",X"C6",X"00",X"8E",
		X"48",X"6A",X"BD",X"7B",X"00",X"8D",X"E4",X"8E",X"25",X"70",X"BD",X"DC",X"3C",X"C6",X"19",X"8E",
		X"CC",X"56",X"31",X"2F",X"A6",X"A0",X"BD",X"D7",X"9A",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",
		X"8A",X"BD",X"D7",X"9A",X"C6",X"88",X"8D",X"C3",X"86",X"34",X"C6",X"22",X"8E",X"48",X"7A",X"BD",
		X"7B",X"00",X"CE",X"DD",X"3B",X"8E",X"CC",X"8A",X"BD",X"D7",X"92",X"8D",X"1F",X"F7",X"BF",X"28",
		X"7F",X"BF",X"1A",X"C6",X"70",X"BD",X"DC",X"1B",X"B6",X"BF",X"28",X"8E",X"CC",X"8A",X"BD",X"D7",
		X"9A",X"86",X"22",X"B7",X"BF",X"1A",X"BD",X"DC",X"1B",X"20",X"DA",X"39",X"B6",X"C8",X"0C",X"85",
		X"02",X"27",X"04",X"32",X"62",X"6E",X"C4",X"B6",X"C8",X"04",X"84",X"0C",X"BD",X"DB",X"E4",X"34",
		X"02",X"B6",X"C8",X"04",X"84",X"0C",X"A1",X"E4",X"35",X"02",X"26",X"E0",X"4D",X"27",X"DD",X"85",
		X"FB",X"26",X"06",X"C1",X"18",X"27",X"D5",X"5A",X"39",X"C1",X"40",X"27",X"CF",X"5C",X"39",X"A6",
		X"84",X"84",X"F0",X"27",X"07",X"CC",X"99",X"99",X"ED",X"81",X"ED",X"81",X"39",X"4F",X"5F",X"33",
		X"A4",X"FD",X"BF",X"1B",X"FD",X"BF",X"1D",X"FD",X"BF",X"1F",X"FD",X"BF",X"21",X"7F",X"BF",X"26",
		X"B6",X"CC",X"05",X"44",X"25",X"03",X"7E",X"00",X"12",X"8E",X"9A",X"73",X"8D",X"D1",X"8E",X"9A",
		X"78",X"8D",X"CC",X"8E",X"9A",X"73",X"BD",X"E0",X"E4",X"24",X"26",X"7C",X"BF",X"26",X"BD",X"00",
		X"03",X"64",X"11",X"E0",X"5E",X"86",X"10",X"9B",X"04",X"A7",X"24",X"4F",X"A7",X"A8",X"35",X"8E",
		X"9A",X"73",X"AF",X"A8",X"31",X"8E",X"DD",X"E9",X"AF",X"C8",X"38",X"6F",X"C8",X"36",X"7E",X"DE",
		X"50",X"8E",X"9A",X"73",X"AF",X"C8",X"31",X"4F",X"BD",X"DE",X"8A",X"8E",X"DD",X"E9",X"AF",X"C8",
		X"38",X"86",X"40",X"A7",X"C8",X"36",X"7E",X"DE",X"50",X"7D",X"C8",X"06",X"2A",X"0E",X"BD",X"00",
		X"2A",X"B6",X"BF",X"FF",X"8A",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"8E",X"9A",X"78",X"BD",
		X"E0",X"E4",X"24",X"27",X"7C",X"BF",X"26",X"BD",X"00",X"03",X"64",X"11",X"E0",X"5E",X"86",X"10",
		X"9B",X"04",X"A7",X"24",X"86",X"01",X"A7",X"A8",X"35",X"8E",X"9A",X"78",X"AF",X"A8",X"31",X"8E",
		X"DE",X"42",X"AF",X"C8",X"38",X"6F",X"C8",X"36",X"7E",X"DE",X"50",X"8E",X"9A",X"78",X"AF",X"C8",
		X"31",X"86",X"01",X"8D",X"55",X"8E",X"DE",X"42",X"AF",X"C8",X"38",X"86",X"40",X"A7",X"C8",X"36",
		X"20",X"0E",X"B6",X"BF",X"FF",X"84",X"FD",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"7E",X"00",X"12",
		X"86",X"11",X"BD",X"00",X"0C",X"26",X"29",X"BD",X"00",X"2A",X"8E",X"2B",X"68",X"86",X"58",X"C6",
		X"11",X"BD",X"7B",X"03",X"86",X"29",X"BD",X"7B",X"15",X"BD",X"00",X"0F",X"0D",X"86",X"1E",X"BD",
		X"00",X"09",X"33",X"A4",X"6A",X"C8",X"36",X"27",X"0A",X"86",X"11",X"BD",X"00",X"0C",X"27",X"ED",
		X"6E",X"D8",X"38",X"86",X"11",X"BD",X"00",X"06",X"20",X"F6",X"BD",X"E0",X"EA",X"24",X"1E",X"7C",
		X"BF",X"26",X"34",X"02",X"BD",X"00",X"03",X"64",X"11",X"DE",X"D0",X"86",X"10",X"9B",X"04",X"A7",
		X"24",X"35",X"02",X"A7",X"A8",X"35",X"AE",X"C8",X"31",X"AF",X"A8",X"31",X"39",X"BD",X"E1",X"07",
		X"24",X"1D",X"7C",X"BF",X"26",X"34",X"02",X"BD",X"00",X"03",X"64",X"11",X"DE",X"D0",X"86",X"08",
		X"9B",X"04",X"A7",X"24",X"35",X"02",X"A7",X"A8",X"35",X"AE",X"C8",X"31",X"AF",X"A8",X"31",X"39",
		X"DE",X"08",X"6F",X"C8",X"30",X"E6",X"C8",X"35",X"26",X"09",X"C6",X"3C",X"34",X"04",X"CC",X"5E",
		X"11",X"20",X"0E",X"C6",X"3C",X"7D",X"C8",X"06",X"2A",X"02",X"C6",X"34",X"34",X"04",X"CC",X"5F",
		X"11",X"8E",X"24",X"B0",X"BD",X"7B",X"03",X"30",X"89",X"03",X"00",X"86",X"57",X"BD",X"7B",X"03",
		X"1F",X"98",X"31",X"4B",X"35",X"04",X"E7",X"24",X"8E",X"DF",X"13",X"AF",X"2C",X"8E",X"44",X"78",
		X"BD",X"E1",X"59",X"BD",X"E0",X"EA",X"24",X"15",X"8E",X"CF",X"EA",X"BD",X"E0",X"0B",X"6D",X"C8",
		X"35",X"26",X"06",X"10",X"BF",X"BF",X"1D",X"20",X"04",X"10",X"BF",X"BF",X"21",X"BD",X"E1",X"07",
		X"24",X"19",X"6D",X"C8",X"30",X"27",X"1D",X"30",X"4B",X"30",X"0F",X"10",X"8E",X"CD",X"66",X"C6",
		X"03",X"BD",X"D2",X"54",X"BD",X"D6",X"1B",X"86",X"05",X"8D",X"75",X"24",X"70",X"1F",X"12",X"BD",
		X"D7",X"31",X"20",X"5B",X"30",X"A9",X"32",X"9A",X"26",X"34",X"8E",X"CF",X"96",X"BD",X"E0",X"26",
		X"31",X"26",X"AE",X"C8",X"31",X"C6",X"04",X"BD",X"D2",X"54",X"10",X"8E",X"CD",X"3E",X"6D",X"C8",
		X"35",X"26",X"09",X"10",X"BF",X"BF",X"1B",X"7F",X"BF",X"1F",X"20",X"07",X"10",X"BF",X"BF",X"1F",
		X"7F",X"BF",X"1B",X"30",X"4B",X"30",X"0F",X"C6",X"14",X"BD",X"D2",X"54",X"20",X"A9",X"BD",X"DF",
		X"C4",X"34",X"01",X"34",X"10",X"10",X"AC",X"E1",X"22",X"11",X"8D",X"6F",X"6D",X"C8",X"35",X"26",
		X"06",X"10",X"BF",X"BF",X"1B",X"20",X"04",X"10",X"BF",X"BF",X"1F",X"35",X"01",X"24",X"0E",X"8E",
		X"30",X"A4",X"CC",X"59",X"AA",X"BD",X"7B",X"03",X"86",X"60",X"BD",X"00",X"09",X"7E",X"00",X"00",
		X"34",X"26",X"20",X"0C",X"34",X"26",X"8E",X"CD",X"66",X"8D",X"26",X"86",X"04",X"25",X"01",X"4C",
		X"B7",X"BF",X"06",X"8E",X"CD",X"74",X"8D",X"19",X"24",X"05",X"7A",X"BF",X"06",X"27",X"0E",X"30",
		X"0E",X"8C",X"CF",X"A4",X"25",X"F0",X"8E",X"CF",X"96",X"1C",X"FE",X"35",X"A6",X"1A",X"01",X"35",
		X"A6",X"34",X"10",X"31",X"4B",X"31",X"2F",X"C6",X"03",X"BD",X"D7",X"81",X"A1",X"A0",X"26",X"07",
		X"5A",X"26",X"F6",X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",X"34",X"20",X"BD",X"E0",X"26",
		X"30",X"4B",X"30",X"0F",X"C6",X"03",X"BD",X"D2",X"54",X"AE",X"C8",X"31",X"C6",X"04",X"BD",X"D2",
		X"54",X"35",X"20",X"7E",X"D6",X"3A",X"34",X"30",X"1F",X"12",X"10",X"BC",X"BF",X"1B",X"26",X"05",
		X"30",X"2E",X"BF",X"BF",X"1B",X"BC",X"BF",X"1D",X"26",X"05",X"30",X"2E",X"BF",X"BF",X"1D",X"10",
		X"AC",X"62",X"27",X"0B",X"30",X"32",X"86",X"0E",X"BD",X"D7",X"51",X"31",X"32",X"20",X"DB",X"30",
		X"A8",X"D8",X"BC",X"BF",X"1B",X"26",X"05",X"30",X"2E",X"BF",X"BF",X"1B",X"35",X"B0",X"DE",X"08",
		X"6C",X"C8",X"30",X"31",X"4B",X"A6",X"C8",X"35",X"26",X"09",X"86",X"3C",X"A7",X"24",X"CC",X"5E",
		X"11",X"20",X"0E",X"86",X"3C",X"7D",X"C8",X"06",X"2A",X"02",X"86",X"34",X"A7",X"24",X"CC",X"5F",
		X"11",X"8E",X"10",X"5B",X"BD",X"7B",X"03",X"86",X"56",X"30",X"89",X"03",X"00",X"BD",X"7B",X"03",
		X"1F",X"98",X"8E",X"E0",X"9A",X"AF",X"2C",X"7E",X"E1",X"4B",X"30",X"2F",X"10",X"8E",X"CD",X"3E",
		X"C6",X"14",X"BD",X"D2",X"54",X"10",X"8E",X"CD",X"66",X"8E",X"CF",X"96",X"BD",X"E0",X"26",X"10",
		X"8E",X"CD",X"74",X"BD",X"D6",X"3A",X"AE",X"C8",X"31",X"10",X"8E",X"CD",X"6C",X"C6",X"04",X"BD",
		X"D2",X"54",X"8E",X"D6",X"08",X"10",X"8E",X"CD",X"66",X"C6",X"03",X"BD",X"D2",X"54",X"BD",X"D6",
		X"1B",X"8E",X"CD",X"3E",X"A6",X"C8",X"35",X"26",X"05",X"BF",X"BF",X"1B",X"20",X"03",X"BF",X"BF",
		X"1F",X"7E",X"DE",X"D5",X"10",X"8E",X"CD",X"6C",X"20",X"36",X"34",X"12",X"10",X"8E",X"CF",X"AA",
		X"AE",X"C8",X"31",X"8D",X"2B",X"25",X"0C",X"31",X"2E",X"10",X"8C",X"CF",X"F8",X"25",X"F4",X"1C",
		X"FE",X"35",X"92",X"31",X"3A",X"35",X"92",X"34",X"12",X"10",X"8E",X"CD",X"6C",X"AE",X"C8",X"31",
		X"8D",X"0E",X"25",X"EF",X"31",X"2E",X"10",X"8C",X"CF",X"96",X"25",X"F4",X"1C",X"FE",X"35",X"92",
		X"34",X"36",X"1E",X"12",X"C6",X"04",X"8D",X"17",X"C1",X"04",X"26",X"02",X"84",X"0F",X"A1",X"A0",
		X"22",X"05",X"25",X"07",X"5A",X"26",X"EF",X"1C",X"FE",X"35",X"B6",X"1A",X"01",X"35",X"B6",X"8C",
		X"C0",X"00",X"25",X"04",X"BD",X"D7",X"81",X"39",X"A6",X"80",X"39",X"8E",X"CC",X"16",X"BD",X"D7",
		X"92",X"BD",X"DA",X"53",X"8E",X"26",X"43",X"20",X"02",X"C6",X"03",X"A7",X"25",X"E7",X"A4",X"86",
		X"02",X"A7",X"2E",X"AF",X"28",X"C6",X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",X"5A",X"26",X"FB",
		X"8E",X"DA",X"D2",X"AF",X"26",X"C6",X"0A",X"6F",X"21",X"E7",X"22",X"86",X"25",X"A7",X"23",X"AD",
		X"B8",X"06",X"25",X"17",X"10",X"AF",X"C8",X"3A",X"ED",X"C8",X"36",X"86",X"03",X"BD",X"00",X"09",
		X"33",X"A4",X"10",X"AE",X"C8",X"3A",X"EC",X"C8",X"36",X"20",X"E4",X"6E",X"B8",X"0C",X"42",X"55",
		X"42",X"42",X"4C",X"45",X"53",X"2D",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"7E",X"E2",X"03",X"31",X"A8",X"1B",X"8E",X"9C",X"22",X"AF",X"2F",X"34",X"10",X"CE",X"75",X"A0",
		X"5F",X"A6",X"C5",X"A7",X"85",X"5C",X"C1",X"78",X"26",X"F7",X"AE",X"E4",X"30",X"89",X"01",X"00",
		X"4F",X"5F",X"A7",X"80",X"5C",X"26",X"FB",X"AE",X"E4",X"30",X"89",X"02",X"00",X"CE",X"CC",X"CC",
		X"34",X"10",X"4F",X"EF",X"81",X"4C",X"81",X"07",X"27",X"36",X"81",X"38",X"10",X"27",X"00",X"59",
		X"81",X"62",X"10",X"27",X"00",X"83",X"81",X"6B",X"26",X"E9",X"1F",X"30",X"81",X"FF",X"26",X"05",
		X"CC",X"BB",X"BB",X"20",X"10",X"C3",X"11",X"11",X"81",X"CC",X"10",X"27",X"00",X"99",X"81",X"DD",
		X"26",X"03",X"C3",X"11",X"11",X"1F",X"03",X"35",X"10",X"30",X"89",X"01",X"00",X"7E",X"E2",X"30",
		X"34",X"02",X"1F",X"30",X"5C",X"26",X"04",X"CB",X"FB",X"20",X"05",X"C1",X"CD",X"26",X"01",X"5C",
		X"1F",X"03",X"EF",X"81",X"5A",X"C1",X"CD",X"26",X"03",X"5A",X"20",X"06",X"C1",X"FA",X"26",X"02",
		X"CB",X"05",X"1F",X"03",X"35",X"02",X"7E",X"E2",X"35",X"34",X"02",X"1F",X"30",X"C1",X"FF",X"26",
		X"05",X"83",X"04",X"40",X"20",X"0A",X"C3",X"01",X"10",X"81",X"CD",X"26",X"03",X"C3",X"01",X"10",
		X"1F",X"03",X"EF",X"81",X"83",X"01",X"10",X"81",X"CD",X"26",X"05",X"83",X"01",X"10",X"20",X"D2",
		X"81",X"FA",X"26",X"CE",X"C3",X"05",X"50",X"20",X"C9",X"34",X"02",X"1F",X"30",X"C1",X"FF",X"26",
		X"04",X"C4",X"BF",X"20",X"08",X"CB",X"10",X"C1",X"DC",X"26",X"02",X"CB",X"10",X"1F",X"03",X"EF",
		X"81",X"C0",X"10",X"C1",X"DC",X"26",X"05",X"C0",X"10",X"7E",X"E2",X"92",X"C1",X"AF",X"10",X"26",
		X"FF",X"A0",X"CB",X"50",X"7E",X"E2",X"92",X"35",X"10",X"FC",X"99",X"FC",X"ED",X"30",X"FC",X"99",
		X"FF",X"ED",X"32",X"BD",X"76",X"8D",X"6F",X"24",X"6F",X"34",X"BD",X"E3",X"26",X"BD",X"E3",X"3E",
		X"6F",X"3F",X"BD",X"E3",X"59",X"35",X"10",X"8E",X"75",X"A0",X"BD",X"E3",X"28",X"96",X"00",X"84",
		X"FB",X"97",X"00",X"7E",X"00",X"00",X"AE",X"62",X"AF",X"39",X"CC",X"0A",X"0C",X"ED",X"35",X"CC",
		X"45",X"8F",X"ED",X"37",X"BD",X"76",X"38",X"BD",X"76",X"8D",X"BD",X"76",X"70",X"39",X"EC",X"37",
		X"8B",X"05",X"C0",X"03",X"ED",X"37",X"AE",X"62",X"30",X"89",X"02",X"00",X"AF",X"62",X"CC",X"03",
		X"03",X"ED",X"35",X"CC",X"06",X"07",X"ED",X"3D",X"39",X"AF",X"39",X"86",X"03",X"A7",X"36",X"E6",
		X"34",X"C1",X"22",X"10",X"26",X"00",X"A6",X"EC",X"37",X"C3",X"3A",X"19",X"ED",X"37",X"33",X"88",
		X"10",X"EF",X"39",X"CC",X"04",X"01",X"ED",X"35",X"86",X"03",X"34",X"02",X"BD",X"76",X"38",X"6C",
		X"37",X"6C",X"38",X"35",X"02",X"4A",X"26",X"F2",X"86",X"03",X"34",X"02",X"6A",X"35",X"BD",X"76",
		X"38",X"6C",X"37",X"6C",X"38",X"35",X"02",X"4A",X"26",X"F0",X"6A",X"37",X"A6",X"38",X"8B",X"A0",
		X"A7",X"38",X"BD",X"76",X"38",X"6A",X"37",X"6C",X"38",X"6C",X"35",X"BD",X"76",X"38",X"6C",X"35",
		X"86",X"04",X"34",X"02",X"6A",X"37",X"6C",X"38",X"BD",X"76",X"38",X"35",X"02",X"4A",X"26",X"F2",
		X"A6",X"37",X"80",X"77",X"A7",X"37",X"86",X"04",X"34",X"02",X"BD",X"76",X"38",X"6A",X"37",X"6A",
		X"38",X"35",X"02",X"4A",X"26",X"F2",X"6C",X"37",X"6A",X"35",X"BD",X"76",X"38",X"6A",X"38",X"6A",
		X"35",X"BD",X"76",X"38",X"A6",X"38",X"80",X"A1",X"A7",X"38",X"86",X"03",X"34",X"02",X"BD",X"76",
		X"38",X"6A",X"38",X"6C",X"35",X"35",X"02",X"4A",X"26",X"F2",X"86",X"03",X"34",X"02",X"BD",X"76",
		X"38",X"6C",X"37",X"6A",X"38",X"35",X"02",X"4A",X"26",X"F2",X"7E",X"EC",X"C6",X"C1",X"1C",X"25",
		X"57",X"C0",X"1B",X"34",X"04",X"86",X"04",X"3D",X"CB",X"1E",X"E7",X"A4",X"E6",X"E4",X"86",X"03",
		X"3D",X"CB",X"04",X"E7",X"21",X"EC",X"37",X"AB",X"A4",X"EB",X"21",X"ED",X"37",X"CC",X"02",X"01",
		X"ED",X"35",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",X"6C",X"37",X"6C",X"36",X"BD",X"76",
		X"38",X"6A",X"38",X"6C",X"36",X"E6",X"E4",X"5C",X"86",X"03",X"3D",X"E7",X"3B",X"35",X"02",X"4C",
		X"81",X"04",X"25",X"09",X"80",X"03",X"C6",X"02",X"3D",X"EB",X"3B",X"E7",X"3B",X"A6",X"34",X"A0",
		X"3B",X"8B",X"03",X"34",X"02",X"7E",X"E5",X"8D",X"54",X"25",X"0A",X"E7",X"3C",X"86",X"0D",X"A0",
		X"3C",X"33",X"86",X"20",X"03",X"33",X"88",X"10",X"EF",X"39",X"A6",X"34",X"81",X"1A",X"26",X"0E",
		X"33",X"88",X"10",X"EF",X"39",X"CC",X"10",X"02",X"ED",X"35",X"6C",X"38",X"20",X"0B",X"81",X"1B",
		X"27",X"0A",X"4D",X"26",X"04",X"86",X"02",X"A7",X"3B",X"BD",X"76",X"38",X"E6",X"34",X"86",X"01",
		X"4C",X"C0",X"04",X"24",X"FB",X"CB",X"04",X"C1",X"02",X"26",X"01",X"4C",X"A7",X"35",X"5D",X"27",
		X"14",X"C1",X"03",X"27",X"10",X"80",X"02",X"A7",X"3C",X"86",X"0E",X"A0",X"3C",X"A7",X"3B",X"33",
		X"86",X"EF",X"39",X"20",X"05",X"33",X"88",X"10",X"EF",X"39",X"A6",X"34",X"27",X"06",X"4A",X"44",
		X"8B",X"03",X"A7",X"3B",X"A6",X"37",X"AB",X"3B",X"A7",X"37",X"6C",X"38",X"A6",X"34",X"81",X"1A",
		X"26",X"08",X"6A",X"38",X"86",X"03",X"A7",X"36",X"20",X"04",X"81",X"1B",X"27",X"03",X"BD",X"76",
		X"38",X"33",X"88",X"10",X"EF",X"39",X"86",X"01",X"A7",X"3B",X"A6",X"34",X"80",X"02",X"25",X"7B",
		X"27",X"53",X"6C",X"3B",X"80",X"04",X"27",X"4D",X"22",X"F8",X"EC",X"37",X"AB",X"3B",X"5C",X"ED",
		X"37",X"A6",X"34",X"81",X"1B",X"26",X"08",X"86",X"01",X"A7",X"36",X"6C",X"38",X"6C",X"38",X"BD",
		X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"34",X"80",X"04",X"25",X"4E",X"44",X"44",X"8B",
		X"02",X"A7",X"3B",X"EC",X"37",X"AB",X"3B",X"5C",X"ED",X"37",X"A6",X"34",X"81",X"1B",X"26",X"04",
		X"6A",X"38",X"6A",X"36",X"BD",X"76",X"38",X"A6",X"34",X"81",X"1B",X"10",X"26",X"00",X"2C",X"6C",
		X"36",X"6A",X"38",X"20",X"26",X"6A",X"35",X"6C",X"3B",X"EC",X"37",X"AB",X"3B",X"5C",X"ED",X"37",
		X"BD",X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"3B",X"81",X"02",X"27",X"0D",X"4A",X"A7",
		X"3B",X"EC",X"37",X"AB",X"3B",X"5C",X"ED",X"37",X"BD",X"76",X"38",X"C6",X"02",X"A6",X"34",X"27",
		X"0A",X"81",X"03",X"22",X"08",X"5C",X"81",X"03",X"26",X"01",X"5C",X"1F",X"98",X"34",X"02",X"6C",
		X"37",X"6C",X"38",X"BD",X"76",X"38",X"35",X"02",X"4A",X"26",X"F2",X"A6",X"34",X"81",X"1D",X"25",
		X"47",X"EC",X"37",X"4C",X"CB",X"03",X"ED",X"37",X"6A",X"35",X"6A",X"36",X"A6",X"34",X"81",X"1D",
		X"27",X"02",X"6A",X"36",X"BD",X"76",X"38",X"86",X"08",X"E6",X"34",X"C0",X"1C",X"3D",X"E7",X"3B",
		X"86",X"70",X"AB",X"3B",X"E6",X"34",X"C1",X"1D",X"27",X"01",X"4C",X"A7",X"22",X"A6",X"38",X"AB",
		X"22",X"A7",X"38",X"BD",X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"34",X"81",X"1D",X"26",
		X"02",X"6C",X"38",X"A6",X"E4",X"7E",X"E7",X"2B",X"33",X"0E",X"EF",X"39",X"6C",X"37",X"6C",X"38",
		X"BD",X"76",X"38",X"A6",X"34",X"10",X"27",X"00",X"6C",X"81",X"17",X"25",X"13",X"80",X"16",X"34",
		X"02",X"C6",X"02",X"3D",X"E7",X"3B",X"86",X"0E",X"A0",X"3B",X"A7",X"3B",X"34",X"02",X"A6",X"34",
		X"4A",X"34",X"02",X"33",X"88",X"10",X"EF",X"39",X"6C",X"38",X"BD",X"76",X"38",X"6C",X"37",X"6C",
		X"38",X"A6",X"34",X"81",X"17",X"25",X"31",X"6A",X"3B",X"26",X"2D",X"81",X"17",X"26",X"04",X"6A",
		X"35",X"20",X"29",X"35",X"02",X"CC",X"01",X"04",X"ED",X"35",X"BD",X"76",X"38",X"A6",X"61",X"C6",
		X"0C",X"3D",X"E7",X"3B",X"A6",X"38",X"8B",X"26",X"AB",X"3B",X"A7",X"38",X"BD",X"76",X"38",X"6C",
		X"38",X"A6",X"E4",X"A7",X"3B",X"7E",X"E6",X"C6",X"33",X"0E",X"EF",X"39",X"BD",X"76",X"38",X"35",
		X"02",X"80",X"02",X"24",X"AC",X"A6",X"34",X"44",X"25",X"2A",X"86",X"02",X"A7",X"3B",X"A6",X"38",
		X"AB",X"3B",X"A7",X"38",X"CC",X"03",X"01",X"ED",X"35",X"33",X"0D",X"EF",X"39",X"A6",X"3D",X"34",
		X"02",X"BD",X"76",X"38",X"6C",X"38",X"35",X"02",X"4A",X"26",X"F4",X"CC",X"02",X"03",X"ED",X"35",
		X"6A",X"38",X"20",X"24",X"33",X"88",X"10",X"EF",X"39",X"A6",X"3E",X"80",X"03",X"23",X"0F",X"E6",
		X"38",X"CB",X"03",X"E7",X"38",X"34",X"02",X"BD",X"76",X"38",X"35",X"02",X"20",X"ED",X"8B",X"03",
		X"A7",X"3B",X"A6",X"38",X"AB",X"3B",X"A7",X"38",X"A6",X"34",X"81",X"17",X"27",X"05",X"33",X"88",
		X"6B",X"EF",X"39",X"BD",X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"34",X"27",X"2D",X"4A",
		X"6A",X"37",X"6C",X"38",X"33",X"88",X"10",X"EF",X"39",X"34",X"02",X"BD",X"76",X"38",X"6C",X"38",
		X"33",X"88",X"6B",X"EF",X"39",X"BD",X"76",X"38",X"A6",X"34",X"81",X"18",X"25",X"08",X"6A",X"3B",
		X"26",X"04",X"35",X"02",X"20",X"06",X"35",X"02",X"80",X"02",X"24",X"D4",X"33",X"88",X"10",X"EF",
		X"39",X"A6",X"34",X"81",X"1C",X"25",X"04",X"A6",X"62",X"20",X"20",X"81",X"03",X"22",X"12",X"C6",
		X"03",X"E7",X"3C",X"81",X"02",X"25",X"12",X"6C",X"3C",X"81",X"03",X"26",X"0C",X"6C",X"3C",X"20",
		X"08",X"A7",X"3C",X"81",X"1B",X"27",X"02",X"6C",X"3C",X"A6",X"3C",X"6A",X"37",X"6C",X"38",X"34",
		X"02",X"BD",X"76",X"38",X"35",X"02",X"4A",X"26",X"F2",X"A6",X"34",X"81",X"1B",X"25",X"50",X"22",
		X"0D",X"6A",X"37",X"6C",X"38",X"6A",X"36",X"BD",X"76",X"38",X"6C",X"36",X"20",X"41",X"6A",X"37",
		X"6C",X"38",X"6A",X"35",X"6A",X"36",X"BD",X"76",X"38",X"6A",X"37",X"6C",X"38",X"6A",X"36",X"BD",
		X"76",X"38",X"A6",X"37",X"A0",X"A4",X"A0",X"A4",X"4A",X"A7",X"37",X"BD",X"76",X"38",X"6C",X"36",
		X"6A",X"37",X"6A",X"38",X"BD",X"76",X"38",X"6A",X"37",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"34",
		X"81",X"1D",X"25",X"04",X"A6",X"E4",X"20",X"02",X"A6",X"62",X"A7",X"3C",X"7E",X"EA",X"22",X"A6",
		X"34",X"81",X"04",X"10",X"24",X"00",X"69",X"44",X"24",X"3C",X"26",X"20",X"33",X"88",X"6B",X"EF",
		X"39",X"6A",X"37",X"6C",X"38",X"BD",X"76",X"38",X"EC",X"37",X"80",X"03",X"5C",X"ED",X"37",X"33",
		X"88",X"10",X"EF",X"39",X"6C",X"35",X"BD",X"76",X"38",X"7E",X"E8",X"E6",X"6A",X"37",X"6A",X"37",
		X"6C",X"38",X"BD",X"76",X"38",X"6C",X"35",X"6C",X"35",X"EC",X"37",X"80",X"04",X"5C",X"ED",X"37",
		X"BD",X"76",X"38",X"7E",X"E8",X"E6",X"6C",X"35",X"33",X"88",X"68",X"EF",X"39",X"6A",X"37",X"6A",
		X"37",X"6C",X"38",X"BD",X"76",X"38",X"A6",X"34",X"10",X"27",X"00",X"FA",X"33",X"88",X"65",X"EF",
		X"39",X"6C",X"35",X"EC",X"37",X"80",X"03",X"5C",X"ED",X"37",X"BD",X"76",X"38",X"7E",X"E8",X"E6",
		X"80",X"04",X"C6",X"01",X"E7",X"3B",X"6F",X"3C",X"6C",X"3B",X"6C",X"35",X"80",X"02",X"25",X"06",
		X"6C",X"3C",X"80",X"02",X"24",X"F0",X"8B",X"02",X"34",X"02",X"EC",X"37",X"A0",X"3B",X"5C",X"ED",
		X"37",X"A6",X"34",X"81",X"1B",X"26",X"26",X"35",X"02",X"6A",X"36",X"6A",X"36",X"BD",X"76",X"38",
		X"A6",X"37",X"80",X"38",X"A7",X"37",X"BD",X"76",X"38",X"6A",X"37",X"6A",X"38",X"CC",X"02",X"02",
		X"ED",X"35",X"BD",X"76",X"38",X"6C",X"36",X"A6",X"34",X"4A",X"7E",X"EA",X"1E",X"BD",X"76",X"38",
		X"EC",X"37",X"A0",X"3B",X"A0",X"3C",X"5C",X"ED",X"37",X"35",X"02",X"E6",X"3C",X"26",X"40",X"81",
		X"00",X"27",X"20",X"BD",X"76",X"18",X"BD",X"76",X"38",X"A6",X"35",X"AB",X"3B",X"A7",X"35",X"A7",
		X"3B",X"EC",X"37",X"A0",X"3B",X"5C",X"ED",X"37",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",
		X"7E",X"E8",X"E6",X"BD",X"76",X"38",X"A6",X"35",X"AB",X"3B",X"A7",X"35",X"4A",X"A7",X"3B",X"EC",
		X"37",X"A0",X"3B",X"5C",X"ED",X"37",X"BD",X"76",X"18",X"BD",X"76",X"38",X"7E",X"E8",X"E6",X"81",
		X"00",X"27",X"18",X"BD",X"76",X"38",X"A6",X"3B",X"4C",X"48",X"A7",X"35",X"A7",X"3B",X"EC",X"37",
		X"A0",X"3B",X"5C",X"ED",X"37",X"BD",X"76",X"38",X"7E",X"E8",X"E6",X"6C",X"35",X"BD",X"76",X"18",
		X"BD",X"76",X"38",X"A6",X"35",X"AB",X"3B",X"A7",X"35",X"4A",X"A7",X"3B",X"EC",X"37",X"A0",X"3B",
		X"5C",X"ED",X"37",X"BD",X"76",X"18",X"A6",X"34",X"81",X"1A",X"26",X"07",X"6A",X"36",X"33",X"88",
		X"10",X"EF",X"39",X"BD",X"76",X"38",X"86",X"02",X"A7",X"3B",X"A6",X"34",X"6C",X"3B",X"80",X"02",
		X"24",X"FA",X"A6",X"37",X"A0",X"3B",X"A7",X"37",X"A6",X"34",X"44",X"25",X"1F",X"A6",X"35",X"80",
		X"02",X"C6",X"02",X"3D",X"E7",X"3C",X"C6",X"C1",X"E0",X"3C",X"1F",X"13",X"3A",X"AF",X"39",X"1F",
		X"31",X"A6",X"34",X"81",X"1A",X"26",X"05",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",X"86",
		X"03",X"A7",X"36",X"A6",X"34",X"10",X"27",X"00",X"D9",X"81",X"04",X"24",X"53",X"81",X"02",X"27",
		X"32",X"6A",X"35",X"C6",X"02",X"E7",X"3B",X"4A",X"27",X"04",X"6A",X"35",X"20",X"06",X"33",X"89",
		X"00",X"C1",X"EF",X"39",X"EC",X"37",X"A0",X"3B",X"5A",X"ED",X"37",X"BD",X"76",X"38",X"A6",X"34",
		X"81",X"03",X"10",X"26",X"00",X"AC",X"EC",X"37",X"A0",X"3B",X"5A",X"ED",X"37",X"BD",X"76",X"38",
		X"7E",X"EA",X"02",X"6A",X"35",X"6A",X"37",X"6A",X"37",X"6A",X"38",X"6A",X"3C",X"6A",X"3C",X"C6",
		X"C1",X"E0",X"3C",X"1F",X"13",X"3A",X"AF",X"39",X"1F",X"31",X"BD",X"76",X"38",X"7E",X"EA",X"02",
		X"C6",X"02",X"E7",X"3C",X"80",X"04",X"6C",X"3C",X"80",X"04",X"24",X"FA",X"8B",X"04",X"81",X"02",
		X"26",X"02",X"6C",X"3C",X"E6",X"3C",X"E7",X"35",X"81",X"00",X"27",X"04",X"81",X"02",X"26",X"01",
		X"5A",X"E7",X"3B",X"34",X"02",X"EC",X"37",X"A0",X"3B",X"5A",X"ED",X"37",X"35",X"02",X"81",X"01",
		X"27",X"1F",X"81",X"02",X"26",X"06",X"86",X"C1",X"A7",X"3C",X"20",X"19",X"33",X"88",X"10",X"EF",
		X"39",X"BD",X"76",X"38",X"EC",X"37",X"A0",X"3B",X"5A",X"ED",X"37",X"BD",X"76",X"38",X"7E",X"EA",
		X"02",X"86",X"C3",X"A7",X"3C",X"A6",X"34",X"44",X"44",X"4C",X"C6",X"02",X"3D",X"E7",X"23",X"E6",
		X"3C",X"E0",X"23",X"1F",X"13",X"3A",X"AF",X"39",X"1F",X"31",X"BD",X"76",X"38",X"A6",X"3B",X"A7",
		X"35",X"6A",X"3B",X"EC",X"37",X"A0",X"3B",X"5A",X"ED",X"37",X"33",X"88",X"10",X"EF",X"39",X"BD",
		X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"33",X"88",X"10",X"EF",X"39",X"A6",X"34",X"81",X"03",
		X"24",X"0C",X"C6",X"03",X"E7",X"3C",X"81",X"02",X"26",X"08",X"6C",X"3C",X"20",X"04",X"A7",X"3C",
		X"6C",X"3C",X"6A",X"37",X"6A",X"38",X"BD",X"76",X"38",X"6A",X"3C",X"26",X"F5",X"A6",X"34",X"81",
		X"1D",X"25",X"2E",X"6A",X"38",X"6A",X"35",X"6A",X"36",X"81",X"1D",X"26",X"04",X"6A",X"38",X"20",
		X"02",X"6A",X"36",X"BD",X"76",X"38",X"A6",X"38",X"A0",X"22",X"A7",X"38",X"BD",X"76",X"38",X"6A",
		X"37",X"6A",X"38",X"6A",X"38",X"CC",X"02",X"03",X"ED",X"35",X"35",X"02",X"A7",X"3C",X"7E",X"EB",
		X"D7",X"6A",X"37",X"6A",X"38",X"1F",X"13",X"C6",X"C1",X"3A",X"AF",X"39",X"1F",X"31",X"BD",X"76",
		X"38",X"A6",X"34",X"10",X"27",X"00",X"69",X"81",X"17",X"25",X"04",X"E6",X"E4",X"E7",X"3B",X"4A",
		X"6A",X"38",X"33",X"88",X"10",X"EF",X"39",X"34",X"02",X"BD",X"76",X"38",X"6A",X"38",X"A6",X"34",
		X"81",X"17",X"25",X"38",X"6A",X"3B",X"26",X"34",X"81",X"17",X"26",X"04",X"6A",X"35",X"20",X"37",
		X"35",X"02",X"CC",X"01",X"04",X"ED",X"35",X"6A",X"38",X"BD",X"76",X"38",X"A6",X"61",X"C6",X"0C",
		X"3D",X"E7",X"3B",X"A6",X"38",X"80",X"26",X"A0",X"3B",X"A7",X"38",X"BD",X"76",X"38",X"6A",X"37",
		X"CC",X"02",X"03",X"ED",X"35",X"35",X"06",X"A7",X"3B",X"7E",X"EB",X"0B",X"6A",X"37",X"1F",X"13",
		X"C6",X"C1",X"3A",X"AF",X"39",X"1F",X"31",X"BD",X"76",X"38",X"35",X"02",X"80",X"02",X"24",X"A0",
		X"A6",X"34",X"44",X"25",X"5C",X"CC",X"03",X"01",X"ED",X"35",X"6A",X"37",X"33",X"88",X"71",X"EF",
		X"39",X"A6",X"3D",X"34",X"02",X"BD",X"76",X"38",X"6A",X"38",X"35",X"02",X"4A",X"26",X"F4",X"6C",
		X"37",X"6A",X"38",X"CC",X"02",X"03",X"ED",X"35",X"BD",X"76",X"38",X"A6",X"34",X"10",X"27",X"00",
		X"92",X"44",X"34",X"02",X"6C",X"37",X"6A",X"38",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",
		X"6A",X"38",X"33",X"88",X"71",X"EF",X"39",X"BD",X"76",X"38",X"A6",X"34",X"81",X"18",X"25",X"09",
		X"6A",X"3B",X"26",X"05",X"35",X"02",X"7E",X"EB",X"A3",X"35",X"02",X"4A",X"26",X"D4",X"7E",X"EB",
		X"A3",X"33",X"88",X"10",X"EF",X"39",X"A6",X"3E",X"80",X"03",X"23",X"0F",X"34",X"02",X"A6",X"38",
		X"80",X"03",X"A7",X"38",X"BD",X"76",X"38",X"35",X"02",X"20",X"ED",X"8B",X"03",X"A7",X"3B",X"A6",
		X"38",X"A0",X"3B",X"A7",X"38",X"A6",X"34",X"81",X"17",X"27",X"05",X"33",X"88",X"71",X"EF",X"39",
		X"BD",X"76",X"38",X"CC",X"02",X"03",X"ED",X"35",X"A6",X"34",X"81",X"17",X"26",X"06",X"6A",X"37",
		X"35",X"04",X"35",X"04",X"4A",X"34",X"02",X"33",X"88",X"10",X"EF",X"39",X"6C",X"37",X"6A",X"38",
		X"BD",X"76",X"38",X"33",X"88",X"71",X"EF",X"39",X"6A",X"38",X"BD",X"76",X"38",X"35",X"02",X"80",
		X"02",X"24",X"E2",X"A6",X"34",X"81",X"1C",X"25",X"0B",X"33",X"88",X"10",X"EF",X"39",X"35",X"02",
		X"A7",X"3C",X"20",X"23",X"81",X"04",X"24",X"12",X"C6",X"03",X"E7",X"3C",X"81",X"02",X"25",X"12",
		X"6C",X"3C",X"81",X"02",X"27",X"0C",X"6C",X"3C",X"20",X"08",X"A7",X"3C",X"81",X"1B",X"27",X"02",
		X"6C",X"3C",X"33",X"88",X"10",X"EF",X"39",X"6C",X"37",X"6A",X"38",X"BD",X"76",X"38",X"6A",X"3C",
		X"26",X"F5",X"A6",X"34",X"81",X"1B",X"25",X"27",X"22",X"14",X"6C",X"37",X"6A",X"36",X"BD",X"76",
		X"38",X"CC",X"08",X"01",X"ED",X"35",X"6C",X"37",X"BD",X"76",X"38",X"7E",X"EC",X"C6",X"6C",X"37",
		X"6A",X"36",X"BD",X"76",X"38",X"6C",X"37",X"6A",X"36",X"BD",X"76",X"38",X"7E",X"EC",X"C6",X"A6",
		X"34",X"81",X"04",X"24",X"3D",X"81",X"03",X"26",X"04",X"6C",X"37",X"20",X"05",X"33",X"88",X"71",
		X"EF",X"39",X"6C",X"37",X"6A",X"38",X"44",X"25",X"02",X"6C",X"35",X"BD",X"76",X"38",X"A6",X"34",
		X"10",X"27",X"00",X"92",X"6C",X"37",X"6C",X"37",X"6A",X"38",X"C6",X"03",X"E7",X"35",X"81",X"02",
		X"25",X"02",X"6C",X"35",X"44",X"24",X"05",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",X"7E",
		X"EC",X"C6",X"6C",X"37",X"6A",X"38",X"80",X"04",X"C6",X"01",X"E7",X"3B",X"6C",X"35",X"6C",X"3B",
		X"80",X"04",X"24",X"F8",X"8B",X"04",X"34",X"02",X"BD",X"76",X"38",X"35",X"02",X"81",X"03",X"26",
		X"02",X"6C",X"3B",X"81",X"02",X"26",X"02",X"6C",X"35",X"81",X"00",X"27",X"09",X"81",X"03",X"27",
		X"05",X"33",X"88",X"71",X"EF",X"39",X"34",X"02",X"EC",X"37",X"AB",X"3B",X"5A",X"ED",X"37",X"BD",
		X"76",X"38",X"35",X"02",X"81",X"02",X"27",X"05",X"33",X"88",X"10",X"EF",X"39",X"E6",X"35",X"EB",
		X"3B",X"E7",X"35",X"81",X"00",X"27",X"06",X"81",X"03",X"27",X"02",X"6C",X"3B",X"EC",X"37",X"AB",
		X"3B",X"5A",X"ED",X"37",X"A6",X"34",X"81",X"1A",X"26",X"09",X"6C",X"38",X"6A",X"36",X"33",X"88",
		X"10",X"EF",X"39",X"BD",X"76",X"38",X"A6",X"24",X"10",X"27",X"01",X"8A",X"BD",X"EF",X"6D",X"BD",
		X"76",X"5C",X"6A",X"34",X"A6",X"34",X"D6",X"8D",X"2B",X"15",X"0D",X"00",X"2A",X"33",X"81",X"11",
		X"26",X"2C",X"34",X"20",X"BD",X"00",X"03",X"64",X"17",X"00",X"27",X"35",X"20",X"20",X"1F",X"81",
		X"13",X"22",X"1B",X"27",X"16",X"81",X"10",X"26",X"09",X"34",X"32",X"86",X"2A",X"BD",X"7B",X"12",
		X"35",X"32",X"BD",X"00",X"21",X"D6",X"37",X"CB",X"03",X"D7",X"37",X"BD",X"00",X"24",X"7E",X"EE",
		X"21",X"81",X"FF",X"27",X"06",X"81",X"14",X"10",X"22",X"01",X"06",X"EC",X"35",X"34",X"7F",X"CC",
		X"02",X"01",X"ED",X"35",X"6F",X"2D",X"A6",X"34",X"81",X"14",X"27",X"44",X"81",X"0D",X"27",X"4E",
		X"81",X"06",X"27",X"53",X"81",X"FF",X"27",X"0A",X"81",X"05",X"10",X"22",X"00",X"7F",X"27",X"4C",
		X"20",X"58",X"EE",X"25",X"BD",X"ED",X"CF",X"EE",X"27",X"BD",X"ED",X"CF",X"CC",X"44",X"A5",X"ED",
		X"29",X"ED",X"2B",X"CE",X"77",X"0E",X"86",X"07",X"34",X"02",X"BD",X"ED",X"CF",X"BD",X"EE",X"10",
		X"6C",X"29",X"6C",X"29",X"6C",X"2B",X"6C",X"2B",X"35",X"02",X"4A",X"26",X"EB",X"7E",X"EE",X"1D",
		X"CE",X"77",X"0E",X"EF",X"25",X"CC",X"0E",X"87",X"ED",X"29",X"86",X"85",X"20",X"3D",X"CC",X"1F",
		X"91",X"ED",X"29",X"86",X"74",X"20",X"34",X"CC",X"64",X"9B",X"20",X"2F",X"CC",X"32",X"9B",X"ED",
		X"29",X"EE",X"25",X"EF",X"27",X"CE",X"77",X"0E",X"EF",X"25",X"EE",X"25",X"BD",X"ED",X"CF",X"34",
		X"40",X"EE",X"27",X"BD",X"ED",X"CF",X"EE",X"25",X"EF",X"27",X"35",X"40",X"BD",X"EE",X"10",X"EF",
		X"25",X"6C",X"29",X"6C",X"29",X"6A",X"2B",X"6A",X"2B",X"20",X"62",X"ED",X"2B",X"EE",X"25",X"BD",
		X"ED",X"CF",X"BD",X"ED",X"CF",X"6C",X"29",X"6C",X"29",X"6A",X"2B",X"6A",X"2B",X"20",X"4E",X"6F",
		X"24",X"6D",X"2D",X"26",X"06",X"EC",X"29",X"6C",X"2D",X"20",X"04",X"EC",X"2B",X"6F",X"2D",X"ED",
		X"37",X"6F",X"2E",X"EC",X"C1",X"34",X"02",X"AB",X"2E",X"A7",X"2E",X"58",X"34",X"04",X"8E",X"76",
		X"9A",X"30",X"85",X"AF",X"39",X"BD",X"76",X"38",X"6C",X"38",X"35",X"04",X"35",X"02",X"4A",X"34",
		X"02",X"26",X"E9",X"32",X"61",X"A6",X"2E",X"81",X"31",X"26",X"D8",X"6C",X"24",X"EF",X"25",X"39",
		X"6F",X"2E",X"A6",X"C1",X"AB",X"2E",X"A7",X"2E",X"81",X"31",X"26",X"F6",X"39",X"35",X"7F",X"ED",
		X"35",X"A6",X"34",X"44",X"24",X"08",X"A6",X"3E",X"80",X"04",X"A7",X"3E",X"20",X"06",X"A6",X"3D",
		X"80",X"04",X"A7",X"3D",X"86",X"4A",X"A7",X"37",X"86",X"21",X"A0",X"34",X"C6",X"03",X"3D",X"E7",
		X"22",X"86",X"29",X"AB",X"22",X"A7",X"38",X"A6",X"34",X"81",X"FF",X"10",X"26",X"F5",X"0A",X"39",
		X"57",X"D8",X"58",X"0E",X"58",X"44",X"A6",X"34",X"81",X"15",X"26",X"03",X"BD",X"00",X"1E",X"81",
		X"22",X"26",X"15",X"BD",X"00",X"0F",X"14",X"BD",X"EE",X"E4",X"6C",X"24",X"86",X"4A",X"A7",X"37",
		X"AE",X"62",X"BD",X"76",X"2A",X"7E",X"E3",X"59",X"80",X"03",X"24",X"FC",X"8E",X"EE",X"56",X"48",
		X"AE",X"86",X"CC",X"47",X"3E",X"1A",X"FF",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"8E",X"02",X"0D",
		X"BF",X"CA",X"06",X"86",X"2A",X"B7",X"CA",X"00",X"8E",X"00",X"09",X"CB",X"09",X"F7",X"CA",X"05",
		X"B7",X"CA",X"00",X"30",X"1F",X"26",X"F4",X"1C",X"00",X"AE",X"62",X"A6",X"3F",X"4C",X"84",X"03",
		X"5F",X"A7",X"3F",X"30",X"8B",X"86",X"4A",X"A7",X"37",X"A6",X"34",X"4C",X"BD",X"76",X"2C",X"6C",
		X"34",X"A6",X"34",X"44",X"8B",X"03",X"A7",X"35",X"A6",X"34",X"44",X"25",X"08",X"A6",X"3E",X"8B",
		X"04",X"A7",X"3E",X"20",X"06",X"A6",X"3D",X"8B",X"04",X"A7",X"3D",X"BD",X"76",X"8D",X"BD",X"76",
		X"70",X"7E",X"E3",X"59",X"AE",X"64",X"A6",X"3F",X"5F",X"30",X"8B",X"86",X"1A",X"A7",X"23",X"A6",
		X"23",X"44",X"8B",X"03",X"A7",X"3B",X"A7",X"35",X"86",X"4A",X"A0",X"3B",X"A7",X"37",X"A6",X"23",
		X"C6",X"03",X"E7",X"36",X"3D",X"E7",X"3B",X"86",X"8C",X"A0",X"3B",X"A7",X"38",X"A6",X"23",X"81",
		X"1A",X"26",X"06",X"6C",X"38",X"6A",X"36",X"20",X"08",X"44",X"25",X"05",X"33",X"88",X"71",X"20",
		X"03",X"33",X"88",X"10",X"EF",X"39",X"BD",X"76",X"38",X"86",X"4A",X"A7",X"37",X"A6",X"23",X"81",
		X"1A",X"27",X"0B",X"44",X"25",X"08",X"86",X"10",X"A0",X"35",X"33",X"86",X"EF",X"39",X"BD",X"76",
		X"38",X"AE",X"64",X"A6",X"3F",X"4A",X"84",X"03",X"5F",X"A7",X"3F",X"30",X"8B",X"6A",X"23",X"2A",
		X"9E",X"8E",X"75",X"A0",X"BD",X"E3",X"28",X"AE",X"64",X"30",X"89",X"FF",X"00",X"8E",X"47",X"3E",
		X"86",X"88",X"A7",X"84",X"30",X"89",X"01",X"00",X"8C",X"4E",X"3E",X"26",X"F5",X"34",X"10",X"4F",
		X"BD",X"00",X"09",X"31",X"A8",X"1B",X"35",X"90",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"D0",X"11",X"3F",X"3F",X"3F",X"3F",X"D0",X"26",
		X"7E",X"F0",X"1F",X"7E",X"F3",X"3E",X"7E",X"F4",X"6F",X"7E",X"F9",X"5F",X"7E",X"FF",X"21",X"00",
		X"F9",X"07",X"28",X"2F",X"00",X"A4",X"15",X"C7",X"FF",X"38",X"17",X"CC",X"81",X"81",X"2F",X"1A",
		X"FF",X"10",X"CE",X"BF",X"00",X"7F",X"C8",X"0D",X"7F",X"C8",X"0C",X"86",X"3C",X"B7",X"C8",X"0D",
		X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",X"B7",X"C8",X"0F",X"86",X"C0",X"B7",
		X"C8",X"0E",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"F0",X"0F",X"10",X"8E",X"C0",X"00",X"EC",X"81",
		X"ED",X"A1",X"8C",X"F0",X"1F",X"25",X"F7",X"86",X"02",X"10",X"8E",X"F0",X"62",X"8E",X"00",X"00",
		X"20",X"3A",X"10",X"8E",X"F0",X"69",X"7E",X"F2",X"8A",X"86",X"34",X"B7",X"C8",X"0D",X"B7",X"C8",
		X"0F",X"7F",X"C8",X"0E",X"86",X"BF",X"1F",X"8B",X"10",X"CE",X"BF",X"00",X"BD",X"D2",X"1E",X"86",
		X"05",X"8E",X"30",X"70",X"C6",X"99",X"BD",X"7B",X"03",X"86",X"06",X"8E",X"3A",X"90",X"C6",X"99",
		X"BD",X"7B",X"03",X"10",X"8E",X"D2",X"00",X"86",X"07",X"7E",X"F1",X"CA",X"1A",X"3F",X"7F",X"C9",
		X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",
		X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"ED",
		X"81",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",X"26",
		X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",X"00",
		X"26",X"C8",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",
		X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"10",X"A3",X"81",X"26",
		X"43",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",X"26",
		X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",X"00",
		X"26",X"C5",X"1F",X"03",X"1F",X"B8",X"81",X"FF",X"26",X"05",X"1F",X"30",X"7E",X"F0",X"A7",X"4A",
		X"1F",X"8B",X"81",X"80",X"27",X"07",X"4D",X"1F",X"30",X"10",X"26",X"FF",X"6A",X"C6",X"01",X"F7",
		X"C9",X"00",X"6E",X"A4",X"30",X"1E",X"A8",X"84",X"E8",X"01",X"4D",X"26",X"07",X"5D",X"26",X"04",
		X"30",X"02",X"20",X"AD",X"CE",X"00",X"30",X"1E",X"10",X"5F",X"1E",X"10",X"8C",X"00",X"00",X"27",
		X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",X"10",X"11",X"83",X"00",X"30",X"23",X"EE",X"CE",X"00",
		X"10",X"20",X"E9",X"33",X"41",X"47",X"25",X"05",X"57",X"25",X"02",X"20",X"F6",X"1F",X"30",X"86",
		X"01",X"B7",X"C9",X"00",X"10",X"CE",X"F1",X"8A",X"20",X"54",X"86",X"BF",X"1F",X"8B",X"1F",X"A8",
		X"43",X"10",X"CE",X"BF",X"00",X"BD",X"D2",X"1E",X"85",X"C0",X"26",X"0A",X"86",X"05",X"8E",X"30",
		X"70",X"C6",X"22",X"BD",X"7B",X"03",X"86",X"07",X"8E",X"40",X"90",X"C6",X"22",X"BD",X"7B",X"03",
		X"1F",X"30",X"1F",X"98",X"C6",X"22",X"BD",X"7B",X"06",X"1F",X"A8",X"85",X"40",X"26",X"03",X"7E",
		X"F8",X"F1",X"10",X"8E",X"D2",X"00",X"20",X"00",X"86",X"20",X"8E",X"58",X"00",X"30",X"1F",X"C6",
		X"39",X"F7",X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",X"EE",X"6E",X"A4",X"1F",X"03",
		X"86",X"02",X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"F1",X"ED",X"7E",X"F2",X"68",X"86",X"02",X"10",
		X"8E",X"F1",X"F5",X"20",X"D5",X"10",X"8E",X"F1",X"FB",X"20",X"5D",X"86",X"01",X"10",X"8E",X"F2",
		X"03",X"20",X"C7",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",X"8E",X"F2",X"11",X"20",
		X"57",X"86",X"02",X"10",X"8E",X"F2",X"19",X"20",X"B1",X"10",X"8E",X"F2",X"1F",X"20",X"39",X"86",
		X"01",X"10",X"8E",X"F2",X"27",X"20",X"A3",X"1F",X"30",X"1F",X"98",X"10",X"8E",X"F2",X"31",X"20",
		X"37",X"86",X"02",X"10",X"8E",X"F2",X"39",X"20",X"91",X"10",X"8E",X"F2",X"3F",X"20",X"19",X"86",
		X"05",X"10",X"8E",X"F2",X"47",X"20",X"83",X"1F",X"B8",X"4A",X"1F",X"8B",X"26",X"96",X"10",X"8E",
		X"F2",X"54",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",
		X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",X"46",X"46",X"46",X"84",X"C0",X"B7",
		X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0F",X"86",X"34",X"C5",
		X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",X"1A",X"3F",X"8E",X"F3",X"1C",X"8C",
		X"F3",X"3C",X"26",X"02",X"6E",X"A4",X"A6",X"01",X"27",X"18",X"A6",X"84",X"5F",X"1F",X"03",X"86",
		X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",X"1E",X"03",X"26",X"F3",X"E1",X"01",
		X"26",X"04",X"30",X"02",X"20",X"D9",X"A6",X"84",X"44",X"44",X"44",X"44",X"81",X"0D",X"25",X"02",
		X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",X"CE",X"F2",X"D0",X"7E",X"F1",X"DE",
		X"86",X"BF",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"BF",X"00",X"BD",X"D2",X"1E",
		X"1F",X"A8",X"43",X"F7",X"BF",X"06",X"85",X"C0",X"26",X"0A",X"86",X"05",X"8E",X"30",X"70",X"C6",
		X"22",X"BD",X"7B",X"03",X"86",X"08",X"8E",X"40",X"90",X"C6",X"22",X"BD",X"7B",X"03",X"B6",X"BF",
		X"06",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"C6",X"22",X"BD",X"7B",X"06",X"1F",X"A9",X"C5",X"40",
		X"26",X"03",X"7E",X"F8",X"F6",X"10",X"8E",X"D2",X"00",X"7E",X"F1",X"C8",X"00",X"22",X"10",X"98",
		X"20",X"FB",X"30",X"AA",X"40",X"99",X"50",X"19",X"60",X"04",X"70",X"70",X"80",X"5A",X"90",X"00",
		X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",X"D9",X"E0",X"8F",X"F0",X"77",X"00",X"F8",X"10",X"CE",
		X"BF",X"00",X"86",X"04",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",
		X"86",X"FF",X"B7",X"BF",X"09",X"BD",X"F4",X"5E",X"B6",X"C8",X"0C",X"46",X"10",X"25",X"06",X"0F",
		X"BD",X"D2",X"1E",X"1A",X"BF",X"10",X"8E",X"F3",X"6C",X"7E",X"F2",X"58",X"86",X"39",X"B7",X"CB",
		X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"10",X"8E",X"F3",X"7F",X"7E",X"F2",X"8A",X"86",
		X"BF",X"1F",X"8B",X"BD",X"D2",X"1E",X"86",X"00",X"BD",X"7B",X"12",X"C6",X"03",X"8E",X"70",X"00",
		X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"16",X"30",X"1F",X"8C",X"00",
		X"00",X"26",X"ED",X"5A",X"26",X"E7",X"10",X"8E",X"F3",X"B2",X"8E",X"00",X"00",X"86",X"FF",X"7E",
		X"F0",X"9C",X"86",X"01",X"B7",X"C9",X"00",X"86",X"BF",X"1F",X"8B",X"BD",X"D2",X"1E",X"86",X"01",
		X"BD",X"7B",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"8E",
		X"9C",X"00",X"6F",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",X"01",X"26",X"F4",X"CC",X"A5",
		X"5A",X"FD",X"BF",X"0B",X"B7",X"BF",X"09",X"8D",X"68",X"BD",X"F9",X"2F",X"BD",X"FE",X"BA",X"86",
		X"02",X"24",X"24",X"C6",X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",X"10",X"CE",X"F4",X"05",
		X"86",X"03",X"7E",X"F1",X"DE",X"10",X"CE",X"BF",X"00",X"8D",X"46",X"86",X"BF",X"1F",X"8B",X"86",
		X"03",X"C1",X"1F",X"22",X"02",X"86",X"04",X"BD",X"D2",X"1E",X"BD",X"7B",X"12",X"BD",X"F9",X"2F",
		X"7F",X"BF",X"08",X"BD",X"FE",X"3A",X"BD",X"FE",X"44",X"BD",X"F9",X"52",X"24",X"F8",X"86",X"3F",
		X"B7",X"C8",X"0E",X"4F",X"BD",X"F9",X"5F",X"4F",X"B7",X"C8",X"0E",X"BD",X"F9",X"2F",X"BD",X"F7",
		X"80",X"BD",X"F9",X"2F",X"BD",X"F6",X"E4",X"BD",X"F9",X"52",X"24",X"03",X"BD",X"F9",X"2F",X"20",
		X"75",X"7F",X"C8",X"0E",X"86",X"34",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"39",X"8E",X"F0",
		X"0F",X"10",X"8E",X"C0",X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"1F",X"25",X"F7",X"39",X"86",
		X"3C",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",X"3F",X"1F",
		X"8A",X"86",X"8F",X"BE",X"C5",X"01",X"30",X"89",X"12",X"34",X"10",X"8E",X"F4",X"91",X"7E",X"F0",
		X"9C",X"10",X"8E",X"F4",X"98",X"7E",X"F2",X"8A",X"86",X"BF",X"1F",X"8B",X"10",X"CE",X"BF",X"00",
		X"BD",X"FE",X"BA",X"24",X"16",X"86",X"04",X"8C",X"CD",X"00",X"23",X"02",X"86",X"03",X"BD",X"D2",
		X"1E",X"BD",X"7B",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"F9",X"8D",X"31",X"10",X"8E",X"F4",
		X"6F",X"86",X"04",X"7E",X"F1",X"CA",X"8D",X"78",X"BD",X"F9",X"2F",X"BD",X"D2",X"1E",X"86",X"07",
		X"B7",X"C0",X"00",X"BD",X"F9",X"2F",X"86",X"38",X"B7",X"C0",X"00",X"BD",X"F9",X"2F",X"86",X"C0",
		X"B7",X"C0",X"00",X"BD",X"F9",X"2F",X"8D",X"06",X"BD",X"F9",X"2F",X"7E",X"F9",X"6F",X"8E",X"C0",
		X"00",X"10",X"8E",X"F5",X"30",X"EC",X"A1",X"ED",X"81",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"C0",
		X"10",X"25",X"F2",X"CC",X"00",X"00",X"8E",X"00",X"00",X"BF",X"BF",X"06",X"30",X"89",X"0F",X"00",
		X"ED",X"83",X"34",X"02",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"02",X"BC",X"BF",X"06",X"26",X"F0",
		X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",X"DA",X"39",
		X"05",X"05",X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",
		X"BD",X"D2",X"1E",X"4F",X"BD",X"F7",X"75",X"7F",X"C9",X"00",X"86",X"FF",X"B7",X"C0",X"01",X"86",
		X"C0",X"B7",X"C0",X"02",X"86",X"38",X"B7",X"C0",X"03",X"86",X"07",X"B7",X"C0",X"04",X"10",X"8E",
		X"F6",X"6C",X"CC",X"01",X"01",X"AE",X"A4",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"01",X"ED",X"81",
		X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"F6",X"94",X"26",X"E9",X"86",X"11",X"10",X"8E",
		X"F6",X"4C",X"AE",X"A4",X"BF",X"BF",X"06",X"A7",X"84",X"7C",X"BF",X"06",X"C6",X"39",X"F7",X"CB",
		X"FF",X"BE",X"BF",X"06",X"AC",X"22",X"26",X"EF",X"31",X"24",X"10",X"8C",X"F6",X"6C",X"26",X"E2",
		X"10",X"8E",X"F6",X"94",X"AE",X"A4",X"BF",X"BF",X"06",X"A6",X"24",X"A7",X"84",X"7C",X"BF",X"06",
		X"C6",X"39",X"F7",X"CB",X"FF",X"BE",X"BF",X"06",X"AC",X"22",X"26",X"EF",X"31",X"25",X"10",X"8C",
		X"F6",X"D0",X"26",X"E0",X"10",X"8E",X"F6",X"D0",X"AE",X"A4",X"A6",X"24",X"A7",X"80",X"C6",X"39",
		X"F7",X"CB",X"FF",X"AC",X"22",X"26",X"F5",X"31",X"25",X"10",X"8C",X"F6",X"E4",X"26",X"E9",X"86",
		X"21",X"B7",X"43",X"7E",X"86",X"20",X"B7",X"93",X"7E",X"8E",X"4B",X"0A",X"A6",X"84",X"84",X"F0",
		X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",X"6D",X"26",X"EE",X"8E",X"4B",
		X"90",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",
		X"F3",X"26",X"EE",X"8E",X"0B",X"18",X"BF",X"BF",X"06",X"BE",X"BF",X"06",X"A6",X"84",X"84",X"F0",
		X"8A",X"01",X"A7",X"84",X"F6",X"BF",X"07",X"CB",X"22",X"25",X"05",X"F7",X"BF",X"07",X"20",X"E9",
		X"C6",X"18",X"F7",X"BF",X"07",X"F6",X"BF",X"06",X"CB",X"10",X"F7",X"BF",X"06",X"C1",X"9B",X"26",
		X"D8",X"C6",X"01",X"F7",X"C9",X"00",X"C6",X"39",X"F7",X"CB",X"FF",X"39",X"04",X"07",X"94",X"07",
		X"04",X"29",X"94",X"29",X"04",X"4B",X"94",X"4B",X"04",X"6D",X"94",X"6D",X"04",X"8F",X"94",X"8F",
		X"04",X"B1",X"94",X"B1",X"04",X"D3",X"94",X"D3",X"04",X"F5",X"94",X"F5",X"03",X"07",X"03",X"F5",
		X"13",X"07",X"13",X"F5",X"23",X"07",X"23",X"F5",X"33",X"07",X"33",X"F5",X"43",X"07",X"43",X"F5",
		X"53",X"07",X"53",X"F5",X"63",X"07",X"63",X"F5",X"73",X"07",X"73",X"F5",X"83",X"07",X"83",X"F5",
		X"93",X"07",X"93",X"F5",X"45",X"05",X"52",X"05",X"44",X"45",X"06",X"52",X"06",X"44",X"45",X"07",
		X"52",X"07",X"00",X"45",X"08",X"52",X"08",X"33",X"45",X"09",X"52",X"09",X"33",X"45",X"F3",X"52",
		X"F3",X"33",X"45",X"F4",X"52",X"F4",X"33",X"45",X"F5",X"52",X"F5",X"00",X"45",X"F6",X"52",X"F6",
		X"44",X"45",X"F7",X"52",X"F7",X"44",X"04",X"7E",X"43",X"7E",X"22",X"54",X"7E",X"93",X"7E",X"22",
		X"02",X"6F",X"02",X"8E",X"04",X"03",X"6F",X"03",X"8E",X"30",X"93",X"6F",X"93",X"8E",X"00",X"94",
		X"6F",X"94",X"8E",X"34",X"BD",X"D2",X"1E",X"86",X"05",X"BD",X"7B",X"12",X"86",X"80",X"B7",X"BF",
		X"28",X"4F",X"BD",X"F9",X"5F",X"BD",X"F9",X"52",X"25",X"33",X"7A",X"BF",X"28",X"26",X"F2",X"B6",
		X"F7",X"5D",X"8D",X"71",X"8D",X"28",X"8E",X"F7",X"5D",X"A6",X"80",X"BF",X"BF",X"06",X"8D",X"65",
		X"86",X"80",X"B7",X"BF",X"28",X"4F",X"BD",X"F9",X"5F",X"BD",X"F9",X"52",X"25",X"0F",X"7A",X"BF",
		X"28",X"26",X"F2",X"BE",X"BF",X"06",X"8C",X"F7",X"65",X"25",X"DE",X"20",X"D9",X"39",X"8E",X"00",
		X"00",X"10",X"8E",X"F7",X"65",X"BF",X"BF",X"06",X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",
		X"ED",X"83",X"C6",X"39",X"F7",X"CB",X"FF",X"BC",X"BF",X"06",X"26",X"F2",X"30",X"89",X"09",X"00",
		X"4D",X"26",X"03",X"8E",X"0D",X"00",X"10",X"8C",X"F7",X"75",X"26",X"D9",X"39",X"02",X"03",X"04",
		X"10",X"18",X"20",X"40",X"80",X"00",X"FF",X"11",X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",
		X"AA",X"66",X"99",X"77",X"88",X"8E",X"C0",X"00",X"A7",X"80",X"8C",X"C0",X"10",X"25",X"F9",X"39",
		X"86",X"0A",X"B7",X"BF",X"06",X"BD",X"D2",X"1E",X"86",X"06",X"BD",X"7B",X"12",X"C6",X"39",X"F7",
		X"CB",X"FF",X"CE",X"BF",X"28",X"6F",X"C0",X"11",X"83",X"BF",X"31",X"23",X"F8",X"CE",X"F8",X"61",
		X"8D",X"29",X"86",X"34",X"B7",X"C8",X"07",X"C6",X"39",X"F7",X"CB",X"FF",X"8D",X"1D",X"86",X"3C",
		X"B7",X"C8",X"07",X"8D",X"26",X"BD",X"F9",X"52",X"24",X"0A",X"C6",X"39",X"F7",X"CB",X"FF",X"7A",
		X"BF",X"06",X"27",X"06",X"4F",X"BD",X"F9",X"5F",X"20",X"D3",X"39",X"AE",X"C1",X"27",X"0B",X"10",
		X"AE",X"C1",X"A6",X"84",X"A8",X"A4",X"A7",X"21",X"20",X"F1",X"39",X"CE",X"F8",X"79",X"10",X"8E",
		X"BF",X"28",X"C6",X"01",X"E5",X"21",X"27",X"02",X"8D",X"15",X"33",X"43",X"58",X"24",X"F5",X"C6",
		X"39",X"F7",X"CB",X"FF",X"31",X"22",X"10",X"8C",X"BF",X"31",X"22",X"02",X"20",X"E4",X"39",X"34",
		X"14",X"86",X"3F",X"B7",X"C8",X"0E",X"E8",X"A4",X"E7",X"A4",X"E6",X"E4",X"E5",X"A4",X"26",X"2A",
		X"E6",X"42",X"27",X"4B",X"86",X"40",X"1F",X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"CC",X"44",X"02",
		X"FD",X"CA",X"06",X"BF",X"CA",X"04",X"BF",X"CA",X"04",X"C6",X"00",X"F7",X"CA",X"01",X"C6",X"12",
		X"F7",X"CA",X"00",X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"94",X"E6",X"42",X"27",X"21",X"86",X"40",
		X"1F",X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"A6",X"C4",X"BD",X"7B",X"0C",X"A6",X"41",
		X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"BD",X"7B",X"0F",X"86",X"3C",X"B7",X"C8",X"0E",X"35",
		X"94",X"C8",X"0C",X"BF",X"28",X"C8",X"04",X"BF",X"2A",X"C8",X"06",X"BF",X"2C",X"00",X"00",X"C8",
		X"04",X"BF",X"2E",X"C8",X"06",X"BF",X"30",X"00",X"00",X"16",X"FF",X"2C",X"17",X"FF",X"33",X"18",
		X"FF",X"3A",X"19",X"FF",X"41",X"1A",X"FF",X"48",X"1B",X"FF",X"4F",X"1C",X"FF",X"56",X"00",X"00",
		X"00",X"21",X"F1",X"5D",X"6D",X"F1",X"64",X"1F",X"F1",X"6B",X"20",X"F1",X"72",X"1E",X"FF",X"79",
		X"1D",X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"21",X"F2",X"87",X"6D",X"F2",X"8E",X"1F",X"F2",X"95",X"20",X"F2",X"9C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CE",X"F3",X"CF",X"20",X"03",X"CE",X"F3",X"A6",X"10",X"CE",X"BF",X"00",X"10",X"8E",X"F9",
		X"06",X"86",X"01",X"7E",X"F1",X"CA",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"10",X"8E",X"F9",
		X"16",X"86",X"01",X"7E",X"F1",X"CA",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F0",X"10",X"8E",X"F9",
		X"26",X"86",X"01",X"7E",X"F1",X"CA",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"6E",X"C4",X"B6",
		X"C8",X"0C",X"85",X"02",X"26",X"06",X"86",X"01",X"8D",X"25",X"20",X"F3",X"7F",X"C0",X"00",X"BD",
		X"D2",X"1E",X"20",X"07",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"06",X"86",X"01",X"8D",X"10",X"20",
		X"F3",X"39",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"03",X"1A",X"01",X"39",X"1C",X"FE",X"39",X"C6",
		X"39",X"8E",X"03",X"00",X"F7",X"CB",X"FF",X"30",X"1F",X"26",X"F9",X"4A",X"2A",X"F1",X"39",X"86",
		X"BF",X"1F",X"8B",X"BD",X"F4",X"5E",X"8D",X"DA",X"24",X"02",X"8D",X"B3",X"86",X"07",X"BD",X"7B",
		X"12",X"CE",X"CD",X"02",X"8E",X"1A",X"30",X"86",X"24",X"34",X"12",X"C6",X"88",X"BD",X"7B",X"03",
		X"1E",X"31",X"BD",X"D2",X"24",X"C5",X"F0",X"26",X"08",X"CA",X"F0",X"C5",X"0F",X"26",X"02",X"CA",
		X"0F",X"1F",X"98",X"43",X"34",X"06",X"BD",X"D2",X"27",X"6D",X"E0",X"26",X"12",X"85",X"F0",X"26",
		X"0E",X"8A",X"F0",X"85",X"0F",X"26",X"08",X"8A",X"0F",X"C5",X"F0",X"26",X"02",X"CA",X"F0",X"1F",
		X"02",X"1E",X"31",X"1F",X"10",X"86",X"6A",X"1F",X"01",X"35",X"02",X"C6",X"88",X"BD",X"7B",X"06",
		X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"20",X"34",X"04",X"C6",X"88",X"BD",X"7B",X"06",X"35",X"02",
		X"BD",X"7B",X"06",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"12",X"30",X"88",X"10",X"4C",X"11",X"83",
		X"CD",X"38",X"23",X"95",X"86",X"2E",X"C6",X"88",X"BD",X"7B",X"03",X"1F",X"10",X"86",X"6E",X"1F",
		X"01",X"1E",X"31",X"8E",X"CD",X"20",X"BD",X"D2",X"24",X"F7",X"BF",X"10",X"BD",X"D2",X"27",X"FD",
		X"BF",X"11",X"8E",X"CD",X"38",X"BD",X"D2",X"24",X"F7",X"BF",X"13",X"BD",X"D2",X"27",X"FD",X"BF",
		X"14",X"1E",X"31",X"8D",X"21",X"C6",X"88",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",X"7B",X"06",
		X"86",X"32",X"BD",X"7B",X"00",X"B6",X"BF",X"12",X"BD",X"7B",X"06",X"86",X"39",X"B7",X"CB",X"FF",
		X"BD",X"F9",X"2F",X"7E",X"FB",X"47",X"34",X"30",X"8D",X"7A",X"FC",X"BF",X"10",X"27",X"0F",X"86",
		X"99",X"34",X"02",X"B7",X"BF",X"12",X"7F",X"BF",X"11",X"7F",X"BF",X"10",X"20",X"4C",X"B6",X"BF",
		X"12",X"34",X"02",X"FC",X"BF",X"0D",X"FD",X"BF",X"10",X"B6",X"BF",X"0F",X"B7",X"BF",X"12",X"CC",
		X"00",X"00",X"FD",X"BF",X"0D",X"B7",X"BF",X"0F",X"86",X"04",X"78",X"BF",X"12",X"79",X"BF",X"11",
		X"79",X"BF",X"10",X"79",X"BF",X"0F",X"4A",X"26",X"F1",X"8E",X"BF",X"13",X"10",X"8E",X"BF",X"13",
		X"CE",X"BF",X"13",X"8D",X"17",X"FC",X"BF",X"0F",X"FD",X"BF",X"16",X"FC",X"BF",X"11",X"FD",X"BF",
		X"18",X"8E",X"BF",X"1A",X"8D",X"06",X"8D",X"04",X"8D",X"23",X"35",X"B2",X"34",X"70",X"C6",X"04",
		X"20",X"04",X"34",X"70",X"C6",X"03",X"1C",X"FE",X"A6",X"82",X"A9",X"A2",X"19",X"A7",X"C2",X"5A",
		X"26",X"F6",X"35",X"F0",X"CC",X"00",X"00",X"FD",X"BF",X"0D",X"B7",X"BF",X"0F",X"FC",X"BF",X"13",
		X"26",X"0F",X"B6",X"BF",X"15",X"26",X"0A",X"CC",X"00",X"00",X"FD",X"BF",X"10",X"B7",X"BF",X"12",
		X"39",X"86",X"07",X"B7",X"BF",X"16",X"8E",X"BF",X"10",X"10",X"8E",X"BF",X"16",X"CE",X"BF",X"1A",
		X"8D",X"35",X"7A",X"BF",X"16",X"26",X"02",X"20",X"2E",X"86",X"04",X"78",X"BF",X"12",X"79",X"BF",
		X"11",X"79",X"BF",X"10",X"79",X"BF",X"0F",X"79",X"BF",X"0E",X"79",X"BF",X"0D",X"4A",X"26",X"EB",
		X"8D",X"A0",X"25",X"02",X"20",X"DC",X"FC",X"BF",X"17",X"FD",X"BF",X"0D",X"B6",X"BF",X"19",X"B7",
		X"BF",X"0F",X"7C",X"BF",X"12",X"20",X"E9",X"34",X"20",X"C6",X"03",X"86",X"99",X"A0",X"A2",X"A7",
		X"A4",X"5A",X"26",X"F7",X"10",X"AE",X"E4",X"C6",X"03",X"1A",X"01",X"A6",X"3F",X"89",X"00",X"19",
		X"A7",X"A2",X"5A",X"26",X"F6",X"35",X"A0",X"8E",X"CC",X"18",X"6F",X"80",X"8C",X"CC",X"24",X"25",
		X"F9",X"BD",X"D2",X"1E",X"BD",X"F9",X"52",X"24",X"03",X"BD",X"F9",X"2F",X"86",X"08",X"BD",X"7B",
		X"12",X"CE",X"CC",X"00",X"8E",X"1A",X"20",X"86",X"30",X"34",X"12",X"C6",X"22",X"BD",X"7B",X"0C",
		X"F7",X"BF",X"1A",X"F7",X"BF",X"0D",X"1F",X"12",X"BD",X"FD",X"1B",X"33",X"42",X"C6",X"39",X"F7",
		X"CB",X"FF",X"35",X"12",X"30",X"0A",X"4C",X"11",X"83",X"CC",X"24",X"2D",X"DC",X"86",X"09",X"BD",
		X"7B",X"15",X"7F",X"BF",X"0D",X"B6",X"CC",X"07",X"84",X"0F",X"81",X"09",X"26",X"0B",X"86",X"5D",
		X"F6",X"BF",X"1A",X"8E",X"70",X"3E",X"BD",X"7B",X"0C",X"10",X"8E",X"16",X"20",X"CE",X"CC",X"00",
		X"1F",X"21",X"86",X"30",X"C6",X"33",X"FD",X"BF",X"28",X"BD",X"7B",X"09",X"86",X"39",X"B7",X"CB",
		X"FF",X"B6",X"C8",X"04",X"84",X"03",X"27",X"02",X"8D",X"1A",X"B6",X"C8",X"04",X"84",X"30",X"27",
		X"03",X"BD",X"FC",X"77",X"C6",X"3C",X"F7",X"C8",X"07",X"BD",X"F9",X"52",X"24",X"DE",X"BD",X"F9",
		X"2F",X"7E",X"D2",X"09",X"B7",X"BF",X"2C",X"B1",X"BF",X"2A",X"27",X"15",X"7F",X"BF",X"2B",X"B6",
		X"BF",X"2C",X"B7",X"BF",X"2A",X"86",X"02",X"BD",X"F9",X"5F",X"B6",X"C8",X"04",X"84",X"03",X"26",
		X"1D",X"C6",X"05",X"F7",X"BF",X"2D",X"B6",X"C8",X"04",X"84",X"03",X"26",X"04",X"7F",X"BF",X"2A",
		X"39",X"86",X"02",X"BD",X"F9",X"5F",X"7A",X"BF",X"2D",X"26",X"EB",X"B6",X"C8",X"04",X"85",X"02",
		X"26",X"22",X"85",X"01",X"27",X"42",X"10",X"8C",X"16",X"20",X"27",X"3C",X"8D",X"3F",X"31",X"36",
		X"33",X"5E",X"11",X"83",X"CC",X"12",X"26",X"0A",X"7D",X"BF",X"0A",X"27",X"05",X"31",X"A8",X"C4",
		X"33",X"54",X"20",X"1C",X"10",X"8C",X"16",X"CA",X"27",X"1E",X"8D",X"21",X"31",X"2A",X"33",X"42",
		X"11",X"83",X"CC",X"08",X"26",X"0A",X"7D",X"BF",X"0A",X"27",X"05",X"31",X"A8",X"3C",X"33",X"4C",
		X"1F",X"21",X"FC",X"BF",X"28",X"BD",X"7B",X"09",X"4F",X"BD",X"F9",X"5F",X"39",X"1F",X"21",X"B6",
		X"BF",X"28",X"5F",X"BD",X"7B",X"09",X"39",X"B7",X"BF",X"2C",X"B1",X"BF",X"2E",X"27",X"15",X"7F",
		X"BF",X"2F",X"B6",X"BF",X"2C",X"B7",X"BF",X"2E",X"86",X"02",X"BD",X"F9",X"5F",X"B6",X"C8",X"04",
		X"84",X"30",X"26",X"1E",X"C6",X"08",X"F7",X"BF",X"31",X"B6",X"C8",X"04",X"84",X"30",X"26",X"04",
		X"7F",X"BF",X"2F",X"39",X"4F",X"BD",X"F9",X"5F",X"7A",X"BF",X"31",X"26",X"EC",X"B6",X"C8",X"04",
		X"84",X"30",X"34",X"02",X"1F",X"31",X"BD",X"D2",X"21",X"34",X"02",X"5F",X"F7",X"BF",X"1A",X"8D",
		X"5A",X"C6",X"39",X"F7",X"CB",X"FF",X"8E",X"FC",X"F7",X"1F",X"30",X"30",X"85",X"35",X"06",X"C5",
		X"10",X"26",X"0C",X"C5",X"20",X"27",X"14",X"A1",X"84",X"27",X"10",X"8B",X"99",X"20",X"06",X"A1",
		X"01",X"27",X"08",X"8B",X"01",X"19",X"1F",X"31",X"BD",X"D2",X"2A",X"C6",X"22",X"F7",X"BF",X"1A",
		X"BD",X"FD",X"1B",X"4F",X"7E",X"F9",X"5F",X"00",X"99",X"01",X"99",X"00",X"01",X"00",X"09",X"00",
		X"99",X"00",X"99",X"00",X"99",X"01",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"03",X"20",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"1F",X"30",X"54",X"8E",X"FD",
		X"7C",X"30",X"85",X"6D",X"84",X"2B",X"2C",X"1F",X"31",X"BD",X"D2",X"21",X"11",X"83",X"CC",X"06",
		X"26",X"0A",X"B7",X"BF",X"0A",X"7D",X"BF",X"0D",X"26",X"02",X"8D",X"52",X"85",X"F0",X"26",X"02",
		X"8A",X"F0",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"F6",X"BF",X"1A",X"BD",
		X"7B",X"0F",X"39",X"A6",X"84",X"85",X"01",X"26",X"1C",X"1F",X"31",X"BD",X"D2",X"24",X"86",X"0D",
		X"5D",X"27",X"02",X"86",X"44",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"F6",
		X"BF",X"1A",X"7E",X"7B",X"0C",X"8D",X"B0",X"86",X"2F",X"7E",X"7B",X"09",X"81",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"34",X"76",
		X"8E",X"00",X"3C",X"BF",X"CA",X"06",X"8E",X"6A",X"48",X"BF",X"CA",X"04",X"5F",X"F7",X"CA",X"01",
		X"C6",X"12",X"F7",X"CA",X"00",X"8E",X"FD",X"FE",X"81",X"09",X"26",X"0F",X"34",X"12",X"86",X"5D",
		X"F6",X"BF",X"1A",X"8E",X"70",X"3E",X"BD",X"7B",X"0C",X"35",X"12",X"1F",X"89",X"58",X"34",X"04",
		X"58",X"EB",X"E0",X"3A",X"33",X"42",X"1E",X"31",X"8C",X"CC",X"14",X"27",X"2F",X"A6",X"C0",X"BD",
		X"D2",X"2A",X"C6",X"39",X"F7",X"CB",X"FF",X"1E",X"31",X"31",X"2A",X"34",X"10",X"30",X"5E",X"BD",
		X"D2",X"21",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",
		X"35",X"02",X"F6",X"BF",X"1A",X"BD",X"7B",X"0F",X"35",X"10",X"20",X"CA",X"35",X"F6",X"01",X"04",
		X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",X"00",X"00",
		X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",X"01",X"02",
		X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"01",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"D2",X"1E",X"CC",X"FE",X"01",
		X"FD",X"BF",X"29",X"39",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"5F",X"4F",X"B7",
		X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"5F",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",
		X"5F",X"FC",X"BF",X"29",X"84",X"3F",X"B7",X"C8",X"0E",X"C6",X"99",X"8E",X"3A",X"80",X"86",X"22",
		X"BD",X"7B",X"03",X"B6",X"BF",X"2A",X"8A",X"F0",X"C6",X"99",X"BD",X"7B",X"06",X"86",X"40",X"B7",
		X"BF",X"28",X"86",X"01",X"BD",X"F9",X"5F",X"BD",X"F9",X"52",X"25",X"05",X"7A",X"BF",X"28",X"26",
		X"F1",X"B6",X"BF",X"08",X"26",X"06",X"B6",X"C8",X"0C",X"46",X"24",X"1D",X"8E",X"57",X"80",X"B6",
		X"BF",X"2A",X"8A",X"F0",X"C6",X"00",X"BD",X"7B",X"06",X"FC",X"BF",X"29",X"1A",X"01",X"49",X"5C",
		X"C1",X"07",X"25",X"02",X"8D",X"87",X"FD",X"BF",X"29",X"39",X"8E",X"CC",X"00",X"10",X"8E",X"9C",
		X"00",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",X"C6",X"06",X"FE",X"BF",X"0B",X"10",
		X"BE",X"BF",X"0A",X"8E",X"CC",X"00",X"BD",X"FF",X"21",X"A7",X"80",X"86",X"39",X"B7",X"CB",X"FF",
		X"8C",X"D0",X"00",X"26",X"F1",X"10",X"BF",X"BF",X"0A",X"FF",X"BF",X"0B",X"8E",X"CC",X"00",X"BD",
		X"FF",X"21",X"A8",X"80",X"84",X"0F",X"26",X"24",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",X"00",
		X"26",X"ED",X"5A",X"26",X"C7",X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"9C",X"00",X"10",X"8E",X"CC",
		X"00",X"A6",X"C0",X"A7",X"A0",X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",X"8D",X"EC",X"1A",X"01",
		X"39",X"34",X"04",X"F6",X"BF",X"0A",X"86",X"03",X"3D",X"CB",X"11",X"B6",X"BF",X"0C",X"44",X"44",
		X"44",X"B8",X"BF",X"0C",X"44",X"76",X"BF",X"0B",X"76",X"BF",X"0C",X"FB",X"BF",X"0C",X"F9",X"BF",
		X"0B",X"F7",X"BF",X"0A",X"B6",X"BF",X"0A",X"35",X"84",X"20",X"42",X"55",X"42",X"42",X"4C",X"45",
		X"53",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"28",
		X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",
		X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",
		X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",
		X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"6E",X"9F",X"EF",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"97",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"7E",X"00",X"89",X"7E",X"00",X"AD",X"7E",X"00",X"EE",X"7E",X"00",X"5C",X"7E",X"01",X"13",X"7E",
		X"07",X"1B",X"7E",X"12",X"E8",X"7E",X"01",X"63",X"7E",X"37",X"25",X"7E",X"01",X"AB",X"7E",X"3A",
		X"69",X"7E",X"23",X"0B",X"7E",X"05",X"0F",X"7E",X"13",X"C0",X"7E",X"38",X"2A",X"34",X"51",X"AE",
		X"22",X"EE",X"A4",X"EF",X"84",X"AF",X"42",X"1F",X"03",X"AE",X"42",X"10",X"AF",X"84",X"AF",X"22",
		X"EF",X"A4",X"10",X"AF",X"42",X"35",X"D1",X"34",X"51",X"1A",X"50",X"AE",X"A4",X"EE",X"22",X"AF",
		X"C4",X"EF",X"02",X"35",X"D1",X"10",X"9E",X"08",X"20",X"09",X"86",X"FF",X"9B",X"04",X"10",X"9E",
		X"08",X"A7",X"24",X"10",X"EF",X"27",X"1A",X"50",X"10",X"AE",X"A4",X"10",X"9F",X"08",X"1C",X"EF",
		X"EC",X"24",X"91",X"04",X"2A",X"F0",X"10",X"EE",X"27",X"C5",X"01",X"27",X"04",X"C5",X"02",X"27",
		X"01",X"39",X"C4",X"FE",X"E7",X"25",X"AD",X"B8",X"09",X"10",X"9E",X"08",X"BD",X"00",X"47",X"30",
		X"A4",X"BD",X"01",X"AB",X"20",X"D2",X"35",X"40",X"A6",X"C0",X"34",X"42",X"BD",X"00",X"5A",X"6A",
		X"E4",X"26",X"F9",X"35",X"82",X"34",X"57",X"EE",X"67",X"37",X"20",X"20",X"08",X"34",X"57",X"EE",
		X"67",X"10",X"8E",X"00",X"8C",X"37",X"04",X"4F",X"BD",X"01",X"63",X"10",X"AF",X"09",X"34",X"10",
		X"AF",X"84",X"AF",X"02",X"30",X"8B",X"30",X"1C",X"37",X"24",X"EF",X"69",X"10",X"AF",X"84",X"35",
		X"20",X"AF",X"27",X"ED",X"25",X"96",X"04",X"4A",X"A7",X"24",X"CC",X"9B",X"DC",X"BD",X"00",X"2D",
		X"35",X"D7",X"34",X"03",X"20",X"02",X"8D",X"06",X"A6",X"C0",X"26",X"FA",X"35",X"83",X"34",X"15",
		X"8E",X"9B",X"DC",X"AE",X"84",X"8C",X"9B",X"DC",X"26",X"02",X"35",X"95",X"A1",X"06",X"26",X"F3",
		X"8D",X"02",X"20",X"EF",X"34",X"05",X"E6",X"05",X"CA",X"01",X"E7",X"05",X"D6",X"04",X"5A",X"E7",
		X"04",X"35",X"85",X"8E",X"9B",X"DC",X"AE",X"84",X"8C",X"9B",X"DC",X"26",X"05",X"8E",X"00",X"00",
		X"4D",X"39",X"A1",X"06",X"26",X"F0",X"39",X"34",X"63",X"96",X"04",X"4A",X"A7",X"04",X"10",X"AE",
		X"84",X"EE",X"02",X"10",X"AF",X"C4",X"EF",X"22",X"10",X"9E",X"08",X"EE",X"A4",X"AF",X"42",X"EF",
		X"84",X"AF",X"A4",X"10",X"AF",X"02",X"35",X"E3",X"34",X"77",X"44",X"34",X"02",X"24",X"05",X"86",
		X"3B",X"BD",X"00",X"5C",X"6A",X"E4",X"2B",X"07",X"86",X"77",X"BD",X"00",X"5C",X"20",X"F5",X"32",
		X"61",X"35",X"F7",X"34",X"06",X"8E",X"A5",X"71",X"EC",X"84",X"2B",X"09",X"27",X"04",X"30",X"8B",
		X"20",X"F6",X"BD",X"01",X"C1",X"88",X"80",X"6D",X"8B",X"2A",X"06",X"E3",X"8B",X"8B",X"80",X"20",
		X"F6",X"10",X"A3",X"E4",X"24",X"08",X"88",X"80",X"ED",X"84",X"88",X"80",X"20",X"E0",X"A3",X"E4",
		X"10",X"83",X"00",X"14",X"2C",X"06",X"E3",X"E4",X"ED",X"81",X"35",X"86",X"88",X"80",X"ED",X"84",
		X"88",X"80",X"30",X"8B",X"35",X"06",X"ED",X"81",X"39",X"30",X"A4",X"34",X"03",X"A6",X"1E",X"8A",
		X"80",X"A7",X"1E",X"35",X"83",X"34",X"07",X"1A",X"50",X"DC",X"0C",X"ED",X"C4",X"DF",X"0C",X"35",
		X"87",X"3F",X"39",X"34",X"57",X"EE",X"67",X"37",X"04",X"4F",X"BD",X"01",X"63",X"31",X"84",X"37",
		X"16",X"EF",X"67",X"33",X"A6",X"86",X"04",X"1A",X"50",X"FF",X"CA",X"04",X"BF",X"CA",X"02",X"FD",
		X"CA",X"06",X"7F",X"CA",X"00",X"35",X"D7",X"10",X"DF",X"20",X"F6",X"C8",X"0E",X"4F",X"F6",X"CB",
		X"00",X"58",X"49",X"58",X"49",X"48",X"26",X"23",X"DC",X"03",X"C3",X"00",X"01",X"DD",X"03",X"F6",
		X"CB",X"00",X"C4",X"FC",X"26",X"14",X"CE",X"99",X"F9",X"37",X"76",X"CE",X"C0",X"10",X"36",X"76",
		X"CE",X"99",X"F1",X"37",X"76",X"CE",X"C0",X"08",X"36",X"76",X"4F",X"8E",X"02",X"2E",X"D6",X"96",
		X"27",X"02",X"88",X"06",X"4D",X"26",X"03",X"8E",X"98",X"0A",X"10",X"CE",X"99",X"E2",X"6E",X"96",
		X"05",X"D8",X"05",X"FB",X"06",X"BF",X"BD",X"15",X"B9",X"BD",X"01",X"48",X"AD",X"B8",X"0B",X"86",
		X"1E",X"BD",X"00",X"5C",X"CE",X"39",X"97",X"BD",X"08",X"38",X"7E",X"00",X"89",X"34",X"07",X"6F",
		X"E2",X"1A",X"50",X"F6",X"BF",X"FF",X"B6",X"C8",X"06",X"2A",X"0C",X"96",X"01",X"27",X"08",X"6C",
		X"E4",X"CA",X"02",X"86",X"34",X"20",X"04",X"C4",X"FD",X"86",X"3C",X"B7",X"C8",X"07",X"35",X"02",
		X"91",X"96",X"27",X"0D",X"97",X"96",X"F7",X"BF",X"FF",X"F7",X"C9",X"00",X"1C",X"EF",X"BD",X"38",
		X"2A",X"35",X"87",X"0D",X"22",X"26",X"02",X"D7",X"22",X"39",X"B6",X"C8",X"04",X"44",X"D6",X"25",
		X"2B",X"0F",X"24",X"14",X"5C",X"C1",X"03",X"2D",X"10",X"C6",X"03",X"8D",X"E6",X"C6",X"FF",X"20",
		X"08",X"25",X"FA",X"5A",X"C1",X"FC",X"2E",X"01",X"5F",X"D7",X"25",X"44",X"D6",X"26",X"2B",X"0F",
		X"24",X"14",X"5C",X"C1",X"03",X"2D",X"10",X"C6",X"04",X"8D",X"C8",X"C6",X"FF",X"20",X"08",X"25",
		X"FA",X"5A",X"C1",X"FC",X"2E",X"01",X"5F",X"D7",X"26",X"44",X"44",X"44",X"D6",X"24",X"2B",X"0F",
		X"24",X"14",X"5C",X"C1",X"03",X"2D",X"10",X"C6",X"02",X"8D",X"A8",X"C6",X"FF",X"20",X"08",X"25",
		X"FA",X"5A",X"C1",X"FC",X"2E",X"01",X"5F",X"D7",X"24",X"44",X"D6",X"23",X"2B",X"0F",X"24",X"14",
		X"5C",X"C1",X"03",X"2D",X"10",X"C6",X"01",X"8D",X"8A",X"C6",X"FF",X"20",X"08",X"25",X"FA",X"5A",
		X"C1",X"FC",X"2E",X"01",X"5F",X"D7",X"23",X"7E",X"D0",X"1C",X"B6",X"C8",X"04",X"44",X"24",X"0B",
		X"D6",X"4E",X"5C",X"C1",X"03",X"2D",X"05",X"C6",X"EC",X"D7",X"4D",X"5F",X"D7",X"4E",X"44",X"24",
		X"0B",X"D6",X"4F",X"5C",X"C1",X"03",X"2D",X"05",X"C6",X"14",X"D7",X"4D",X"5F",X"D7",X"4F",X"44",
		X"24",X"0B",X"D6",X"50",X"5C",X"C1",X"03",X"2D",X"05",X"C6",X"EC",X"D7",X"4C",X"5F",X"D7",X"50",
		X"44",X"24",X"0B",X"D6",X"51",X"5C",X"C1",X"03",X"2D",X"05",X"C6",X"14",X"D7",X"4C",X"5F",X"D7",
		X"51",X"7E",X"D0",X"1C",X"96",X"3E",X"2A",X"01",X"40",X"A7",X"E2",X"96",X"40",X"2A",X"01",X"40",
		X"A1",X"E4",X"24",X"02",X"A6",X"E4",X"8B",X"02",X"A7",X"E4",X"DC",X"4C",X"4D",X"27",X"0F",X"5D",
		X"27",X"0C",X"80",X"06",X"2A",X"02",X"8B",X"0C",X"C0",X"06",X"2A",X"02",X"CB",X"0C",X"DD",X"4C",
		X"27",X"2F",X"9E",X"52",X"26",X"44",X"A6",X"E4",X"81",X"04",X"24",X"3E",X"8E",X"02",X"00",X"5D",
		X"2E",X"09",X"8E",X"00",X"00",X"5D",X"27",X"03",X"8E",X"FD",X"FF",X"9F",X"40",X"8E",X"02",X"00",
		X"96",X"4C",X"2E",X"09",X"8E",X"00",X"00",X"4D",X"27",X"03",X"8E",X"FD",X"FF",X"9F",X"3E",X"20",
		X"19",X"9E",X"52",X"27",X"15",X"A6",X"E4",X"8B",X"06",X"81",X"10",X"24",X"0D",X"BD",X"1F",X"69",
		X"A7",X"E2",X"1D",X"DD",X"40",X"E6",X"E0",X"1D",X"DD",X"3E",X"DC",X"4C",X"5D",X"27",X"13",X"D8",
		X"40",X"57",X"59",X"D8",X"40",X"24",X"0B",X"86",X"F0",X"58",X"58",X"3D",X"2A",X"02",X"80",X"F0",
		X"1F",X"89",X"86",X"11",X"5D",X"3D",X"2A",X"02",X"80",X"11",X"D3",X"40",X"DD",X"40",X"A6",X"E4",
		X"81",X"04",X"25",X"16",X"96",X"40",X"43",X"50",X"82",X"FF",X"47",X"56",X"47",X"56",X"47",X"56",
		X"47",X"56",X"47",X"56",X"47",X"56",X"D3",X"40",X"DD",X"40",X"D6",X"4C",X"27",X"13",X"D8",X"3E",
		X"57",X"59",X"D8",X"3E",X"24",X"0B",X"86",X"F0",X"58",X"58",X"3D",X"2A",X"02",X"80",X"F0",X"1F",
		X"89",X"86",X"11",X"5D",X"3D",X"2A",X"02",X"80",X"11",X"D3",X"3E",X"DD",X"3E",X"A6",X"E4",X"81",
		X"04",X"25",X"16",X"96",X"3E",X"43",X"50",X"82",X"FF",X"47",X"56",X"47",X"56",X"47",X"56",X"47",
		X"56",X"47",X"56",X"47",X"56",X"D3",X"3E",X"DD",X"3E",X"9E",X"4C",X"9F",X"52",X"8E",X"00",X"00",
		X"96",X"00",X"2A",X"02",X"9F",X"4C",X"A6",X"E4",X"81",X"04",X"24",X"04",X"4F",X"5F",X"20",X"0C",
		X"0F",X"54",X"DC",X"40",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"D3",X"3C",X"81",X"3F",
		X"22",X"0A",X"96",X"40",X"2A",X"02",X"9F",X"40",X"86",X"3F",X"0C",X"54",X"9B",X"45",X"25",X"04",
		X"81",X"EA",X"25",X"0A",X"96",X"40",X"2B",X"02",X"9F",X"40",X"86",X"EA",X"0C",X"54",X"97",X"39",
		X"90",X"45",X"97",X"37",X"DD",X"3C",X"A6",X"E4",X"81",X"04",X"24",X"04",X"4F",X"5F",X"20",X"0A",
		X"DC",X"3E",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"D3",X"3A",X"D7",X"3B",X"D6",X"36",
		X"C1",X"08",X"22",X"0E",X"4D",X"2E",X"12",X"4F",X"0C",X"54",X"D6",X"3E",X"2A",X"0B",X"9F",X"3E",
		X"20",X"07",X"C1",X"F6",X"25",X"03",X"4D",X"2A",X"08",X"9B",X"44",X"25",X"04",X"81",X"FE",X"25",
		X"0A",X"86",X"FE",X"0C",X"54",X"D6",X"3E",X"2B",X"02",X"9F",X"3E",X"97",X"38",X"90",X"44",X"97",
		X"36",X"97",X"3A",X"BD",X"23",X"0B",X"8D",X"27",X"D6",X"1C",X"D7",X"1A",X"10",X"CE",X"9A",X"13",
		X"B6",X"9A",X"0F",X"32",X"E6",X"86",X"18",X"B7",X"9A",X"0F",X"11",X"8C",X"9A",X"2B",X"10",X"2C",
		X"CB",X"1A",X"35",X"36",X"BD",X"0A",X"4E",X"A6",X"2B",X"84",X"7F",X"A7",X"2B",X"20",X"EB",X"34",
		X"57",X"1A",X"50",X"96",X"00",X"85",X"08",X"27",X"5A",X"CE",X"99",X"F1",X"9E",X"42",X"DC",X"5A",
		X"2A",X"07",X"9B",X"36",X"25",X"07",X"4F",X"20",X"04",X"9B",X"36",X"25",X"08",X"AB",X"1C",X"25",
		X"04",X"81",X"FE",X"23",X"02",X"86",X"FE",X"97",X"5E",X"A0",X"1C",X"5D",X"2A",X"0A",X"DB",X"37",
		X"C1",X"3F",X"24",X"02",X"C6",X"3F",X"20",X"02",X"DB",X"37",X"EB",X"1D",X"C1",X"EA",X"23",X"02",
		X"C6",X"EA",X"D7",X"5F",X"E0",X"1D",X"DD",X"5C",X"8B",X"15",X"46",X"FD",X"CA",X"04",X"36",X"06",
		X"BF",X"CA",X"02",X"EC",X"1E",X"FD",X"CA",X"06",X"86",X"0A",X"24",X"02",X"8A",X"20",X"36",X"12",
		X"B7",X"CA",X"00",X"CE",X"99",X"EC",X"DC",X"36",X"D3",X"56",X"8B",X"15",X"46",X"FD",X"CA",X"04",
		X"36",X"06",X"9E",X"46",X"BF",X"CA",X"02",X"EC",X"1E",X"FD",X"CA",X"06",X"86",X"0A",X"24",X"02",
		X"8A",X"20",X"36",X"12",X"B7",X"CA",X"00",X"DC",X"36",X"D3",X"58",X"8B",X"15",X"46",X"FD",X"CA",
		X"04",X"36",X"06",X"9E",X"48",X"BF",X"CA",X"02",X"EC",X"1E",X"FD",X"CA",X"06",X"86",X"0A",X"24",
		X"02",X"8A",X"20",X"36",X"12",X"B7",X"CA",X"00",X"9E",X"4A",X"BF",X"CA",X"02",X"AE",X"1E",X"BF",
		X"CA",X"06",X"DC",X"36",X"D3",X"56",X"C3",X"16",X"01",X"46",X"FD",X"CA",X"04",X"86",X"0A",X"24",
		X"02",X"8A",X"20",X"B7",X"CA",X"00",X"35",X"D7",X"10",X"CE",X"9A",X"2B",X"B6",X"9A",X"10",X"32",
		X"E6",X"86",X"18",X"B7",X"9A",X"10",X"11",X"8C",X"9A",X"43",X"10",X"2C",X"92",X"22",X"35",X"36",
		X"BD",X"0A",X"4E",X"A6",X"2B",X"84",X"7F",X"A7",X"2B",X"20",X"EB",X"96",X"00",X"84",X"80",X"27",
		X"11",X"DC",X"17",X"83",X"00",X"01",X"2E",X"08",X"C6",X"06",X"BD",X"D2",X"1B",X"CC",X"0E",X"10",
		X"DD",X"17",X"96",X"88",X"27",X"02",X"0A",X"88",X"DC",X"83",X"DD",X"84",X"DC",X"81",X"DD",X"82",
		X"DC",X"7F",X"DD",X"80",X"DC",X"7D",X"DD",X"7E",X"FC",X"C8",X"0C",X"97",X"7D",X"85",X"40",X"27",
		X"04",X"C6",X"78",X"D7",X"88",X"D6",X"7D",X"DA",X"7E",X"DA",X"7F",X"DA",X"80",X"DA",X"81",X"DA",
		X"82",X"DA",X"83",X"DA",X"84",X"DA",X"85",X"D4",X"86",X"D7",X"87",X"94",X"7E",X"9A",X"87",X"D6",
		X"86",X"97",X"86",X"53",X"D4",X"86",X"C4",X"3E",X"27",X"36",X"54",X"34",X"04",X"64",X"E4",X"24",
		X"03",X"7E",X"F0",X"03",X"96",X"88",X"26",X"09",X"64",X"E4",X"24",X"05",X"8D",X"4A",X"BD",X"D2",
		X"3F",X"64",X"E4",X"24",X"03",X"BD",X"D2",X"15",X"96",X"88",X"26",X"12",X"64",X"E4",X"24",X"05",
		X"8D",X"36",X"BD",X"D2",X"39",X"64",X"E4",X"24",X"05",X"8D",X"2D",X"BD",X"D2",X"3C",X"35",X"04",
		X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"9A",X"43",X"B6",X"9A",X"11",X"32",X"E6",X"86",X"18",
		X"B7",X"9A",X"11",X"11",X"8C",X"9A",X"5B",X"10",X"2C",X"91",X"65",X"35",X"36",X"BD",X"0A",X"4E",
		X"A6",X"2B",X"84",X"7F",X"A7",X"2B",X"20",X"EB",X"34",X"17",X"C6",X"17",X"7E",X"07",X"29",X"9E",
		X"13",X"DC",X"27",X"26",X"1A",X"30",X"03",X"A6",X"84",X"27",X"04",X"9F",X"13",X"20",X"18",X"96",
		X"97",X"97",X"29",X"27",X"06",X"9E",X"98",X"0F",X"97",X"20",X"EA",X"C6",X"13",X"20",X"0F",X"5A",
		X"D7",X"28",X"26",X"14",X"4A",X"27",X"DE",X"E6",X"01",X"5C",X"DD",X"27",X"E6",X"02",X"86",X"3F",
		X"B7",X"C8",X"0E",X"C8",X"3F",X"F7",X"C8",X"0E",X"10",X"CE",X"9A",X"5B",X"B6",X"9A",X"12",X"32",
		X"E6",X"86",X"18",X"B7",X"9A",X"12",X"11",X"8C",X"9A",X"73",X"10",X"2C",X"91",X"02",X"35",X"36",
		X"BD",X"0A",X"4E",X"A6",X"2B",X"84",X"7F",X"A7",X"2B",X"20",X"EB",X"34",X"17",X"1A",X"50",X"AE",
		X"65",X"E6",X"80",X"AF",X"65",X"96",X"00",X"2A",X"1E",X"58",X"8E",X"07",X"55",X"AE",X"85",X"A6",
		X"02",X"84",X"7F",X"91",X"29",X"24",X"12",X"D6",X"97",X"C4",X"7F",X"E7",X"E2",X"A1",X"E0",X"25",
		X"06",X"A6",X"02",X"97",X"97",X"9F",X"98",X"35",X"97",X"A6",X"02",X"97",X"29",X"4F",X"5F",X"DD",
		X"27",X"9F",X"13",X"35",X"97",X"07",X"83",X"07",X"88",X"07",X"8D",X"07",X"92",X"07",X"9A",X"07",
		X"9F",X"07",X"A4",X"07",X"AF",X"07",X"B4",X"07",X"B9",X"07",X"C1",X"07",X"C6",X"07",X"D1",X"07",
		X"D6",X"07",X"DB",X"07",X"E0",X"07",X"E5",X"07",X"EA",X"07",X"EF",X"07",X"F7",X"07",X"FC",X"08",
		X"04",X"08",X"09",X"08",X"0E",X"7F",X"01",X"90",X"14",X"00",X"14",X"01",X"32",X"02",X"00",X"14",
		X"01",X"46",X"08",X"00",X"1E",X"02",X"0B",X"04",X"01",X"14",X"04",X"00",X"1E",X"01",X"28",X"07",
		X"00",X"14",X"01",X"0A",X"09",X"00",X"7E",X"03",X"0A",X"0A",X"01",X"1E",X"09",X"01",X"01",X"13",
		X"00",X"70",X"08",X"0A",X"0E",X"00",X"1E",X"01",X"28",X"0D",X"00",X"7D",X"01",X"30",X"0C",X"01",
		X"28",X"0E",X"00",X"7F",X"01",X"01",X"13",X"00",X"FF",X"01",X"77",X"15",X"01",X"30",X"0B",X"01",
		X"01",X"13",X"00",X"29",X"01",X"50",X"04",X"00",X"7F",X"01",X"32",X"19",X"00",X"72",X"01",X"2D",
		X"0E",X"00",X"29",X"01",X"0A",X"08",X"00",X"72",X"01",X"FA",X"11",X"00",X"6A",X"01",X"1E",X"18",
		X"00",X"50",X"01",X"1E",X"1D",X"01",X"01",X"13",X"00",X"76",X"01",X"FA",X"11",X"00",X"7A",X"01",
		X"28",X"12",X"01",X"01",X"10",X"00",X"1E",X"01",X"02",X"05",X"00",X"7E",X"01",X"90",X"10",X"00",
		X"FF",X"01",X"40",X"04",X"00",X"34",X"53",X"9B",X"04",X"A7",X"2A",X"20",X"02",X"34",X"53",X"8E",
		X"9A",X"01",X"A6",X"25",X"AE",X"84",X"A1",X"05",X"22",X"FA",X"AF",X"A4",X"EE",X"02",X"EF",X"22",
		X"10",X"AF",X"02",X"10",X"AF",X"C4",X"35",X"D3",X"34",X"36",X"34",X"01",X"1A",X"50",X"EC",X"C1",
		X"27",X"1E",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"37",X"36",X"10",X"BF",X"CA",X"04",X"BF",
		X"CA",X"02",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"5F",X"F7",X"CA",X"01",X"35",X"01",X"20",X"DA",
		X"35",X"B7",X"34",X"57",X"86",X"0A",X"20",X"04",X"34",X"57",X"86",X"1A",X"AE",X"28",X"1A",X"50",
		X"A7",X"E2",X"EC",X"24",X"8B",X"15",X"46",X"BF",X"CA",X"02",X"EE",X"1E",X"FF",X"CA",X"06",X"FD",
		X"CA",X"04",X"A6",X"E0",X"24",X"02",X"8A",X"20",X"8C",X"90",X"00",X"25",X"02",X"8A",X"04",X"B7",
		X"CA",X"00",X"35",X"D7",X"96",X"04",X"4C",X"A7",X"2A",X"AD",X"B8",X"0E",X"AE",X"28",X"EC",X"24",
		X"39",X"A7",X"24",X"BD",X"18",X"4D",X"AD",X"B8",X"10",X"A6",X"24",X"81",X"08",X"22",X"08",X"8D",
		X"E3",X"2A",X"1E",X"86",X"FF",X"20",X"EA",X"A6",X"26",X"81",X"F6",X"25",X"12",X"8D",X"D5",X"AB",
		X"1C",X"25",X"06",X"81",X"FF",X"A6",X"24",X"25",X"08",X"86",X"FF",X"A0",X"1C",X"20",X"D2",X"8D",
		X"C3",X"C1",X"3F",X"25",X"CC",X"EB",X"1D",X"25",X"C8",X"C1",X"EA",X"22",X"C4",X"AB",X"1C",X"ED",
		X"26",X"96",X"96",X"27",X"21",X"AE",X"22",X"E6",X"25",X"E1",X"05",X"24",X"18",X"EE",X"A4",X"EF",
		X"84",X"AF",X"42",X"AE",X"02",X"E1",X"05",X"25",X"FA",X"EE",X"84",X"10",X"AF",X"84",X"AF",X"22",
		X"EF",X"A4",X"10",X"AF",X"42",X"39",X"E6",X"25",X"AE",X"A4",X"E1",X"05",X"23",X"18",X"EE",X"22",
		X"AF",X"C4",X"EF",X"02",X"AE",X"84",X"E1",X"05",X"22",X"FA",X"AF",X"A4",X"EE",X"02",X"10",X"AF",
		X"02",X"10",X"AF",X"C4",X"EF",X"22",X"39",X"BD",X"00",X"5A",X"96",X"95",X"26",X"F9",X"96",X"96",
		X"10",X"26",X"00",X"9B",X"BE",X"9A",X"09",X"9F",X"2A",X"1C",X"EF",X"10",X"9E",X"2A",X"AE",X"22",
		X"8C",X"9A",X"07",X"27",X"E2",X"9F",X"2A",X"F6",X"CB",X"00",X"CB",X"0C",X"E1",X"25",X"24",X"27",
		X"EC",X"2A",X"91",X"04",X"2A",X"03",X"5D",X"27",X"05",X"BD",X"09",X"06",X"20",X"DB",X"EC",X"24",
		X"AE",X"28",X"34",X"16",X"BD",X"08",X"A9",X"F6",X"CB",X"00",X"CB",X"0C",X"E1",X"25",X"24",X"25",
		X"35",X"16",X"BD",X"0A",X"4C",X"20",X"C2",X"EC",X"2A",X"90",X"04",X"4A",X"2A",X"DB",X"5D",X"26",
		X"D8",X"EC",X"24",X"AE",X"28",X"34",X"16",X"BD",X"08",X"A9",X"6C",X"2A",X"F6",X"CB",X"00",X"E1",
		X"27",X"24",X"DD",X"20",X"02",X"6C",X"2A",X"E6",X"27",X"CB",X"40",X"4F",X"58",X"49",X"58",X"49",
		X"26",X"01",X"4C",X"8D",X"05",X"27",X"C9",X"7E",X"09",X"39",X"CE",X"9A",X"0F",X"1A",X"50",X"E6",
		X"C6",X"27",X"17",X"C0",X"06",X"E7",X"C6",X"8E",X"09",X"CB",X"EB",X"86",X"33",X"C5",X"86",X"80",
		X"A7",X"2B",X"36",X"20",X"35",X"36",X"36",X"30",X"34",X"06",X"39",X"0A",X"22",X"3A",X"52",X"BE",
		X"9A",X"01",X"9F",X"2A",X"1C",X"EF",X"10",X"9E",X"2A",X"AE",X"A4",X"8C",X"9A",X"01",X"10",X"27",
		X"FF",X"45",X"9F",X"2A",X"F6",X"CB",X"00",X"CB",X"0C",X"53",X"E1",X"27",X"23",X"28",X"EC",X"2A",
		X"91",X"04",X"2A",X"03",X"5D",X"27",X"05",X"BD",X"08",X"E5",X"20",X"D8",X"EC",X"24",X"AE",X"28",
		X"34",X"16",X"BD",X"08",X"A9",X"F6",X"CB",X"00",X"CB",X"0C",X"53",X"E1",X"27",X"23",X"26",X"35",
		X"16",X"BD",X"0A",X"4C",X"20",X"BE",X"EC",X"2A",X"90",X"04",X"4A",X"2A",X"DA",X"5D",X"26",X"D7",
		X"EC",X"24",X"AE",X"28",X"34",X"16",X"BD",X"08",X"A9",X"6C",X"2A",X"F6",X"CB",X"00",X"53",X"E1",
		X"25",X"23",X"DC",X"20",X"02",X"6C",X"2A",X"E6",X"25",X"C0",X"40",X"4F",X"58",X"49",X"58",X"49",
		X"26",X"02",X"86",X"03",X"BD",X"09",X"AA",X"27",X"C6",X"7E",X"09",X"D4",X"1A",X"50",X"BF",X"CA",
		X"02",X"EE",X"1E",X"FF",X"CA",X"06",X"8B",X"15",X"46",X"FD",X"CA",X"04",X"86",X"1A",X"24",X"02",
		X"8A",X"20",X"8C",X"90",X"00",X"25",X"02",X"8A",X"04",X"B7",X"CA",X"00",X"AE",X"28",X"BF",X"CA",
		X"02",X"EE",X"1E",X"FF",X"CA",X"06",X"EC",X"24",X"8B",X"15",X"46",X"FD",X"CA",X"04",X"86",X"0A",
		X"24",X"02",X"8A",X"20",X"8C",X"90",X"00",X"25",X"02",X"8A",X"04",X"B7",X"CA",X"00",X"39",X"86",
		X"02",X"BD",X"00",X"5C",X"96",X"95",X"26",X"F7",X"CE",X"9A",X"07",X"AE",X"42",X"8C",X"9A",X"01",
		X"27",X"ED",X"CE",X"1B",X"B8",X"A6",X"0C",X"48",X"10",X"AE",X"C6",X"33",X"84",X"AE",X"84",X"EC",
		X"04",X"E1",X"47",X"22",X"E6",X"A1",X"46",X"22",X"F4",X"EC",X"0C",X"A6",X"A6",X"27",X"EE",X"E4",
		X"4D",X"27",X"EA",X"EC",X"06",X"A1",X"44",X"25",X"E4",X"E1",X"47",X"23",X"02",X"E6",X"47",X"E0",
		X"05",X"D7",X"2B",X"EC",X"04",X"A3",X"44",X"97",X"2A",X"58",X"34",X"50",X"EE",X"48",X"EE",X"5A",
		X"33",X"C5",X"AE",X"08",X"AE",X"1A",X"EC",X"81",X"DB",X"2A",X"E1",X"C1",X"2D",X"06",X"9B",X"2A",
		X"A1",X"5F",X"2F",X"08",X"0A",X"2B",X"2A",X"EE",X"35",X"50",X"20",X"B1",X"35",X"10",X"10",X"AE",
		X"E4",X"A6",X"2C",X"A1",X"0C",X"23",X"02",X"1E",X"12",X"BD",X"0C",X"64",X"35",X"40",X"7E",X"0A",
		X"9B",X"32",X"66",X"BD",X"00",X"5A",X"1A",X"50",X"DC",X"36",X"9E",X"38",X"DE",X"19",X"34",X"56",
		X"DC",X"5C",X"9E",X"5E",X"1C",X"EF",X"34",X"16",X"96",X"00",X"84",X"08",X"27",X"77",X"8E",X"9A",
		X"01",X"AE",X"84",X"EC",X"04",X"E1",X"63",X"22",X"6C",X"A1",X"62",X"22",X"F4",X"EC",X"06",X"E1",
		X"61",X"25",X"EE",X"A1",X"E4",X"25",X"EA",X"A6",X"0D",X"84",X"03",X"27",X"E4",X"CE",X"0C",X"0E",
		X"5F",X"A6",X"0C",X"5A",X"A1",X"C5",X"27",X"06",X"C1",X"FC",X"2E",X"F7",X"20",X"D3",X"D7",X"30",
		X"A6",X"E4",X"E6",X"62",X"A0",X"04",X"E0",X"04",X"DD",X"2C",X"E6",X"63",X"E1",X"07",X"23",X"02",
		X"E6",X"07",X"EE",X"08",X"EE",X"5A",X"A6",X"61",X"A0",X"05",X"25",X"07",X"48",X"33",X"C6",X"E0",
		X"61",X"20",X"02",X"E0",X"05",X"D7",X"2E",X"EC",X"C1",X"D1",X"2C",X"2D",X"04",X"91",X"2D",X"2F",
		X"06",X"0A",X"2E",X"2A",X"F2",X"20",X"9A",X"10",X"8E",X"9A",X"99",X"96",X"30",X"4C",X"A7",X"0C",
		X"BD",X"0C",X"64",X"20",X"8C",X"32",X"64",X"8E",X"9A",X"01",X"AE",X"84",X"EC",X"06",X"E1",X"61",
		X"25",X"F8",X"A1",X"E4",X"25",X"F4",X"EC",X"04",X"E1",X"63",X"10",X"22",X"FF",X"53",X"A1",X"62",
		X"22",X"E8",X"A0",X"E4",X"97",X"2C",X"A6",X"0D",X"84",X"03",X"27",X"DE",X"10",X"AE",X"64",X"EE",
		X"08",X"EE",X"5A",X"A6",X"07",X"A1",X"63",X"23",X"02",X"A6",X"63",X"E0",X"61",X"58",X"25",X"06",
		X"31",X"A5",X"A0",X"05",X"20",X"05",X"50",X"33",X"C5",X"A0",X"61",X"97",X"2E",X"37",X"06",X"DB",
		X"2C",X"E1",X"A1",X"2D",X"06",X"9B",X"2C",X"A1",X"3F",X"2F",X"06",X"0A",X"2E",X"2A",X"EE",X"20",
		X"A9",X"10",X"8E",X"9A",X"99",X"BD",X"0C",X"64",X"20",X"A0",X"09",X"07",X"08",X"04",X"20",X"42",
		X"55",X"42",X"42",X"4C",X"45",X"53",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",
		X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",
		X"4F",X"4E",X"49",X"43",X"53",X"20",X"31",X"39",X"38",X"33",X"34",X"77",X"1A",X"50",X"A6",X"2B",
		X"85",X"80",X"27",X"1E",X"84",X"7F",X"A7",X"2B",X"CE",X"9A",X"13",X"37",X"36",X"10",X"AC",X"65",
		X"26",X"F9",X"34",X"40",X"BD",X"0A",X"4E",X"35",X"40",X"8E",X"0D",X"A5",X"10",X"8E",X"D0",X"97",
		X"36",X"36",X"35",X"F7",X"34",X"30",X"8D",X"D2",X"1E",X"12",X"8D",X"CE",X"1E",X"12",X"E6",X"2C",
		X"CE",X"1B",X"D0",X"58",X"EE",X"C5",X"E6",X"0C",X"E0",X"2C",X"58",X"AD",X"D5",X"35",X"B0",X"8E",
		X"0D",X"49",X"4F",X"5F",X"ED",X"98",X"08",X"EE",X"81",X"EF",X"98",X"06",X"8C",X"0D",X"51",X"26",
		X"F3",X"8E",X"97",X"FF",X"86",X"39",X"B7",X"CB",X"FF",X"6F",X"80",X"8C",X"BF",X"7F",X"23",X"F6",
		X"86",X"98",X"1F",X"8B",X"7F",X"CA",X"01",X"10",X"CE",X"9C",X"22",X"CE",X"0D",X"2F",X"BD",X"08",
		X"38",X"8E",X"9B",X"DC",X"BF",X"9B",X"DC",X"BF",X"9B",X"DE",X"CC",X"02",X"08",X"FD",X"9B",X"E1",
		X"CC",X"99",X"8D",X"FD",X"A5",X"71",X"8E",X"9B",X"D6",X"AF",X"1A",X"30",X"1A",X"8C",X"9A",X"B0",
		X"26",X"F7",X"1C",X"EF",X"BD",X"00",X"AD",X"2F",X"03",X"1A",X"41",X"8E",X"CC",X"00",X"BD",X"D2",
		X"21",X"97",X"1D",X"8E",X"CD",X"00",X"BD",X"D2",X"24",X"1F",X"98",X"81",X"20",X"22",X"06",X"84",
		X"0F",X"81",X"09",X"23",X"07",X"5F",X"8E",X"CD",X"00",X"BD",X"D2",X"2D",X"F7",X"BF",X"23",X"8E",
		X"CC",X"14",X"BD",X"D2",X"21",X"C6",X"19",X"3D",X"D7",X"1E",X"50",X"D7",X"1F",X"BD",X"38",X"2A",
		X"BD",X"31",X"E6",X"BD",X"00",X"5A",X"BD",X"15",X"BD",X"96",X"22",X"27",X"F6",X"8E",X"0D",X"25",
		X"48",X"AD",X"96",X"0F",X"22",X"20",X"EC",X"0D",X"F5",X"0D",X"E6",X"31",X"C4",X"31",X"CB",X"00",
		X"17",X"00",X"00",X"0D",X"59",X"98",X"06",X"00",X"31",X"00",X"00",X"0D",X"70",X"99",X"E2",X"00",
		X"04",X"00",X"00",X"0D",X"AC",X"98",X"62",X"00",X"00",X"00",X"34",X"FF",X"35",X"00",X"34",X"00",
		X"3C",X"C8",X"0C",X"C8",X"0E",X"C8",X"04",X"C8",X"06",X"A5",X"5A",X"9B",X"DC",X"04",X"EC",X"9A",
		X"B0",X"C8",X"04",X"7E",X"02",X"8A",X"07",X"C1",X"FF",X"FF",X"0E",X"10",X"99",X"00",X"99",X"00",
		X"C0",X"0D",X"A5",X"00",X"00",X"C0",X"0D",X"A5",X"00",X"00",X"C0",X"0D",X"A5",X"00",X"00",X"C9",
		X"FF",X"2F",X"1F",X"06",X"0A",X"DA",X"AC",X"80",X"00",X"F0",X"C5",X"53",X"92",X"A6",X"00",X"9A",
		X"07",X"9A",X"07",X"00",X"00",X"9A",X"01",X"9A",X"01",X"00",X"FF",X"FF",X"FF",X"18",X"18",X"18",
		X"18",X"00",X"00",X"04",X"05",X"00",X"98",X"19",X"19",X"CF",X"9A",X"78",X"19",X"91",X"9A",X"73",
		X"03",X"0C",X"00",X"01",X"00",X"8E",X"CC",X"06",X"BD",X"D2",X"21",X"81",X"09",X"27",X"26",X"F1",
		X"BF",X"23",X"23",X"02",X"35",X"86",X"B6",X"BF",X"23",X"5A",X"27",X"08",X"C6",X"0A",X"BD",X"D2",
		X"1B",X"8B",X"99",X"19",X"C6",X"0A",X"BD",X"D2",X"1B",X"8B",X"99",X"19",X"B7",X"BF",X"23",X"8E",
		X"CD",X"00",X"BD",X"D2",X"2A",X"39",X"C6",X"02",X"D7",X"02",X"8D",X"C9",X"C6",X"09",X"BD",X"D2",
		X"1B",X"86",X"C0",X"20",X"0E",X"C6",X"FF",X"D7",X"02",X"50",X"8D",X"B9",X"C6",X"08",X"BD",X"D2",
		X"1B",X"86",X"80",X"97",X"00",X"97",X"93",X"97",X"94",X"97",X"96",X"BD",X"00",X"AD",X"4D",X"1A",
		X"02",X"36",X"7F",X"BF",X"25",X"0F",X"01",X"BD",X"07",X"1B",X"00",X"8E",X"03",X"0A",X"9F",X"11",
		X"CE",X"0E",X"9B",X"BD",X"08",X"38",X"96",X"1D",X"97",X"6B",X"B7",X"9A",X"90",X"8E",X"CC",X"02",
		X"BD",X"D2",X"24",X"BD",X"D2",X"45",X"F7",X"9A",X"7D",X"F7",X"9A",X"8B",X"5A",X"D7",X"66",X"CE",
		X"14",X"59",X"BD",X"00",X"E2",X"37",X"16",X"ED",X"2B",X"BD",X"02",X"4D",X"BD",X"00",X"5A",X"96",
		X"90",X"26",X"F9",X"BD",X"38",X"2A",X"BD",X"30",X"46",X"BD",X"1A",X"C5",X"7A",X"9A",X"7D",X"BD",
		X"00",X"AD",X"4D",X"06",X"13",X"43",X"BD",X"00",X"AD",X"43",X"04",X"45",X"C1",X"BD",X"00",X"A5",
		X"3A",X"CB",X"39",X"10",X"39",X"A1",X"BD",X"00",X"AD",X"2F",X"19",X"31",X"0E",X"7F",X"9A",X"98",
		X"7E",X"11",X"FC",X"78",X"45",X"84",X"51",X"78",X"00",X"45",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"A5",X"78",X"45",X"84",X"51",X"0D",X"AC",X"00",X"10",X"01",X"FE",X"00",X"09",X"00",X"00",X"0D",
		X"AC",X"98",X"62",X"00",X"05",X"00",X"00",X"0D",X"B0",X"98",X"66",X"00",X"05",X"00",X"00",X"0D",
		X"B0",X"9A",X"7D",X"00",X"05",X"00",X"00",X"0D",X"B0",X"9A",X"8B",X"00",X"0A",X"10",X"00",X"00",
		X"00",X"9A",X"73",X"00",X"0A",X"00",X"00",X"0E",X"91",X"9A",X"9D",X"00",X"0E",X"00",X"00",X"0E",
		X"83",X"98",X"36",X"00",X"11",X"00",X"00",X"0D",X"70",X"99",X"E2",X"00",X"00",X"01",X"00",X"01",
		X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"10",X"7C",X"02",X"00",X"00",X"00",X"00",
		X"00",X"28",X"F6",X"00",X"00",X"0C",X"FA",X"10",X"65",X"02",X"00",X"00",X"00",X"00",X"00",X"28",
		X"FA",X"01",X"00",X"0C",X"FA",X"10",X"65",X"03",X"00",X"00",X"00",X"14",X"F8",X"14",X"FA",X"01",
		X"00",X"0C",X"FA",X"10",X"65",X"03",X"00",X"02",X"00",X"14",X"F8",X"14",X"FA",X"01",X"00",X"0C",
		X"FA",X"10",X"65",X"00",X"00",X"00",X"00",X"1E",X"F2",X"00",X"00",X"06",X"00",X"0C",X"FA",X"10",
		X"69",X"03",X"00",X"03",X"00",X"14",X"F8",X"14",X"FA",X"02",X"02",X"0C",X"FA",X"10",X"69",X"06",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"03",X"00",X"0C",X"FA",X"10",X"69",X"00",X"00",X"06",
		X"00",X"14",X"00",X"14",X"00",X"02",X"02",X"0C",X"FA",X"10",X"69",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"28",X"F1",X"10",X"6D",X"04",X"00",X"03",X"00",X"00",X"00",X"28",
		X"F3",X"02",X"04",X"11",X"F8",X"10",X"72",X"02",X"02",X"04",X"02",X"14",X"00",X"14",X"00",X"03",
		X"00",X"11",X"F8",X"10",X"72",X"03",X"02",X"03",X"02",X"1E",X"F6",X"14",X"F6",X"04",X"00",X"11",
		X"F8",X"10",X"72",X"00",X"00",X"00",X"00",X"30",X"EC",X"00",X"00",X"06",X"08",X"14",X"F6",X"10",
		X"72",X"05",X"02",X"04",X"02",X"19",X"F6",X"19",X"F6",X"00",X"00",X"13",X"F8",X"10",X"72",X"00",
		X"00",X"04",X"08",X"14",X"00",X"14",X"00",X"03",X"03",X"13",X"F8",X"10",X"76",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"F1",X"10",X"6D",X"05",X"02",X"05",X"02",X"19",
		X"F6",X"19",X"F6",X"03",X"03",X"0F",X"F8",X"10",X"76",X"07",X"05",X"00",X"00",X"14",X"00",X"14",
		X"00",X"03",X"03",X"14",X"F8",X"10",X"76",X"05",X"05",X"02",X"04",X"00",X"00",X"32",X"F1",X"04",
		X"06",X"14",X"F6",X"10",X"7A",X"00",X"00",X"00",X"00",X"2D",X"EC",X"00",X"00",X"0A",X"0A",X"14",
		X"F6",X"10",X"7A",X"05",X"02",X"05",X"02",X"19",X"F6",X"23",X"F6",X"04",X"03",X"28",X"EE",X"10",
		X"7C",X"04",X"07",X"04",X"06",X"1E",X"F6",X"19",X"F6",X"00",X"00",X"14",X"F6",X"10",X"7A",X"00",
		X"00",X"06",X"08",X"14",X"00",X"14",X"00",X"03",X"08",X"1E",X"F2",X"10",X"7A",X"04",X"05",X"03",
		X"06",X"19",X"F6",X"19",X"F6",X"04",X"08",X"19",X"F6",X"10",X"7A",X"0A",X"08",X"00",X"00",X"14",
		X"00",X"14",X"00",X"05",X"08",X"19",X"F6",X"10",X"7A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"28",X"F1",X"10",X"7D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"06",X"32",X"E7",X"10",X"7A",X"14",X"93",X"A4",X"00",X"13",X"A3",X"94",X"00",X"22",X"B2",X"22",
		X"B2",X"00",X"13",X"A2",X"93",X"00",X"13",X"A2",X"A3",X"00",X"12",X"C2",X"00",X"B1",X"21",X"A2",
		X"22",X"A2",X"00",X"0C",X"14",X"1E",X"06",X"00",X"02",X"00",X"08",X"00",X"0B",X"11",X"0C",X"0C",
		X"0D",X"37",X"0D",X"03",X"12",X"14",X"1E",X"07",X"02",X"04",X"02",X"09",X"04",X"09",X"0E",X"0C",
		X"14",X"0E",X"2D",X"0F",X"04",X"14",X"1E",X"19",X"08",X"03",X"05",X"03",X"0A",X"04",X"07",X"0B",
		X"10",X"14",X"0C",X"23",X"12",X"04",X"14",X"1E",X"14",X"08",X"04",X"05",X"05",X"0A",X"04",X"06",
		X"09",X"14",X"14",X"0B",X"1E",X"14",X"05",X"14",X"1E",X"14",X"09",X"0F",X"0A",X"0A",X"04",X"04",
		X"05",X"08",X"14",X"19",X"0A",X"1E",X"18",X"05",X"14",X"1E",X"0F",X"09",X"04",X"06",X"03",X"07",
		X"0A",X"06",X"09",X"14",X"1E",X"0A",X"1E",X"1C",X"04",X"19",X"1E",X"0F",X"09",X"04",X"06",X"06",
		X"0A",X"04",X"06",X"09",X"19",X"1E",X"09",X"19",X"1E",X"04",X"19",X"1E",X"0F",X"09",X"14",X"0A",
		X"0A",X"04",X"04",X"04",X"07",X"19",X"1E",X"09",X"19",X"20",X"05",X"1E",X"1E",X"0E",X"0A",X"02",
		X"05",X"05",X"0A",X"04",X"05",X"08",X"1E",X"1E",X"09",X"19",X"22",X"05",X"1E",X"1E",X"0C",X"0B",
		X"06",X"06",X"09",X"08",X"07",X"05",X"08",X"1E",X"1E",X"08",X"19",X"26",X"05",X"1E",X"1E",X"0A",
		X"0C",X"08",X"06",X"09",X"08",X"0C",X"03",X"05",X"1E",X"1E",X"07",X"19",X"28",X"03",X"1E",X"1E",
		X"08",X"0D",X"08",X"09",X"05",X"06",X"08",X"02",X"04",X"1E",X"1E",X"07",X"19",X"28",X"04",X"1E",
		X"1E",X"0C",X"0E",X"09",X"06",X"03",X"08",X"07",X"04",X"06",X"1E",X"1E",X"06",X"19",X"23",X"07",
		X"1E",X"1E",X"04",X"0F",X"0A",X"0F",X"0A",X"04",X"03",X"02",X"04",X"1E",X"1E",X"06",X"19",X"23",
		X"06",X"1E",X"1E",X"02",X"10",X"0A",X"07",X"04",X"08",X"09",X"03",X"05",X"1E",X"1E",X"06",X"14",
		X"2D",X"06",X"1E",X"1E",X"02",X"11",X"0A",X"07",X"04",X"08",X"0A",X"02",X"04",X"1E",X"1E",X"05",
		X"14",X"28",X"04",X"1E",X"1E",X"06",X"14",X"0A",X"08",X"04",X"04",X"0A",X"06",X"09",X"1E",X"1E",
		X"05",X"14",X"23",X"05",X"34",X"77",X"20",X"03",X"BD",X"00",X"5A",X"96",X"00",X"84",X"20",X"27",
		X"F7",X"AE",X"69",X"EE",X"81",X"AF",X"69",X"BD",X"15",X"AE",X"35",X"F7",X"BD",X"1A",X"C5",X"CE",
		X"0E",X"C3",X"BD",X"08",X"38",X"BD",X"00",X"5A",X"BD",X"00",X"AD",X"39",X"05",X"20",X"04",X"BD",
		X"00",X"AD",X"57",X"01",X"0A",X"8F",X"BD",X"00",X"AD",X"57",X"09",X"0B",X"13",X"96",X"73",X"27",
		X"06",X"96",X"00",X"8A",X"08",X"97",X"00",X"86",X"02",X"BD",X"00",X"5C",X"BD",X"18",X"34",X"39",
		X"0C",X"69",X"27",X"FC",X"BD",X"07",X"1B",X"06",X"86",X"0C",X"97",X"67",X"0F",X"73",X"BD",X"37",
		X"64",X"4F",X"5F",X"BD",X"1E",X"E5",X"BD",X"00",X"AD",X"7F",X"1A",X"44",X"10",X"CE",X"0E",X"DD",
		X"D6",X"1E",X"D7",X"30",X"D6",X"69",X"C1",X"14",X"23",X"0D",X"C0",X"14",X"D7",X"30",X"C0",X"09",
		X"24",X"FC",X"CB",X"09",X"CE",X"0F",X"E7",X"86",X"0E",X"3D",X"8E",X"98",X"6C",X"33",X"CB",X"DF",
		X"7B",X"D6",X"30",X"A6",X"41",X"3D",X"2A",X"02",X"90",X"30",X"AB",X"C1",X"A7",X"80",X"8C",X"98",
		X"72",X"26",X"EE",X"96",X"6E",X"9B",X"6F",X"97",X"72",X"BD",X"00",X"5A",X"BD",X"2F",X"10",X"BD",
		X"11",X"BC",X"D6",X"69",X"54",X"C1",X"09",X"23",X"06",X"C0",X"07",X"24",X"FC",X"CB",X"11",X"CE",
		X"10",X"83",X"86",X"11",X"3D",X"33",X"CB",X"DF",X"79",X"A6",X"C8",X"10",X"97",X"8E",X"EC",X"C1",
		X"DD",X"74",X"96",X"6C",X"BD",X"24",X"0E",X"33",X"47",X"96",X"6D",X"BD",X"26",X"11",X"96",X"6E",
		X"E6",X"C0",X"BD",X"28",X"5A",X"96",X"6F",X"E6",X"C0",X"BD",X"27",X"34",X"96",X"70",X"BD",X"30",
		X"13",X"BD",X"00",X"AD",X"39",X"0C",X"29",X"29",X"86",X"01",X"BD",X"01",X"48",X"96",X"00",X"8A",
		X"20",X"97",X"00",X"BD",X"00",X"AD",X"39",X"18",X"29",X"EE",X"BD",X"00",X"AD",X"39",X"02",X"09",
		X"27",X"39",X"BD",X"07",X"1B",X"0B",X"BD",X"14",X"85",X"86",X"04",X"BD",X"00",X"5C",X"CE",X"14",
		X"52",X"BD",X"00",X"E2",X"96",X"00",X"84",X"7F",X"97",X"00",X"86",X"FF",X"97",X"8F",X"8E",X"02",
		X"8A",X"9F",X"11",X"BD",X"37",X"12",X"0F",X"01",X"BD",X"02",X"4D",X"BD",X"00",X"AD",X"7F",X"12",
		X"12",X"E5",X"7E",X"00",X"89",X"7E",X"D2",X"51",X"0F",X"8F",X"BD",X"02",X"4D",X"CE",X"32",X"3D",
		X"BD",X"31",X"E1",X"7E",X"00",X"89",X"BD",X"14",X"85",X"96",X"00",X"85",X"40",X"27",X"3A",X"96",
		X"02",X"26",X"15",X"0A",X"02",X"96",X"01",X"88",X"01",X"8B",X"12",X"34",X"02",X"BD",X"7B",X"12",
		X"BD",X"37",X"12",X"35",X"02",X"BD",X"7B",X"1A",X"BD",X"02",X"4D",X"96",X"01",X"8B",X"12",X"BD",
		X"7B",X"12",X"86",X"02",X"D6",X"02",X"2B",X"05",X"F6",X"C8",X"06",X"2A",X"02",X"86",X"01",X"BD",
		X"01",X"48",X"96",X"01",X"8B",X"12",X"BD",X"7B",X"1A",X"0A",X"66",X"9E",X"62",X"6A",X"98",X"F6",
		X"BD",X"11",X"FE",X"BD",X"00",X"5A",X"96",X"71",X"27",X"F9",X"BD",X"00",X"5A",X"BD",X"18",X"46",
		X"81",X"05",X"22",X"F6",X"BD",X"00",X"AD",X"25",X"15",X"3A",X"1C",X"BD",X"15",X"BD",X"86",X"14",
		X"3D",X"8B",X"06",X"A7",X"2B",X"BD",X"18",X"46",X"27",X"0D",X"4F",X"BD",X"00",X"5C",X"6A",X"2B",
		X"26",X"F3",X"BD",X"31",X"23",X"20",X"E4",X"BD",X"1F",X"61",X"86",X"01",X"BD",X"00",X"5C",X"C6",
		X"01",X"96",X"67",X"81",X"12",X"24",X"01",X"50",X"D7",X"8D",X"BD",X"31",X"3D",X"96",X"8D",X"2A",
		X"19",X"BD",X"00",X"AD",X"4D",X"14",X"14",X"F3",X"30",X"A4",X"BD",X"01",X"27",X"B6",X"13",X"9D",
		X"BD",X"00",X"5C",X"20",X"F8",X"0F",X"8D",X"BD",X"31",X"3D",X"BD",X"00",X"5A",X"86",X"17",X"BD",
		X"01",X"13",X"27",X"F6",X"BD",X"18",X"28",X"BD",X"23",X"0B",X"BD",X"11",X"F0",X"7E",X"13",X"43",
		X"4F",X"5F",X"DD",X"56",X"DD",X"58",X"CC",X"24",X"52",X"0D",X"8D",X"26",X"03",X"CC",X"25",X"10",
		X"34",X"06",X"BD",X"1E",X"D9",X"BD",X"14",X"25",X"BD",X"18",X"23",X"86",X"02",X"BD",X"00",X"5C",
		X"A6",X"E4",X"BD",X"7B",X"12",X"BD",X"07",X"1B",X"16",X"96",X"67",X"80",X"11",X"2F",X"2A",X"8E",
		X"51",X"51",X"34",X"12",X"C6",X"DD",X"BD",X"7B",X"00",X"BD",X"14",X"25",X"A6",X"64",X"D6",X"8D",
		X"26",X"05",X"BD",X"19",X"1B",X"20",X"03",X"BD",X"19",X"24",X"86",X"0A",X"BD",X"00",X"5C",X"35",
		X"12",X"5F",X"BD",X"7B",X"00",X"0A",X"67",X"20",X"D0",X"A6",X"E1",X"BD",X"7B",X"1A",X"BD",X"07",
		X"1B",X"0A",X"7E",X"00",X"89",X"D6",X"67",X"C0",X"0C",X"58",X"8E",X"23",X"9A",X"3A",X"EC",X"84",
		X"DD",X"48",X"EC",X"06",X"DD",X"46",X"EC",X"88",X"20",X"DD",X"4A",X"CC",X"19",X"53",X"0D",X"01",
		X"27",X"02",X"86",X"CC",X"7E",X"1F",X"41",X"0D",X"0E",X"0F",X"0C",X"09",X"01",X"0A",X"18",X"15",
		X"05",X"00",X"10",X"07",X"16",X"15",X"19",X"04",X"00",X"1B",X"0B",X"11",X"12",X"06",X"14",X"00",
		X"23",X"66",X"96",X"00",X"84",X"C7",X"97",X"00",X"BD",X"22",X"F4",X"CE",X"14",X"47",X"BD",X"00",
		X"E2",X"86",X"0D",X"BD",X"01",X"13",X"26",X"03",X"BD",X"01",X"27",X"7E",X"18",X"28",X"A6",X"2A",
		X"8B",X"04",X"A7",X"2A",X"39",X"8E",X"9A",X"01",X"CE",X"14",X"7E",X"AE",X"84",X"8C",X"9A",X"07",
		X"27",X"04",X"EF",X"0E",X"20",X"F5",X"8D",X"CA",X"BD",X"22",X"99",X"86",X"02",X"BD",X"00",X"EE",
		X"BD",X"00",X"5A",X"BE",X"9A",X"0F",X"8C",X"18",X"18",X"26",X"F5",X"BE",X"9A",X"11",X"8C",X"18",
		X"18",X"26",X"ED",X"8E",X"9A",X"01",X"AE",X"84",X"8C",X"9A",X"07",X"26",X"0D",X"0F",X"89",X"0F",
		X"8A",X"BE",X"99",X"B2",X"2A",X"03",X"7F",X"99",X"B2",X"39",X"8C",X"A5",X"71",X"23",X"E7",X"A6",
		X"0B",X"84",X"10",X"26",X"E1",X"31",X"84",X"96",X"90",X"81",X"0E",X"27",X"03",X"BD",X"08",X"68",
		X"BD",X"00",X"47",X"BD",X"01",X"A9",X"20",X"CE",X"BD",X"12",X"AA",X"CC",X"7D",X"90",X"DD",X"60",
		X"7E",X"23",X"0B",X"96",X"00",X"8A",X"20",X"97",X"00",X"8D",X"ED",X"BD",X"1F",X"41",X"BD",X"05",
		X"0F",X"86",X"01",X"BD",X"00",X"5C",X"9E",X"8B",X"A6",X"0C",X"81",X"0A",X"27",X"23",X"BD",X"1F",
		X"2D",X"34",X"06",X"EC",X"04",X"AB",X"06",X"46",X"EB",X"07",X"56",X"A0",X"E4",X"E0",X"61",X"BD",
		X"15",X"DA",X"1F",X"98",X"D6",X"67",X"54",X"54",X"BD",X"16",X"23",X"AB",X"E0",X"EB",X"E0",X"DD",
		X"60",X"BD",X"07",X"1B",X"09",X"DE",X"08",X"86",X"02",X"A7",X"45",X"BD",X"14",X"68",X"96",X"90",
		X"27",X"06",X"CE",X"36",X"6A",X"7E",X"36",X"73",X"C6",X"07",X"BD",X"D2",X"1B",X"96",X"02",X"2B",
		X"51",X"D6",X"66",X"D7",X"02",X"10",X"8E",X"0D",X"AC",X"CE",X"9A",X"7D",X"8E",X"9A",X"8B",X"0A",
		X"01",X"27",X"06",X"31",X"3C",X"1E",X"13",X"00",X"01",X"1A",X"50",X"BF",X"CA",X"04",X"8E",X"98",
		X"66",X"BF",X"CA",X"02",X"CC",X"04",X"0A",X"FD",X"CA",X"06",X"86",X"04",X"B7",X"CA",X"00",X"C6",
		X"00",X"FF",X"CA",X"02",X"BF",X"CA",X"04",X"B7",X"CA",X"00",X"8E",X"98",X"62",X"10",X"BF",X"CA",
		X"02",X"BF",X"CA",X"04",X"F7",X"CA",X"07",X"7F",X"CA",X"00",X"BD",X"11",X"A4",X"12",X"F6",X"7E",
		X"00",X"89",X"96",X"66",X"26",X"F4",X"BD",X"11",X"A4",X"12",X"B2",X"7E",X"00",X"89",X"86",X"06",
		X"BD",X"01",X"13",X"EF",X"98",X"07",X"7E",X"01",X"27",X"8D",X"02",X"1F",X"98",X"34",X"03",X"D6",
		X"05",X"86",X"03",X"3D",X"CB",X"11",X"96",X"07",X"44",X"44",X"44",X"98",X"07",X"44",X"06",X"06",
		X"06",X"07",X"DB",X"07",X"D9",X"06",X"D7",X"05",X"35",X"83",X"34",X"13",X"DD",X"34",X"2A",X"01",
		X"40",X"5D",X"2A",X"01",X"50",X"DD",X"2C",X"5F",X"91",X"2D",X"24",X"02",X"CA",X"20",X"86",X"10",
		X"DD",X"2F",X"8E",X"16",X"47",X"DA",X"2F",X"3A",X"96",X"2D",X"E6",X"88",X"40",X"3D",X"DD",X"32",
		X"96",X"2C",X"E6",X"84",X"3D",X"93",X"32",X"22",X"06",X"D6",X"30",X"DA",X"2F",X"D7",X"30",X"D6",
		X"30",X"04",X"2F",X"24",X"DD",X"96",X"34",X"2A",X"03",X"50",X"CB",X"80",X"96",X"35",X"2A",X"01",
		X"50",X"35",X"93",X"8E",X"16",X"47",X"DD",X"2F",X"84",X"7F",X"A6",X"86",X"3D",X"D6",X"2F",X"2A",
		X"01",X"40",X"97",X"32",X"CB",X"40",X"D7",X"33",X"C4",X"7F",X"E6",X"85",X"96",X"30",X"3D",X"D6",
		X"33",X"2A",X"01",X"40",X"D6",X"32",X"39",X"00",X"06",X"0D",X"13",X"19",X"1F",X"25",X"2C",X"32",
		X"38",X"3E",X"44",X"4A",X"50",X"56",X"5C",X"62",X"67",X"6D",X"72",X"78",X"7E",X"83",X"88",X"8E",
		X"93",X"98",X"9D",X"A2",X"A7",X"AB",X"B0",X"B4",X"B9",X"BD",X"C1",X"C5",X"C9",X"CD",X"D0",X"D4",
		X"D7",X"DB",X"DE",X"E1",X"E4",X"E7",X"E9",X"EC",X"EE",X"F0",X"F2",X"F4",X"F6",X"F7",X"F9",X"FA",
		X"FB",X"FC",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FD",X"FC",X"FB",X"FA",
		X"F9",X"F7",X"F6",X"F4",X"F2",X"F0",X"EE",X"EC",X"E9",X"E7",X"E4",X"E1",X"DE",X"DB",X"D7",X"D4",
		X"D0",X"CD",X"C9",X"C5",X"C1",X"BD",X"B9",X"B4",X"B0",X"AB",X"A7",X"A2",X"9D",X"98",X"93",X"8E",
		X"88",X"83",X"7E",X"78",X"72",X"6D",X"67",X"62",X"5C",X"56",X"50",X"4A",X"44",X"3E",X"38",X"32",
		X"2C",X"25",X"1F",X"19",X"13",X"0D",X"06",X"34",X"15",X"DD",X"2C",X"27",X"3D",X"48",X"29",X"06",
		X"58",X"28",X"FA",X"56",X"47",X"49",X"46",X"DD",X"2C",X"D6",X"2C",X"2A",X"02",X"40",X"50",X"3D",
		X"DD",X"2E",X"96",X"2D",X"D6",X"2D",X"2A",X"02",X"40",X"50",X"3D",X"D3",X"2E",X"2A",X"02",X"86",
		X"7F",X"8E",X"16",X"FC",X"30",X"86",X"A6",X"84",X"D6",X"2D",X"3D",X"2A",X"02",X"A0",X"84",X"A7",
		X"61",X"A6",X"84",X"D6",X"2C",X"3D",X"2A",X"02",X"A0",X"84",X"35",X"95",X"FF",X"FB",X"F3",X"EC",
		X"E5",X"DF",X"D9",X"D6",X"D1",X"CC",X"C9",X"C4",X"C2",X"BD",X"BB",X"B7",X"B5",X"B3",X"AF",X"AD",
		X"AA",X"A8",X"A6",X"A4",X"A1",X"A0",X"9E",X"9C",X"99",X"98",X"97",X"95",X"94",X"91",X"90",X"8F",
		X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"86",X"85",X"84",X"83",X"82",X"81",X"7F",X"7F",X"7E",X"7D",
		X"7C",X"7B",X"7A",X"79",X"78",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"72",X"71",X"71",X"70",
		X"6F",X"6F",X"6E",X"6D",X"6C",X"6C",X"6C",X"6B",X"6A",X"69",X"69",X"69",X"68",X"67",X"67",X"66",
		X"66",X"66",X"65",X"64",X"64",X"64",X"63",X"62",X"62",X"61",X"61",X"61",X"60",X"60",X"60",X"5F",
		X"5E",X"5E",X"5E",X"5D",X"5D",X"5C",X"5C",X"5C",X"5B",X"5B",X"5B",X"5A",X"34",X"57",X"4F",X"5F",
		X"ED",X"63",X"43",X"53",X"DD",X"2E",X"8E",X"9A",X"01",X"AE",X"84",X"8C",X"9A",X"01",X"26",X"02",
		X"35",X"D7",X"EE",X"65",X"A6",X"C0",X"27",X"F1",X"A1",X"0C",X"26",X"F8",X"A6",X"04",X"A0",X"61",
		X"46",X"2A",X"01",X"40",X"1F",X"89",X"3D",X"DD",X"2C",X"A6",X"05",X"A0",X"62",X"46",X"2A",X"01",
		X"40",X"1F",X"89",X"3D",X"D3",X"2C",X"10",X"93",X"2E",X"24",X"CE",X"DD",X"2E",X"AF",X"63",X"20",
		X"C8",X"31",X"84",X"8E",X"6B",X"84",X"CC",X"92",X"A2",X"20",X"0E",X"34",X"16",X"8E",X"64",X"31",
		X"CC",X"98",X"59",X"9B",X"67",X"DB",X"67",X"20",X"02",X"34",X"16",X"A1",X"24",X"25",X"12",X"E1",
		X"25",X"25",X"0E",X"1F",X"10",X"A1",X"26",X"22",X"0A",X"E1",X"27",X"22",X"06",X"1A",X"01",X"35",
		X"96",X"1C",X"FE",X"35",X"96",X"34",X"17",X"AE",X"28",X"BD",X"15",X"BD",X"E7",X"24",X"EB",X"1C",
		X"25",X"F7",X"E7",X"26",X"C1",X"FE",X"24",X"F1",X"BD",X"15",X"BD",X"86",X"AB",X"3D",X"8B",X"3F",
		X"A7",X"25",X"AB",X"1D",X"25",X"F2",X"A7",X"27",X"81",X"EA",X"24",X"EC",X"BD",X"17",X"C3",X"25",
		X"D6",X"35",X"97",X"CC",X"04",X"E3",X"20",X"03",X"CC",X"04",X"EC",X"DD",X"0A",X"4F",X"5F",X"DD",
		X"3E",X"DD",X"40",X"39",X"CC",X"03",X"0A",X"0D",X"90",X"27",X"03",X"CC",X"02",X"8A",X"DD",X"11",
		X"CC",X"03",X"54",X"DD",X"0A",X"39",X"96",X"6E",X"9B",X"6F",X"9B",X"71",X"39",X"CE",X"00",X"00",
		X"EC",X"24",X"81",X"FE",X"25",X"03",X"33",X"41",X"4F",X"AB",X"1C",X"25",X"04",X"81",X"FE",X"23",
		X"1C",X"33",X"43",X"86",X"FE",X"C1",X"3F",X"24",X"02",X"C6",X"3F",X"C1",X"47",X"22",X"02",X"33",
		X"44",X"EB",X"1D",X"C1",X"EA",X"22",X"14",X"C1",X"E2",X"23",X"14",X"20",X"10",X"C1",X"3F",X"24",
		X"04",X"C6",X"3F",X"33",X"44",X"EB",X"1D",X"C1",X"EA",X"23",X"04",X"C6",X"EA",X"33",X"4C",X"ED",
		X"26",X"A0",X"1C",X"E0",X"1D",X"ED",X"24",X"1F",X"30",X"5D",X"39",X"AC",X"C1",X"26",X"FC",X"6F",
		X"C2",X"6F",X"C2",X"39",X"34",X"07",X"EC",X"1A",X"AF",X"3A",X"A3",X"3A",X"33",X"AB",X"EF",X"3A",
		X"EC",X"1E",X"ED",X"3E",X"EC",X"1C",X"ED",X"3C",X"34",X"06",X"34",X"02",X"8D",X"14",X"EC",X"E4",
		X"A0",X"01",X"E0",X"81",X"ED",X"A1",X"6A",X"62",X"2A",X"F4",X"32",X"63",X"30",X"06",X"31",X"26",
		X"35",X"87",X"44",X"34",X"06",X"25",X"23",X"30",X"86",X"E6",X"84",X"C4",X"F0",X"E7",X"A4",X"E6",
		X"82",X"C4",X"0F",X"EA",X"A4",X"E7",X"A0",X"4A",X"26",X"EF",X"E6",X"80",X"C4",X"F0",X"E7",X"A0",
		X"A6",X"E4",X"30",X"86",X"6A",X"61",X"2A",X"DF",X"35",X"86",X"E6",X"86",X"58",X"C9",X"00",X"58",
		X"C9",X"00",X"58",X"C9",X"00",X"58",X"C9",X"00",X"E7",X"A0",X"4A",X"2A",X"ED",X"6F",X"A0",X"A6",
		X"E4",X"30",X"86",X"30",X"02",X"6A",X"61",X"2A",X"E1",X"35",X"86",X"34",X"27",X"10",X"9E",X"64",
		X"AB",X"22",X"20",X"14",X"34",X"27",X"10",X"9E",X"64",X"1F",X"89",X"84",X"F0",X"C4",X"0F",X"AB",
		X"23",X"19",X"A7",X"23",X"1F",X"98",X"A9",X"22",X"19",X"A7",X"22",X"86",X"01",X"A7",X"24",X"A6",
		X"21",X"89",X"00",X"19",X"A7",X"21",X"A6",X"A4",X"89",X"00",X"19",X"24",X"02",X"8B",X"10",X"A7",
		X"A4",X"96",X"00",X"2A",X"30",X"96",X"6A",X"27",X"06",X"A8",X"21",X"84",X"F0",X"26",X"26",X"EC",
		X"21",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"D1",X"6B",X"25",X"18",X"BD",X"1B",X"34",
		X"0F",X"6A",X"96",X"6B",X"9B",X"1D",X"19",X"97",X"6B",X"24",X"0A",X"A6",X"21",X"84",X"F0",X"8B",
		X"10",X"19",X"4C",X"97",X"6A",X"35",X"A7",X"9A",X"7D",X"1A",X"FC",X"30",X"1D",X"22",X"20",X"1B",
		X"20",X"9A",X"77",X"1A",X"AA",X"9A",X"73",X"14",X"18",X"1A",X"94",X"9A",X"74",X"17",X"18",X"1A",
		X"90",X"9A",X"74",X"1A",X"18",X"1A",X"94",X"9A",X"75",X"1D",X"18",X"1A",X"90",X"9A",X"75",X"20",
		X"18",X"1A",X"94",X"9A",X"76",X"23",X"18",X"1A",X"90",X"00",X"00",X"FF",X"9A",X"76",X"26",X"18",
		X"1A",X"94",X"00",X"00",X"FF",X"9A",X"8B",X"1B",X"0E",X"5A",X"1D",X"7A",X"20",X"1B",X"2A",X"9A",
		X"7C",X"1A",X"AA",X"9A",X"78",X"6C",X"18",X"1A",X"94",X"9A",X"79",X"6F",X"18",X"1A",X"90",X"9A",
		X"79",X"72",X"18",X"1A",X"94",X"9A",X"7A",X"75",X"18",X"1A",X"90",X"9A",X"7A",X"78",X"18",X"1A",
		X"94",X"9A",X"7B",X"7B",X"18",X"1A",X"90",X"00",X"00",X"FF",X"9A",X"7B",X"7E",X"18",X"1A",X"94",
		X"00",X"00",X"FF",X"9A",X"7D",X"1A",X"FC",X"30",X"1D",X"22",X"20",X"1B",X"20",X"9A",X"AF",X"1A",
		X"AA",X"9A",X"AB",X"14",X"18",X"1A",X"94",X"9A",X"AC",X"17",X"18",X"1A",X"90",X"9A",X"AC",X"1A",
		X"18",X"1A",X"94",X"9A",X"AD",X"1D",X"18",X"1A",X"90",X"9A",X"AD",X"20",X"18",X"1A",X"94",X"9A",
		X"AE",X"23",X"18",X"1A",X"90",X"00",X"00",X"FF",X"9A",X"AE",X"26",X"18",X"1A",X"94",X"00",X"00",
		X"FF",X"9E",X"62",X"30",X"88",X"2B",X"AF",X"2B",X"DE",X"62",X"EE",X"42",X"10",X"AE",X"02",X"2B",
		X"0B",X"E6",X"94",X"AD",X"98",X"04",X"AE",X"2B",X"30",X"06",X"20",X"EA",X"BD",X"00",X"5A",X"9E",
		X"62",X"E6",X"94",X"27",X"F7",X"6F",X"94",X"5D",X"2B",X"D7",X"30",X"04",X"E6",X"94",X"26",X"D6",
		X"30",X"06",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"CC",X"30",X"06",X"20",X"C8",X"30",X"0C",
		X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"BE",X"30",X"06",X"20",X"BA",X"30",X"0C",X"20",X"B6",
		X"56",X"56",X"56",X"56",X"C4",X"0F",X"58",X"BE",X"7B",X"18",X"AE",X"85",X"30",X"02",X"CC",X"07",
		X"03",X"1A",X"50",X"BF",X"CA",X"02",X"FD",X"CA",X"06",X"10",X"BF",X"CA",X"04",X"CC",X"12",X"00",
		X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"1F",X"30",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"4F",X"B7",
		X"CA",X"01",X"7E",X"00",X"5A",X"96",X"00",X"84",X"40",X"27",X"06",X"96",X"90",X"26",X"02",X"8D",
		X"1A",X"9E",X"64",X"63",X"04",X"BD",X"00",X"96",X"02",X"9E",X"64",X"6C",X"04",X"BD",X"00",X"96",
		X"07",X"96",X"00",X"84",X"80",X"27",X"03",X"BD",X"1B",X"50",X"39",X"8D",X"02",X"8D",X"E2",X"DC",
		X"64",X"C8",X"0B",X"DD",X"64",X"DC",X"62",X"C8",X"5E",X"DD",X"62",X"39",X"17",X"0D",X"12",X"00",
		X"00",X"00",X"12",X"20",X"09",X"10",X"12",X"AA",X"00",X"00",X"30",X"1D",X"00",X"00",X"17",X"0D",
		X"12",X"00",X"00",X"00",X"6A",X"20",X"09",X"10",X"12",X"AA",X"00",X"00",X"5A",X"1D",X"00",X"00",
		X"12",X"22",X"16",X"21",X"1A",X"22",X"1E",X"23",X"22",X"22",X"6A",X"22",X"6E",X"21",X"72",X"22",
		X"76",X"23",X"7A",X"22",X"34",X"15",X"BD",X"07",X"1B",X"0D",X"C6",X"05",X"BD",X"D2",X"1B",X"D6",
		X"66",X"CB",X"01",X"C2",X"00",X"D7",X"66",X"9E",X"62",X"E7",X"98",X"F6",X"8D",X"02",X"35",X"95",
		X"34",X"77",X"10",X"9E",X"62",X"EE",X"38",X"BD",X"08",X"38",X"A6",X"B8",X"F6",X"81",X"63",X"23",
		X"02",X"86",X"63",X"81",X"0A",X"25",X"12",X"8E",X"64",X"D1",X"EE",X"3A",X"8D",X"29",X"C6",X"CC",
		X"30",X"C9",X"02",X"05",X"BD",X"37",X"C8",X"86",X"09",X"81",X"05",X"2F",X"09",X"8E",X"63",X"2E",
		X"EE",X"3C",X"8D",X"13",X"80",X"05",X"8E",X"61",X"CB",X"10",X"AE",X"3E",X"4A",X"2B",X"06",X"EE",
		X"A1",X"8D",X"04",X"20",X"F7",X"35",X"F7",X"34",X"45",X"1A",X"50",X"FF",X"CA",X"04",X"EE",X"1E",
		X"FF",X"CA",X"06",X"BF",X"CA",X"02",X"C6",X"0A",X"F7",X"CA",X"00",X"35",X"C5",X"35",X"40",X"A6",
		X"C0",X"BD",X"19",X"24",X"E6",X"C4",X"4F",X"7E",X"1E",X"E5",X"1B",X"E5",X"1C",X"0F",X"1C",X"1F",
		X"1C",X"2F",X"1C",X"47",X"1C",X"59",X"1C",X"69",X"1C",X"77",X"1C",X"85",X"1C",X"93",X"1C",X"A3",
		X"1C",X"AF",X"1B",X"FA",X"1C",X"12",X"1C",X"24",X"1C",X"3C",X"1C",X"50",X"1C",X"64",X"1C",X"70",
		X"1C",X"80",X"1C",X"90",X"1C",X"9E",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"00",X"1C",X"F4",X"1D",X"2F",X"1D",X"4D",X"2C",X"FE",X"01",X"C1",X"26",X"82",X"26",X"82",
		X"1C",X"DC",X"2C",X"10",X"1C",X"E8",X"1D",X"17",X"1D",X"4D",X"1C",X"F4",X"1D",X"F9",X"1C",X"BC",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"1C",X"C6",X"1C",X"CE",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"1C",X"C6",X"1C",X"CE",
		X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"2C",X"AC",X"0A",X"8E",
		X"0A",X"8E",X"1D",X"85",X"1D",X"8B",X"1D",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"00",X"00",X"00",X"2B",X"DB",X"2B",X"ED",X"2B",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"27",X"D6",X"27",X"E4",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"1D",X"87",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"01",X"00",X"00",X"1D",X"8D",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"1D",X"81",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",
		X"1D",X"0D",X"1D",X"A4",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"DC",X"40",X"C3",X"02",
		X"00",X"DD",X"40",X"7E",X"1D",X"0D",X"0A",X"6E",X"BD",X"07",X"1B",X"04",X"20",X"06",X"0A",X"6F",
		X"BD",X"07",X"1B",X"08",X"7E",X"1D",X"73",X"31",X"84",X"7E",X"08",X"62",X"9C",X"9F",X"26",X"01",
		X"39",X"C6",X"0A",X"BD",X"36",X"A3",X"20",X"05",X"C6",X"06",X"BD",X"36",X"A3",X"BD",X"07",X"1B",
		X"0E",X"7E",X"15",X"08",X"BD",X"07",X"1B",X"0C",X"C6",X"03",X"BD",X"36",X"A3",X"8D",X"13",X"BD",
		X"17",X"C1",X"30",X"A4",X"24",X"05",X"8D",X"0A",X"BD",X"37",X"E2",X"0A",X"71",X"31",X"84",X"7E",
		X"1D",X"64",X"BD",X"1B",X"AD",X"51",X"46",X"DC",X"3E",X"47",X"56",X"47",X"56",X"D3",X"3E",X"8D",
		X"74",X"DD",X"3E",X"DC",X"40",X"47",X"56",X"47",X"56",X"D3",X"40",X"8D",X"68",X"DD",X"40",X"BD",
		X"07",X"1B",X"0F",X"C6",X"04",X"BD",X"36",X"A3",X"0A",X"6E",X"8D",X"0C",X"BD",X"17",X"C1",X"24",
		X"23",X"8D",X"05",X"BD",X"37",X"E2",X"20",X"1C",X"BD",X"1B",X"AD",X"02",X"3C",X"BD",X"07",X"1B",
		X"0C",X"C6",X"02",X"BD",X"36",X"A3",X"0A",X"6F",X"8D",X"20",X"BD",X"17",X"C1",X"24",X"05",X"BD",
		X"37",X"E2",X"8D",X"16",X"34",X"10",X"BD",X"08",X"68",X"BD",X"00",X"47",X"30",X"A4",X"BD",X"01",
		X"AB",X"35",X"90",X"1E",X"12",X"8D",X"ED",X"7E",X"1C",X"D7",X"BD",X"1B",X"AD",X"51",X"2D",X"31",
		X"84",X"0A",X"71",X"20",X"0A",X"31",X"84",X"0A",X"6E",X"20",X"04",X"31",X"84",X"0A",X"6F",X"BD",
		X"07",X"1B",X"03",X"20",X"CF",X"81",X"40",X"2D",X"03",X"CC",X"40",X"00",X"81",X"C0",X"2C",X"03",
		X"CC",X"C0",X"00",X"39",X"BD",X"1D",X"0D",X"EC",X"A8",X"10",X"83",X"26",X"5D",X"26",X"07",X"DE",
		X"9C",X"2A",X"03",X"BD",X"18",X"9B",X"0C",X"9E",X"86",X"20",X"BD",X"19",X"1B",X"BD",X"07",X"1B",
		X"03",X"BD",X"00",X"A5",X"1D",X"D4",X"4D",X"01",X"1D",X"E2",X"8E",X"47",X"84",X"AF",X"2B",X"86",
		X"40",X"A7",X"2D",X"39",X"0F",X"9E",X"5F",X"AE",X"2B",X"86",X"20",X"BD",X"7B",X"0F",X"4F",X"7E",
		X"7B",X"0F",X"8D",X"F2",X"6A",X"2D",X"26",X"05",X"8D",X"EA",X"7E",X"00",X"89",X"6A",X"2C",X"C6",
		X"44",X"8D",X"E4",X"4F",X"BD",X"00",X"5C",X"20",X"E9",X"BD",X"1F",X"2D",X"DD",X"32",X"A0",X"04",
		X"10",X"2B",X"00",X"A0",X"81",X"13",X"10",X"22",X"00",X"9A",X"E0",X"05",X"10",X"2B",X"00",X"94",
		X"C1",X"0B",X"10",X"22",X"00",X"8E",X"FE",X"3B",X"E2",X"58",X"33",X"C5",X"A1",X"C4",X"10",X"25",
		X"00",X"82",X"A1",X"41",X"10",X"22",X"00",X"7C",X"96",X"67",X"81",X"12",X"25",X"30",X"BD",X"18",
		X"23",X"BD",X"07",X"1B",X"10",X"86",X"25",X"BD",X"19",X"1B",X"D6",X"90",X"27",X"10",X"CE",X"35",
		X"2E",X"C6",X"0D",X"BD",X"36",X"A3",X"26",X"03",X"CE",X"35",X"7C",X"7E",X"36",X"73",X"0C",X"69",
		X"27",X"FC",X"96",X"15",X"49",X"BD",X"11",X"A4",X"13",X"A5",X"10",X"25",X"E2",X"2B",X"BD",X"07",
		X"1B",X"03",X"BD",X"18",X"23",X"6F",X"E2",X"BD",X"1F",X"2D",X"80",X"7E",X"8B",X"01",X"81",X"02",
		X"25",X"0C",X"49",X"86",X"01",X"25",X"01",X"40",X"9B",X"36",X"97",X"36",X"6C",X"E4",X"C0",X"92",
		X"CB",X"01",X"C1",X"02",X"25",X"0C",X"59",X"C6",X"01",X"25",X"01",X"50",X"DB",X"37",X"D7",X"37",
		X"6C",X"E4",X"6D",X"E0",X"26",X"08",X"C6",X"01",X"BD",X"36",X"A3",X"7E",X"15",X"08",X"4F",X"BD",
		X"00",X"5C",X"20",X"C1",X"CC",X"7E",X"92",X"90",X"32",X"D0",X"33",X"BD",X"16",X"C7",X"A7",X"E2",
		X"86",X"C8",X"58",X"3D",X"2A",X"02",X"80",X"C8",X"E6",X"E4",X"A7",X"E4",X"86",X"C8",X"58",X"3D",
		X"2A",X"02",X"80",X"C8",X"1F",X"89",X"1D",X"D3",X"3E",X"BD",X"1D",X"95",X"DD",X"3E",X"E6",X"E0",
		X"1D",X"D3",X"40",X"BD",X"1D",X"95",X"DD",X"40",X"39",X"86",X"C0",X"B7",X"99",X"E2",X"B7",X"99",
		X"E7",X"B7",X"99",X"EC",X"39",X"34",X"37",X"0F",X"2E",X"DC",X"67",X"81",X"12",X"24",X"02",X"03",
		X"2E",X"E3",X"61",X"81",X"18",X"23",X"02",X"86",X"18",X"81",X"0C",X"24",X"02",X"86",X"0C",X"DD",
		X"67",X"5F",X"81",X"12",X"25",X"0A",X"96",X"2E",X"27",X"04",X"BD",X"07",X"1B",X"12",X"C6",X"21",
		X"D7",X"89",X"35",X"B7",X"86",X"0A",X"BD",X"00",X"5C",X"CC",X"FF",X"00",X"BD",X"1E",X"E5",X"86",
		X"05",X"BD",X"00",X"5C",X"96",X"00",X"84",X"EF",X"97",X"00",X"7E",X"00",X"89",X"34",X"05",X"96",
		X"67",X"44",X"9B",X"37",X"9B",X"57",X"A7",X"61",X"96",X"67",X"44",X"9B",X"36",X"9B",X"56",X"35",
		X"85",X"34",X"07",X"96",X"67",X"5F",X"40",X"47",X"56",X"34",X"06",X"AB",X"63",X"90",X"56",X"1A",
		X"50",X"DD",X"3A",X"97",X"36",X"35",X"06",X"AB",X"62",X"90",X"57",X"DD",X"3C",X"97",X"37",X"35",
		X"87",X"86",X"05",X"BD",X"01",X"13",X"7E",X"01",X"27",X"9E",X"40",X"DC",X"3E",X"26",X"04",X"30",
		X"84",X"27",X"18",X"58",X"49",X"29",X"0F",X"1E",X"10",X"58",X"49",X"29",X"04",X"1E",X"10",X"20",
		X"F2",X"46",X"1E",X"01",X"47",X"49",X"46",X"34",X"10",X"E6",X"E1",X"39",X"8D",X"DB",X"7E",X"16",
		X"C7",X"34",X"50",X"96",X"00",X"85",X"08",X"27",X"5D",X"8D",X"F1",X"DD",X"2C",X"26",X"04",X"C6",
		X"40",X"D7",X"2D",X"C6",X"FE",X"81",X"CE",X"2D",X"18",X"5C",X"81",X"EC",X"2D",X"0D",X"5C",X"81",
		X"14",X"2D",X"08",X"5C",X"81",X"32",X"2D",X"03",X"5C",X"20",X"06",X"96",X"2D",X"2B",X"02",X"CB",
		X"04",X"8E",X"23",X"4E",X"58",X"58",X"30",X"85",X"EE",X"84",X"DF",X"42",X"96",X"67",X"44",X"97",
		X"2F",X"49",X"D6",X"2C",X"3D",X"2A",X"02",X"90",X"67",X"58",X"49",X"9B",X"56",X"9B",X"2F",X"A0",
		X"02",X"97",X"5A",X"96",X"67",X"D6",X"2D",X"3D",X"2A",X"02",X"90",X"67",X"58",X"49",X"9B",X"57",
		X"9B",X"2F",X"A0",X"03",X"97",X"5B",X"1C",X"EF",X"10",X"9E",X"1B",X"35",X"D0",X"32",X"61",X"86",
		X"04",X"BD",X"00",X"5C",X"1A",X"50",X"D6",X"1A",X"C8",X"50",X"D7",X"1C",X"31",X"2B",X"D6",X"67",
		X"8E",X"23",X"88",X"58",X"EE",X"85",X"1C",X"EF",X"DF",X"46",X"CE",X"23",X"A2",X"EE",X"C5",X"DF",
		X"4A",X"CE",X"23",X"14",X"33",X"C5",X"A6",X"C0",X"AE",X"86",X"9F",X"48",X"5F",X"44",X"97",X"55",
		X"90",X"67",X"47",X"56",X"ED",X"28",X"37",X"02",X"A7",X"2A",X"DC",X"3A",X"9B",X"56",X"ED",X"A4",
		X"DC",X"3C",X"9B",X"57",X"ED",X"22",X"DC",X"3E",X"E6",X"2A",X"40",X"3D",X"2A",X"02",X"A0",X"2A",
		X"E3",X"A4",X"A3",X"28",X"ED",X"24",X"DC",X"40",X"E6",X"2A",X"40",X"3D",X"2A",X"02",X"A0",X"2A",
		X"E3",X"22",X"A3",X"28",X"ED",X"26",X"9E",X"48",X"AE",X"1C",X"DE",X"46",X"EE",X"5C",X"A0",X"22",
		X"10",X"22",X"00",X"B9",X"40",X"97",X"57",X"A7",X"E2",X"9B",X"67",X"4A",X"97",X"45",X"A6",X"A4",
		X"97",X"3A",X"A0",X"24",X"23",X"55",X"97",X"56",X"9B",X"67",X"4A",X"97",X"44",X"4F",X"5F",X"DD",
		X"58",X"EC",X"24",X"DD",X"3A",X"BD",X"1F",X"91",X"20",X"04",X"EC",X"81",X"ED",X"A1",X"6A",X"E4",
		X"2A",X"F8",X"96",X"55",X"90",X"57",X"27",X"1A",X"A7",X"E4",X"37",X"06",X"9B",X"56",X"DB",X"56",
		X"A1",X"80",X"23",X"02",X"A6",X"1F",X"E1",X"80",X"24",X"02",X"A6",X"1F",X"ED",X"A1",X"6A",X"E4",
		X"26",X"E8",X"96",X"67",X"9B",X"57",X"90",X"55",X"27",X"0E",X"A7",X"E4",X"37",X"06",X"9B",X"56",
		X"DB",X"56",X"ED",X"A1",X"6A",X"E4",X"26",X"F4",X"7E",X"1F",X"FD",X"40",X"5F",X"D7",X"56",X"DD",
		X"58",X"9B",X"55",X"91",X"67",X"2C",X"02",X"96",X"67",X"4A",X"97",X"44",X"BD",X"1F",X"91",X"20",
		X"08",X"EC",X"81",X"9B",X"58",X"DB",X"58",X"ED",X"A1",X"6A",X"E4",X"2A",X"F4",X"96",X"55",X"90",
		X"57",X"27",X"1A",X"A7",X"E4",X"EC",X"81",X"9B",X"58",X"DB",X"58",X"A1",X"C0",X"23",X"02",X"A6",
		X"5F",X"E1",X"C0",X"24",X"02",X"E6",X"5F",X"ED",X"A1",X"6A",X"E4",X"26",X"E8",X"96",X"67",X"9B",
		X"57",X"90",X"55",X"37",X"10",X"AF",X"A1",X"4A",X"26",X"F9",X"7E",X"1F",X"FD",X"97",X"59",X"A7",
		X"E2",X"9B",X"55",X"91",X"67",X"2C",X"02",X"96",X"67",X"4A",X"97",X"45",X"A6",X"22",X"97",X"3C",
		X"A6",X"A4",X"97",X"3A",X"A0",X"24",X"10",X"23",X"00",X"88",X"97",X"56",X"9B",X"67",X"4A",X"97",
		X"44",X"A6",X"24",X"97",X"3A",X"4F",X"5F",X"DD",X"57",X"BD",X"1F",X"91",X"20",X"08",X"37",X"06",
		X"9B",X"56",X"DB",X"56",X"ED",X"A1",X"6A",X"E4",X"2A",X"F4",X"96",X"67",X"90",X"59",X"91",X"55",
		X"2E",X"2E",X"A7",X"E4",X"27",X"18",X"37",X"06",X"9B",X"56",X"DB",X"56",X"A1",X"80",X"23",X"02",
		X"A6",X"1F",X"E1",X"80",X"24",X"02",X"E6",X"1F",X"ED",X"A1",X"6A",X"E4",X"26",X"E8",X"96",X"55",
		X"9B",X"59",X"90",X"67",X"27",X"07",X"EE",X"81",X"EF",X"A1",X"4A",X"26",X"F9",X"7E",X"1F",X"FD",
		X"96",X"55",X"A7",X"E4",X"37",X"06",X"9B",X"56",X"DB",X"56",X"A1",X"80",X"23",X"02",X"A6",X"1F",
		X"E1",X"80",X"24",X"02",X"E6",X"1F",X"ED",X"A1",X"6A",X"E4",X"26",X"E8",X"96",X"67",X"90",X"55",
		X"90",X"59",X"A7",X"E4",X"37",X"06",X"9B",X"56",X"DB",X"56",X"ED",X"A1",X"6A",X"E4",X"26",X"F4",
		X"20",X"CB",X"40",X"97",X"58",X"9B",X"55",X"91",X"67",X"2C",X"02",X"96",X"67",X"4A",X"97",X"44",
		X"4F",X"5F",X"DD",X"56",X"BD",X"1F",X"91",X"20",X"04",X"37",X"06",X"ED",X"A1",X"6A",X"E4",X"2A",
		X"F8",X"96",X"67",X"90",X"59",X"91",X"55",X"2E",X"33",X"A7",X"E4",X"EC",X"81",X"9B",X"58",X"DB",
		X"58",X"A1",X"C0",X"23",X"02",X"A6",X"5F",X"E1",X"C0",X"24",X"02",X"E6",X"5F",X"ED",X"A1",X"6A",
		X"E4",X"26",X"E8",X"96",X"55",X"9B",X"59",X"90",X"67",X"27",X"0E",X"A7",X"E4",X"EC",X"81",X"9B",
		X"58",X"DB",X"58",X"ED",X"A1",X"6A",X"E4",X"26",X"F4",X"7E",X"1F",X"FD",X"96",X"55",X"A7",X"E4",
		X"EC",X"81",X"9B",X"58",X"DB",X"58",X"A1",X"C0",X"23",X"02",X"A6",X"5F",X"E1",X"C0",X"24",X"02",
		X"E6",X"5F",X"ED",X"A1",X"6A",X"E4",X"26",X"E8",X"96",X"67",X"90",X"55",X"90",X"59",X"37",X"10",
		X"AF",X"A1",X"4A",X"26",X"F9",X"20",X"D2",X"6A",X"A8",X"14",X"10",X"27",X"0E",X"AB",X"6C",X"A8",
		X"13",X"EC",X"A8",X"12",X"BD",X"16",X"23",X"9B",X"60",X"DB",X"61",X"ED",X"24",X"39",X"57",X"31",
		X"57",X"41",X"57",X"4E",X"57",X"5E",X"57",X"6A",X"57",X"7A",X"57",X"86",X"57",X"96",X"57",X"A3",
		X"57",X"B3",X"57",X"C0",X"57",X"D0",X"56",X"F8",X"57",X"08",X"57",X"14",X"57",X"24",X"00",X"00",
		X"00",X"00",X"22",X"57",X"38",X"1D",X"00",X"00",X"1E",X"BD",X"15",X"B9",X"CA",X"01",X"84",X"3F",
		X"34",X"06",X"34",X"02",X"BD",X"01",X"C3",X"17",X"0A",X"0F",X"22",X"8E",X"DC",X"60",X"ED",X"24",
		X"ED",X"26",X"A6",X"E4",X"48",X"48",X"A7",X"A8",X"12",X"E6",X"E4",X"54",X"54",X"C9",X"00",X"C4",
		X"0F",X"58",X"8E",X"22",X"6E",X"AE",X"85",X"AF",X"28",X"BD",X"18",X"4D",X"27",X"05",X"BD",X"01",
		X"A9",X"20",X"04",X"4F",X"BD",X"08",X"15",X"BD",X"00",X"5A",X"A6",X"E4",X"AB",X"62",X"84",X"3F",
		X"A7",X"E4",X"A1",X"61",X"26",X"BE",X"32",X"63",X"96",X"90",X"27",X"01",X"39",X"86",X"1E",X"BD",
		X"00",X"5C",X"20",X"17",X"8D",X"0C",X"96",X"00",X"84",X"F7",X"97",X"00",X"86",X"C0",X"B7",X"99",
		X"EC",X"39",X"34",X"77",X"CE",X"99",X"EC",X"C6",X"01",X"20",X"07",X"34",X"77",X"CE",X"99",X"E2",
		X"C6",X"03",X"1A",X"50",X"37",X"32",X"10",X"BF",X"CA",X"04",X"BF",X"CA",X"02",X"AE",X"1E",X"BF",
		X"CA",X"06",X"8A",X"10",X"B7",X"CA",X"00",X"5A",X"26",X"EA",X"35",X"F7",X"12",X"14",X"14",X"16",
		X"16",X"18",X"18",X"19",X"1A",X"1A",X"1C",X"1B",X"1E",X"1C",X"20",X"1D",X"22",X"1E",X"24",X"1F",
		X"26",X"20",X"28",X"21",X"2A",X"22",X"56",X"C4",X"05",X"02",X"56",X"DC",X"05",X"05",X"56",X"2C",
		X"02",X"05",X"56",X"42",X"01",X"05",X"56",X"5E",X"00",X"02",X"56",X"A8",X"05",X"00",X"56",X"92",
		X"02",X"00",X"56",X"76",X"00",X"00",X"CE",X"23",X"79",X"AE",X"C1",X"EC",X"C1",X"80",X"35",X"88",
		X"5A",X"BD",X"7B",X"00",X"A6",X"C0",X"26",X"F5",X"39",X"10",X"F8",X"A5",X"11",X"8C",X"A6",X"85",
		X"B0",X"7E",X"81",X"81",X"7E",X"86",X"82",X"7C",X"85",X"8A",X"81",X"8A",X"8C",X"79",X"7B",X"78",
		X"77",X"7E",X"8C",X"7C",X"85",X"7E",X"77",X"8C",X"A9",X"00",X"61",X"CB",X"62",X"0E",X"62",X"62",
		X"62",X"BE",X"63",X"2E",X"63",X"A7",X"64",X"37",X"64",X"D1",X"65",X"85",X"66",X"44",X"67",X"20",
		X"68",X"08",X"69",X"10",X"6A",X"25",X"6B",X"5D",X"6C",X"A3",X"6E",X"0D",X"6E",X"4B",X"6E",X"8F",
		X"6E",X"E5",X"6F",X"42",X"6F",X"B4",X"70",X"2E",X"70",X"C0",X"71",X"5B",X"72",X"11",X"72",X"D1",
		X"73",X"AF",X"74",X"98",X"49",X"4A",X"00",X"00",X"02",X"FF",X"24",X"7E",X"2E",X"61",X"BD",X"17",
		X"CB",X"25",X"1B",X"8E",X"70",X"3F",X"CC",X"8C",X"A2",X"BD",X"17",X"D9",X"25",X"10",X"A6",X"25",
		X"90",X"67",X"81",X"49",X"25",X"08",X"A6",X"63",X"BD",X"08",X"15",X"BD",X"08",X"62",X"39",X"BD",
		X"01",X"C3",X"1C",X"08",X"0E",X"23",X"D4",X"6F",X"A8",X"18",X"6F",X"A8",X"19",X"39",X"34",X"77",
		X"E6",X"61",X"27",X"39",X"CB",X"02",X"58",X"4F",X"BD",X"01",X"63",X"9F",X"9C",X"34",X"10",X"BD",
		X"00",X"A5",X"24",X"4F",X"4D",X"0A",X"24",X"54",X"8D",X"D5",X"AE",X"E4",X"10",X"AF",X"81",X"AF",
		X"E4",X"BD",X"17",X"F5",X"5F",X"BD",X"23",X"DE",X"25",X"F7",X"96",X"04",X"A7",X"2A",X"BD",X"15",
		X"B9",X"BD",X"25",X"16",X"6A",X"63",X"26",X"E0",X"CC",X"00",X"01",X"ED",X"F1",X"35",X"F7",X"9E",
		X"9C",X"7E",X"01",X"AB",X"CE",X"FF",X"FF",X"EF",X"2F",X"DE",X"9C",X"EF",X"2D",X"BD",X"00",X"5A",
		X"EE",X"2D",X"AE",X"C1",X"27",X"FC",X"2A",X"0F",X"BD",X"2D",X"99",X"10",X"A3",X"2F",X"24",X"EB",
		X"AF",X"A8",X"11",X"ED",X"2F",X"20",X"E4",X"AE",X"A8",X"11",X"9F",X"9A",X"20",X"D6",X"10",X"9C",
		X"9A",X"26",X"11",X"6A",X"A8",X"19",X"2A",X"0C",X"DC",X"36",X"BD",X"25",X"16",X"DE",X"79",X"A6",
		X"42",X"A7",X"A8",X"19",X"A6",X"A8",X"18",X"6C",X"A8",X"18",X"4D",X"27",X"19",X"2B",X"12",X"90",
		X"8E",X"2B",X"26",X"48",X"8E",X"24",X"A9",X"6E",X"96",X"24",X"C4",X"24",X"E4",X"24",X"F2",X"25",
		X"0D",X"6C",X"A8",X"18",X"20",X"00",X"8E",X"48",X"06",X"A6",X"A8",X"12",X"2A",X"03",X"8E",X"48",
		X"A8",X"AF",X"28",X"39",X"8E",X"49",X"4A",X"AF",X"28",X"A6",X"24",X"E6",X"A8",X"16",X"E3",X"A8",
		X"12",X"A7",X"24",X"E7",X"A8",X"16",X"A6",X"25",X"E6",X"A8",X"17",X"E3",X"A8",X"14",X"A7",X"25",
		X"E7",X"A8",X"17",X"39",X"8E",X"48",X"A8",X"A6",X"A8",X"12",X"2A",X"03",X"8E",X"48",X"06",X"AF",
		X"28",X"39",X"A6",X"24",X"E6",X"A8",X"16",X"A3",X"A8",X"12",X"A7",X"24",X"E7",X"A8",X"16",X"A6",
		X"25",X"E6",X"A8",X"17",X"A3",X"A8",X"14",X"A7",X"25",X"E7",X"A8",X"17",X"39",X"6F",X"A8",X"18",
		X"8E",X"49",X"4A",X"AF",X"28",X"39",X"A0",X"24",X"46",X"97",X"2C",X"2A",X"02",X"03",X"2C",X"E0",
		X"25",X"56",X"2B",X"08",X"D1",X"2C",X"23",X"02",X"D6",X"2C",X"20",X"08",X"53",X"D1",X"2C",X"23",
		X"02",X"D6",X"2C",X"53",X"BD",X"16",X"C7",X"34",X"06",X"96",X"75",X"D6",X"05",X"3D",X"9B",X"74",
		X"97",X"2C",X"E6",X"E0",X"3D",X"2A",X"02",X"90",X"2C",X"47",X"56",X"47",X"56",X"ED",X"A8",X"12",
		X"96",X"2C",X"E6",X"E0",X"3D",X"2A",X"02",X"90",X"2C",X"47",X"56",X"47",X"56",X"ED",X"A8",X"14",
		X"39",X"86",X"7E",X"C5",X"04",X"26",X"05",X"BD",X"15",X"BD",X"20",X"09",X"C5",X"01",X"26",X"03",
		X"BD",X"15",X"B9",X"C6",X"92",X"A0",X"24",X"E0",X"25",X"BD",X"25",X"97",X"40",X"50",X"BD",X"15",
		X"DA",X"E7",X"A8",X"1C",X"EC",X"A8",X"1C",X"BD",X"16",X"23",X"40",X"AB",X"24",X"A7",X"A8",X"17",
		X"50",X"EB",X"25",X"E7",X"A8",X"19",X"39",X"34",X"17",X"BD",X"16",X"C7",X"DD",X"32",X"9E",X"79",
		X"BD",X"15",X"BD",X"96",X"1E",X"3D",X"E6",X"04",X"3D",X"AB",X"03",X"97",X"2F",X"D6",X"32",X"3D",
		X"2A",X"02",X"90",X"2F",X"47",X"56",X"47",X"56",X"ED",X"A8",X"12",X"96",X"2F",X"D6",X"33",X"3D",
		X"2A",X"02",X"90",X"2F",X"47",X"56",X"47",X"56",X"ED",X"A8",X"14",X"35",X"97",X"EC",X"A8",X"17",
		X"E3",X"A8",X"12",X"ED",X"A8",X"17",X"EC",X"A8",X"19",X"E3",X"A8",X"14",X"ED",X"A8",X"19",X"EC",
		X"A8",X"1C",X"AB",X"A8",X"1B",X"A7",X"A8",X"1C",X"BD",X"16",X"23",X"AB",X"A8",X"17",X"EB",X"A8",
		X"19",X"ED",X"24",X"CE",X"49",X"DF",X"E6",X"A8",X"16",X"5C",X"E7",X"A8",X"16",X"C4",X"10",X"27",
		X"03",X"CE",X"4A",X"3D",X"EF",X"28",X"39",X"49",X"DF",X"00",X"00",X"03",X"FF",X"25",X"CD",X"25",
		X"61",X"34",X"77",X"6A",X"61",X"2A",X"02",X"35",X"F7",X"BD",X"01",X"C3",X"20",X"08",X"0E",X"26",
		X"07",X"BD",X"17",X"F5",X"9E",X"79",X"A6",X"06",X"BD",X"15",X"BD",X"3D",X"D6",X"1E",X"3D",X"AB",
		X"05",X"BD",X"15",X"BD",X"5D",X"2A",X"01",X"40",X"A7",X"A8",X"1B",X"A6",X"08",X"BD",X"15",X"BD",
		X"E7",X"A8",X"16",X"3D",X"AB",X"07",X"A7",X"A8",X"1D",X"BD",X"15",X"B9",X"BD",X"25",X"97",X"BD",
		X"15",X"BD",X"BD",X"25",X"81",X"BD",X"23",X"DE",X"25",X"C7",X"7E",X"26",X"13",X"BD",X"15",X"B9",
		X"BD",X"25",X"16",X"C6",X"02",X"8E",X"24",X"7E",X"CE",X"2E",X"61",X"E7",X"2C",X"86",X"FF",X"A7",
		X"2D",X"AF",X"2E",X"EF",X"A8",X"10",X"6E",X"C4",X"8E",X"25",X"CD",X"CE",X"25",X"61",X"C6",X"03",
		X"20",X"E9",X"96",X"00",X"85",X"10",X"26",X"21",X"D6",X"67",X"C1",X"12",X"24",X"10",X"C6",X"07",
		X"A6",X"0C",X"81",X"02",X"27",X"02",X"C6",X"08",X"BD",X"36",X"A3",X"7E",X"1C",X"ED",X"8A",X"10",
		X"97",X"00",X"BD",X"00",X"AD",X"39",X"0F",X"1F",X"14",X"86",X"FC",X"A7",X"0D",X"86",X"30",X"BD",
		X"19",X"24",X"BD",X"07",X"1B",X"11",X"A6",X"0C",X"C6",X"0B",X"BD",X"36",X"A3",X"81",X"02",X"27",
		X"08",X"60",X"88",X"1B",X"CC",X"26",X"78",X"20",X"03",X"CC",X"26",X"5D",X"ED",X"88",X"10",X"BD",
		X"1F",X"2D",X"DD",X"32",X"EC",X"04",X"AB",X"06",X"46",X"EB",X"07",X"56",X"90",X"32",X"D0",X"33",
		X"BD",X"16",X"C7",X"D7",X"2F",X"CE",X"4A",X"3D",X"E6",X"0C",X"C1",X"02",X"26",X"09",X"CE",X"48",
		X"06",X"4D",X"2A",X"03",X"CE",X"48",X"A8",X"31",X"84",X"BD",X"08",X"68",X"EF",X"08",X"5F",X"47",
		X"56",X"47",X"56",X"47",X"56",X"ED",X"88",X"12",X"96",X"2F",X"5F",X"47",X"56",X"47",X"56",X"47",
		X"56",X"ED",X"88",X"14",X"CC",X"24",X"C9",X"ED",X"0E",X"86",X"0C",X"A7",X"0C",X"39",X"4A",X"9D",
		X"00",X"00",X"08",X"FF",X"27",X"2A",X"01",X"C1",X"00",X"80",X"A6",X"A8",X"18",X"AB",X"2A",X"A7",
		X"2A",X"7E",X"24",X"C9",X"34",X"77",X"6A",X"61",X"2B",X"0C",X"BD",X"01",X"C3",X"1B",X"08",X"08",
		X"27",X"1E",X"8D",X"04",X"20",X"F0",X"35",X"F7",X"BD",X"17",X"F5",X"A6",X"63",X"BD",X"08",X"15",
		X"BD",X"08",X"62",X"CC",X"7C",X"90",X"E0",X"25",X"34",X"04",X"2A",X"01",X"50",X"A0",X"24",X"34",
		X"06",X"2A",X"01",X"40",X"34",X"02",X"A1",X"62",X"CC",X"01",X"00",X"24",X"14",X"6D",X"63",X"2A",
		X"01",X"40",X"ED",X"A8",X"14",X"A6",X"68",X"E6",X"62",X"8D",X"19",X"ED",X"A8",X"12",X"32",X"64",
		X"39",X"6D",X"61",X"2A",X"01",X"40",X"ED",X"A8",X"12",X"A6",X"68",X"E6",X"E1",X"8D",X"05",X"ED",
		X"A8",X"14",X"35",X"86",X"34",X"02",X"68",X"63",X"58",X"28",X"FB",X"6F",X"E2",X"86",X"01",X"34",
		X"06",X"CC",X"80",X"00",X"64",X"61",X"66",X"62",X"10",X"A3",X"61",X"25",X"02",X"A3",X"61",X"69",
		X"E4",X"24",X"F1",X"A6",X"E4",X"43",X"32",X"63",X"E6",X"63",X"3D",X"58",X"49",X"E6",X"E4",X"A7",
		X"E2",X"3D",X"C6",X"B0",X"3D",X"AB",X"61",X"A7",X"A8",X"18",X"E6",X"E1",X"4F",X"6D",X"63",X"2A",
		X"04",X"43",X"50",X"82",X"FF",X"39",X"34",X"20",X"BD",X"01",X"C3",X"1B",X"08",X"0E",X"28",X"50",
		X"0C",X"6E",X"20",X"0C",X"34",X"20",X"BD",X"01",X"C3",X"1B",X"08",X"08",X"27",X"1E",X"0C",X"6F",
		X"CC",X"00",X"FD",X"E7",X"0D",X"E7",X"2D",X"E6",X"88",X"18",X"34",X"07",X"EE",X"08",X"EC",X"88",
		X"12",X"47",X"56",X"47",X"56",X"D7",X"2F",X"EC",X"88",X"14",X"47",X"56",X"47",X"56",X"96",X"2F",
		X"BD",X"16",X"C7",X"DD",X"32",X"50",X"8D",X"12",X"31",X"84",X"BD",X"00",X"47",X"BD",X"08",X"68",
		X"DC",X"32",X"40",X"8D",X"05",X"35",X"27",X"7E",X"08",X"62",X"34",X"02",X"86",X"1C",X"5D",X"3D",
		X"2A",X"02",X"80",X"1C",X"AB",X"04",X"A7",X"24",X"AB",X"5C",X"A7",X"26",X"86",X"1C",X"E6",X"E0",
		X"3D",X"2A",X"02",X"80",X"1C",X"AB",X"05",X"A7",X"25",X"AB",X"5D",X"A7",X"27",X"7E",X"27",X"4B",
		X"4A",X"C1",X"00",X"00",X"07",X"FF",X"27",X"2A",X"01",X"C1",X"34",X"77",X"6A",X"61",X"2B",X"0D",
		X"BD",X"01",X"C3",X"1B",X"08",X"0E",X"28",X"50",X"BD",X"27",X"48",X"20",X"EF",X"35",X"F7",X"EC",
		X"24",X"6D",X"A8",X"13",X"26",X"0E",X"81",X"7A",X"25",X"32",X"C1",X"8E",X"C6",X"01",X"25",X"02",
		X"C6",X"03",X"20",X"1A",X"81",X"7A",X"23",X"F2",X"20",X"22",X"A6",X"A8",X"13",X"46",X"46",X"EC",
		X"24",X"25",X"15",X"C1",X"8E",X"25",X"15",X"5F",X"81",X"7A",X"23",X"02",X"C6",X"02",X"E7",X"A8",
		X"13",X"CC",X"28",X"AC",X"ED",X"2E",X"20",X"04",X"C1",X"8E",X"23",X"EB",X"6C",X"A8",X"12",X"EC",
		X"A8",X"12",X"58",X"EB",X"A8",X"13",X"58",X"8E",X"28",X"C8",X"3A",X"84",X"01",X"48",X"EE",X"86",
		X"EF",X"28",X"E6",X"A8",X"14",X"6E",X"98",X"04",X"54",X"9A",X"54",X"D8",X"28",X"E0",X"55",X"16",
		X"55",X"58",X"28",X"F0",X"55",X"9A",X"55",X"D8",X"28",X"E7",X"54",X"16",X"54",X"58",X"28",X"F7",
		X"A6",X"24",X"E3",X"A8",X"15",X"20",X"05",X"A6",X"24",X"A3",X"A8",X"15",X"A7",X"24",X"20",X"0E",
		X"A6",X"25",X"E3",X"A8",X"15",X"20",X"05",X"A6",X"25",X"A3",X"A8",X"15",X"A7",X"25",X"E7",X"A8",
		X"14",X"6A",X"A8",X"17",X"27",X"01",X"39",X"96",X"78",X"26",X"13",X"BD",X"15",X"BD",X"86",X"32",
		X"3D",X"8B",X"0F",X"A7",X"A8",X"17",X"BD",X"15",X"BD",X"C4",X"03",X"E7",X"A8",X"13",X"39",X"54",
		X"16",X"00",X"00",X"09",X"FF",X"28",X"AC",X"29",X"07",X"0F",X"78",X"D6",X"71",X"34",X"04",X"26",
		X"03",X"7E",X"00",X"89",X"BD",X"01",X"C3",X"1A",X"08",X"0E",X"29",X"1F",X"DE",X"79",X"A6",X"4C",
		X"BD",X"15",X"BD",X"3D",X"D6",X"1E",X"3D",X"AB",X"4B",X"44",X"56",X"44",X"56",X"44",X"56",X"44",
		X"56",X"ED",X"A8",X"15",X"8D",X"B1",X"CE",X"29",X"CB",X"58",X"EE",X"C5",X"EF",X"24",X"EF",X"26",
		X"4F",X"BD",X"08",X"15",X"BD",X"15",X"BD",X"54",X"DE",X"79",X"A6",X"4E",X"3D",X"BD",X"15",X"BD",
		X"54",X"24",X"01",X"40",X"AB",X"4E",X"BD",X"00",X"5C",X"6A",X"E4",X"26",X"B7",X"9E",X"79",X"A6",
		X"0D",X"BD",X"01",X"48",X"86",X"01",X"97",X"78",X"8E",X"9A",X"01",X"AE",X"84",X"8C",X"9A",X"07",
		X"27",X"9F",X"A6",X"0C",X"81",X"09",X"26",X"F3",X"CE",X"28",X"8A",X"CC",X"7A",X"8E",X"E0",X"05",
		X"56",X"E7",X"E2",X"2A",X"01",X"50",X"E7",X"E2",X"C6",X"01",X"A0",X"04",X"46",X"97",X"2F",X"2A",
		X"01",X"40",X"A1",X"E0",X"22",X"08",X"96",X"2F",X"A7",X"E4",X"5F",X"CE",X"28",X"6F",X"A6",X"E0",
		X"2A",X"02",X"CA",X"02",X"E7",X"88",X"13",X"EF",X"0E",X"20",X"C0",X"92",X"92",X"7E",X"A2",X"63",
		X"92",X"7E",X"7C",X"7E",X"92",X"00",X"00",X"4D",X"32",X"00",X"00",X"05",X"FF",X"2B",X"1D",X"2B",
		X"93",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"0F",X"76",
		X"0F",X"77",X"BD",X"00",X"A5",X"2D",X"86",X"2F",X"0D",X"2D",X"B4",X"9E",X"7B",X"AE",X"0C",X"A6",
		X"80",X"26",X"03",X"7E",X"00",X"89",X"84",X"7F",X"81",X"10",X"24",X"07",X"84",X"0F",X"BD",X"01",
		X"48",X"20",X"EC",X"1F",X"89",X"CE",X"2A",X"2E",X"6D",X"1F",X"2A",X"03",X"CE",X"2D",X"31",X"84",
		X"0F",X"C4",X"F0",X"BD",X"01",X"48",X"AD",X"C4",X"C0",X"10",X"26",X"F3",X"20",X"D1",X"34",X"77",
		X"BD",X"00",X"A5",X"2A",X"E5",X"39",X"0E",X"2A",X"61",X"33",X"A4",X"BD",X"01",X"C3",X"23",X"04",
		X"1F",X"29",X"D3",X"10",X"AF",X"4B",X"EF",X"A8",X"1F",X"4F",X"BD",X"08",X"15",X"BD",X"15",X"BD",
		X"5D",X"2A",X"05",X"86",X"FE",X"A7",X"A8",X"12",X"BD",X"15",X"BD",X"1D",X"ED",X"A8",X"14",X"35",
		X"F7",X"BD",X"00",X"5A",X"10",X"AE",X"2B",X"A6",X"A8",X"19",X"27",X"F5",X"CE",X"2B",X"12",X"EF",
		X"2E",X"CE",X"2B",X"C5",X"A6",X"24",X"E6",X"27",X"BD",X"17",X"7C",X"30",X"84",X"27",X"35",X"A0",
		X"04",X"46",X"40",X"E0",X"05",X"56",X"50",X"BD",X"16",X"C7",X"97",X"2F",X"1D",X"58",X"49",X"58",
		X"49",X"ED",X"A8",X"14",X"D6",X"2F",X"1D",X"58",X"49",X"58",X"49",X"ED",X"A8",X"12",X"86",X"0F",
		X"BD",X"00",X"5C",X"BD",X"15",X"BD",X"C1",X"08",X"25",X"0A",X"10",X"AE",X"2B",X"E6",X"A8",X"18",
		X"2B",X"EC",X"20",X"BD",X"8E",X"2B",X"1D",X"AF",X"2E",X"CC",X"77",X"8B",X"A0",X"24",X"E0",X"25",
		X"BD",X"16",X"C7",X"97",X"2F",X"1D",X"58",X"49",X"ED",X"A8",X"14",X"D6",X"2F",X"1D",X"58",X"49",
		X"ED",X"A8",X"12",X"86",X"03",X"BD",X"00",X"5C",X"10",X"AE",X"2B",X"EC",X"24",X"83",X"77",X"8B",
		X"26",X"D7",X"10",X"9E",X"08",X"10",X"AE",X"2B",X"BD",X"0C",X"3A",X"BD",X"1D",X"64",X"8D",X"03",
		X"7E",X"00",X"89",X"34",X"17",X"EC",X"24",X"C0",X"05",X"C1",X"3F",X"23",X"13",X"8B",X"15",X"46",
		X"8E",X"0C",X"01",X"1A",X"50",X"BF",X"CA",X"06",X"FD",X"CA",X"04",X"86",X"12",X"B7",X"CA",X"00",
		X"35",X"97",X"6C",X"A8",X"18",X"BD",X"17",X"C3",X"24",X"10",X"6F",X"A8",X"18",X"8E",X"4D",X"32",
		X"A6",X"A8",X"12",X"2A",X"22",X"8E",X"4C",X"68",X"20",X"1D",X"EC",X"A8",X"14",X"2A",X"04",X"43",
		X"50",X"82",X"FF",X"6D",X"A8",X"12",X"2B",X"44",X"A3",X"A8",X"12",X"2E",X"47",X"8E",X"2B",X"B5",
		X"E6",X"A8",X"18",X"C4",X"06",X"AE",X"85",X"AF",X"28",X"8D",X"A8",X"BD",X"24",X"C9",X"BD",X"18",
		X"4D",X"26",X"40",X"EC",X"24",X"C0",X"05",X"C1",X"3F",X"22",X"01",X"39",X"8B",X"15",X"46",X"1F",
		X"01",X"EC",X"A8",X"1D",X"4D",X"26",X"01",X"4A",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",
		X"D7",X"2F",X"C6",X"EE",X"BD",X"7B",X"0F",X"96",X"2F",X"7E",X"7B",X"0F",X"8E",X"2B",X"BD",X"E3",
		X"A8",X"12",X"2B",X"BC",X"8E",X"52",X"B0",X"E6",X"A8",X"18",X"C4",X"04",X"27",X"B9",X"8E",X"53",
		X"6E",X"20",X"B4",X"E7",X"A8",X"19",X"56",X"56",X"2A",X"0B",X"86",X"01",X"24",X"01",X"40",X"A7",
		X"A8",X"12",X"6F",X"A8",X"13",X"56",X"56",X"2A",X"0B",X"86",X"01",X"24",X"01",X"40",X"A7",X"A8",
		X"14",X"6F",X"A8",X"15",X"39",X"50",X"56",X"51",X"14",X"51",X"CE",X"51",X"14",X"4D",X"FC",X"4E",
		X"BA",X"4F",X"74",X"4E",X"BA",X"08",X"07",X"09",X"00",X"35",X"40",X"A6",X"C0",X"AB",X"A8",X"1E",
		X"19",X"A7",X"A8",X"1E",X"24",X"03",X"6C",X"A8",X"1D",X"6E",X"C4",X"A6",X"07",X"A1",X"27",X"24",
		X"01",X"39",X"BD",X"2B",X"C9",X"20",X"0A",X"6E",X"6C",X"A8",X"1A",X"20",X"0F",X"A6",X"07",X"A1",
		X"27",X"25",X"EE",X"BD",X"2B",X"C9",X"15",X"0A",X"6F",X"6C",X"A8",X"1B",X"7E",X"1D",X"0D",X"A6",
		X"07",X"A1",X"27",X"25",X"DC",X"BD",X"2B",X"C9",X"15",X"6C",X"A8",X"1C",X"0A",X"71",X"20",X"EC",
		X"C6",X"09",X"BD",X"36",X"A3",X"BD",X"2D",X"2B",X"20",X"03",X"BD",X"1D",X"7A",X"6A",X"88",X"1B",
		X"2A",X"F8",X"20",X"03",X"BD",X"1D",X"48",X"6A",X"88",X"1A",X"2A",X"F8",X"20",X"03",X"BD",X"1D",
		X"12",X"6A",X"88",X"1C",X"2A",X"F8",X"31",X"84",X"6F",X"2D",X"AE",X"A8",X"1F",X"BD",X"01",X"04",
		X"86",X"20",X"A7",X"2B",X"EE",X"28",X"EC",X"58",X"E3",X"24",X"91",X"36",X"25",X"40",X"D1",X"37",
		X"25",X"3C",X"90",X"36",X"97",X"2F",X"D1",X"39",X"23",X"02",X"D6",X"39",X"D7",X"2E",X"EC",X"56",
		X"E3",X"24",X"D1",X"39",X"22",X"28",X"91",X"38",X"22",X"24",X"90",X"36",X"DD",X"2C",X"96",X"2E",
		X"9E",X"19",X"D0",X"37",X"25",X"06",X"58",X"3A",X"90",X"2D",X"20",X"02",X"90",X"37",X"97",X"2E",
		X"EC",X"81",X"D1",X"2C",X"2D",X"04",X"91",X"2F",X"2F",X"05",X"0A",X"2E",X"2A",X"F2",X"39",X"1A",
		X"50",X"96",X"00",X"8A",X"08",X"97",X"00",X"97",X"73",X"0F",X"5F",X"7E",X"1F",X"91",X"72",X"89",
		X"8A",X"9B",X"0D",X"A5",X"00",X"00",X"04",X"FF",X"2E",X"98",X"2E",X"61",X"A6",X"A8",X"1A",X"AA",
		X"88",X"1A",X"26",X"49",X"A6",X"A8",X"12",X"A8",X"88",X"12",X"2B",X"36",X"A6",X"A8",X"14",X"A8",
		X"88",X"14",X"2B",X"2E",X"EC",X"24",X"6D",X"A8",X"12",X"2A",X"04",X"86",X"FE",X"A0",X"24",X"97",
		X"2F",X"C0",X"3F",X"A6",X"A8",X"14",X"2A",X"04",X"C6",X"EA",X"E0",X"25",X"86",X"1E",X"A7",X"A8",
		X"1A",X"A7",X"88",X"1A",X"D1",X"2F",X"22",X"0B",X"EC",X"A8",X"12",X"43",X"50",X"82",X"FF",X"ED",
		X"A8",X"12",X"39",X"EC",X"A8",X"14",X"43",X"50",X"82",X"FF",X"ED",X"A8",X"14",X"39",X"C6",X"FF",
		X"BD",X"36",X"A3",X"BD",X"22",X"F4",X"0F",X"73",X"BD",X"00",X"A5",X"2F",X"D2",X"39",X"18",X"2F",
		X"5A",X"AF",X"2B",X"31",X"84",X"BD",X"00",X"47",X"BD",X"07",X"1B",X"09",X"8D",X"0B",X"EE",X"A8",
		X"1B",X"31",X"C4",X"BD",X"00",X"47",X"7E",X"01",X"B5",X"8D",X"00",X"BD",X"1B",X"AD",X"05",X"80",
		X"39",X"34",X"77",X"BD",X"07",X"1B",X"07",X"86",X"5A",X"34",X"02",X"4F",X"BD",X"00",X"5C",X"86",
		X"07",X"97",X"8A",X"35",X"02",X"4A",X"26",X"F1",X"BD",X"01",X"C3",X"1F",X"04",X"0A",X"2C",X"9E",
		X"10",X"9F",X"9F",X"BD",X"D0",X"00",X"9E",X"76",X"AF",X"C4",X"2A",X"02",X"EF",X"02",X"DF",X"76",
		X"8E",X"98",X"76",X"AF",X"42",X"10",X"AF",X"44",X"EF",X"A8",X"1B",X"4F",X"A7",X"A8",X"1A",X"BD",
		X"08",X"15",X"BD",X"08",X"62",X"BD",X"15",X"B9",X"BD",X"2D",X"EF",X"86",X"0F",X"BD",X"00",X"5C",
		X"0F",X"9F",X"0F",X"8A",X"35",X"F7",X"9E",X"76",X"2A",X"0C",X"33",X"84",X"AE",X"84",X"BD",X"01",
		X"B5",X"8C",X"00",X"00",X"2B",X"F4",X"0F",X"76",X"39",X"A6",X"04",X"90",X"36",X"46",X"2A",X"01",
		X"40",X"1F",X"89",X"3D",X"ED",X"E3",X"E6",X"05",X"D0",X"37",X"56",X"2A",X"01",X"50",X"1F",X"98",
		X"3D",X"E3",X"E1",X"39",X"BD",X"00",X"5A",X"DE",X"76",X"2A",X"F9",X"CC",X"FF",X"FF",X"DD",X"2F",
		X"AE",X"44",X"8D",X"D5",X"10",X"93",X"2F",X"24",X"04",X"DD",X"2F",X"9F",X"34",X"EE",X"C4",X"2B",
		X"EF",X"10",X"9E",X"34",X"A6",X"A8",X"1A",X"27",X"05",X"BD",X"00",X"5C",X"20",X"D6",X"DC",X"36",
		X"A0",X"24",X"46",X"E0",X"25",X"56",X"8D",X"07",X"86",X"05",X"BD",X"00",X"5C",X"20",X"C5",X"BD",
		X"15",X"DA",X"C1",X"40",X"22",X"0E",X"C1",X"26",X"23",X"02",X"C6",X"26",X"C1",X"1A",X"24",X"02",
		X"C6",X"1A",X"20",X"2F",X"5D",X"2B",X"0E",X"C1",X"66",X"23",X"02",X"C6",X"66",X"C1",X"5A",X"24",
		X"02",X"C6",X"5A",X"20",X"1E",X"C1",X"C0",X"22",X"0E",X"C1",X"A6",X"23",X"02",X"C6",X"A6",X"C1",
		X"9A",X"24",X"02",X"C6",X"9A",X"20",X"0C",X"C1",X"E6",X"23",X"02",X"C6",X"E6",X"C1",X"DA",X"24",
		X"02",X"C6",X"DA",X"D7",X"2F",X"BD",X"15",X"BD",X"DE",X"79",X"A6",X"4F",X"3D",X"AB",X"4F",X"1F",
		X"89",X"96",X"2F",X"BD",X"16",X"23",X"5F",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",
		X"A8",X"12",X"5F",X"96",X"32",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",X"A8",X"14",
		X"39",X"A6",X"24",X"E6",X"A8",X"12",X"2A",X"06",X"81",X"14",X"22",X"10",X"20",X"04",X"81",X"D1",
		X"25",X"0A",X"EC",X"A8",X"12",X"43",X"50",X"82",X"FF",X"ED",X"A8",X"12",X"A6",X"25",X"E6",X"A8",
		X"14",X"2A",X"06",X"81",X"53",X"22",X"10",X"20",X"04",X"81",X"BD",X"25",X"0A",X"EC",X"A8",X"14",
		X"43",X"50",X"82",X"FF",X"ED",X"A8",X"14",X"39",X"A6",X"A8",X"1A",X"27",X"03",X"6A",X"A8",X"1A",
		X"CE",X"2E",X"DC",X"8E",X"2E",X"FC",X"A6",X"A8",X"12",X"2A",X"06",X"8E",X"99",X"A0",X"33",X"C8",
		X"10",X"A6",X"A8",X"14",X"2A",X"04",X"30",X"08",X"33",X"48",X"EC",X"A8",X"18",X"8B",X"64",X"24",
		X"15",X"6C",X"A8",X"19",X"C4",X"03",X"58",X"AE",X"85",X"AF",X"28",X"33",X"C5",X"EC",X"24",X"AB",
		X"C4",X"EB",X"41",X"ED",X"24",X"4F",X"A7",X"A8",X"18",X"7E",X"24",X"C9",X"00",X"FE",X"00",X"01",
		X"01",X"03",X"FF",X"FE",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"00",X"FF",X"FE",X"01",X"01",
		X"00",X"03",X"00",X"FE",X"00",X"00",X"00",X"00",X"01",X"00",X"FF",X"00",X"58",X"80",X"59",X"94",
		X"5A",X"99",X"5B",X"63",X"5C",X"59",X"5D",X"6D",X"5E",X"81",X"5F",X"95",X"60",X"A5",X"61",X"37",
		X"8E",X"9C",X"22",X"31",X"02",X"10",X"BF",X"99",X"B2",X"CE",X"08",X"08",X"EF",X"3E",X"96",X"15",
		X"A8",X"3C",X"A7",X"3C",X"8E",X"61",X"37",X"CC",X"16",X"0B",X"BD",X"18",X"D2",X"EF",X"A1",X"CC",
		X"16",X"0B",X"8E",X"60",X"A5",X"10",X"BF",X"99",X"B0",X"BD",X"18",X"D2",X"31",X"26",X"C6",X"0E",
		X"34",X"24",X"BD",X"00",X"5A",X"35",X"24",X"8E",X"99",X"A0",X"10",X"AF",X"85",X"8E",X"2E",X"FC",
		X"AE",X"85",X"BD",X"18",X"A4",X"C0",X"02",X"2A",X"E7",X"39",X"86",X"1E",X"A7",X"2D",X"10",X"AE",
		X"2B",X"EC",X"24",X"C1",X"44",X"24",X"02",X"C6",X"44",X"C1",X"DF",X"23",X"02",X"C6",X"DF",X"81",
		X"E8",X"23",X"02",X"86",X"E8",X"ED",X"24",X"86",X"01",X"BD",X"00",X"5C",X"6A",X"2D",X"2B",X"24",
		X"E6",X"2D",X"10",X"AE",X"2B",X"BD",X"08",X"68",X"8E",X"2F",X"0C",X"A6",X"A8",X"12",X"2A",X"03",
		X"8E",X"99",X"B0",X"C4",X"01",X"58",X"AE",X"85",X"AF",X"28",X"BD",X"08",X"62",X"C6",X"99",X"BD",
		X"2F",X"E1",X"20",X"D3",X"86",X"78",X"A7",X"2D",X"96",X"00",X"2A",X"03",X"BD",X"D0",X"5F",X"4F",
		X"BD",X"00",X"5C",X"EE",X"2B",X"BD",X"15",X"BD",X"86",X"08",X"3D",X"8B",X"05",X"AB",X"45",X"97",
		X"2F",X"BD",X"15",X"BD",X"86",X"17",X"3D",X"AB",X"44",X"D6",X"2F",X"BD",X"D0",X"36",X"6A",X"2D",
		X"26",X"DD",X"10",X"AE",X"2B",X"5F",X"8D",X"09",X"BD",X"08",X"68",X"BD",X"01",X"A9",X"7E",X"00",
		X"89",X"D7",X"30",X"EC",X"24",X"C0",X"05",X"8B",X"1D",X"46",X"1F",X"01",X"86",X"10",X"D6",X"30",
		X"BD",X"7B",X"0F",X"4F",X"7E",X"7B",X"0F",X"A6",X"2A",X"8B",X"02",X"A7",X"2A",X"CC",X"0D",X"A5",
		X"ED",X"68",X"A6",X"29",X"88",X"E0",X"A7",X"29",X"39",X"4B",X"24",X"00",X"00",X"06",X"02",X"2F",
		X"F7",X"01",X"C1",X"34",X"77",X"6A",X"61",X"2A",X"02",X"35",X"F7",X"BD",X"01",X"C3",X"14",X"08",
		X"0E",X"30",X"09",X"BD",X"17",X"F5",X"8E",X"23",X"60",X"CC",X"DB",X"C9",X"BD",X"17",X"D9",X"24",
		X"F2",X"BD",X"23",X"DE",X"25",X"ED",X"20",X"DD",X"74",X"8C",X"87",X"97",X"3B",X"E8",X"00",X"10",
		X"0A",X"FF",X"01",X"C1",X"01",X"C1",X"BD",X"00",X"A5",X"30",X"E3",X"25",X"07",X"30",X"60",X"6F",
		X"2B",X"BD",X"01",X"C3",X"14",X"04",X"0A",X"30",X"38",X"10",X"9F",X"8B",X"BD",X"08",X"1D",X"39",
		X"7F",X"9A",X"00",X"6F",X"2B",X"86",X"03",X"BD",X"00",X"5C",X"96",X"00",X"85",X"04",X"26",X"F5",
		X"96",X"95",X"26",X"F1",X"6A",X"2B",X"2A",X"0F",X"86",X"03",X"A7",X"2B",X"96",X"89",X"63",X"2C",
		X"2A",X"02",X"96",X"8A",X"B7",X"9A",X"00",X"8D",X"41",X"CE",X"98",X"76",X"EE",X"C4",X"2A",X"07",
		X"10",X"AE",X"44",X"8D",X"2C",X"20",X"F5",X"10",X"9E",X"8B",X"10",X"AE",X"22",X"A6",X"25",X"81",
		X"79",X"23",X"04",X"8D",X"12",X"20",X"F3",X"10",X"9E",X"8B",X"10",X"AE",X"A4",X"A6",X"25",X"81",
		X"9E",X"24",X"B2",X"8D",X"02",X"20",X"F3",X"E6",X"2C",X"C1",X"02",X"27",X"04",X"C1",X"03",X"26",
		X"08",X"BD",X"17",X"C3",X"24",X"03",X"7E",X"08",X"62",X"39",X"8E",X"3B",X"E8",X"EE",X"1E",X"CC",
		X"41",X"86",X"1A",X"50",X"BF",X"CA",X"02",X"FF",X"CA",X"06",X"FD",X"CA",X"04",X"86",X"0A",X"B7",
		X"CA",X"00",X"39",X"7F",X"9A",X"00",X"10",X"9E",X"8B",X"BD",X"00",X"47",X"7E",X"01",X"A9",X"77",
		X"3F",X"77",X"3F",X"4B",X"06",X"00",X"00",X"0B",X"FF",X"31",X"01",X"01",X"C1",X"00",X"00",X"02",
		X"00",X"A6",X"25",X"81",X"90",X"10",X"25",X"F3",X"C0",X"32",X"62",X"7E",X"38",X"1D",X"BD",X"15",
		X"BD",X"86",X"64",X"3D",X"8B",X"10",X"BD",X"00",X"5C",X"96",X"00",X"85",X"20",X"27",X"EF",X"8D",
		X"02",X"20",X"EB",X"BD",X"01",X"C3",X"1A",X"04",X"16",X"30",X"EF",X"BD",X"07",X"1B",X"15",X"BD",
		X"15",X"BD",X"86",X"0A",X"3D",X"AB",X"24",X"A7",X"24",X"4F",X"7E",X"08",X"15",X"BD",X"07",X"1B",
		X"13",X"96",X"00",X"8A",X"04",X"97",X"00",X"BD",X"14",X"62",X"BD",X"14",X"9B",X"CC",X"00",X"03",
		X"DD",X"56",X"CC",X"01",X"00",X"DD",X"59",X"96",X"67",X"40",X"47",X"8B",X"7E",X"C6",X"54",X"D0",
		X"67",X"DD",X"36",X"CC",X"98",X"A8",X"8E",X"F8",X"E0",X"0D",X"8D",X"26",X"06",X"CC",X"7F",X"FF",
		X"8E",X"AD",X"07",X"8D",X"2F",X"BD",X"00",X"A5",X"31",X"AB",X"57",X"14",X"E2",X"00",X"6F",X"A8",
		X"2A",X"BD",X"00",X"5A",X"96",X"00",X"84",X"04",X"26",X"F7",X"96",X"8D",X"2A",X"0A",X"86",X"1E",
		X"BD",X"00",X"5C",X"86",X"2A",X"BD",X"7B",X"1A",X"CE",X"39",X"7D",X"BD",X"08",X"38",X"CC",X"C5",
		X"53",X"8E",X"A6",X"00",X"FD",X"99",X"FC",X"BF",X"99",X"FF",X"39",X"AE",X"A8",X"2A",X"2A",X"00",
		X"96",X"00",X"84",X"FB",X"97",X"00",X"20",X"E0",X"86",X"05",X"BD",X"01",X"48",X"A6",X"2B",X"97",
		X"8F",X"7E",X"00",X"89",X"86",X"01",X"CE",X"32",X"3D",X"20",X"05",X"CE",X"32",X"72",X"86",X"02",
		X"95",X"8F",X"26",X"11",X"C6",X"03",X"D7",X"8F",X"BD",X"00",X"AD",X"2F",X"13",X"31",X"B8",X"A7",
		X"2B",X"8D",X"03",X"EF",X"2B",X"39",X"34",X"40",X"CE",X"32",X"09",X"BD",X"00",X"E2",X"7F",X"9A",
		X"00",X"BD",X"00",X"AD",X"39",X"0B",X"31",X"FF",X"CE",X"32",X"3B",X"EF",X"2B",X"35",X"C0",X"BD",
		X"00",X"5A",X"96",X"90",X"26",X"F9",X"6E",X"B8",X"0B",X"1B",X"14",X"0B",X"00",X"BD",X"31",X"3D",
		X"CE",X"33",X"CB",X"BD",X"08",X"38",X"BD",X"30",X"CA",X"86",X"03",X"BD",X"01",X"48",X"BD",X"D2",
		X"4E",X"86",X"2C",X"BD",X"7B",X"15",X"86",X"03",X"BD",X"01",X"48",X"86",X"2C",X"BD",X"7B",X"1D",
		X"86",X"26",X"BD",X"7B",X"15",X"86",X"03",X"BD",X"01",X"48",X"39",X"8D",X"D0",X"8E",X"CC",X"04",
		X"BD",X"D2",X"21",X"46",X"24",X"2C",X"BD",X"38",X"2A",X"BD",X"D2",X"33",X"86",X"26",X"BD",X"7B",
		X"1D",X"86",X"28",X"BD",X"7B",X"15",X"8E",X"54",X"DC",X"96",X"1D",X"C6",X"AA",X"BD",X"7B",X"0F",
		X"86",X"0A",X"BD",X"01",X"48",X"0F",X"8F",X"86",X"2F",X"BD",X"7B",X"12",X"86",X"01",X"97",X"8D",
		X"8D",X"9B",X"BD",X"38",X"2A",X"86",X"11",X"BD",X"7B",X"12",X"CE",X"33",X"99",X"BD",X"08",X"38",
		X"CC",X"1D",X"05",X"BD",X"33",X"53",X"86",X"16",X"BD",X"7B",X"15",X"CE",X"33",X"71",X"BD",X"08",
		X"38",X"86",X"18",X"BD",X"7B",X"15",X"CE",X"33",X"B7",X"BD",X"08",X"38",X"86",X"17",X"BD",X"7B",
		X"15",X"CE",X"33",X"7B",X"BD",X"08",X"38",X"86",X"1C",X"BD",X"7B",X"15",X"CE",X"33",X"A3",X"BD",
		X"08",X"38",X"86",X"30",X"BD",X"7B",X"15",X"86",X"31",X"BD",X"7B",X"15",X"CC",X"14",X"05",X"BD",
		X"33",X"53",X"86",X"1A",X"BD",X"7B",X"15",X"CE",X"33",X"8F",X"BD",X"08",X"38",X"86",X"19",X"BD",
		X"7B",X"15",X"CE",X"33",X"85",X"BD",X"08",X"38",X"CC",X"15",X"05",X"BD",X"33",X"53",X"CC",X"1E",
		X"05",X"BD",X"33",X"53",X"86",X"1F",X"BD",X"7B",X"15",X"CE",X"33",X"C1",X"BD",X"08",X"38",X"CE",
		X"33",X"AD",X"BD",X"08",X"38",X"CC",X"20",X"05",X"BD",X"33",X"53",X"86",X"7E",X"BD",X"00",X"5C",
		X"86",X"1C",X"BD",X"7B",X"1D",X"86",X"2E",X"BD",X"7B",X"15",X"CE",X"33",X"A3",X"BD",X"08",X"38",
		X"86",X"30",X"BD",X"7B",X"1D",X"86",X"31",X"BD",X"7B",X"1D",X"86",X"21",X"BD",X"7B",X"15",X"CC",
		X"22",X"0F",X"BD",X"7B",X"15",X"C6",X"14",X"BD",X"34",X"C5",X"86",X"02",X"BD",X"01",X"48",X"86",
		X"7F",X"C6",X"00",X"8E",X"32",X"DC",X"BD",X"7B",X"0C",X"86",X"26",X"BD",X"7B",X"15",X"86",X"04",
		X"BD",X"01",X"48",X"0F",X"8F",X"0F",X"15",X"BD",X"00",X"A5",X"36",X"87",X"4D",X"1B",X"34",X"F8",
		X"7E",X"00",X"89",X"34",X"06",X"BD",X"7B",X"15",X"86",X"14",X"BD",X"00",X"5C",X"35",X"06",X"5A",
		X"27",X"0E",X"34",X"06",X"BD",X"7B",X"1D",X"86",X"0E",X"BD",X"00",X"5C",X"35",X"06",X"20",X"E3",
		X"39",X"04",X"06",X"0A",X"00",X"4A",X"9D",X"2C",X"66",X"00",X"00",X"05",X"09",X"0A",X"00",X"4A",
		X"C1",X"30",X"8C",X"00",X"00",X"09",X"08",X"0A",X"00",X"49",X"DF",X"5F",X"7D",X"00",X"00",X"09",
		X"0D",X"0A",X"00",X"49",X"4A",X"61",X"68",X"00",X"00",X"09",X"10",X"0A",X"00",X"70",X"2E",X"45",
		X"6D",X"00",X"00",X"0A",X"0F",X"0A",X"00",X"4D",X"FC",X"2D",X"A8",X"00",X"00",X"0D",X"12",X"0A",
		X"00",X"58",X"80",X"6A",X"A2",X"00",X"00",X"06",X"07",X"0A",X"00",X"54",X"9A",X"2A",X"7B",X"00",
		X"00",X"09",X"0E",X"0A",X"00",X"4B",X"24",X"58",X"8F",X"00",X"00",X"0C",X"16",X"0A",X"00",X"74",
		X"98",X"44",X"65",X"00",X"00",X"81",X"01",X"26",X"0D",X"86",X"1D",X"BD",X"7B",X"15",X"BD",X"34",
		X"0E",X"86",X"1D",X"7E",X"7B",X"1D",X"81",X"05",X"10",X"24",X"00",X"6E",X"8B",X"60",X"8D",X"27",
		X"C5",X"80",X"27",X"04",X"30",X"89",X"E8",X"00",X"34",X"12",X"8D",X"55",X"86",X"60",X"30",X"09",
		X"C5",X"80",X"27",X"04",X"30",X"89",X"E8",X"00",X"8D",X"31",X"35",X"12",X"20",X"3B",X"34",X"16",
		X"86",X"02",X"BD",X"01",X"48",X"35",X"96",X"34",X"02",X"EC",X"04",X"C1",X"80",X"24",X"08",X"CB",
		X"10",X"8D",X"0C",X"C4",X"F0",X"35",X"82",X"C0",X"24",X"8D",X"04",X"CA",X"0F",X"35",X"82",X"8B",
		X"15",X"46",X"1F",X"01",X"5F",X"81",X"46",X"25",X"01",X"5A",X"39",X"8D",X"14",X"30",X"07",X"4C",
		X"8D",X"0F",X"8D",X"CA",X"8D",X"03",X"4A",X"30",X"19",X"34",X"12",X"5F",X"BD",X"7B",X"0C",X"35",
		X"92",X"34",X"16",X"C6",X"11",X"BD",X"7B",X"0C",X"35",X"96",X"26",X"0F",X"BD",X"34",X"17",X"C5",
		X"80",X"27",X"04",X"30",X"89",X"E0",X"00",X"86",X"74",X"20",X"D0",X"81",X"08",X"24",X"15",X"8B",
		X"5F",X"8D",X"A4",X"C5",X"80",X"27",X"04",X"30",X"89",X"EE",X"00",X"34",X"12",X"8D",X"D2",X"86",
		X"77",X"16",X"FF",X"7A",X"26",X"0E",X"8D",X"8F",X"C5",X"80",X"27",X"04",X"30",X"89",X"E0",X"00",
		X"86",X"6F",X"20",X"A7",X"81",X"0A",X"24",X"0F",X"BD",X"34",X"17",X"C5",X"80",X"27",X"04",X"30",
		X"89",X"E0",X"00",X"86",X"67",X"20",X"94",X"26",X"0C",X"86",X"7E",X"8E",X"36",X"AB",X"8D",X"A1",
		X"BD",X"34",X"0E",X"20",X"94",X"81",X"0C",X"24",X"28",X"86",X"22",X"BD",X"7B",X"15",X"86",X"21",
		X"BD",X"7B",X"15",X"C6",X"04",X"34",X"04",X"86",X"21",X"B7",X"9A",X"00",X"86",X"0A",X"BD",X"00",
		X"5C",X"86",X"00",X"B7",X"9A",X"00",X"86",X"05",X"BD",X"00",X"5C",X"35",X"04",X"5A",X"26",X"E5",
		X"39",X"86",X"30",X"BD",X"7B",X"15",X"86",X"31",X"BD",X"7B",X"15",X"BD",X"34",X"0E",X"86",X"30",
		X"BD",X"7B",X"1D",X"86",X"31",X"7E",X"7B",X"1D",X"CE",X"14",X"5A",X"BD",X"00",X"E2",X"C6",X"01",
		X"D7",X"90",X"BD",X"30",X"46",X"8E",X"9A",X"AB",X"9F",X"64",X"4F",X"5F",X"ED",X"84",X"ED",X"02",
		X"A7",X"04",X"8E",X"1A",X"0D",X"9F",X"62",X"BD",X"00",X"A5",X"3A",X"CB",X"39",X"10",X"39",X"A1",
		X"BD",X"00",X"AD",X"2F",X"19",X"31",X"0E",X"0F",X"93",X"0F",X"94",X"BD",X"38",X"2A",X"4F",X"5F",
		X"DD",X"4C",X"CE",X"14",X"47",X"BD",X"00",X"E2",X"BD",X"14",X"9B",X"86",X"0C",X"D6",X"90",X"C1",
		X"0A",X"25",X"02",X"86",X"15",X"97",X"67",X"86",X"04",X"C1",X"05",X"26",X"01",X"4F",X"97",X"69",
		X"C1",X"0B",X"26",X"25",X"0F",X"9C",X"BD",X"11",X"BC",X"BD",X"23",X"FF",X"CC",X"74",X"74",X"ED",
		X"24",X"CC",X"88",X"7E",X"ED",X"26",X"97",X"9E",X"CC",X"0A",X"8E",X"ED",X"2E",X"4F",X"BD",X"08",
		X"15",X"BD",X"08",X"62",X"BD",X"12",X"AA",X"20",X"03",X"BD",X"11",X"FE",X"D6",X"90",X"5A",X"27",
		X"14",X"C1",X"0A",X"23",X"20",X"C1",X"0B",X"27",X"46",X"C1",X"0C",X"27",X"08",X"0F",X"8D",X"BD",
		X"31",X"E6",X"7E",X"36",X"87",X"CC",X"78",X"8C",X"7E",X"36",X"2B",X"08",X"09",X"07",X"F6",X"06",
		X"02",X"03",X"05",X"04",X"02",X"8E",X"35",X"9A",X"A6",X"85",X"5F",X"DD",X"91",X"2A",X"20",X"BD",
		X"18",X"46",X"26",X"1B",X"C6",X"05",X"BD",X"36",X"A3",X"86",X"FF",X"97",X"8D",X"BD",X"31",X"3D",
		X"BD",X"14",X"E8",X"7E",X"36",X"6A",X"BD",X"18",X"28",X"BD",X"23",X"0B",X"7E",X"35",X"2E",X"CE",
		X"36",X"64",X"10",X"8E",X"36",X"5F",X"96",X"00",X"85",X"08",X"26",X"04",X"33",X"41",X"31",X"3F",
		X"DC",X"36",X"BD",X"17",X"7C",X"A6",X"0C",X"91",X"91",X"27",X"3E",X"96",X"36",X"DE",X"2E",X"11",
		X"83",X"01",X"00",X"24",X"07",X"A0",X"04",X"46",X"E0",X"05",X"20",X"34",X"0D",X"91",X"2B",X"24",
		X"CE",X"98",X"91",X"DC",X"36",X"BD",X"17",X"7C",X"30",X"84",X"26",X"1D",X"86",X"18",X"BD",X"01",
		X"13",X"27",X"11",X"96",X"9E",X"27",X"AF",X"4F",X"5F",X"DD",X"4C",X"DD",X"3E",X"DD",X"40",X"BD",
		X"00",X"5A",X"20",X"EF",X"33",X"A4",X"BD",X"17",X"7C",X"EC",X"04",X"90",X"36",X"46",X"D0",X"37",
		X"56",X"BD",X"15",X"DA",X"54",X"54",X"54",X"54",X"54",X"C9",X"00",X"58",X"8E",X"36",X"4E",X"AE",
		X"85",X"9F",X"4C",X"4F",X"BD",X"00",X"5C",X"96",X"95",X"26",X"F8",X"7E",X"35",X"7C",X"14",X"00",
		X"14",X"14",X"00",X"14",X"EC",X"14",X"EC",X"00",X"EC",X"EC",X"00",X"EC",X"14",X"EC",X"04",X"08",
		X"05",X"07",X"09",X"00",X"04",X"02",X"03",X"0A",X"06",X"00",X"BD",X"14",X"62",X"BD",X"14",X"85",
		X"7E",X"35",X"2E",X"86",X"1B",X"BD",X"01",X"13",X"27",X"01",X"3F",X"EF",X"98",X"07",X"BD",X"18",
		X"28",X"BD",X"23",X"0B",X"7E",X"00",X"89",X"8E",X"9A",X"73",X"9F",X"64",X"8E",X"19",X"91",X"9F",
		X"62",X"BD",X"14",X"62",X"CE",X"14",X"52",X"BD",X"00",X"E2",X"BD",X"14",X"9B",X"0F",X"90",X"0F",
		X"95",X"20",X"DB",X"34",X"76",X"5D",X"2A",X"12",X"CE",X"98",X"93",X"5C",X"26",X"02",X"33",X"41",
		X"A6",X"C4",X"34",X"01",X"26",X"3B",X"63",X"C4",X"20",X"1B",X"D1",X"90",X"34",X"01",X"26",X"31",
		X"0C",X"90",X"C1",X"0B",X"26",X"0F",X"BD",X"00",X"AD",X"2F",X"1C",X"37",X"04",X"C6",X"07",X"81",
		X"02",X"27",X"02",X"C6",X"08",X"86",X"FF",X"97",X"95",X"34",X"04",X"BD",X"18",X"28",X"E6",X"E4",
		X"CE",X"36",X"F6",X"A6",X"C5",X"BD",X"33",X"D5",X"35",X"04",X"C1",X"0D",X"27",X"05",X"BD",X"18",
		X"34",X"0F",X"95",X"35",X"F7",X"0A",X"08",X"01",X"02",X"03",X"04",X"0C",X"05",X"06",X"07",X"09",
		X"08",X"01",X"01",X"0B",X"86",X"05",X"BD",X"01",X"48",X"D6",X"90",X"27",X"02",X"0C",X"90",X"7E",
		X"00",X"89",X"34",X"77",X"86",X"23",X"BD",X"7B",X"12",X"86",X"64",X"BD",X"00",X"5C",X"86",X"23",
		X"BD",X"7B",X"1A",X"35",X"F7",X"34",X"77",X"B6",X"BF",X"23",X"27",X"24",X"8E",X"CC",X"06",X"BD",
		X"D2",X"21",X"81",X"09",X"27",X"1A",X"86",X"27",X"BD",X"7B",X"15",X"34",X"10",X"CC",X"31",X"AA",
		X"BD",X"7B",X"09",X"BD",X"7B",X"09",X"35",X"10",X"C6",X"DD",X"B6",X"BF",X"23",X"BD",X"7B",X"0F",
		X"35",X"F7",X"09",X"0D",X"12",X"AA",X"00",X"00",X"07",X"20",X"09",X"0D",X"12",X"AA",X"00",X"00",
		X"85",X"20",X"00",X"00",X"34",X"57",X"CE",X"37",X"52",X"BD",X"08",X"38",X"CC",X"76",X"DD",X"8E",
		X"07",X"20",X"BD",X"7B",X"0C",X"96",X"00",X"2A",X"21",X"84",X"40",X"27",X"1D",X"86",X"76",X"8E",
		X"85",X"20",X"BD",X"7B",X"0C",X"D6",X"69",X"96",X"01",X"26",X"03",X"F6",X"9A",X"8E",X"8D",X"13",
		X"88",X"28",X"DD",X"F6",X"9A",X"80",X"96",X"01",X"26",X"02",X"D6",X"69",X"8D",X"05",X"0C",X"28",
		X"DD",X"35",X"D7",X"EE",X"E1",X"37",X"10",X"4F",X"C1",X"64",X"25",X"0A",X"C0",X"64",X"4C",X"C1",
		X"64",X"25",X"03",X"C0",X"64",X"4C",X"D7",X"2F",X"E6",X"C0",X"4D",X"27",X"05",X"8A",X"F0",X"BD",
		X"7B",X"0F",X"96",X"2F",X"8D",X"02",X"6E",X"C4",X"BD",X"D2",X"48",X"7E",X"7B",X"0F",X"56",X"14",
		X"00",X"00",X"00",X"00",X"37",X"D8",X"38",X"1D",X"6A",X"A8",X"18",X"10",X"27",X"F9",X"2A",X"7E",
		X"24",X"C9",X"34",X"30",X"C6",X"FE",X"BD",X"36",X"A3",X"BD",X"01",X"C3",X"1B",X"08",X"0E",X"37",
		X"CE",X"86",X"3C",X"A7",X"A8",X"18",X"AE",X"62",X"EC",X"04",X"ED",X"24",X"ED",X"26",X"BD",X"15",
		X"B9",X"BD",X"16",X"C7",X"97",X"2F",X"1D",X"58",X"49",X"58",X"49",X"ED",X"A8",X"12",X"D6",X"2F",
		X"1D",X"58",X"49",X"58",X"49",X"ED",X"A8",X"14",X"BD",X"08",X"15",X"35",X"B0",X"BD",X"00",X"47",
		X"8E",X"D0",X"97",X"1E",X"12",X"32",X"62",X"7E",X"01",X"AB",X"34",X"40",X"86",X"C9",X"8E",X"99",
		X"F1",X"A7",X"89",X"26",X"0F",X"A7",X"80",X"8C",X"9A",X"01",X"25",X"F5",X"BD",X"D2",X"1E",X"CE",
		X"38",X"9D",X"BD",X"08",X"38",X"10",X"8E",X"38",X"78",X"8D",X"1C",X"8E",X"99",X"F1",X"CE",X"0D",
		X"7F",X"37",X"06",X"ED",X"81",X"8C",X"9A",X"01",X"25",X"F7",X"BD",X"37",X"25",X"96",X"90",X"26",
		X"03",X"BD",X"1A",X"C5",X"35",X"40",X"39",X"A6",X"A4",X"81",X"FF",X"27",X"F9",X"EE",X"A1",X"AE",
		X"A1",X"EC",X"A1",X"BD",X"D0",X"A1",X"20",X"EF",X"07",X"2F",X"8C",X"2F",X"0A",X"19",X"07",X"DF",
		X"8C",X"DF",X"09",X"0E",X"10",X"13",X"29",X"13",X"04",X"08",X"10",X"29",X"29",X"29",X"04",X"08",
		X"10",X"13",X"81",X"13",X"04",X"08",X"10",X"29",X"81",X"29",X"04",X"08",X"FF",X"97",X"3F",X"12",
		X"AA",X"00",X"00",X"00",X"00",X"10",X"C0",X"12",X"AA",X"00",X"00",X"00",X"3F",X"0B",X"C0",X"12",
		X"AA",X"00",X"00",X"8C",X"3F",X"7C",X"12",X"12",X"AA",X"00",X"00",X"10",X"ED",X"80",X"AE",X"12",
		X"00",X"00",X"00",X"0A",X"3F",X"19",X"17",X"12",X"00",X"00",X"00",X"11",X"16",X"19",X"17",X"12",
		X"00",X"00",X"00",X"69",X"16",X"7C",X"0F",X"12",X"88",X"00",X"00",X"10",X"30",X"02",X"97",X"12",
		X"88",X"00",X"00",X"08",X"48",X"02",X"97",X"12",X"88",X"00",X"00",X"8A",X"48",X"01",X"97",X"12",
		X"88",X"00",X"00",X"07",X"48",X"01",X"97",X"12",X"88",X"00",X"00",X"8C",X"48",X"76",X"02",X"12",
		X"88",X"00",X"00",X"0F",X"EB",X"0A",X"19",X"02",X"00",X"3A",X"D0",X"07",X"30",X"09",X"0E",X"02",
		X"00",X"3D",X"AA",X"07",X"DF",X"12",X"18",X"0A",X"00",X"3B",X"E8",X"41",X"86",X"04",X"08",X"0A",
		X"00",X"44",X"4F",X"10",X"13",X"04",X"05",X"0A",X"00",X"45",X"AD",X"10",X"29",X"04",X"08",X"0A",
		X"00",X"44",X"4F",X"68",X"13",X"04",X"05",X"0A",X"00",X"45",X"AD",X"68",X"29",X"15",X"04",X"12",
		X"88",X"00",X"00",X"13",X"13",X"15",X"04",X"12",X"88",X"00",X"00",X"6B",X"13",X"14",X"01",X"12",
		X"88",X"00",X"00",X"13",X"2D",X"14",X"01",X"12",X"88",X"00",X"00",X"6B",X"2D",X"01",X"0F",X"12",
		X"88",X"00",X"00",X"10",X"1A",X"01",X"0F",X"12",X"88",X"00",X"00",X"68",X"1A",X"01",X"0F",X"12",
		X"88",X"00",X"00",X"29",X"1A",X"01",X"0F",X"12",X"88",X"00",X"00",X"81",X"1A",X"13",X"1B",X"0A",
		X"00",X"3E",X"28",X"41",X"0A",X"12",X"0B",X"2A",X"00",X"44",X"6F",X"41",X"25",X"08",X"0F",X"0A",
		X"00",X"45",X"35",X"47",X"30",X"00",X"00",X"70",X"08",X"12",X"00",X"00",X"00",X"00",X"F8",X"00",
		X"00",X"CC",X"01",X"7A",X"BD",X"01",X"63",X"AF",X"2B",X"31",X"84",X"CC",X"11",X"18",X"8E",X"3A",
		X"D0",X"BD",X"18",X"D2",X"CC",X"10",X"0D",X"8E",X"3D",X"AA",X"BD",X"18",X"D2",X"BD",X"00",X"5A",
		X"8E",X"3A",X"D0",X"10",X"8E",X"07",X"30",X"CC",X"0A",X"19",X"8D",X"31",X"BD",X"00",X"5A",X"8E",
		X"3D",X"AA",X"10",X"8E",X"07",X"DF",X"CC",X"09",X"0E",X"8D",X"22",X"BD",X"00",X"5A",X"AE",X"2B",
		X"10",X"8E",X"84",X"30",X"CC",X"0A",X"19",X"8D",X"14",X"BD",X"00",X"5A",X"AE",X"2B",X"30",X"89",
		X"00",X"FA",X"10",X"8E",X"84",X"DF",X"CC",X"09",X"0E",X"8D",X"02",X"20",X"C0",X"34",X"01",X"1A",
		X"50",X"10",X"BF",X"CA",X"04",X"BF",X"CA",X"02",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"D6",
		X"54",X"C1",X"02",X"2C",X"05",X"86",X"0E",X"B7",X"CA",X"00",X"35",X"81",X"8E",X"40",X"29",X"8D",
		X"18",X"86",X"0A",X"BD",X"00",X"5C",X"8D",X"51",X"86",X"0A",X"BD",X"00",X"5C",X"8E",X"3E",X"28",
		X"8D",X"07",X"86",X"0A",X"BD",X"00",X"5C",X"20",X"E3",X"10",X"8E",X"41",X"0A",X"CC",X"13",X"1B",
		X"20",X"70",X"86",X"05",X"A7",X"2B",X"8D",X"31",X"86",X"03",X"BD",X"00",X"5C",X"8E",X"40",X"29",
		X"8D",X"E7",X"86",X"03",X"BD",X"00",X"5C",X"6A",X"2B",X"10",X"27",X"C6",X"2C",X"8E",X"3E",X"28",
		X"8D",X"D7",X"86",X"03",X"BD",X"00",X"5C",X"20",X"DD",X"34",X"20",X"86",X"15",X"BD",X"00",X"EE",
		X"BD",X"00",X"AD",X"25",X"16",X"3A",X"42",X"35",X"A0",X"CE",X"3A",X"8B",X"BD",X"08",X"38",X"8E",
		X"42",X"2A",X"10",X"8E",X"41",X"0A",X"CC",X"12",X"1B",X"20",X"27",X"14",X"1B",X"12",X"AA",X"00",
		X"00",X"41",X"0A",X"00",X"00",X"8E",X"40",X"29",X"8D",X"9F",X"86",X"0F",X"BD",X"00",X"5C",X"8D",
		X"D8",X"86",X"0F",X"BD",X"00",X"5C",X"8E",X"3E",X"28",X"8D",X"8E",X"86",X"0F",X"BD",X"00",X"5C",
		X"20",X"E3",X"34",X"01",X"1A",X"50",X"10",X"BF",X"CA",X"04",X"BF",X"CA",X"02",X"88",X"04",X"C8",
		X"04",X"FD",X"CA",X"06",X"86",X"02",X"B7",X"CA",X"00",X"35",X"81",X"AE",X"2B",X"7E",X"01",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AD",X"08",X"88",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"D8",
		X"88",X"88",X"88",X"88",X"AA",X"AA",X"AA",X"AA",X"D8",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",
		X"AA",X"D8",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AA",X"AD",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"AA",X"AA",X"D8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"AD",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"A8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"AA",X"D8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"AA",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"AD",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"A8",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"A8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"D8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"08",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",
		X"80",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"88",X"88",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"80",X"00",X"00",X"00",
		X"00",X"00",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0C",X"04",X"0F",X"02",X"11",
		X"01",X"12",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"01",X"12",X"02",X"11",X"04",X"0F",
		X"06",X"0D",X"3B",X"CA",X"23",X"18",X"16",X"1D",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",
		X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",
		X"66",X"DD",X"DD",X"66",X"DD",X"66",X"DD",X"DD",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"66",X"DD",X"DD",X"DD",X"D6",X"DD",X"6D",X"DD",X"DD",X"DD",X"66",X"60",X"00",X"00",X"00",
		X"00",X"00",X"66",X"DD",X"6D",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D6",X"DD",X"66",X"00",
		X"00",X"00",X"00",X"06",X"68",X"6D",X"DA",X"D6",X"66",X"66",X"66",X"66",X"66",X"6D",X"AD",X"D6",
		X"86",X"60",X"00",X"00",X"00",X"66",X"D6",X"DD",X"DD",X"66",X"6D",X"88",X"88",X"88",X"D6",X"66",
		X"DD",X"DD",X"6D",X"66",X"00",X"00",X"06",X"6D",X"66",X"68",X"66",X"68",X"88",X"88",X"80",X"80",
		X"80",X"06",X"66",X"86",X"66",X"D6",X"60",X"00",X"66",X"D6",X"66",X"86",X"68",X"88",X"88",X"08",
		X"80",X"80",X"80",X"00",X"06",X"68",X"66",X"6D",X"66",X"00",X"6D",X"66",X"A8",X"66",X"88",X"88",
		X"88",X"08",X"80",X"80",X"80",X"08",X"00",X"66",X"8A",X"66",X"D6",X"00",X"6D",X"DD",X"DD",X"68",
		X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"08",X"00",X"0A",X"DD",X"DD",X"D6",X"00",X"6D",X"D6",
		X"AD",X"A8",X"88",X"80",X"0F",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"0A",X"DA",X"6D",X"D6",X"00",
		X"6D",X"DD",X"DD",X"A8",X"88",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"0A",X"DD",X"DD",
		X"D6",X"00",X"6D",X"DD",X"DD",X"A8",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0A",
		X"DD",X"DD",X"D6",X"00",X"6D",X"66",X"A8",X"6A",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"A6",X"8A",X"66",X"D6",X"00",X"66",X"D6",X"66",X"86",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FA",X"68",X"66",X"6D",X"66",X"00",X"06",X"6D",X"66",X"A8",X"6A",X"6F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"F6",X"A6",X"8A",X"66",X"D6",X"60",X"00",X"08",X"6A",X"D6",X"DD",X"DD",X"6A",
		X"6F",X"FF",X"FF",X"FF",X"F6",X"A6",X"DD",X"DD",X"6D",X"66",X"80",X"00",X"00",X"86",X"6D",X"6D",
		X"DA",X"D6",X"AA",X"AA",X"AA",X"AA",X"AA",X"6D",X"AD",X"D6",X"8A",X"68",X"00",X"00",X"00",X"08",
		X"6A",X"DD",X"6D",X"DD",X"DD",X"8D",X"DD",X"D8",X"DD",X"DD",X"D6",X"DD",X"66",X"80",X"00",X"00",
		X"00",X"00",X"86",X"A6",X"DD",X"DD",X"DD",X"DA",X"DD",X"AD",X"DD",X"DD",X"DD",X"6A",X"68",X"00",
		X"00",X"00",X"00",X"00",X"08",X"D6",X"A6",X"DD",X"DD",X"66",X"DD",X"66",X"DD",X"DD",X"6A",X"6D",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"D6",X"A6",X"DD",X"DD",X"DD",X"DD",X"DD",X"6A",
		X"6D",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"D6",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"6D",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"D8",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"D8",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"88",
		X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"A0",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"AA",X"D8",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"AD",X"88",X"88",X"80",X"00",X"00",X"00",X"00",X"AA",X"AA",X"D8",X"88",X"88",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"AD",X"88",X"88",X"80",X"00",X"00",X"00",X"AA",X"AA",X"AA",
		X"AD",X"88",X"88",X"80",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AD",X"88",X"88",X"88",X"88",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AD",X"08",X"88",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"66",X"66",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"61",X"11",X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"D1",X"11",X"11",X"1D",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"D1",X"11",X"11",X"1D",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"66",X"11",
		X"11",X"66",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D1",X"16",X"66",X"66",X"61",X"1D",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"66",X"A6",X"66",X"66",X"66",X"81",X"18",X"66",X"66",X"66",X"6A",X"66",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"6A",X"11",X"11",X"11",X"11",X"86",X"1D",X"D1",X"68",X"11",X"11",X"11",X"11",X"A6",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"11",X"11",X"11",X"11",X"66",X"D6",X"81",X"18",X"6D",X"66",X"11",
		X"11",X"11",X"11",X"A6",X"AA",X"AA",X"A6",X"11",X"17",X"17",X"17",X"18",X"11",X"68",X"66",X"66",
		X"86",X"11",X"81",X"71",X"71",X"71",X"11",X"6A",X"AA",X"61",X"A7",X"A6",X"A6",X"AD",X"A8",X"11",
		X"18",X"88",X"88",X"81",X"11",X"8A",X"DA",X"6A",X"6A",X"7A",X"16",X"AA",X"AA",X"A6",X"AD",X"AD",
		X"AD",X"A8",X"81",X"81",X"1D",X"D1",X"18",X"18",X"8A",X"DA",X"DA",X"DA",X"6A",X"AA",X"AA",X"66",
		X"AD",X"AD",X"AD",X"A8",X"A8",X"68",X"D1",X"17",X"71",X"1D",X"86",X"8A",X"8A",X"DA",X"DA",X"DA",
		X"66",X"AA",X"6D",X"A8",X"A8",X"A8",X"A8",X"A8",X"6D",X"81",X"11",X"11",X"18",X"D6",X"8A",X"8A",
		X"8A",X"8A",X"8A",X"D6",X"AA",X"D8",X"68",X"68",X"68",X"68",X"68",X"6D",X"81",X"11",X"11",X"18",
		X"D6",X"86",X"86",X"86",X"86",X"86",X"8D",X"AA",X"A8",X"88",X"88",X"88",X"88",X"88",X"6D",X"81",
		X"11",X"11",X"18",X"D6",X"88",X"88",X"88",X"88",X"88",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"6D",X"81",X"11",X"11",X"18",X"D6",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"8D",X"81",X"11",X"11",X"18",X"D8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"81",X"11",X"11",X"18",X"8A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"81",X"11",X"11",X"18",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"81",X"11",
		X"11",X"18",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"61",X"81",X"77",X"77",X"18",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"61",X"16",X"87",X"76",X"67",X"78",X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"6D",X"87",X"66",X"66",X"78",X"D8",X"88",X"88",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"1A",X"DD",X"88",X"66",X"66",X"88",X"DD",X"88",
		X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"AD",X"DD",X"D8",X"88",X"88",
		X"8D",X"DD",X"68",X"88",X"88",X"86",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"66",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"66",X"61",X"11",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"11",X"11",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"A6",X"11",X"11",X"11",X"1D",X"66",X"6A",
		X"AA",X"66",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"AD",X"A6",X"11",X"11",
		X"16",X"11",X"6D",X"66",X"11",X"11",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"6D",
		X"AD",X"A6",X"6D",X"66",X"66",X"D6",X"11",X"11",X"11",X"11",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"88",X"AD",X"61",X"66",X"11",X"81",X"66",X"A1",X"11",X"11",X"1A",X"16",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"68",X"11",X"86",X"8D",X"D8",X"68",X"66",X"1A",X"6A",X"6A",
		X"6A",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"88",X"66",X"D6",X"18",X"11",X"6D",X"16",
		X"6A",X"DA",X"DA",X"DA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"11",X"D8",X"66",
		X"66",X"86",X"16",X"DA",X"DA",X"DA",X"86",X"8A",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"11",
		X"16",X"66",X"88",X"88",X"68",X"A8",X"DA",X"DA",X"86",X"88",X"DA",X"AA",X"AA",X"AA",X"AA",X"61",
		X"11",X"11",X"11",X"DA",X"11",X"16",X"D1",X"11",X"88",X"D6",X"88",X"88",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"11",X"11",X"11",X"6A",X"88",X"11",X"16",X"11",X"11",X"11",X"88",X"86",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"1A",X"DA",X"86",X"88",X"8D",X"A1",X"11",X"11",X"16",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"6A",X"DA",X"86",X"6D",X"D8",X"A7",
		X"11",X"11",X"11",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"11",X"11",X"1A",X"DA",X"8A",X"86",
		X"6D",X"D8",X"A6",X"A1",X"11",X"11",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"16",X"71",X"6A",
		X"DA",X"86",X"86",X"6D",X"D8",X"AD",X"A7",X"11",X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"66",X"61",X"DA",X"86",X"88",X"8D",X"6D",X"D8",X"AD",X"A6",X"11",X"11",X"11",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"A8",X"66",X"6A",X"D6",X"88",X"DA",X"AD",X"8D",X"D8",X"68",X"AD",X"A1",X"11",X"11",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"66",X"88",X"DA",X"AA",X"A6",X"D8",X"88",X"88",X"6D",
		X"A7",X"17",X"77",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"DA",X"AA",X"AA",X"A6",X"AA",
		X"AD",X"D8",X"88",X"A6",X"17",X"66",X"76",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"61",X"DA",X"66",X"D8",X"88",X"6D",X"A6",X"66",X"68",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A6",X"61",X"1D",X"D8",X"88",X"88",X"8D",X"8D",X"66",X"66",X"86",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"DD",X"88",X"6A",X"66",X"88",X"68",X"88",X"88",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",X"11",X"1D",X"DD",X"8A",X"A6",X"66",X"68",X"D6",
		X"88",X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"6D",X"DD",X"8A",X"66",
		X"66",X"68",X"DD",X"68",X"88",X"88",X"86",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"66",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"11",X"17",X"67",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"11",X"11",X"11",X"16",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"66",X"AA",X"A6",X"66",X"D1",X"11",X"11",X"11",X"7A",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"11",X"11",X"66",X"D1",X"11",X"61",X"11",X"11",
		X"7A",X"6A",X"DA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"11",X"11",X"11",X"11",X"66",X"66",X"66",
		X"6A",X"66",X"6A",X"D6",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"A1",X"11",X"11",X"11",X"16",
		X"18",X"18",X"6D",X"16",X"DA",X"86",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"A6",X"A6",X"A7",X"A1",
		X"16",X"D6",X"1D",X"D1",X"68",X"61",X"86",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AD",X"AD",
		X"A6",X"A6",X"61",X"D6",X"81",X"81",X"6D",X"66",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",
		X"68",X"AD",X"AD",X"AD",X"61",X"68",X"66",X"66",X"8D",X"11",X"11",X"16",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"88",X"68",X"AD",X"AD",X"8A",X"86",X"88",X"88",X"6A",X"61",X"11",X"11",X"16",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"68",X"1D",X"D8",X"11",X"16",X"D1",X"11",X"1D",X"11",X"11",
		X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"88",X"11",X"11",X"11",X"61",X"11",X"8D",
		X"A7",X"11",X"11",X"11",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"61",X"11",X"11",X"1A",X"D8",
		X"88",X"68",X"A6",X"A1",X"11",X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"11",X"11",X"11",
		X"7A",X"8D",X"DD",X"68",X"AD",X"A7",X"11",X"11",X"16",X"AA",X"AA",X"AA",X"AA",X"AA",X"A1",X"11",
		X"11",X"1A",X"6A",X"8D",X"DD",X"68",X"AD",X"A6",X"A1",X"17",X"71",X"6A",X"AA",X"AA",X"AA",X"AA",
		X"61",X"11",X"11",X"7A",X"DA",X"8D",X"DD",X"68",X"68",X"AD",X"A7",X"17",X"67",X"6A",X"AA",X"AA",
		X"AA",X"A6",X"11",X"11",X"1A",X"6A",X"DA",X"8D",X"DD",X"88",X"88",X"6D",X"AD",X"76",X"66",X"6A",
		X"AA",X"AA",X"AA",X"A1",X"17",X"11",X"1A",X"DA",X"86",X"8D",X"D8",X"6A",X"A8",X"88",X"6D",X"76",
		X"66",X"8A",X"AA",X"AA",X"AA",X"61",X"76",X"11",X"7A",X"D6",X"88",X"88",X"88",X"8A",X"AA",X"A8",
		X"88",X"A6",X"88",X"AA",X"AA",X"AA",X"AA",X"66",X"66",X"61",X"6A",X"88",X"8A",X"66",X"68",X"8A",
		X"AA",X"AA",X"A8",X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"66",X"67",X"D6",X"86",X"A6",X"66",
		X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"66",X"66",X"D8",X"68",
		X"88",X"88",X"8D",X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"88",X"D8",
		X"86",X"88",X"6A",X"66",X"88",X"D8",X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"61",
		X"11",X"1A",X"6D",X"8A",X"A6",X"66",X"68",X"DD",X"88",X"88",X"88",X"6A",X"AA",X"AA",X"AA",X"AA",
		X"61",X"11",X"11",X"A6",X"DD",X"8A",X"66",X"66",X"68",X"DD",X"D8",X"88",X"88",X"86",X"AA",X"AA",
		X"96",X"00",X"10",X"2A",X"BC",X"73",X"CC",X"00",X"0B",X"33",X"A5",X"8E",X"D0",X"DB",X"1E",X"01",
		X"9F",X"15",X"30",X"89",X"0C",X"03",X"34",X"46",X"34",X"10",X"8E",X"02",X"1E",X"1E",X"13",X"34",
		X"50",X"CE",X"44",X"3F",X"C6",X"0F",X"A6",X"C5",X"43",X"A7",X"85",X"5A",X"2A",X"F8",X"39",X"CA",
		X"D9",X"1F",X"5F",X"7D",X"FF",X"DB",X"05",X"A3",X"D8",X"FB",X"79",X"7F",X"68",X"EA",X"C6",X"AD",
		X"88",X"88",X"00",X"D8",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",X"88",X"88",X"00",X"88",
		X"80",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"AA",
		X"A6",X"11",X"11",X"A6",X"DD",X"8A",X"6A",X"66",X"66",X"68",X"DD",X"68",X"88",X"88",X"8A",X"AA",
		X"00",X"AA",X"61",X"11",X"1A",X"6D",X"D8",X"6A",X"6A",X"6A",X"66",X"66",X"8D",X"D6",X"88",X"88",
		X"86",X"AA",X"00",X"AA",X"61",X"11",X"A6",X"DD",X"D8",X"AA",X"6A",X"6A",X"66",X"66",X"8D",X"DD",
		X"68",X"88",X"88",X"AA",X"00",X"A6",X"11",X"1A",X"6D",X"DD",X"D8",X"AA",X"61",X"6A",X"6A",X"66",
		X"8D",X"DD",X"D6",X"88",X"88",X"6A",X"00",X"A6",X"11",X"A6",X"DD",X"DD",X"D8",X"AA",X"61",X"66",
		X"6A",X"66",X"8D",X"DD",X"DD",X"68",X"88",X"8A",X"00",X"61",X"1A",X"6D",X"DD",X"DD",X"D8",X"AA",
		X"61",X"16",X"AA",X"66",X"8D",X"DD",X"DD",X"D6",X"88",X"86",X"00",X"61",X"A6",X"DD",X"DD",X"DD",
		X"D8",X"AA",X"AA",X"11",X"AA",X"A6",X"8D",X"DD",X"DD",X"DD",X"68",X"88",X"00",X"6A",X"AA",X"A6",
		X"A6",X"D6",X"68",X"AA",X"11",X"1A",X"AA",X"A6",X"8D",X"66",X"DD",X"66",X"6A",X"88",X"00",X"88",
		X"88",X"88",X"88",X"88",X"88",X"AA",X"1A",X"66",X"6D",X"D6",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"A6",X"99",X"99",X"99",X"99",X"98",X"A1",X"A1",X"11",X"A6",X"D8",X"89",X"99",X"99",X"99",
		X"99",X"6A",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"11",X"A1",X"1A",X"A6",X"68",X"8A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"00",X"8D",X"1A",X"A1",X"1A",X"A6",X"6D",X"88",X"00",X"8D",X"1A",X"A1",
		X"AA",X"A6",X"6D",X"88",X"00",X"8D",X"1A",X"A1",X"A6",X"A6",X"6D",X"88",X"00",X"8D",X"1A",X"A1",
		X"AA",X"A6",X"6D",X"88",X"00",X"8D",X"1A",X"A1",X"A6",X"A6",X"6D",X"88",X"00",X"86",X"1A",X"A1",
		X"A6",X"A8",X"6D",X"D8",X"00",X"68",X"1A",X"A1",X"A6",X"A6",X"6D",X"DD",X"00",X"A8",X"1A",X"A1",
		X"A6",X"A8",X"6D",X"86",X"00",X"A8",X"1A",X"61",X"A6",X"18",X"6D",X"86",X"00",X"A6",X"81",X"61",
		X"AD",X"A8",X"68",X"66",X"00",X"61",X"68",X"61",X"A6",X"68",X"86",X"AD",X"00",X"DD",X"11",X"68",
		X"88",X"86",X"AA",X"DD",X"00",X"8D",X"6A",X"11",X"11",X"11",X"AD",X"D8",X"00",X"88",X"DD",X"66",
		X"AA",X"66",X"DD",X"88",X"00",X"88",X"80",X"DD",X"DD",X"DD",X"08",X"88",X"00",X"88",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"D8",X"00",X"00",X"00",X"AD",X"88",X"88",
		X"00",X"CE",X"46",X"28",X"8D",X"50",X"26",X"F9",X"A6",X"41",X"27",X"08",X"8D",X"48",X"27",X"FC",
		X"33",X"41",X"20",X"F0",X"1A",X"FF",X"BD",X"D2",X"1E",X"CC",X"00",X"FF",X"FD",X"C0",X"00",X"10",
		X"8E",X"46",X"2D",X"8E",X"10",X"30",X"34",X"10",X"C6",X"11",X"A6",X"A0",X"88",X"9B",X"80",X"35",
		X"2B",X"10",X"27",X"05",X"BD",X"7B",X"00",X"20",X"F1",X"AE",X"E4",X"30",X"88",X"10",X"AF",X"E4",
		X"20",X"E8",X"8E",X"1B",X"E6",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"13",X"27",X"F4",X"30",X"1F",
		X"26",X"F3",X"6E",X"9F",X"FF",X"FE",X"34",X"40",X"86",X"1E",X"BD",X"00",X"09",X"35",X"40",X"A6",
		X"9F",X"98",X"0E",X"A0",X"C4",X"91",X"31",X"39",X"15",X"32",X"26",X"18",X"00",X"C8",X"DC",X"D3",
		X"C9",X"A4",X"D3",X"C9",X"A4",X"DA",X"CF",X"DA",X"DA",X"D0",X"DF",X"C9",X"AE",X"D8",X"DF",X"C9",
		X"D3",X"DD",X"D6",X"DF",X"D8",X"A4",X"DA",X"C3",X"A4",X"CD",X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",
		X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",
		X"D9",X"F8",X"AE",X"C4",X"D9",X"FB",X"A4",X"AD",X"A5",X"A6",X"A3",X"A4",X"CD",X"D3",X"D0",X"D0",
		X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",
		X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",X"DB",X"D0",X"D0",X"A4",X"CA",X"D3",X"DD",X"DC",X"C8",X"C9",
		X"A4",X"CA",X"DF",X"C9",X"DF",X"CA",X"CE",X"DF",X"D8",X"2E",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"48",X"88",X"12",X"0C",X"0E",X"09",X"00",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"CC",X"B3",X"C3",X"BC",X"C0",X"00",X"00",X"00",X"00",X"0C",X"C1",X"1B",X"CB",
		X"11",X"CC",X"00",X"00",X"00",X"0C",X"CC",X"C1",X"49",X"11",X"49",X"CC",X"CC",X"00",X"00",X"33",
		X"3C",X"CC",X"11",X"81",X"1C",X"CC",X"33",X"30",X"00",X"55",X"33",X"3C",X"CC",X"CC",X"CC",X"33",
		X"35",X"50",X"00",X"39",X"55",X"33",X"3C",X"CC",X"33",X"35",X"59",X"C0",X"02",X"09",X"39",X"55",
		X"33",X"C3",X"35",X"59",X"C9",X"E0",X"A0",X"92",X"09",X"39",X"55",X"25",X"59",X"C9",X"E9",X"00",
		X"09",X"A0",X"92",X"09",X"39",X"59",X"C9",X"E9",X"90",X"00",X"00",X"09",X"A0",X"92",X"49",X"39",
		X"E9",X"90",X"00",X"00",X"00",X"00",X"09",X"A0",X"92",X"9E",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"A9",X"00",X"00",X"00",X"00",X"00",X"09",X"0B",X"06",X"0E",X"05",X"0F",X"03",X"11",
		X"02",X"12",X"02",X"12",X"02",X"12",X"01",X"12",X"00",X"11",X"01",X"10",X"03",X"0E",X"05",X"0C",
		X"07",X"09",X"49",X"2A",X"12",X"0C",X"0E",X"09",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"B3",X"C3",X"BC",X"C0",X"00",X"00",X"00",X"00",X"0C",X"C1",X"1B",
		X"CB",X"11",X"CC",X"00",X"00",X"00",X"0C",X"CC",X"C9",X"41",X"19",X"41",X"CC",X"CC",X"00",X"00",
		X"33",X"3C",X"CC",X"11",X"81",X"1C",X"CC",X"33",X"30",X"00",X"55",X"33",X"3C",X"CC",X"CC",X"CC",
		X"33",X"35",X"50",X"00",X"39",X"55",X"33",X"3C",X"CC",X"33",X"35",X"59",X"C0",X"00",X"29",X"39",
		X"55",X"33",X"C3",X"35",X"59",X"C9",X"0E",X"00",X"09",X"29",X"39",X"55",X"25",X"59",X"C9",X"0E",
		X"90",X"A0",X"00",X"99",X"29",X"39",X"59",X"C9",X"0E",X"90",X"A9",X"00",X"00",X"00",X"99",X"29",
		X"39",X"0E",X"90",X"A9",X"00",X"00",X"00",X"00",X"00",X"93",X"9E",X"90",X"A9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"A9",X"00",X"00",X"00",X"00",X"07",X"09",X"04",X"0C",X"03",X"0D",
		X"01",X"0F",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"01",X"12",X"02",X"11",X"04",X"0F",
		X"06",X"0D",X"09",X"0B",X"49",X"BF",X"10",X"0C",X"0D",X"09",X"00",X"00",X"00",X"0C",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"CC",X"B3",X"C3",X"BC",X"C0",X"00",X"00",X"00",X"0C",X"C1",X"1B",
		X"CB",X"11",X"CC",X"00",X"00",X"0C",X"CC",X"C1",X"99",X"19",X"91",X"CC",X"CC",X"00",X"33",X"3C",
		X"CC",X"11",X"81",X"1C",X"CC",X"33",X"30",X"55",X"33",X"3C",X"CC",X"CC",X"CC",X"33",X"35",X"50",
		X"39",X"55",X"33",X"3C",X"CC",X"33",X"35",X"59",X"C0",X"29",X"39",X"55",X"33",X"C3",X"35",X"59",
		X"C9",X"C0",X"29",X"29",X"39",X"55",X"25",X"59",X"C9",X"C9",X"E0",X"19",X"29",X"29",X"39",X"59",
		X"C9",X"C9",X"E9",X"E0",X"09",X"19",X"29",X"29",X"39",X"C9",X"E9",X"E9",X"00",X"00",X"09",X"19",
		X"29",X"29",X"E9",X"79",X"00",X"00",X"00",X"00",X"09",X"19",X"19",X"79",X"00",X"00",X"00",X"07",
		X"09",X"04",X"0C",X"03",X"0D",X"01",X"0F",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",
		X"10",X"00",X"10",X"01",X"0F",X"03",X"0D",X"05",X"0B",X"4A",X"27",X"10",X"07",X"0D",X"0C",X"00",
		X"00",X"C3",X"32",X"32",X"33",X"C0",X"00",X"00",X"00",X"C3",X"34",X"34",X"44",X"34",X"33",X"C0",
		X"00",X"03",X"54",X"11",X"99",X"19",X"91",X"15",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",
		X"33",X"43",X"30",X"39",X"34",X"55",X"55",X"55",X"55",X"54",X"39",X"30",X"0E",X"39",X"53",X"22",
		X"22",X"23",X"59",X"33",X"00",X"00",X"43",X"34",X"3C",X"CC",X"34",X"33",X"C0",X"00",X"00",X"00",
		X"43",X"35",X"93",X"43",X"C0",X"00",X"00",X"04",X"0C",X"02",X"0E",X"01",X"0F",X"00",X"10",X"00",
		X"10",X"01",X"0F",X"02",X"0E",X"04",X"0C",X"4A",X"85",X"0E",X"08",X"0C",X"0D",X"00",X"00",X"33",
		X"43",X"43",X"30",X"00",X"00",X"00",X"33",X"11",X"D4",X"D1",X"13",X"30",X"00",X"03",X"C1",X"19",
		X"51",X"59",X"11",X"33",X"00",X"33",X"34",X"11",X"15",X"11",X"14",X"53",X"30",X"35",X"33",X"39",
		X"99",X"99",X"33",X"E4",X"30",X"33",X"43",X"99",X"99",X"99",X"93",X"43",X"30",X"49",X"33",X"99",
		X"94",X"99",X"93",X"39",X"30",X"0E",X"C3",X"32",X"33",X"24",X"34",X"3C",X"00",X"00",X"03",X"43",
		X"59",X"33",X"43",X"C0",X"00",X"04",X"0A",X"02",X"0C",X"01",X"0D",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"01",X"0D",X"03",X"0C",X"4A",X"B1",X"06",X"04",X"00",X"01",X"00",X"06",X"7D",
		X"00",X"D2",X"51",X"B1",X"D0",X"72",X"31",X"36",X"10",X"20",X"7B",X"32",X"30",X"01",X"CC",X"A6",
		X"B0",X"03",X"05",X"00",X"06",X"00",X"06",X"00",X"06",X"01",X"06",X"4A",X"EE",X"08",X"08",X"01",
		X"0D",X"00",X"00",X"55",X"50",X"00",X"05",X"50",X"55",X"55",X"00",X"55",X"58",X"55",X"58",X"00",
		X"55",X"55",X"58",X"00",X"00",X"09",X"55",X"55",X"88",X"00",X"55",X"59",X"85",X"55",X"80",X"08",
		X"80",X"08",X"55",X"80",X"00",X"05",X"50",X"88",X"00",X"00",X"08",X"80",X"00",X"00",X"04",X"06",
		X"01",X"07",X"00",X"07",X"00",X"05",X"01",X"07",X"00",X"08",X"01",X"08",X"03",X"07",X"03",X"04",
		X"4B",X"12",X"02",X"05",X"06",X"02",X"0D",X"00",X"06",X"00",X"06",X"00",X"DA",X"D0",X"D6",X"D0",
		X"0D",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"02",X"00",X"02",X"01",X"01",X"4B",X"A2",
		X"0F",X"0D",X"0D",X"0A",X"00",X"D6",X"86",X"A0",X"00",X"00",X"00",X"00",X"00",X"06",X"6D",X"6D",
		X"61",X"00",X"00",X"00",X"00",X"00",X"D6",X"D6",X"66",X"D6",X"A0",X"00",X"00",X"00",X"00",X"0D",
		X"66",X"88",X"6D",X"61",X"00",X"00",X"00",X"00",X"16",X"D6",X"88",X"66",X"D6",X"A0",X"00",X"00",
		X"00",X"0A",X"6D",X"66",X"86",X"6D",X"6A",X"00",X"00",X"00",X"00",X"A6",X"D6",X"68",X"86",X"D6",
		X"A0",X"00",X"00",X"00",X"0A",X"6D",X"68",X"86",X"6D",X"6A",X"00",X"00",X"00",X"00",X"A6",X"D6",
		X"68",X"66",X"D6",X"A0",X"00",X"00",X"00",X"01",X"6D",X"66",X"88",X"6D",X"61",X"00",X"00",X"00",
		X"00",X"A6",X"D6",X"88",X"66",X"60",X"00",X"00",X"00",X"00",X"0A",X"6D",X"66",X"6D",X"66",X"00",
		X"00",X"00",X"00",X"00",X"16",X"D6",X"D6",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"68",X"6D",
		X"00",X"00",X"02",X"06",X"01",X"07",X"00",X"08",X"01",X"09",X"00",X"0A",X"01",X"0B",X"02",X"0C",
		X"03",X"0D",X"04",X"0E",X"05",X"0F",X"06",X"0E",X"07",X"0F",X"08",X"0E",X"09",X"0D",X"4C",X"42",
		X"0F",X"0D",X"0D",X"0A",X"00",X"D6",X"86",X"10",X"00",X"00",X"00",X"00",X"00",X"06",X"6D",X"6D",
		X"6A",X"00",X"00",X"00",X"00",X"00",X"D6",X"D6",X"66",X"D6",X"10",X"00",X"00",X"00",X"00",X"0D",
		X"66",X"88",X"6D",X"6A",X"00",X"00",X"00",X"00",X"A6",X"D6",X"88",X"66",X"D6",X"A0",X"00",X"00",
		X"00",X"0A",X"6D",X"66",X"86",X"6D",X"6A",X"00",X"00",X"00",X"00",X"A6",X"D6",X"68",X"86",X"D6",
		X"10",X"00",X"00",X"00",X"01",X"6D",X"68",X"86",X"6D",X"6A",X"00",X"00",X"00",X"00",X"A6",X"D6",
		X"68",X"66",X"D6",X"A0",X"00",X"00",X"00",X"0A",X"6D",X"66",X"88",X"6D",X"6A",X"00",X"00",X"00",
		X"00",X"A6",X"D6",X"88",X"66",X"60",X"00",X"00",X"00",X"00",X"01",X"6D",X"66",X"6D",X"66",X"00",
		X"00",X"00",X"00",X"00",X"A6",X"D6",X"D6",X"60",X"00",X"00",X"00",X"00",X"00",X"01",X"68",X"6D",
		X"00",X"00",X"02",X"06",X"01",X"07",X"00",X"08",X"01",X"09",X"00",X"0A",X"01",X"0B",X"02",X"0C",
		X"03",X"0D",X"04",X"0E",X"05",X"0F",X"06",X"0E",X"07",X"0F",X"08",X"0E",X"09",X"0D",X"00",X"09",
		X"11",X"0F",X"4D",X"08",X"11",X"0F",X"0E",X"14",X"00",X"70",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"BB",X"BB",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"E3",X"EE",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"83",X"8E",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"3E",X"EE",X"66",X"DC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"34",X"E3",X"54",X"BB",X"CC",X"00",X"00",X"00",X"00",X"00",X"53",
		X"35",X"5E",X"EB",X"4C",X"00",X"00",X"00",X"00",X"00",X"EC",X"55",X"4E",X"E4",X"44",X"00",X"00",
		X"00",X"00",X"0C",X"E0",X"04",X"EE",X"44",X"44",X"00",X"00",X"21",X"00",X"EE",X"00",X"0E",X"E4",
		X"44",X"45",X"00",X"C2",X"4C",X"00",X"E9",X"99",X"EE",X"99",X"44",X"49",X"99",X"24",X"27",X"00",
		X"00",X"00",X"EE",X"04",X"94",X"44",X"00",X"C2",X"4C",X"00",X"00",X"00",X"00",X"09",X"90",X"49",
		X"90",X"00",X"21",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"02",X"05",X"03",X"04",X"01",X"06",X"01",X"07",
		X"00",X"07",X"01",X"0A",X"02",X"0B",X"02",X"0B",X"02",X"0B",X"01",X"11",X"00",X"11",X"00",X"11",
		X"04",X"11",X"07",X"11",X"06",X"0B",X"09",X"0A",X"00",X"09",X"11",X"0F",X"4D",X"D2",X"11",X"0F",
		X"0E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"BB",X"BB",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AB",X"EE",X"3E",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",
		X"E8",X"E8",X"E6",X"00",X"00",X"00",X"00",X"0C",X"CD",X"66",X"EE",X"E3",X"E0",X"00",X"00",X"00",
		X"00",X"CC",X"BB",X"45",X"3E",X"43",X"00",X"00",X"00",X"00",X"00",X"C4",X"BE",X"E5",X"53",X"35",
		X"00",X"00",X"00",X"00",X"00",X"44",X"4E",X"E4",X"55",X"CE",X"00",X"00",X"12",X"00",X"00",X"44",
		X"44",X"EE",X"40",X"0E",X"C0",X"00",X"C4",X"2C",X"00",X"54",X"44",X"4E",X"E0",X"00",X"EE",X"00",
		X"72",X"42",X"99",X"94",X"44",X"99",X"EE",X"99",X"9E",X"00",X"C4",X"2C",X"00",X"44",X"49",X"00",
		X"EE",X"00",X"00",X"00",X"12",X"00",X"09",X"94",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"0F",X"0D",X"0E",X"0B",X"10",X"0A",X"10",X"0A",X"11",X"07",X"10",X"06",X"0F",
		X"06",X"0F",X"06",X"0F",X"00",X"10",X"00",X"11",X"00",X"11",X"00",X"0D",X"00",X"0A",X"06",X"0B",
		X"07",X"08",X"00",X"00",X"04",X"0E",X"4E",X"92",X"11",X"0E",X"0E",X"0B",X"0D",X"EE",X"00",X"70",
		X"07",X"00",X"00",X"00",X"00",X"00",X"0E",X"9E",X"D0",X"07",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"E0",X"BB",X"BB",X"A0",X"00",X"00",X"00",X"00",X"00",X"90",X"0B",X"E3",X"EE",X"BA",
		X"00",X"00",X"00",X"00",X"00",X"90",X"0E",X"8E",X"8E",X"BA",X"00",X"00",X"00",X"00",X"00",X"90",
		X"0E",X"3E",X"EE",X"E5",X"4C",X"CC",X"00",X"00",X"00",X"9D",X"00",X"33",X"33",X"4B",X"B4",X"4C",
		X"C0",X"00",X"0E",X"EE",X"00",X"04",X"55",X"EE",X"B4",X"44",X"C0",X"00",X"0E",X"EE",X"EE",X"EE",
		X"EE",X"E4",X"54",X"44",X"C0",X"00",X"00",X"90",X"CC",X"CC",X"CC",X"55",X"44",X"44",X"49",X"00",
		X"00",X"90",X"00",X"00",X"55",X"5C",X"44",X"40",X"99",X"00",X"0C",X"2C",X"00",X"00",X"0C",X"44",
		X"44",X"09",X"90",X"00",X"02",X"42",X"00",X"99",X"99",X"44",X"40",X"00",X"00",X"00",X"24",X"24",
		X"20",X"09",X"99",X"54",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"01",X"09",X"01",X"08",X"02",X"0A",X"02",X"0B",X"02",X"0B",X"02",X"0F",X"02",X"10",
		X"01",X"10",X"01",X"10",X"02",X"11",X"02",X"11",X"01",X"10",X"01",X"0C",X"00",X"0B",X"00",X"0A",
		X"00",X"05",X"08",X"0F",X"4F",X"4A",X"10",X"0F",X"0D",X"14",X"00",X"00",X"00",X"70",X"07",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"BB",X"A0",X"00",X"00",X"00",X"EE",X"D0",X"0B",X"E3",X"EE",X"BA",X"00",X"00",X"00",X"E9",X"EE",
		X"CE",X"83",X"8E",X"BA",X"00",X"00",X"00",X"09",X"00",X"0E",X"3E",X"EE",X"65",X"4C",X"CC",X"00",
		X"00",X"90",X"00",X"39",X"E3",X"5B",X"B4",X"CC",X"C0",X"00",X"90",X"00",X"03",X"35",X"EE",X"B4",
		X"44",X"C0",X"00",X"09",X"00",X"00",X"5E",X"E3",X"54",X"44",X"C0",X"00",X"0D",X"EE",X"CC",X"EE",
		X"35",X"54",X"44",X"40",X"00",X"0E",X"DE",X"EE",X"E3",X"55",X"5C",X"44",X"40",X"00",X"00",X"90",
		X"00",X"00",X"09",X"5C",X"44",X"00",X"00",X"00",X"02",X"00",X"09",X"99",X"54",X"44",X"00",X"00",
		X"00",X"64",X"20",X"00",X"00",X"04",X"44",X"40",X"00",X"00",X"24",X"42",X"00",X"00",X"05",X"59",
		X"90",X"00",X"00",X"10",X"20",X"10",X"09",X"99",X"90",X"90",X"06",X"09",X"07",X"08",X"06",X"0A",
		X"00",X"0B",X"00",X"0B",X"01",X"0F",X"02",X"10",X"02",X"10",X"03",X"10",X"03",X"10",X"03",X"10",
		X"04",X"0F",X"05",X"0F",X"04",X"10",X"04",X"10",X"04",X"10",X"00",X"08",X"0E",X"11",X"50",X"28",
		X"12",X"11",X"0E",X"16",X"00",X"00",X"70",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"E3",X"EE",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"8E",X"8E",
		X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"3E",X"EE",X"65",X"BC",X"CC",X"00",X"00",X"00",
		X"0D",X"ED",X"39",X"9E",X"4E",X"EB",X"4C",X"C0",X"00",X"00",X"EE",X"D0",X"03",X"83",X"4E",X"EB",
		X"44",X"CC",X"00",X"00",X"29",X"00",X"00",X"34",X"4E",X"E5",X"44",X"4C",X"00",X"00",X"0C",X"90",
		X"00",X"55",X"4E",X"E5",X"44",X"4C",X"00",X"00",X"00",X"09",X"00",X"44",X"EE",X"55",X"44",X"4C",
		X"00",X"00",X"00",X"00",X"90",X"92",X"E5",X"55",X"54",X"44",X"40",X"00",X"00",X"00",X"0E",X"1E",
		X"99",X"55",X"55",X"44",X"49",X"00",X"00",X"00",X"01",X"90",X"00",X"00",X"05",X"54",X"49",X"90",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"23",X"60",
		X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"02",X"42",X"24",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"16",X"26",X"10",X"00",X"00",X"04",X"07",X"05",X"06",X"04",X"08",X"03",X"09",
		X"03",X"09",X"03",X"0D",X"01",X"0E",X"00",X"0F",X"00",X"0F",X"01",X"0F",X"03",X"0F",X"04",X"10",
		X"05",X"11",X"05",X"12",X"07",X"11",X"08",X"11",X"09",X"0D",X"0A",X"0E",X"0C",X"00",X"11",X"0E",
		X"50",X"EC",X"11",X"0E",X"0E",X"0B",X"00",X"00",X"00",X"00",X"70",X"07",X"00",X"EE",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"06",X"70",X"0D",X"E9",X"E0",X"00",X"00",X"00",X"00",X"0A",X"BB",X"BB",
		X"0E",X"09",X"00",X"00",X"00",X"00",X"00",X"AB",X"EE",X"3E",X"B0",X"09",X"00",X"00",X"00",X"00",
		X"00",X"AB",X"E8",X"E8",X"E0",X"09",X"00",X"00",X"00",X"CC",X"C4",X"5E",X"EE",X"E3",X"E0",X"09",
		X"00",X"00",X"0C",X"C4",X"4B",X"B4",X"33",X"33",X"00",X"D9",X"00",X"00",X"0C",X"44",X"4B",X"EE",
		X"55",X"40",X"00",X"EE",X"E0",X"00",X"0C",X"44",X"45",X"4E",X"EE",X"EE",X"EE",X"EE",X"E0",X"00",
		X"94",X"44",X"44",X"55",X"CC",X"CC",X"CC",X"09",X"00",X"00",X"99",X"04",X"44",X"C5",X"55",X"00",
		X"00",X"09",X"00",X"00",X"09",X"90",X"44",X"44",X"C0",X"00",X"00",X"C2",X"C0",X"00",X"00",X"00",
		X"04",X"44",X"99",X"99",X"00",X"24",X"20",X"00",X"00",X"00",X"00",X"45",X"99",X"90",X"02",X"42",
		X"42",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"01",X"07",X"01",X"00",X"08",X"10",X"09",X"10",
		X"07",X"0F",X"06",X"0F",X"06",X"0F",X"02",X"0F",X"01",X"0F",X"01",X"10",X"01",X"10",X"00",X"0F",
		X"00",X"0F",X"01",X"10",X"05",X"10",X"06",X"11",X"07",X"11",X"08",X"03",X"0F",X"10",X"51",X"A4",
		X"10",X"0F",X"0D",X"14",X"00",X"00",X"00",X"07",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"BB",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"BE",X"E3",X"EB",X"00",X"DE",X"E0",X"00",X"00",X"0A",X"BE",X"83",X"8E",X"CE",X"E9",
		X"E0",X"0C",X"CC",X"45",X"6E",X"EE",X"3E",X"00",X"09",X"00",X"CC",X"C4",X"BB",X"53",X"E9",X"30",
		X"00",X"90",X"00",X"C4",X"44",X"BE",X"E5",X"33",X"00",X"00",X"90",X"00",X"C4",X"44",X"53",X"EE",
		X"50",X"00",X"09",X"00",X"00",X"44",X"44",X"55",X"3E",X"EC",X"CE",X"ED",X"00",X"00",X"44",X"4C",
		X"55",X"53",X"EE",X"EE",X"DE",X"00",X"00",X"04",X"4C",X"59",X"00",X"00",X"00",X"90",X"00",X"00",
		X"04",X"44",X"59",X"99",X"00",X"02",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"24",X"60",
		X"00",X"00",X"99",X"55",X"00",X"00",X"02",X"44",X"20",X"00",X"00",X"90",X"99",X"99",X"00",X"10",
		X"20",X"10",X"00",X"00",X"07",X"0A",X"08",X"09",X"06",X"0A",X"05",X"10",X"05",X"10",X"01",X"0F",
		X"00",X"0E",X"00",X"0E",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"01",X"0C",X"01",X"0B",X"00",X"0C",
		X"00",X"0C",X"00",X"0C",X"04",X"07",X"10",X"12",X"52",X"82",X"12",X"11",X"0E",X"16",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"BB",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"BE",X"E3",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"BE",X"8E",X"8E",X"00",X"00",
		X"00",X"00",X"0C",X"CC",X"B5",X"6E",X"EE",X"32",X"00",X"00",X"00",X"00",X"CC",X"4B",X"EE",X"4E",
		X"99",X"3D",X"ED",X"00",X"00",X"0C",X"C4",X"4B",X"EE",X"43",X"83",X"00",X"DE",X"E0",X"00",X"0C",
		X"44",X"45",X"EE",X"44",X"30",X"00",X"09",X"20",X"00",X"0C",X"44",X"45",X"EE",X"45",X"50",X"00",
		X"9C",X"00",X"00",X"0C",X"44",X"45",X"5E",X"E4",X"40",X"09",X"00",X"00",X"00",X"44",X"44",X"55",
		X"55",X"E2",X"90",X"90",X"00",X"00",X"09",X"44",X"45",X"55",X"59",X"9E",X"1E",X"00",X"00",X"00",
		X"99",X"44",X"55",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"63",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"22",X"42",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"26",X"10",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"0E",X"0C",X"0D",X"0A",X"0E",X"09",X"0F",X"09",X"0F",X"05",X"0F",X"04",X"11",
		X"03",X"12",X"03",X"12",X"03",X"11",X"03",X"0F",X"02",X"0E",X"01",X"0D",X"00",X"0D",X"01",X"0B",
		X"01",X"0A",X"05",X"09",X"04",X"08",X"00",X"00",X"04",X"11",X"53",X"40",X"0F",X"11",X"0C",X"16",
		X"00",X"00",X"00",X"07",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"BB",X"BA",X"00",X"00",X"00",X"00",X"00",X"BE",X"3E",X"EB",X"A0",X"00",
		X"00",X"09",X"00",X"E8",X"E8",X"EB",X"A0",X"00",X"00",X"EE",X"00",X"E3",X"EE",X"E6",X"C0",X"00",
		X"00",X"E9",X"ED",X"E3",X"99",X"34",X"D0",X"00",X"00",X"09",X"00",X"4E",X"38",X"34",X"4D",X"00",
		X"00",X"09",X"04",X"44",X"33",X"45",X"EE",X"00",X"00",X"09",X"04",X"44",X"45",X"5E",X"EE",X"00",
		X"00",X"39",X"C0",X"55",X"5E",X"EE",X"E4",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"E4",X"54",X"00",
		X"00",X"09",X"04",X"44",X"44",X"55",X"54",X"00",X"00",X"09",X"00",X"44",X"44",X"45",X"54",X"00",
		X"00",X"C2",X"C0",X"59",X"94",X"44",X"54",X"00",X"00",X"24",X"20",X"99",X"00",X"44",X"44",X"00",
		X"02",X"43",X"20",X"00",X"00",X"09",X"99",X"00",X"10",X"10",X"20",X"00",X"00",X"00",X"99",X"00",
		X"07",X"0A",X"08",X"09",X"07",X"0B",X"06",X"0C",X"03",X"0C",X"02",X"0C",X"02",X"0C",X"03",X"0D",
		X"03",X"0D",X"03",X"0D",X"02",X"0D",X"02",X"0D",X"03",X"0D",X"03",X"0D",X"02",X"0D",X"02",X"0D",
		X"01",X"0D",X"00",X"0D",X"00",X"09",X"0C",X"11",X"53",X"EC",X"0F",X"11",X"03",X"16",X"00",X"00",
		X"60",X"06",X"00",X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",X"AB",X"BB",
		X"00",X"00",X"00",X"00",X"0A",X"E3",X"EE",X"30",X"00",X"00",X"00",X"AB",X"E8",X"38",X"EB",X"00",
		X"00",X"00",X"AB",X"3E",X"EE",X"E0",X"00",X"00",X"00",X"0E",X"33",X"93",X"54",X"00",X"00",X"DD",
		X"E5",X"E3",X"E3",X"5E",X"E0",X"00",X"EE",X"44",X"44",X"55",X"5E",X"EE",X"00",X"E9",X"04",X"44",
		X"45",X"55",X"EE",X"00",X"00",X"94",X"44",X"44",X"45",X"EE",X"00",X"00",X"49",X"44",X"45",X"5E",
		X"EE",X"00",X"00",X"44",X"9D",X"EE",X"EE",X"ED",X"00",X"00",X"44",X"4E",X"EE",X"44",X"80",X"00",
		X"00",X"44",X"4E",X"90",X"09",X"99",X"00",X"00",X"44",X"55",X"02",X"20",X"00",X"00",X"00",X"99",
		X"90",X"00",X"34",X"20",X"00",X"00",X"99",X"00",X"00",X"20",X"30",X"20",X"04",X"07",X"05",X"06",
		X"04",X"07",X"03",X"08",X"02",X"09",X"02",X"08",X"03",X"09",X"00",X"0A",X"00",X"0B",X"00",X"0B",
		X"02",X"0B",X"02",X"0B",X"02",X"0B",X"02",X"0A",X"02",X"0B",X"02",X"08",X"02",X"0A",X"02",X"0C",
		X"54",X"3E",X"06",X"09",X"00",X"0E",X"80",X"50",X"50",X"00",X"08",X"05",X"00",X"00",X"08",X"09",
		X"08",X"00",X"00",X"89",X"80",X"80",X"00",X"05",X"00",X"00",X"00",X"99",X"98",X"80",X"08",X"09",
		X"08",X"00",X"08",X"00",X"00",X"80",X"08",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"04",
		X"01",X"03",X"01",X"05",X"02",X"06",X"03",X"03",X"02",X"06",X"01",X"05",X"01",X"06",X"01",X"01",
		X"00",X"00",X"54",X"80",X"06",X"09",X"00",X"0E",X"00",X"50",X"50",X"80",X"00",X"05",X"08",X"00",
		X"08",X"09",X"08",X"00",X"80",X"89",X"80",X"00",X"00",X"05",X"00",X"00",X"88",X"99",X"90",X"00",
		X"08",X"09",X"08",X"00",X"80",X"00",X"08",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"80",
		X"02",X"06",X"03",X"05",X"01",X"05",X"00",X"04",X"03",X"03",X"00",X"04",X"01",X"05",X"00",X"05",
		X"05",X"05",X"06",X"06",X"54",X"C4",X"09",X"06",X"02",X"03",X"80",X"00",X"00",X"00",X"08",X"00",
		X"08",X"88",X"00",X"08",X"80",X"00",X"00",X"00",X"90",X"80",X"05",X"00",X"00",X"09",X"95",X"99",
		X"50",X"00",X"00",X"00",X"90",X"80",X"05",X"00",X"00",X"08",X"80",X"08",X"00",X"00",X"00",X"80",
		X"80",X"80",X"00",X"00",X"00",X"09",X"01",X"08",X"04",X"09",X"03",X"08",X"04",X"09",X"03",X"07",
		X"02",X"06",X"55",X"02",X"09",X"06",X"02",X"03",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"08",
		X"80",X"08",X"00",X"00",X"00",X"00",X"90",X"80",X"05",X"00",X"00",X"09",X"95",X"99",X"50",X"00",
		X"00",X"00",X"90",X"80",X"05",X"00",X"08",X"88",X"00",X"08",X"80",X"00",X"80",X"00",X"00",X"00",
		X"08",X"00",X"02",X"06",X"03",X"07",X"04",X"09",X"03",X"08",X"04",X"09",X"01",X"08",X"00",X"09",
		X"55",X"3E",X"06",X"09",X"00",X"0E",X"80",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"08",X"00",
		X"00",X"80",X"08",X"09",X"08",X"00",X"00",X"99",X"98",X"80",X"00",X"05",X"00",X"00",X"00",X"89",
		X"80",X"80",X"08",X"09",X"08",X"00",X"08",X"05",X"00",X"00",X"80",X"50",X"50",X"00",X"00",X"00",
		X"01",X"01",X"01",X"06",X"01",X"05",X"02",X"06",X"03",X"03",X"02",X"06",X"01",X"05",X"01",X"03",
		X"00",X"04",X"55",X"80",X"06",X"09",X"00",X"0E",X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"00",
		X"80",X"00",X"08",X"00",X"08",X"09",X"08",X"00",X"88",X"99",X"90",X"00",X"00",X"05",X"00",X"00",
		X"80",X"89",X"80",X"00",X"08",X"09",X"08",X"00",X"00",X"05",X"08",X"00",X"00",X"50",X"50",X"80",
		X"06",X"06",X"05",X"05",X"00",X"05",X"01",X"05",X"00",X"04",X"03",X"03",X"00",X"04",X"01",X"05",
		X"03",X"05",X"02",X"06",X"55",X"C4",X"09",X"06",X"02",X"03",X"80",X"00",X"00",X"00",X"08",X"00",
		X"08",X"80",X"00",X"88",X"80",X"00",X"50",X"08",X"09",X"00",X"00",X"00",X"05",X"99",X"59",X"90",
		X"00",X"00",X"50",X"08",X"09",X"00",X"00",X"00",X"00",X"80",X"08",X"80",X"00",X"00",X"00",X"08",
		X"08",X"08",X"00",X"00",X"00",X"09",X"01",X"08",X"00",X"05",X"01",X"06",X"00",X"05",X"02",X"06",
		X"03",X"07",X"56",X"02",X"09",X"06",X"02",X"03",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"80",
		X"08",X"80",X"00",X"00",X"50",X"08",X"09",X"00",X"00",X"00",X"05",X"99",X"59",X"90",X"00",X"00",
		X"50",X"08",X"09",X"00",X"00",X"00",X"08",X"80",X"00",X"88",X"80",X"00",X"80",X"00",X"00",X"00",
		X"08",X"00",X"03",X"07",X"02",X"06",X"00",X"05",X"01",X"06",X"00",X"05",X"01",X"08",X"00",X"09",
		X"06",X"04",X"00",X"01",X"44",X"40",X"00",X"00",X"00",X"40",X"40",X"40",X"04",X"40",X"04",X"00",
		X"40",X"00",X"40",X"40",X"44",X"40",X"00",X"00",X"04",X"05",X"07",X"02",X"10",X"70",X"10",X"24",
		X"24",X"20",X"02",X"42",X"00",X"0C",X"2C",X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"05",X"05",
		X"00",X"02",X"00",X"10",X"00",X"00",X"0E",X"00",X"00",X"00",X"02",X"42",X"00",X"00",X"0C",X"64",
		X"01",X"00",X"02",X"C2",X"E0",X"00",X"90",X"00",X"00",X"00",X"05",X"04",X"00",X"01",X"00",X"00",
		X"21",X"00",X"00",X"C2",X"40",X"00",X"99",X"24",X"27",X"00",X"00",X"C2",X"40",X"00",X"00",X"00",
		X"21",X"00",X"05",X"05",X"00",X"02",X"90",X"00",X"00",X"00",X"02",X"C2",X"E0",X"00",X"0C",X"64",
		X"01",X"00",X"02",X"42",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"04",X"05",
		X"07",X"02",X"00",X"90",X"00",X"00",X"90",X"00",X"0C",X"2C",X"00",X"02",X"42",X"00",X"24",X"24",
		X"20",X"10",X"70",X"10",X"05",X"05",X"00",X"02",X"00",X"00",X"09",X"00",X"0E",X"2C",X"20",X"00",
		X"10",X"46",X"C0",X"00",X"00",X"24",X"20",X"00",X"00",X"00",X"E0",X"00",X"00",X"01",X"00",X"00",
		X"05",X"04",X"00",X"01",X"12",X"00",X"00",X"00",X"04",X"2C",X"00",X"00",X"72",X"42",X"99",X"00",
		X"04",X"2C",X"00",X"00",X"12",X"00",X"00",X"00",X"05",X"05",X"00",X"02",X"00",X"01",X"00",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"24",X"20",X"00",X"10",X"46",X"C0",X"00",X"0E",X"2C",X"20",X"00",
		X"00",X"00",X"09",X"00",X"02",X"05",X"06",X"02",X"0D",X"00",X"D6",X"D0",X"DA",X"D0",X"06",X"00",
		X"06",X"00",X"0D",X"00",X"02",X"03",X"06",X"00",X"0D",X"60",X"0A",X"D0",X"D6",X"00",X"D0",X"00",
		X"03",X"03",X"07",X"00",X"00",X"D6",X"00",X"0D",X"AD",X"00",X"06",X"D0",X"00",X"D0",X"00",X"00",
		X"03",X"02",X"07",X"07",X"00",X"D6",X"00",X"06",X"AD",X"00",X"DD",X"00",X"00",X"05",X"02",X"00",
		X"07",X"00",X"0D",X"D0",X"00",X"D6",X"6A",X"6D",X"00",X"00",X"0D",X"D0",X"00",X"03",X"02",X"07",
		X"07",X"DD",X"00",X"00",X"06",X"AD",X"00",X"00",X"D6",X"00",X"03",X"03",X"07",X"00",X"D0",X"00",
		X"00",X"06",X"D0",X"00",X"0D",X"AD",X"00",X"00",X"D6",X"00",X"02",X"03",X"06",X"00",X"D0",X"00",
		X"D6",X"00",X"0A",X"D0",X"0D",X"60",X"02",X"05",X"06",X"02",X"0D",X"00",X"06",X"00",X"06",X"00",
		X"DA",X"D0",X"D6",X"D0",X"0D",X"00",X"02",X"03",X"06",X"00",X"00",X"D0",X"06",X"D0",X"DA",X"00",
		X"6D",X"00",X"03",X"03",X"07",X"00",X"00",X"0D",X"00",X"0D",X"60",X"00",X"DA",X"D0",X"00",X"6D",
		X"00",X"00",X"03",X"02",X"07",X"07",X"00",X"DD",X"00",X"DA",X"60",X"00",X"6D",X"00",X"00",X"05",
		X"02",X"00",X"07",X"0D",X"D0",X"00",X"00",X"D6",X"A6",X"6D",X"00",X"0D",X"D0",X"00",X"00",X"03",
		X"02",X"07",X"07",X"6D",X"00",X"00",X"DA",X"60",X"00",X"00",X"DD",X"00",X"03",X"03",X"07",X"00",
		X"6D",X"00",X"00",X"DA",X"D0",X"00",X"0D",X"60",X"00",X"00",X"0D",X"00",X"02",X"03",X"06",X"00",
		X"6D",X"00",X"DA",X"00",X"06",X"D0",X"00",X"D0",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",
		X"6A",X"AA",X"86",X"00",X"A6",X"16",X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",
		X"61",X"61",X"6A",X"AA",X"86",X"00",X"A6",X"16",X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",
		X"A6",X"00",X"61",X"61",X"6A",X"AA",X"86",X"00",X"A6",X"16",X"A0",X"A6",X"A8",X"00",X"A6",X"16",
		X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",X"6A",X"AA",X"86",X"00",
		X"A6",X"16",X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",X"6A",X"AA",
		X"86",X"00",X"A6",X"16",X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",
		X"6A",X"AA",X"86",X"00",X"61",X"61",X"6A",X"AA",X"86",X"00",X"A6",X"16",X"A0",X"A6",X"A8",X"00",
		X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",X"6A",X"AA",X"86",X"00",X"A6",X"16",X"A0",X"A6",
		X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"61",X"61",X"6A",X"AA",X"86",X"00",X"A6",X"16",
		X"A0",X"A6",X"A8",X"00",X"A1",X"16",X"AA",X"D6",X"A6",X"00",X"59",X"6A",X"18",X"11",X"09",X"16",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"99",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"90",X"90",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"90",X"08",X"98",X"98",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"08",X"89",X"59",X"89",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"88",X"95",X"98",X"99",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"98",X"89",X"59",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"80",X"95",X"55",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"99",X"99",X"55",X"88",X"89",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"58",X"85",X"58",X"08",X"90",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"99",X"85",X"99",X"40",X"09",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"08",
		X"90",X"05",X"49",X"98",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"98",
		X"90",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"00",X"00",X"07",X"07",X"08",X"08",X"00",X"0C",
		X"01",X"0C",X"02",X"0D",X"05",X"0E",X"06",X"13",X"07",X"14",X"08",X"11",X"0B",X"12",X"08",X"15",
		X"08",X"16",X"07",X"17",X"06",X"18",X"05",X"18",X"0E",X"16",X"0F",X"16",X"10",X"14",X"5A",X"71",
		X"17",X"10",X"09",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"90",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"08",X"95",X"98",X"90",
		X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"09",X"90",X"08",X"89",X"89",X"88",X"99",X"99",X"00",
		X"00",X"00",X"09",X"90",X"00",X"99",X"99",X"88",X"95",X"90",X"90",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"08",X"99",X"98",X"09",X"59",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"88",X"95",X"55",X"80",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"55",X"88",X"89",X"80",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"80",X"00",X"58",X"85",X"58",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"85",X"99",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"90",X"05",X"49",X"98",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"09",X"00",X"00",X"90",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"98",X"00",
		X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",
		X"00",X"0D",X"0D",X"0C",X"0C",X"07",X"0D",X"08",X"0E",X"04",X"0E",X"00",X"13",X"01",X"14",X"07",
		X"11",X"0B",X"15",X"0A",X"16",X"09",X"17",X"09",X"14",X"09",X"15",X"09",X"16",X"08",X"16",X"0D",
		X"16",X"0D",X"14",X"5B",X"41",X"16",X"0D",X"08",X"0A",X"00",X"00",X"00",X"09",X"09",X"00",X"00",
		X"09",X"98",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"58",X"89",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"95",X"90",X"80",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"88",X"98",X"09",X"89",X"89",X"90",X"09",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"88",X"95",
		X"98",X"80",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"98",X"89",X"55",X"58",X"08",X"99",
		X"00",X"00",X"90",X"00",X"08",X"99",X"99",X"95",X"58",X"88",X"99",X"08",X"00",X"99",X"00",X"00",
		X"09",X"00",X"00",X"05",X"88",X"55",X"80",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",
		X"98",X"59",X"99",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"09",X"80",X"00",X"59",X"99",X"80",
		X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"08",X"89",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"89",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"07",X"11",X"08",X"0E",X"08",X"12",X"06",X"13",X"04",X"10",X"03",X"15",X"02",X"15",X"00",
		X"12",X"06",X"13",X"05",X"14",X"04",X"15",X"0A",X"16",X"08",X"10",X"10",X"10",X"5C",X"33",X"17",
		X"0F",X"09",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"90",X"89",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"08",X"95",
		X"90",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"90",X"08",X"09",X"59",X"80",X"00",
		X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"88",X"95",X"98",X"99",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"89",X"98",X"89",X"89",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"95",X"55",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"99",X"99",X"55",X"88",X"89",X"00",X"90",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"58",
		X"85",X"58",X"00",X"09",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"99",X"85",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",X"05",X"99",X"98",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"88",X"80",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"09",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"0D",X"0E",X"07",X"0C",X"08",X"13",X"04",X"11",X"03",X"12",X"00",X"12",X"07",
		X"11",X"0C",X"15",X"08",X"16",X"06",X"17",X"03",X"14",X"0D",X"15",X"0D",X"16",X"0D",X"17",X"0C",
		X"11",X"11",X"11",X"5D",X"43",X"17",X"11",X"09",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"49",X"90",X"09",X"00",X"00",X"00",X"00",X"00",
		X"98",X"99",X"00",X"89",X"55",X"99",X"49",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"85",
		X"58",X"85",X"59",X"80",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"55",X"88",X"50",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"09",X"98",X"95",X"98",X"58",X"99",X"99",X"90",X"00",
		X"00",X"00",X"00",X"09",X"99",X"89",X"59",X"08",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"08",X"95",X"98",X"89",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"89",
		X"88",X"90",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"90",X"98",X"89",X"90",X"00",
		X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"09",X"90",X"00",X"00",X"09",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"89",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"12",X"0E",X"11",X"0D",X"16",X"0D",X"15",X"06",X"17",X"09",X"16",X"09",
		X"15",X"07",X"14",X"05",X"0E",X"04",X"10",X"03",X"11",X"02",X"12",X"01",X"13",X"00",X"14",X"09",
		X"0A",X"08",X"08",X"07",X"07",X"06",X"06",X"5E",X"57",X"17",X"11",X"09",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"90",X"09",X"80",X"00",X"90",
		X"09",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"49",X"90",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"89",X"55",X"99",X"49",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"85",X"58",X"85",X"59",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"89",X"55",X"88",X"85",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"95",X"98",X"58",
		X"99",X"99",X"99",X"00",X"00",X"00",X"09",X"00",X"89",X"89",X"59",X"88",X"90",X"00",X"00",X"00",
		X"98",X"00",X"00",X"90",X"00",X"08",X"98",X"90",X"89",X"99",X"99",X"99",X"80",X"00",X"00",X"09",
		X"00",X"00",X"09",X"59",X"88",X"98",X"00",X"00",X"00",X"09",X"00",X"00",X"90",X"00",X"00",X"90",
		X"98",X"89",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"90",X"00",X"89",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"98",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"12",X"0B",X"11",X"07",X"16",X"09",X"15",X"09",
		X"14",X"09",X"12",X"09",X"11",X"04",X"15",X"03",X"17",X"02",X"14",X"01",X"15",X"00",X"0D",X"05",
		X"0E",X"07",X"0F",X"0D",X"0D",X"0C",X"0C",X"0B",X"0B",X"0A",X"0A",X"5F",X"6B",X"17",X"11",X"09",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"98",X"00",
		X"09",X"99",X"00",X"08",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"08",X"95",X"59",X"99",X"80",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"98",X"55",X"88",X"55",X"98",X"89",X"90",X"00",X"00",
		X"09",X"09",X"98",X"00",X"88",X"95",X"58",X"88",X"50",X"00",X"00",X"00",X"00",X"90",X"00",X"99",
		X"98",X"89",X"59",X"85",X"89",X"98",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"90",X"98",X"98",
		X"89",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"59",X"88",X"99",X"99",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"95",X"90",X"89",X"90",X"00",X"90",X"09",X"00",X"00",
		X"00",X"00",X"00",X"09",X"09",X"88",X"89",X"99",X"80",X"09",X"00",X"98",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"08",X"99",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"00",X"00",X"00",X"11",X"11",X"10",X"10",X"0A",
		X"10",X"06",X"17",X"07",X"17",X"04",X"16",X"03",X"12",X"02",X"13",X"00",X"13",X"08",X"14",X"08",
		X"15",X"07",X"17",X"09",X"14",X"11",X"15",X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"13",X"60",
		X"7F",X"17",X"11",X"09",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"80",X"08",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"99",X"90",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",
		X"55",X"99",X"98",X"00",X"90",X"00",X"00",X"00",X"08",X"98",X"98",X"05",X"58",X"85",X"59",X"88",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"89",X"55",X"88",X"85",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"98",X"98",X"98",X"58",X"99",X"99",X"98",X"00",X"00",X"00",X"09",X"00",
		X"89",X"89",X"59",X"88",X"90",X"00",X"00",X"00",X"98",X"00",X"00",X"90",X"00",X"00",X"95",X"98",
		X"89",X"98",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"09",X"59",X"88",X"98",X"09",X"80",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"90",X"90",X"89",X"99",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"90",X"00",X"89",X"90",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"00",X"00",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"10",X"0B",X"0F",X"0B",X"13",X"0C",X"16",X"0C",X"16",X"05",X"15",X"09",X"11",X"04",X"15",X"03",
		X"17",X"02",X"0F",X"01",X"10",X"00",X"10",X"05",X"11",X"07",X"11",X"0D",X"11",X"0C",X"0C",X"0B",
		X"0B",X"0A",X"0A",X"08",X"08",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",
		X"90",X"00",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"90",X"09",X"00",X"09",X"09",
		X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"90",X"09",X"00",X"90",X"00",X"90",X"00",X"90",X"00",
		X"00",X"09",X"00",X"09",X"00",X"90",X"90",X"00",X"90",X"09",X"00",X"09",X"00",X"00",X"99",X"00",
		X"90",X"90",X"90",X"00",X"90",X"09",X"09",X"00",X"90",X"00",X"09",X"90",X"90",X"90",X"50",X"09",
		X"00",X"90",X"00",X"90",X"90",X"09",X"00",X"99",X"98",X"95",X"89",X"98",X"88",X"50",X"09",X"00",
		X"90",X"00",X"98",X"89",X"99",X"58",X"89",X"98",X"85",X"88",X"99",X"99",X"00",X"00",X"89",X"99",
		X"99",X"85",X"99",X"99",X"85",X"99",X"94",X"90",X"00",X"00",X"08",X"88",X"88",X"80",X"88",X"88",
		X"00",X"08",X"80",X"00",X"00",X"08",X"08",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"09",X"09",X"00",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"90",
		X"90",X"90",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"90",X"00",X"90",X"90",X"09",X"00",X"00",
		X"90",X"00",X"00",X"09",X"00",X"09",X"00",X"90",X"90",X"00",X"90",X"09",X"00",X"00",X"90",X"00",
		X"99",X"00",X"90",X"90",X"90",X"00",X"90",X"09",X"00",X"90",X"90",X"00",X"09",X"90",X"90",X"90",
		X"50",X"09",X"00",X"90",X"00",X"90",X"90",X"90",X"00",X"99",X"98",X"95",X"89",X"98",X"88",X"50",
		X"09",X"00",X"90",X"09",X"98",X"89",X"99",X"58",X"89",X"98",X"85",X"88",X"99",X"99",X"00",X"00",
		X"89",X"99",X"99",X"85",X"99",X"99",X"85",X"99",X"99",X"90",X"00",X"00",X"08",X"89",X"98",X"80",
		X"89",X"88",X"00",X"08",X"80",X"00",X"00",X"61",X"F8",X"01",X"0D",X"00",X"6A",X"AA",X"60",X"00",
		X"0A",X"A1",X"11",X"AA",X"00",X"6A",X"11",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"60",X"A1",
		X"AA",X"AA",X"AA",X"60",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",X"AA",X"60",X"06",X"AA",
		X"AA",X"A6",X"00",X"00",X"66",X"66",X"60",X"00",X"02",X"06",X"01",X"07",X"00",X"08",X"00",X"08",
		X"00",X"08",X"00",X"08",X"00",X"08",X"01",X"07",X"02",X"06",X"62",X"4A",X"02",X"0E",X"00",X"6A",
		X"AA",X"A6",X"00",X"00",X"0A",X"A1",X"11",X"1A",X"A0",X"00",X"6A",X"11",X"AA",X"AA",X"A6",X"00",
		X"A1",X"1A",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",
		X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"AA",X"AA",X"A6",X"00",X"06",X"AA",
		X"AA",X"AA",X"60",X"00",X"00",X"66",X"66",X"66",X"00",X"00",X"02",X"07",X"01",X"08",X"00",X"09",
		X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"00",X"09",X"01",X"08",X"02",X"07",X"62",X"A4",
		X"02",X"0F",X"00",X"06",X"AA",X"A6",X"00",X"00",X"00",X"AA",X"11",X"1A",X"A0",X"00",X"0A",X"11",
		X"1A",X"AA",X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"60",X"A1",X"1A",X"AA",X"AA",X"AA",X"60",
		X"A1",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"60",X"0A",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"6A",X"AA",X"AA",X"60",X"00",X"00",X"00",
		X"66",X"60",X"00",X"00",X"03",X"07",X"02",X"08",X"01",X"09",X"00",X"0A",X"00",X"0A",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"01",X"09",X"02",X"08",X"04",X"06",X"63",X"12",X"03",X"08",X"00",X"06",
		X"AA",X"AA",X"60",X"00",X"00",X"00",X"AA",X"11",X"11",X"AA",X"00",X"00",X"0A",X"11",X"1A",X"AA",
		X"AA",X"A0",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"A6",
		X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"06",X"AA",X"AA",
		X"AA",X"AA",X"60",X"00",X"00",X"6A",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"06",X"66",X"66",X"60",
		X"00",X"00",X"03",X"08",X"02",X"09",X"01",X"0A",X"00",X"0B",X"00",X"0B",X"00",X"0B",X"00",X"0B",
		X"00",X"0B",X"00",X"0B",X"01",X"0A",X"02",X"09",X"03",X"08",X"63",X"89",X"03",X"09",X"00",X"00",
		X"6A",X"AA",X"60",X"00",X"00",X"00",X"0A",X"A1",X"11",X"AA",X"00",X"00",X"00",X"A1",X"11",X"AA",
		X"AA",X"A0",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",
		X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"A6",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"06",X"AA",X"AA",X"A6",
		X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"04",X"08",X"03",X"09",X"02",X"0A",X"01",
		X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"01",X"0B",X"02",X"0A",X"03",
		X"09",X"05",X"07",X"64",X"17",X"0C",X"0A",X"00",X"00",X"6A",X"AA",X"A6",X"00",X"00",X"00",X"00",
		X"0A",X"A1",X"11",X"1A",X"A0",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"00",X"00",X"0A",
		X"11",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",
		X"6A",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"06",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",
		X"00",X"06",X"66",X"66",X"00",X"00",X"00",X"04",X"09",X"03",X"0A",X"02",X"0B",X"01",X"0C",X"00",
		X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"00",X"0D",X"01",X"0C",X"02",X"0B",X"03",
		X"0A",X"05",X"09",X"64",X"AF",X"0C",X"0B",X"00",X"00",X"6A",X"AA",X"AA",X"60",X"00",X"00",X"00",
		X"0A",X"A1",X"11",X"1A",X"AA",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",
		X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",
		X"06",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"00",X"00",X"00",X"04",
		X"0A",X"03",X"0B",X"02",X"0C",X"01",X"0D",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
		X"0E",X"00",X"0E",X"00",X"0E",X"01",X"0D",X"02",X"0C",X"03",X"0B",X"05",X"09",X"65",X"61",X"0D",
		X"14",X"00",X"00",X"6A",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",X"0A",X"A1",X"11",X"11",X"AA",
		X"A0",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"11",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"1A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",
		X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"00",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",
		X"06",X"6A",X"AA",X"AA",X"A6",X"60",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"60",X"00",X"00",
		X"00",X"04",X"0B",X"03",X"0C",X"02",X"0D",X"01",X"0E",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"01",X"0E",X"02",X"0D",X"03",X"0C",X"05",
		X"0A",X"66",X"1E",X"0D",X"15",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"0A",
		X"A1",X"11",X"11",X"1A",X"AA",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"0A",X"11",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"6A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"60",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"1A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"60",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"60",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"06",X"6A",X"AA",
		X"AA",X"AA",X"66",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"00",X"00",X"00",X"04",X"0C",
		X"03",X"0D",X"02",X"0E",X"01",X"0F",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",
		X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"01",X"0F",X"02",X"0E",X"03",X"0D",X"05",X"0B",
		X"66",X"F8",X"0E",X"16",X"00",X"00",X"06",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"11",X"11",X"1A",X"AA",X"00",X"00",X"00",X"00",X"DA",X"11",X"1A",X"AA",X"AA",X"AA",X"AD",
		X"00",X"00",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"11",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",
		X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"66",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",
		X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"D6",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"6D",X"00",X"00",X"00",X"00",X"66",X"AA",X"AA",X"AA",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"05",X"0C",X"04",X"0D",X"02",X"0F",X"02",X"0F",
		X"01",X"10",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",
		X"00",X"11",X"01",X"10",X"02",X"0F",X"02",X"0F",X"04",X"0D",X"06",X"0B",X"67",X"DE",X"0E",X"17",
		X"00",X"00",X"06",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",X"00",X"AA",X"11",X"11",X"1A",
		X"AA",X"A0",X"00",X"00",X"00",X"DA",X"11",X"1A",X"AA",X"AA",X"AA",X"AA",X"D0",X"00",X"00",X"A1",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"1A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",
		X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"60",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"60",X"06",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",
		X"00",X"D6",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"D0",X"00",X"00",X"00",X"66",X"AA",X"AA",X"AA",
		X"A6",X"60",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"05",X"0D",
		X"04",X"0E",X"02",X"10",X"02",X"10",X"01",X"11",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",
		X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"01",X"11",X"02",X"10",X"02",X"10",
		X"04",X"0E",X"06",X"0C",X"68",X"E4",X"0F",X"10",X"00",X"00",X"06",X"AA",X"AA",X"AA",X"AA",X"60",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"11",X"11",X"11",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0A",
		X"11",X"1A",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"6A",
		X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",
		X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"00",X"06",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"00",X"00",X"00",X"06",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",
		X"66",X"AA",X"AA",X"AA",X"AA",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"66",
		X"00",X"00",X"00",X"00",X"05",X"0E",X"04",X"0F",X"03",X"10",X"02",X"11",X"01",X"12",X"00",X"13",
		X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",
		X"01",X"13",X"01",X"12",X"02",X"11",X"03",X"10",X"04",X"0F",X"06",X"0D",X"69",X"F7",X"0F",X"11",
		X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"A1",X"11",
		X"11",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"00",X"00",X"01",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"A1",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"1A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"60",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",
		X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"0A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",
		X"00",X"00",X"00",X"06",X"6A",X"AA",X"AA",X"AA",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",
		X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"06",X"0E",X"05",X"0F",X"04",X"10",X"03",X"11",X"02",
		X"12",X"01",X"13",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"00",
		X"14",X"00",X"14",X"00",X"14",X"01",X"13",X"02",X"12",X"03",X"11",X"04",X"10",X"05",X"0F",X"07",
		X"0D",X"6B",X"2D",X"08",X"12",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"A1",X"11",X"11",X"1A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"A1",
		X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"00",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",
		X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"6A",X"1A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",
		X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",
		X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"06",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"00",X"00",X"00",X"00",X"00",X"06",X"6A",X"AA",X"AA",X"AA",X"A6",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"06",X"0F",X"05",
		X"10",X"04",X"11",X"03",X"12",X"02",X"13",X"01",X"14",X"00",X"15",X"00",X"15",X"00",X"15",X"00",
		X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"01",X"14",X"02",
		X"13",X"03",X"12",X"04",X"11",X"05",X"10",X"07",X"0E",X"6C",X"71",X"08",X"13",X"00",X"00",X"00",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",X"00",X"0A",X"A1",X"11",X"11",X"11",
		X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"A1",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",
		X"00",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"A1",X"1A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"60",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"60",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",
		X"00",X"00",X"06",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",X"6A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"00",X"00",X"06",X"6A",X"AA",X"AA",X"AA",
		X"AA",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"66",X"66",X"66",X"00",X"00",X"00",
		X"00",X"06",X"10",X"05",X"11",X"04",X"12",X"03",X"13",X"02",X"14",X"01",X"15",X"00",X"16",X"00",
		X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",
		X"16",X"00",X"16",X"01",X"15",X"02",X"14",X"03",X"13",X"04",X"12",X"05",X"11",X"07",X"0F",X"6D",
		X"DB",X"09",X"1C",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"A1",X"11",X"11",X"11",X"1A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"A1",
		X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0A",X"11",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"A1",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"00",X"00",X"0A",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",
		X"00",X"6A",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"1A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"A1",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A6",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"06",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"60",X"00",X"00",X"00",X"00",X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",
		X"00",X"00",X"00",X"06",X"6A",X"AA",X"AA",X"AA",X"AA",X"A6",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"66",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"00",X"06",X"11",X"05",X"12",X"04",
		X"13",X"03",X"14",X"02",X"15",X"01",X"16",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",
		X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"01",
		X"16",X"02",X"15",X"03",X"14",X"04",X"13",X"05",X"12",X"07",X"10",X"02",X"0E",X"00",X"01",X"11",
		X"10",X"00",X"00",X"01",X"11",X"AA",X"AA",X"A0",X"00",X"01",X"AA",X"AA",X"AA",X"A0",X"00",X"1A",
		X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"AA",X"AA",
		X"AA",X"A0",X"00",X"00",X"0A",X"AA",X"A0",X"00",X"00",X"02",X"0F",X"00",X"00",X"11",X"10",X"00",
		X"00",X"00",X"11",X"1A",X"AA",X"A0",X"00",X"01",X"1A",X"AA",X"AA",X"AA",X"00",X"01",X"AA",X"AA",
		X"AA",X"AA",X"00",X"1A",X"11",X"1A",X"11",X"1A",X"A0",X"1A",X"19",X"81",X"19",X"81",X"A0",X"1A",
		X"11",X"1A",X"11",X"1A",X"A0",X"0A",X"AA",X"A6",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",
		X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"03",X"08",X"00",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"00",X"00",X"01",X"1A",X"AA",
		X"AA",X"AA",X"A0",X"00",X"01",X"A1",X"AA",X"AA",X"1A",X"A0",X"00",X"11",X"11",X"11",X"A1",X"11",
		X"1A",X"00",X"1A",X"18",X"91",X"A1",X"98",X"1A",X"00",X"1A",X"11",X"11",X"A1",X"11",X"1A",X"00",
		X"1A",X"AA",X"A6",X"A6",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"00",X"00",X"00",X"03",X"09",X"00",X"00",X"11",X"11",X"A0",X"00",X"00",X"00",X"11",X"1A",X"AA",
		X"AA",X"A0",X"00",X"01",X"1A",X"AA",X"AA",X"AA",X"AA",X"00",X"01",X"AA",X"1A",X"AA",X"1A",X"AA",
		X"00",X"11",X"11",X"11",X"A1",X"11",X"1A",X"A0",X"1A",X"18",X"91",X"A1",X"98",X"1A",X"A0",X"1A",
		X"11",X"11",X"A1",X"11",X"1A",X"A0",X"1A",X"AA",X"A6",X"A6",X"AA",X"AA",X"A0",X"1A",X"AA",X"AA",
		X"6A",X"AA",X"AA",X"A0",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"00",
		X"0C",X"0A",X"00",X"00",X"11",X"11",X"1A",X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"AA",
		X"00",X"00",X"01",X"1A",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"01",X"AA",X"1A",X"AA",X"A1",X"AA",
		X"A0",X"00",X"11",X"11",X"11",X"A6",X"11",X"11",X"AA",X"00",X"1A",X"18",X"91",X"AA",X"19",X"81",
		X"AA",X"00",X"16",X"11",X"11",X"AA",X"11",X"11",X"6A",X"00",X"1A",X"AA",X"A6",X"AA",X"6A",X"AA",
		X"AA",X"00",X"1A",X"AA",X"AA",X"66",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"00",
		X"00",X"00",X"0C",X"0B",X"00",X"00",X"11",X"11",X"11",X"A0",X"00",X"00",X"00",X"11",X"1A",X"AA",
		X"AA",X"AA",X"A0",X"00",X"01",X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"01",X"1A",X"11",X"AA",
		X"61",X"1A",X"AA",X"00",X"11",X"A1",X"11",X"1A",X"11",X"11",X"AA",X"A0",X"11",X"A1",X"89",X"1A",
		X"19",X"81",X"AA",X"A0",X"1A",X"61",X"11",X"1A",X"11",X"11",X"6A",X"A0",X"1A",X"AA",X"AA",X"61",
		X"A6",X"AA",X"AA",X"A0",X"1A",X"A6",X"6A",X"A6",X"6A",X"A6",X"AA",X"A0",X"1A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"0A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"0D",X"14",X"00",X"00",
		X"01",X"11",X"11",X"A0",X"00",X"00",X"00",X"00",X"01",X"11",X"AA",X"AA",X"A1",X"A0",X"00",X"00",
		X"00",X"11",X"AA",X"AA",X"AA",X"AA",X"1A",X"00",X"00",X"01",X"1A",X"11",X"1A",X"61",X"11",X"1A",
		X"A0",X"00",X"01",X"A1",X"89",X"1A",X"A1",X"98",X"1A",X"A0",X"00",X"11",X"61",X"11",X"1A",X"A1",
		X"11",X"16",X"AA",X"00",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"1A",X"6A",X"AA",
		X"61",X"A6",X"AA",X"A6",X"AA",X"00",X"18",X"AA",X"6A",X"A6",X"6A",X"A6",X"AA",X"8A",X"00",X"1A",
		X"0A",X"AA",X"AA",X"AA",X"AA",X"A0",X"AA",X"00",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"0A",X"AA",
		X"00",X"0A",X"A6",X"06",X"AA",X"AA",X"60",X"6A",X"A0",X"00",X"0A",X"AA",X"66",X"88",X"88",X"66",
		X"AA",X"A0",X"00",X"00",X"AA",X"A6",X"66",X"66",X"6A",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"66",
		X"66",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"0D",X"15",
		X"00",X"00",X"01",X"11",X"11",X"AA",X"00",X"00",X"00",X"00",X"01",X"11",X"AA",X"AA",X"A1",X"1A",
		X"00",X"00",X"00",X"11",X"AA",X"AA",X"AA",X"AA",X"A1",X"A0",X"00",X"01",X"1A",X"61",X"11",X"61",
		X"11",X"6A",X"AA",X"00",X"01",X"A6",X"18",X"91",X"A1",X"98",X"16",X"AA",X"00",X"11",X"A6",X"11",
		X"11",X"A1",X"11",X"16",X"AA",X"A0",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"1A",
		X"66",X"AA",X"61",X"1A",X"6A",X"A6",X"6A",X"A0",X"18",X"AA",X"66",X"A6",X"66",X"A6",X"6A",X"A8",
		X"A0",X"1A",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"0A",X"A0",X"A6",X"A0",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"A6",X"A0",X"AA",X"A6",X"06",X"AA",X"AA",X"A6",X"06",X"AA",X"A0",X"0A",X"AA",X"66",X"08",
		X"88",X"06",X"6A",X"AA",X"00",X"0A",X"AA",X"A6",X"66",X"16",X"66",X"AA",X"AA",X"00",X"00",X"AA",
		X"AA",X"66",X"66",X"6A",X"AA",X"A0",X"00",X"00",X"0A",X"AA",X"A6",X"66",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"0E",X"16",X"00",X"00",X"01",X"11",X"11",
		X"1A",X"A0",X"00",X"00",X"00",X"00",X"01",X"11",X"1A",X"AA",X"AA",X"11",X"A0",X"00",X"00",X"00",
		X"11",X"AA",X"AA",X"AA",X"AA",X"AA",X"1A",X"00",X"00",X"01",X"1A",X"61",X"11",X"A6",X"11",X"16",
		X"AA",X"A0",X"00",X"01",X"A6",X"18",X"91",X"AA",X"19",X"81",X"6A",X"A0",X"00",X"11",X"A6",X"11",
		X"11",X"AA",X"11",X"11",X"6A",X"AA",X"00",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"00",X"1A",X"66",X"AA",X"A6",X"11",X"6A",X"AA",X"66",X"AA",X"00",X"18",X"AA",X"66",X"6A",X"66",
		X"A6",X"66",X"AA",X"8A",X"00",X"1A",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"00",X"16",
		X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"6A",X"00",X"AA",X"AA",X"86",X"AA",X"AA",X"AA",X"68",
		X"AA",X"AA",X"00",X"AA",X"A6",X"A6",X"88",X"88",X"88",X"6A",X"6A",X"AA",X"00",X"0A",X"AA",X"6A",
		X"A6",X"88",X"6A",X"A6",X"AA",X"A0",X"00",X"0A",X"AA",X"A6",X"AA",X"11",X"AA",X"6A",X"AA",X"A0",
		X"00",X"00",X"AA",X"AA",X"66",X"66",X"66",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"A6",X"66",
		X"6A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"0E",
		X"17",X"00",X"00",X"00",X"11",X"11",X"1A",X"A0",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",
		X"AA",X"11",X"A0",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"AA",X"AA",X"1A",X"A0",X"00",X"00",
		X"11",X"AA",X"11",X"6A",X"61",X"1A",X"A1",X"A0",X"00",X"01",X"1A",X"A1",X"11",X"16",X"11",X"11",
		X"AA",X"AA",X"00",X"01",X"AA",X"61",X"89",X"1A",X"19",X"81",X"6A",X"AA",X"00",X"11",X"A6",X"61",
		X"11",X"1A",X"11",X"11",X"66",X"AA",X"A0",X"1A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A0",X"1A",X"66",X"AA",X"A6",X"11",X"A6",X"AA",X"A6",X"6A",X"A0",X"18",X"AA",X"66",X"6A",X"66",
		X"6A",X"66",X"6A",X"A8",X"A0",X"1A",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"A0",X"A6",
		X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"A6",X"A0",X"AA",X"AA",X"06",X"AA",X"AA",X"AA",X"A6",
		X"0A",X"AA",X"A0",X"0A",X"A6",X"A6",X"88",X"88",X"88",X"86",X"A6",X"AA",X"00",X"0A",X"AA",X"6A",
		X"66",X"88",X"86",X"6A",X"6A",X"AA",X"00",X"00",X"AA",X"A6",X"AA",X"11",X"1A",X"A6",X"AA",X"A0",
		X"00",X"00",X"AA",X"AA",X"66",X"66",X"66",X"6A",X"AA",X"A0",X"00",X"00",X"00",X"AA",X"AA",X"60",
		X"6A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"0F",
		X"10",X"00",X"00",X"00",X"11",X"11",X"11",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",
		X"AA",X"AA",X"A1",X"1A",X"00",X"00",X"00",X"00",X"01",X"1A",X"6A",X"AA",X"AA",X"A6",X"A1",X"A0",
		X"00",X"00",X"00",X"11",X"AA",X"11",X"AA",X"AA",X"11",X"AA",X"1A",X"00",X"00",X"01",X"1A",X"A1",
		X"A1",X"1A",X"61",X"1A",X"1A",X"AA",X"A0",X"00",X"01",X"AA",X"61",X"89",X"1A",X"A1",X"98",X"16",
		X"AA",X"A0",X"00",X"11",X"A6",X"61",X"11",X"1A",X"A1",X"11",X"16",X"6A",X"AA",X"00",X"1A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"11",X"66",X"A1",X"A6",X"61",X"16",X"6A",
		X"1A",X"66",X"1A",X"00",X"18",X"AA",X"66",X"6A",X"A6",X"6A",X"A6",X"66",X"AA",X"8A",X"00",X"1A",
		X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"00",X"16",X"A8",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"8A",X"6A",X"00",X"AA",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"A8",X"AA",X"AA",X"00",
		X"AA",X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"AA",X"00",X"0A",X"AA",X"6A",X"68",X"88",
		X"88",X"86",X"A6",X"AA",X"A0",X"00",X"0A",X"AA",X"A6",X"AA",X"88",X"88",X"AA",X"6A",X"AA",X"A0",
		X"00",X"00",X"AA",X"AA",X"6A",X"A1",X"1A",X"A6",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"A6",
		X"66",X"66",X"6A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"60",X"06",X"AA",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"0F",X"11",X"00",
		X"00",X"00",X"11",X"11",X"11",X"1A",X"A0",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",
		X"AA",X"11",X"A0",X"00",X"00",X"00",X"01",X"1A",X"A6",X"AA",X"AA",X"A6",X"AA",X"1A",X"00",X"00",
		X"00",X"11",X"AA",X"A1",X"1A",X"AA",X"11",X"AA",X"A1",X"A0",X"00",X"01",X"1A",X"A6",X"1A",X"11",
		X"61",X"1A",X"16",X"AA",X"AA",X"00",X"01",X"A6",X"61",X"18",X"91",X"A1",X"98",X"11",X"66",X"AA",
		X"00",X"11",X"AA",X"AA",X"11",X"11",X"A1",X"11",X"AA",X"AA",X"AA",X"A0",X"1A",X"AA",X"AA",X"AA",
		X"A6",X"A6",X"AA",X"AA",X"AA",X"AA",X"A0",X"11",X"66",X"A1",X"A6",X"61",X"1A",X"66",X"A1",X"A6",
		X"61",X"A0",X"18",X"AA",X"66",X"6A",X"A6",X"66",X"AA",X"66",X"6A",X"A8",X"A0",X"1A",X"8A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"A0",X"16",X"A8",X"AA",X"AA",X"AA",X"6A",X"AA",X"AA",
		X"A8",X"A6",X"A0",X"1A",X"AA",X"8A",X"AA",X"AA",X"AA",X"AA",X"AA",X"8A",X"AA",X"A0",X"AA",X"AA",
		X"A8",X"6A",X"AA",X"AA",X"AA",X"68",X"AA",X"AA",X"A0",X"AA",X"AA",X"AA",X"68",X"88",X"88",X"88",
		X"6A",X"AA",X"AA",X"A0",X"0A",X"AA",X"6A",X"A6",X"A1",X"11",X"A6",X"AA",X"6A",X"AA",X"00",X"0A",
		X"AA",X"A6",X"AA",X"68",X"88",X"6A",X"A6",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"6A",X"AA",X"AA",
		X"AA",X"6A",X"AA",X"A0",X"00",X"00",X"0A",X"AA",X"A6",X"AA",X"11",X"A6",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"AA",X"AA",X"66",X"66",X"6A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"A0",X"00",X"00",X"00",X"08",X"12",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"1A",X"AA",X"AA",X"AA",X"A1",X"1A",X"00",X"00",X"00",
		X"00",X"01",X"1A",X"AA",X"6A",X"AA",X"A6",X"AA",X"A1",X"A0",X"00",X"00",X"00",X"11",X"AA",X"A1",
		X"1A",X"AA",X"A1",X"1A",X"AA",X"1A",X"00",X"00",X"01",X"1A",X"A6",X"1A",X"11",X"A6",X"11",X"A1",
		X"6A",X"AA",X"A0",X"00",X"01",X"A6",X"61",X"10",X"91",X"AA",X"19",X"01",X"16",X"6A",X"A0",X"00",
		X"11",X"AA",X"AA",X"A1",X"11",X"AA",X"11",X"1A",X"AA",X"AA",X"AA",X"00",X"11",X"66",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"1A",X"00",X"16",X"AA",X"6A",X"1A",X"66",X"11",X"66",X"A1",
		X"A6",X"AA",X"6A",X"00",X"1A",X"8A",X"A6",X"66",X"AA",X"66",X"AA",X"66",X"6A",X"A8",X"AA",X"00",
		X"1A",X"68",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"86",X"AA",X"00",X"16",X"A9",X"06",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"60",X"9A",X"6A",X"00",X"1A",X"AA",X"90",X"06",X"AA",X"AA",X"AA",X"60",
		X"09",X"AA",X"AA",X"00",X"1A",X"AA",X"A9",X"10",X"66",X"66",X"66",X"01",X"9A",X"AA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"91",X"11",X"11",X"11",X"19",X"AA",X"AA",X"AA",X"00",X"AA",X"AA",X"6A",X"A9",
		X"A1",X"11",X"1A",X"9A",X"A6",X"AA",X"AA",X"00",X"0A",X"AA",X"A6",X"AA",X"99",X"99",X"99",X"AA",
		X"6A",X"AA",X"A0",X"00",X"0A",X"AA",X"AA",X"6A",X"A6",X"99",X"6A",X"A6",X"AA",X"AA",X"A0",X"00",
		X"00",X"AA",X"AA",X"66",X"AA",X"AA",X"AA",X"66",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"A6",
		X"66",X"11",X"66",X"6A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"66",X"66",X"66",X"AA",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",X"CB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"CB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"00",X"00",X"A6",X"35",X"80",X"02",X"C6",X"03",X"3D",X"E7",
		X"3C",X"86",X"6B",X"A0",X"3C",X"33",X"86",X"EF",X"39",X"39",X"A6",X"34",X"C6",X"03",X"3D",X"E7",
		X"3C",X"86",X"8C",X"A0",X"3C",X"A7",X"38",X"39",X"34",X"01",X"1A",X"50",X"EC",X"35",X"88",X"04",
		X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"39",X"FD",X"CA",X"02",X"EC",X"37",X"FD",X"CA",X"04",X"86",
		X"1E",X"E6",X"24",X"26",X"02",X"86",X"0E",X"B7",X"CA",X"00",X"35",X"81",X"EC",X"30",X"1E",X"89",
		X"ED",X"30",X"EC",X"31",X"1E",X"89",X"ED",X"31",X"EC",X"32",X"1E",X"89",X"ED",X"32",X"20",X"12",
		X"EC",X"32",X"1E",X"89",X"ED",X"32",X"EC",X"31",X"1E",X"89",X"ED",X"31",X"EC",X"30",X"1E",X"89",
		X"ED",X"30",X"EC",X"30",X"FD",X"99",X"FC",X"EC",X"32",X"FD",X"99",X"FF",X"39",X"BD",X"EF",X"6D",
		X"CC",X"12",X"00",X"5A",X"26",X"FD",X"4A",X"26",X"FA",X"39",X"00",X"00",X"00",X"01",X"00",X"11",
		X"01",X"11",X"09",X"91",X"09",X"11",X"09",X"99",X"00",X"08",X"08",X"88",X"08",X"00",X"00",X"98",
		X"00",X"88",X"00",X"99",X"00",X"09",X"00",X"90",X"10",X"00",X"11",X"00",X"11",X"10",X"11",X"11",
		X"11",X"19",X"11",X"18",X"11",X"88",X"18",X"88",X"11",X"99",X"19",X"00",X"19",X"99",X"19",X"88",
		X"19",X"89",X"19",X"98",X"11",X"89",X"89",X"99",X"88",X"99",X"88",X"09",X"88",X"00",X"80",X"00",
		X"80",X"01",X"80",X"99",X"88",X"80",X"88",X"88",X"88",X"89",X"88",X"11",X"88",X"81",X"81",X"11",
		X"88",X"91",X"89",X"91",X"80",X"11",X"99",X"91",X"99",X"99",X"91",X"11",X"99",X"00",X"90",X"00",
		X"99",X"90",X"99",X"11",X"98",X"91",X"99",X"88",X"99",X"98",X"99",X"10",X"91",X"10",X"07",X"00",
		X"03",X"01",X"05",X"02",X"05",X"03",X"0B",X"12",X"05",X"03",X"04",X"02",X"04",X"01",X"05",X"00",
		X"05",X"00",X"02",X"0F",X"02",X"10",X"03",X"11",X"01",X"12",X"01",X"28",X"01",X"29",X"01",X"26",
		X"01",X"25",X"01",X"09",X"05",X"00",X"01",X"0F",X"01",X"10",X"02",X"11",X"0B",X"12",X"02",X"11",
		X"02",X"10",X"02",X"0F",X"05",X"00",X"01",X"01",X"02",X"02",X"02",X"03",X"29",X"12",X"01",X"03",
		X"01",X"02",X"01",X"01",X"01",X"00",X"01",X"0F",X"01",X"10",X"01",X"11",X"07",X"12",X"01",X"28",
		X"03",X"26",X"01",X"08",X"01",X"07",X"03",X"00",X"01",X"10",X"01",X"11",X"17",X"12",X"01",X"11",
		X"01",X"10",X"02",X"00",X"06",X"12",X"01",X"13",X"02",X"14",X"04",X"15",X"05",X"16",X"09",X"12",
		X"09",X"16",X"04",X"15",X"02",X"14",X"07",X"12",X"01",X"11",X"04",X"12",X"01",X"30",X"01",X"34",
		X"01",X"2E",X"02",X"2F",X"02",X"06",X"02",X"0A",X"01",X"0B",X"03",X"00",X"01",X"10",X"0A",X"12",
		X"01",X"03",X"01",X"05",X"01",X"04",X"03",X"0C",X"01",X"06",X"03",X"2F",X"02",X"2E",X"01",X"30",
		X"06",X"12",X"01",X"10",X"01",X"10",X"05",X"12",X"01",X"2E",X"01",X"2F",X"02",X"1E",X"01",X"1F",
		X"01",X"20",X"01",X"21",X"04",X"22",X"01",X"23",X"09",X"12",X"01",X"2D",X"06",X"22",X"01",X"21",
		X"01",X"20",X"02",X"1E",X"02",X"2F",X"01",X"2E",X"01",X"30",X"07",X"12",X"05",X"12",X"01",X"19",
		X"03",X"2F",X"01",X"31",X"05",X"32",X"01",X"31",X"01",X"18",X"01",X"11",X"08",X"12",X"01",X"03",
		X"01",X"01",X"03",X"00",X"04",X"32",X"01",X"31",X"05",X"2F",X"01",X"19",X"07",X"12",X"01",X"00",
		X"01",X"0F",X"05",X"12",X"01",X"30",X"01",X"34",X"04",X"2E",X"02",X"04",X"01",X"05",X"01",X"03",
		X"0C",X"12",X"01",X"34",X"01",X"04",X"03",X"06",X"03",X"2F",X"01",X"2E",X"01",X"34",X"01",X"30",
		X"07",X"12",X"01",X"11",X"01",X"0F",X"01",X"00",X"01",X"02",X"05",X"12",X"01",X"13",X"05",X"17",
		X"02",X"13",X"09",X"12",X"01",X"03",X"01",X"01",X"03",X"00",X"01",X"22",X"01",X"25",X"02",X"26",
		X"02",X"27",X"03",X"17",X"02",X"13",X"06",X"12",X"01",X"03",X"01",X"02",X"01",X"00",X"03",X"00",
		X"01",X"0F",X"01",X"11",X"10",X"12",X"02",X"11",X"15",X"12",X"01",X"11",X"01",X"10",X"01",X"0F",
		X"02",X"00",X"03",X"00",X"01",X"01",X"01",X"02",X"01",X"03",X"0F",X"12",X"01",X"03",X"01",X"02",
		X"01",X"01",X"03",X"00",X"01",X"09",X"01",X"25",X"04",X"26",X"01",X"15",X"08",X"12",X"01",X"03",
		X"01",X"02",X"01",X"01",X"04",X"00",X"06",X"00",X"02",X"0F",X"02",X"10",X"08",X"11",X"02",X"10",
		X"01",X"0F",X"03",X"00",X"01",X"0F",X"01",X"10",X"02",X"11",X"0A",X"12",X"02",X"11",X"02",X"10",
		X"01",X"0F",X"06",X"00",X"08",X"00",X"02",X"01",X"08",X"02",X"02",X"01",X"08",X"00",X"01",X"07",
		X"01",X"08",X"01",X"16",X"01",X"15",X"01",X"12",X"03",X"03",X"02",X"02",X"02",X"01",X"09",X"00",
		X"08",X"00",X"03",X"01",X"03",X"02",X"05",X"03",X"0A",X"12",X"04",X"03",X"03",X"02",X"02",X"01",
		X"0B",X"00",X"07",X"00",X"01",X"0F",X"02",X"10",X"01",X"38",X"01",X"33",X"01",X"31",X"16",X"00",
		X"01",X"32",X"01",X"33",X"01",X"2F",X"01",X"2E",X"01",X"39",X"01",X"11",X"01",X"10",X"02",X"0F",
		X"05",X"00",X"02",X"00",X"01",X"01",X"01",X"02",X"02",X"03",X"22",X"12",X"02",X"03",X"01",X"02",
		X"01",X"01",X"05",X"00",X"02",X"00",X"01",X"0F",X"01",X"10",X"01",X"11",X"03",X"12",X"01",X"34",
		X"05",X"2F",X"01",X"0E",X"04",X"00",X"01",X"31",X"01",X"33",X"08",X"11",X"05",X"00",X"01",X"0D",
		X"01",X"06",X"04",X"2F",X"01",X"2E",X"04",X"12",X"01",X"11",X"01",X"10",X"01",X"0F",X"01",X"00",
		X"01",X"03",X"03",X"12",X"05",X"14",X"04",X"15",X"02",X"1A",X"01",X"1B",X"02",X"1A",X"01",X"1C",
		X"01",X"1B",X"01",X"1C",X"01",X"19",X"01",X"1C",X"09",X"19",X"03",X"17",X"02",X"13",X"08",X"12",
		X"01",X"03",X"01",X"02",X"01",X"01",X"01",X"00",X"01",X"10",X"07",X"12",X"05",X"2F",X"05",X"00",
		X"01",X"32",X"02",X"2F",X"08",X"12",X"07",X"00",X"05",X"2F",X"07",X"12",X"01",X"11",X"04",X"22",
		X"06",X"21",X"07",X"22",X"01",X"32",X"01",X"22",X"02",X"32",X"01",X"22",X"05",X"32",X"03",X"31",
		X"01",X"33",X"07",X"2F",X"01",X"19",X"01",X"17",X"08",X"12",X"01",X"03",X"08",X"12",X"05",X"2F",
		X"02",X"22",X"03",X"00",X"01",X"06",X"01",X"2F",X"01",X"13",X"08",X"12",X"02",X"00",X"03",X"22",
		X"02",X"21",X"02",X"1E",X"03",X"2F",X"08",X"12",X"04",X"07",X"06",X"0B",X"07",X"07",X"01",X"0D",
		X"01",X"07",X"02",X"0D",X"01",X"07",X"05",X"0D",X"03",X"0C",X"01",X"06",X"07",X"2F",X"01",X"2E",
		X"01",X"34",X"08",X"12",X"01",X"11",X"08",X"12",X"03",X"1D",X"08",X"15",X"01",X"17",X"09",X"12",
		X"0C",X"14",X"07",X"12",X"01",X"03",X"01",X"11",X"03",X"12",X"05",X"2A",X"04",X"28",X"02",X"2B",
		X"01",X"35",X"02",X"2B",X"01",X"2C",X"01",X"35",X"01",X"2C",X"01",X"2E",X"01",X"2C",X"09",X"2E",
		X"03",X"34",X"02",X"30",X"08",X"12",X"01",X"11",X"01",X"10",X"01",X"0F",X"01",X"00",X"01",X"00",
		X"02",X"01",X"01",X"02",X"02",X"03",X"22",X"12",X"02",X"03",X"02",X"02",X"02",X"01",X"03",X"00",
		X"02",X"00",X"01",X"0F",X"01",X"10",X"02",X"11",X"22",X"12",X"02",X"11",X"01",X"10",X"01",X"0F",
		X"05",X"00",X"08",X"00",X"02",X"01",X"02",X"02",X"03",X"03",X"0E",X"12",X"04",X"03",X"03",X"02",
		X"02",X"01",X"0B",X"00",X"08",X"00",X"03",X"0F",X"03",X"10",X"05",X"11",X"0A",X"12",X"04",X"11",
		X"03",X"10",X"02",X"0F",X"0B",X"00",X"1D",X"00",X"01",X"31",X"01",X"2F",X"01",X"2E",X"01",X"30",
		X"03",X"11",X"02",X"10",X"02",X"0F",X"09",X"00",X"1C",X"00",X"01",X"33",X"04",X"2F",X"01",X"2E",
		X"01",X"30",X"07",X"12",X"02",X"11",X"01",X"10",X"01",X"0F",X"03",X"00",X"1D",X"00",X"01",X"0C",
		X"01",X"2F",X"01",X"1E",X"01",X"1F",X"01",X"27",X"05",X"26",X"02",X"29",X"01",X"2D",X"01",X"2A",
		X"04",X"12",X"01",X"11",X"01",X"10",X"21",X"00",X"02",X"07",X"02",X"36",X"02",X"37",X"04",X"2F",
		X"06",X"12",X"04",X"21",X"03",X"25",X"03",X"21",X"05",X"22",X"10",X"00",X"03",X"22",X"01",X"21",
		X"02",X"1F",X"01",X"24",X"01",X"1E",X"02",X"06",X"02",X"2F",X"06",X"12",X"03",X"12",X"02",X"14",
		X"03",X"15",X"04",X"16",X"15",X"26",X"04",X"16",X"04",X"15",X"02",X"14",X"05",X"12",X"01",X"03",
		X"01",X"00",X"02",X"01",X"01",X"02",X"02",X"03",X"22",X"12",X"02",X"03",X"02",X"02",X"02",X"01",
		X"03",X"00",X"08",X"00",X"02",X"01",X"02",X"02",X"03",X"03",X"0E",X"12",X"04",X"03",X"03",X"02",
		X"02",X"01",X"0B",X"00",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"7E",X"7B",X"2A",X"7E",X"7B",X"74",X"7E",X"7B",X"9C",X"7E",X"7B",X"22",X"7E",X"7B",X"6D",X"7E",
		X"7B",X"95",X"7E",X"7B",X"CA",X"7E",X"7B",X"BD",X"7B",X"EF",X"7E",X"7B",X"C5",X"7E",X"7B",X"B8",
		X"7C",X"59",X"34",X"67",X"10",X"8E",X"7C",X"59",X"20",X"06",X"34",X"67",X"10",X"8E",X"7B",X"EF",
		X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"11",X"7F",X"CA",X"01",X"35",X"E7",X"84",X"0F",X"81",X"0A",
		X"2F",X"02",X"86",X"0A",X"10",X"BE",X"BF",X"02",X"BF",X"CA",X"04",X"48",X"81",X"6A",X"25",X"02",
		X"86",X"5C",X"10",X"AE",X"A6",X"EC",X"A1",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"10",X"BF",
		X"CA",X"02",X"C6",X"1A",X"F7",X"CA",X"00",X"88",X"04",X"5F",X"30",X"8B",X"39",X"34",X"67",X"CE",
		X"7C",X"59",X"20",X"05",X"34",X"67",X"CE",X"7B",X"EF",X"1A",X"FF",X"FF",X"BF",X"02",X"F7",X"CA",
		X"01",X"CE",X"83",X"B6",X"33",X"C6",X"EE",X"C6",X"A6",X"C4",X"8D",X"B8",X"A6",X"C0",X"2A",X"F8",
		X"7F",X"CA",X"01",X"35",X"E7",X"34",X"67",X"CE",X"7C",X"59",X"20",X"05",X"34",X"67",X"CE",X"7B",
		X"EF",X"1A",X"FF",X"FF",X"BF",X"02",X"F7",X"CA",X"01",X"44",X"44",X"44",X"44",X"8D",X"8D",X"A6",
		X"61",X"8D",X"89",X"7F",X"CA",X"01",X"35",X"E7",X"7C",X"BF",X"27",X"20",X"03",X"7F",X"BF",X"27",
		X"CE",X"7B",X"0C",X"20",X"0B",X"7C",X"BF",X"27",X"20",X"03",X"7F",X"BF",X"27",X"CE",X"7B",X"03",
		X"10",X"8E",X"8D",X"83",X"48",X"31",X"B6",X"AE",X"A1",X"E6",X"A0",X"7D",X"BF",X"27",X"27",X"01",
		X"5F",X"A6",X"A4",X"84",X"7F",X"AD",X"C4",X"A6",X"A0",X"2A",X"EC",X"7F",X"CA",X"01",X"39",X"7C",
		X"C3",X"7C",X"DA",X"7C",X"F1",X"7D",X"08",X"7D",X"1F",X"7D",X"36",X"7D",X"4D",X"7D",X"64",X"7D",
		X"7B",X"7D",X"92",X"7D",X"A9",X"7D",X"C0",X"7D",X"D7",X"7D",X"EE",X"7E",X"05",X"7E",X"1C",X"7E",
		X"33",X"7E",X"4A",X"7E",X"61",X"7E",X"78",X"7E",X"88",X"7E",X"9F",X"7E",X"B6",X"7E",X"CD",X"7E",
		X"EB",X"7F",X"02",X"7F",X"19",X"7F",X"30",X"7F",X"47",X"7F",X"5E",X"7F",X"75",X"7F",X"8C",X"7F",
		X"A3",X"7F",X"BA",X"7F",X"D8",X"7F",X"EF",X"80",X"06",X"80",X"1D",X"80",X"31",X"80",X"42",X"80",
		X"50",X"80",X"67",X"80",X"70",X"80",X"80",X"80",X"90",X"80",X"94",X"80",X"A4",X"80",X"AD",X"80",
		X"C4",X"80",X"DB",X"80",X"E1",X"80",X"F1",X"81",X"0B",X"81",X"22",X"81",X"2E",X"81",X"3A",X"81",
		X"46",X"81",X"52",X"81",X"5E",X"81",X"6A",X"81",X"76",X"81",X"82",X"81",X"8E",X"81",X"9A",X"81",
		X"A6",X"81",X"B2",X"81",X"BE",X"81",X"CA",X"81",X"D6",X"81",X"E2",X"81",X"EE",X"81",X"FA",X"82",
		X"06",X"82",X"12",X"82",X"1E",X"82",X"2A",X"82",X"36",X"82",X"47",X"81",X"22",X"82",X"53",X"82",
		X"5F",X"82",X"6B",X"81",X"5E",X"82",X"77",X"82",X"83",X"82",X"8F",X"82",X"E9",X"82",X"FA",X"83",
		X"06",X"83",X"12",X"83",X"1E",X"83",X"2A",X"83",X"34",X"83",X"3C",X"83",X"48",X"83",X"4F",X"83",
		X"5B",X"83",X"67",X"83",X"6B",X"83",X"72",X"83",X"79",X"83",X"99",X"83",X"AA",X"83",X"72",X"83",
		X"72",X"83",X"72",X"03",X"07",X"11",X"11",X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"10",X"01",
		X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"03",X"07",X"00",X"11",X"10",X"01",
		X"11",X"10",X"11",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",
		X"10",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"11",X"00",X"01",
		X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"10",
		X"00",X"01",X"10",X"01",X"11",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"11",X"11",X"10",X"03",
		X"07",X"00",X"01",X"10",X"00",X"11",X"10",X"01",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",
		X"00",X"01",X"10",X"00",X"01",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"11",
		X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",
		X"10",X"11",X"11",X"10",X"03",X"07",X"01",X"11",X"10",X"00",X"01",X"10",X"00",X"11",X"00",X"01",
		X"10",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"03",X"07",X"11",X"11",X"10",
		X"11",X"00",X"10",X"11",X"00",X"10",X"01",X"11",X"00",X"11",X"00",X"10",X"11",X"00",X"10",X"11",
		X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",
		X"00",X"00",X"10",X"00",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"11",X"11",X"10",X"11",X"11",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"10",X"01",
		X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"03",X"07",X"11",X"11",X"00",X"11",X"01",X"10",X"11",
		X"01",X"10",X"11",X"11",X"00",X"11",X"01",X"10",X"11",X"01",X"10",X"11",X"11",X"00",X"03",X"07",
		X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",
		X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"00",X"10",X"01",X"10",X"10",X"01",X"10",
		X"10",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"11",X"11",X"00",X"03",X"07",X"11",X"11",
		X"10",X"11",X"00",X"00",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",
		X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"11",X"00",X"11",X"00",
		X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"03",X"07",X"11",X"11",X"10",X"11",
		X"01",X"10",X"11",X"00",X"00",X"11",X"01",X"10",X"11",X"00",X"10",X"11",X"11",X"10",X"11",X"11",
		X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",X"11",
		X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"02",X"07",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"03",X"07",X"00",X"01",X"10",X"00",X"01",X"10",
		X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"03",
		X"07",X"11",X"00",X"10",X"11",X"01",X"00",X"11",X"10",X"00",X"11",X"10",X"00",X"11",X"11",X"00",
		X"11",X"01",X"10",X"11",X"00",X"10",X"03",X"07",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"10",X"11",X"11",X"10",X"04",X"07",X"11",
		X"11",X"11",X"10",X"11",X"00",X"10",X"10",X"11",X"00",X"10",X"10",X"11",X"00",X"10",X"10",X"11",
		X"00",X"10",X"10",X"11",X"00",X"00",X"10",X"11",X"00",X"00",X"10",X"03",X"07",X"11",X"11",X"10",
		X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",
		X"00",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",
		X"11",X"00",X"10",X"11",X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",
		X"10",X"11",X"11",X"10",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",
		X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"10",
		X"10",X"11",X"01",X"00",X"11",X"10",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",
		X"11",X"10",X"11",X"10",X"00",X"11",X"11",X"00",X"11",X"01",X"10",X"11",X"00",X"10",X"03",X"07",
		X"11",X"11",X"10",X"10",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"11",
		X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"01",X"10",X"00",X"01",X"10",X"00",
		X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"03",X"07",X"11",X"00",
		X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",
		X"11",X"11",X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",
		X"10",X"01",X"01",X"00",X"01",X"11",X"00",X"00",X"11",X"00",X"04",X"07",X"11",X"00",X"00",X"10",
		X"11",X"00",X"00",X"10",X"11",X"00",X"00",X"10",X"11",X"01",X"00",X"10",X"11",X"01",X"00",X"10",
		X"11",X"01",X"00",X"10",X"11",X"11",X"11",X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",
		X"01",X"11",X"00",X"00",X"10",X"00",X"01",X"01",X"00",X"11",X"00",X"10",X"11",X"00",X"10",X"03",
		X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"01",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"00",X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"10",X"11",X"11",X"10",X"03",X"06",X"00",
		X"00",X"00",X"00",X"10",X"00",X"01",X"10",X"00",X"11",X"11",X"10",X"01",X"10",X"00",X"00",X"10",
		X"00",X"03",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"11",
		X"11",X"10",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",
		X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"07",X"10",X"10",X"10",X"10",X"10",X"00",X"10",
		X"02",X"07",X"00",X"10",X"01",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",
		X"02",X"07",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"01",X"00",X"10",X"00",
		X"01",X"02",X"10",X"10",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"11",X"00",X"01",X"00",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"03",X"07",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"00",X"03",X"07",X"01",X"00",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"01",
		X"00",X"00",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"10",X"10",X"02",X"02",X"10",X"10",X"10",
		X"10",X"02",X"07",X"00",X"00",X"11",X"10",X"11",X"10",X"00",X"00",X"00",X"00",X"11",X"10",X"11",
		X"10",X"03",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"00",X"10",X"00",
		X"01",X"11",X"00",X"11",X"11",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",
		X"10",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"10",X"02",X"05",
		X"01",X"00",X"11",X"00",X"01",X"00",X"01",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",
		X"11",X"10",X"10",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"11",X"10",X"00",X"10",
		X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"02",X"05",
		X"11",X"10",X"10",X"00",X"11",X"10",X"00",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",
		X"11",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"01",X"00",
		X"01",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",X"02",X"05",
		X"11",X"10",X"10",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"02",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",
		X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"11",X"10",X"02",X"05",
		X"11",X"10",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"10",X"02",X"05",X"11",X"00",X"10",X"10",
		X"10",X"10",X"10",X"10",X"11",X"00",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"00",X"10",X"00",
		X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"00",X"10",X"00",X"10",X"00",X"02",X"05",
		X"11",X"10",X"10",X"00",X"10",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",
		X"11",X"10",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",X"00",X"01",X"00",X"01",X"00",
		X"11",X"10",X"02",X"05",X"00",X"10",X"00",X"10",X"00",X"10",X"10",X"10",X"11",X"10",X"02",X"05",
		X"10",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"10",X"00",X"10",X"00",
		X"10",X"00",X"10",X"00",X"11",X"10",X"03",X"05",X"11",X"11",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"00",X"10",X"00",X"02",
		X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"00",X"10",X"02",X"05",X"11",X"10",X"10",
		X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",X"00",X"01",X"00",X"01",
		X"00",X"01",X"00",X"02",X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"10",X"02",
		X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"00",X"20",X"42",X"55",X"42",X"42",
		X"4C",X"45",X"53",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",
		X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",
		X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"03",X"05",X"10",X"00",X"10",X"10",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",
		X"01",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"10",X"01",X"00",
		X"01",X"00",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"11",X"10",X"02",X"05",
		X"00",X"10",X"01",X"00",X"11",X"10",X"01",X"00",X"00",X"10",X"02",X"04",X"00",X"00",X"11",X"10",
		X"00",X"00",X"11",X"10",X"02",X"03",X"00",X"00",X"00",X"00",X"11",X"10",X"02",X"05",X"11",X"10",
		X"00",X"10",X"01",X"10",X"00",X"00",X"01",X"00",X"01",X"05",X"10",X"10",X"10",X"00",X"10",X"02",
		X"05",X"00",X"10",X"01",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"02",X"05",X"10",X"00",X"01",
		X"00",X"00",X"10",X"01",X"00",X"10",X"00",X"01",X"02",X"10",X"10",X"01",X"05",X"00",X"00",X"00",
		X"10",X"10",X"01",X"05",X"00",X"00",X"00",X"00",X"10",X"06",X"05",X"11",X"10",X"11",X"10",X"11",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"03",X"05",X"00",X"10",X"00",X"00",X"11",
		X"00",X"11",X"11",X"10",X"00",X"11",X"00",X"00",X"10",X"00",X"02",X"05",X"11",X"10",X"11",X"10",
		X"11",X"10",X"11",X"10",X"11",X"10",X"85",X"09",X"84",X"B6",X"84",X"D4",X"84",X"EF",X"84",X"FB",
		X"85",X"13",X"85",X"29",X"85",X"37",X"85",X"41",X"85",X"4B",X"85",X"56",X"85",X"66",X"85",X"7B",
		X"85",X"8F",X"85",X"91",X"85",X"98",X"85",X"A6",X"85",X"BD",X"85",X"D9",X"85",X"F1",X"85",X"FF",
		X"86",X"1B",X"86",X"26",X"86",X"2D",X"86",X"34",X"86",X"3E",X"86",X"4E",X"86",X"57",X"86",X"62",
		X"86",X"6D",X"86",X"7D",X"86",X"8D",X"86",X"96",X"86",X"A0",X"86",X"B0",X"86",X"BA",X"86",X"CC",
		X"86",X"DB",X"86",X"EC",X"86",X"FC",X"87",X"08",X"87",X"10",X"87",X"25",X"87",X"35",X"87",X"48",
		X"87",X"58",X"87",X"6C",X"87",X"83",X"87",X"93",X"87",X"A2",X"87",X"B7",X"87",X"D1",X"87",X"E2",
		X"87",X"F5",X"88",X"0A",X"88",X"1E",X"88",X"3B",X"88",X"5E",X"88",X"7E",X"88",X"90",X"88",X"A9",
		X"88",X"C1",X"88",X"D9",X"88",X"EF",X"88",X"F9",X"89",X"11",X"89",X"27",X"89",X"3C",X"89",X"64",
		X"89",X"67",X"89",X"71",X"89",X"77",X"89",X"91",X"89",X"99",X"89",X"B2",X"89",X"D4",X"89",X"EF",
		X"89",X"F7",X"8A",X"0D",X"8A",X"21",X"8A",X"2E",X"8A",X"36",X"8A",X"4A",X"8B",X"2B",X"8B",X"3B",
		X"8B",X"60",X"8A",X"68",X"8A",X"86",X"8A",X"99",X"8A",X"AE",X"8A",X"BE",X"8A",X"FE",X"85",X"09",
		X"8B",X"20",X"8B",X"73",X"8B",X"7B",X"8D",X"13",X"8B",X"83",X"8B",X"B4",X"8B",X"CB",X"8B",X"BE",
		X"8B",X"DA",X"8B",X"D4",X"8B",X"F0",X"8B",X"DF",X"8B",X"FD",X"8B",X"FF",X"8C",X"0F",X"8C",X"19",
		X"86",X"A7",X"8C",X"C5",X"8C",X"40",X"8C",X"55",X"8C",X"66",X"8C",X"7D",X"8C",X"95",X"8C",X"A2",
		X"8C",X"B2",X"8C",X"C1",X"8B",X"9B",X"8C",X"29",X"8C",X"F4",X"8A",X"E2",X"8C",X"DB",X"8D",X"26",
		X"8D",X"41",X"8D",X"57",X"8D",X"6C",X"1D",X"13",X"18",X"15",X"0A",X"0F",X"18",X"0E",X"1D",X"0A",
		X"21",X"12",X"0F",X"18",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"1D",X"0A",X"0B",X"1C",X"0F",X"0A",
		X"11",X"19",X"18",X"8F",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"0A",X"13",X"1D",X"0A",X"21",X"0B",
		X"1D",X"12",X"0F",X"0E",X"0A",X"0E",X"19",X"21",X"18",X"0A",X"0E",X"1C",X"0B",X"13",X"98",X"1E",
		X"19",X"0A",X"11",X"0F",X"1E",X"0A",X"0C",X"1C",X"19",X"19",X"97",X"1E",X"19",X"1F",X"0D",X"12",
		X"0A",X"13",X"1E",X"0A",X"10",X"13",X"1C",X"1D",X"9E",X"11",X"0B",X"17",X"0F",X"0A",X"19",X"20",
		X"0F",X"1C",X"8A",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"0A",X"1E",X"0F",X"1D",X"1E",X"1D",
		X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",X"8F",X"0B",X"16",X"16",X"0A",X"1D",X"23",X"1D",
		X"1E",X"0F",X"17",X"1D",X"0A",X"11",X"99",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",
		X"8A",X"1C",X"19",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"0B",X"16",X"16",X"0A",X"1C",
		X"19",X"17",X"1D",X"0A",X"19",X"95",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",
		X"19",X"16",X"16",X"19",X"21",X"9D",X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",
		X"18",X"0D",X"0F",X"0A",X"1E",X"19",X"0A",X"0F",X"22",X"13",X"9E",X"0A",X"1C",X"0B",X"17",X"0A",
		X"0F",X"1C",X"1C",X"19",X"1C",X"1D",X"0A",X"0E",X"0F",X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",
		X"99",X"18",X"19",X"0A",X"0D",X"17",X"19",X"9D",X"0D",X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",
		X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",
		X"0A",X"17",X"1F",X"1D",X"1E",X"0A",X"0C",X"0F",X"0A",X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",
		X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"1A",X"0A",X"1C",X"0B",X"1D",X"13",X"0F",X"0E",
		X"0A",X"10",X"19",X"1C",X"0A",X"1E",X"0F",X"1D",X"9E",X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",
		X"0F",X"0A",X"1A",X"1C",X"19",X"1E",X"0F",X"0D",X"1E",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",
		X"8F",X"0D",X"19",X"16",X"19",X"1C",X"0A",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"9E",X"20",
		X"0F",X"1C",X"1E",X"13",X"0D",X"0B",X"16",X"0A",X"0C",X"0B",X"1C",X"1D",X"0A",X"13",X"18",X"0E",
		X"13",X"0D",X"0B",X"1E",X"0F",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"1D",X"21",X"13",X"1E",X"0D",
		X"12",X"0A",X"1E",X"0F",X"1D",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",
		X"0B",X"18",X"0D",X"8F",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",
		X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",
		X"10",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",
		X"13",X"98",X"1D",X"16",X"0B",X"17",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"17",X"19",X"20",
		X"0F",X"0A",X"16",X"0F",X"10",X"9E",X"17",X"19",X"20",X"0F",X"0A",X"1C",X"13",X"11",X"12",X"9E",
		X"17",X"19",X"20",X"0F",X"0A",X"1F",X"9A",X"17",X"19",X"20",X"0F",X"0A",X"0E",X"19",X"21",X"98",
		X"1D",X"19",X"1F",X"18",X"0E",X"0A",X"16",X"13",X"18",X"8F",X"0C",X"19",X"19",X"15",X"15",X"0F",
		X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"16",X"0F",X"10",X"1E",
		X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",
		X"1C",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1C",X"13",X"11",X"12",
		X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1A",X"0B",X"13",X"0E",
		X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"9D",X"10",X"1C",X"0F",X"0F",X"0A",X"17",X"0F",X"98",
		X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"13",X"18",X"0A",X"17",X"13",
		X"18",X"1F",X"1E",X"0F",X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"17",X"0F",X"18",X"0A",X"1A",
		X"16",X"0B",X"23",X"0F",X"8E",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1D",X"13",X"18",X"11",X"16",
		X"0F",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1E",X"21",
		X"19",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",
		X"0F",X"0E",X"13",X"1E",X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",
		X"0B",X"11",X"0F",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"9E",X"11",X"0B",X"17",X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",
		X"18",X"1E",X"9D",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"17",X"0B",X"18",X"0A",X"0F",X"20",X"0F",
		X"1C",X"A3",X"17",X"0F",X"18",X"0A",X"10",X"19",X"1C",X"0A",X"01",X"0A",X"0D",X"1C",X"0F",X"0E",
		X"13",X"1E",X"0A",X"11",X"0B",X"17",X"8F",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",
		X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0B",X"1E",X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",X"0F",
		X"8E",X"1A",X"1C",X"13",X"0D",X"13",X"18",X"11",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"13",
		X"19",X"98",X"0A",X"0A",X"0A",X"0A",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",
		X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1C",X"13",
		X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",
		X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",
		X"0A",X"10",X"19",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"1F",
		X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",
		X"1C",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",
		X"0A",X"0A",X"17",X"13",X"18",X"13",X"17",X"1F",X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",
		X"10",X"19",X"1C",X"0A",X"0B",X"18",X"23",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0E",X"13",
		X"10",X"10",X"13",X"0D",X"1F",X"16",X"1E",X"23",X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",
		X"16",X"0F",X"1E",X"1E",X"0F",X"1C",X"1D",X"0A",X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",
		X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",X"1C",X"8F",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",
		X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",
		X"9D",X"0D",X"16",X"0F",X"0B",X"1C",X"0A",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",
		X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",
		X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"0B",
		X"1F",X"1E",X"19",X"0A",X"0D",X"23",X"0D",X"16",X"8F",X"1D",X"0F",X"1E",X"0A",X"0B",X"1E",X"1E",
		X"1C",X"0B",X"0D",X"1E",X"0A",X"17",X"19",X"0E",X"0F",X"0A",X"17",X"0F",X"1D",X"1D",X"0B",X"11",
		X"8F",X"1D",X"0F",X"1E",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",
		X"1C",X"0F",X"0A",X"18",X"0B",X"17",X"8F",X"1F",X"1D",X"0F",X"0A",X"2C",X"17",X"19",X"20",X"0F",
		X"2C",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"8A",X"1F",X"1D",X"0F",X"0A",
		X"2C",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"2C",X"0A",X"0C",X"19",X"1E",X"1E",X"19",X"18",X"1D",
		X"0A",X"1E",X"19",X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"20",
		X"0B",X"16",X"1F",X"8F",X"23",X"0F",X"9D",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",
		X"9E",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"17",X"19",X"20",X"0F",X"0A",X"0E",X"19",X"21",X"18",
		X"0A",X"10",X"19",X"1C",X"0A",X"13",X"18",X"1D",X"1E",X"1C",X"1F",X"0D",X"1E",X"13",X"19",X"18",
		X"9D",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",
		X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"1D",X"0A",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",
		X"0F",X"8E",X"0C",X"23",X"0A",X"19",X"1A",X"0F",X"18",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",
		X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",
		X"0A",X"1E",X"19",X"9A",X"0B",X"18",X"0E",X"0A",X"1E",X"1F",X"1C",X"18",X"13",X"18",X"11",X"0A",
		X"11",X"0B",X"17",X"0F",X"0A",X"19",X"18",X"0A",X"0B",X"18",X"0E",X"0A",X"19",X"10",X"90",X"0A",
		X"0D",X"16",X"0F",X"0B",X"1C",X"0F",X"8E",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",
		X"0F",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"1E",X"19",X"0E",
		X"0B",X"23",X"2C",X"1D",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",
		X"9D",X"0C",X"0F",X"1D",X"1E",X"0A",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"9D",X"0D",X"1C",
		X"0F",X"0E",X"13",X"1E",X"1D",X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"17",X"19",X"20",X"0F",X"2C",
		X"0A",X"1E",X"19",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"9C",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"16",X"13",X"18",X"0F",X"0A",X"0C",X"23",X"0A",X"1A",X"1C",X"0F",X"1D",X"1D",X"13",X"18",X"11",
		X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",X"23",X"19",X"1F",X"2C",X"1C",X"0F",X"0A",X"1E",
		X"12",X"0F",X"0A",X"0C",X"0F",X"1D",X"1E",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"1D",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"1C",
		X"0A",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"9D",X"23",X"19",X"1F",X"0A",X"0B",X"1C",X"0F",
		X"0A",X"0B",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"1D",X"0A",X"1A",X"1C",X"99",X"17",X"0B",
		X"22",X"13",X"17",X"1F",X"17",X"0A",X"05",X"0A",X"0F",X"18",X"1E",X"1C",X"23",X"9D",X"1F",X"1D",
		X"0F",X"0A",X"27",X"17",X"19",X"20",X"0F",X"0A",X"1F",X"1A",X"2D",X"0A",X"0E",X"19",X"21",X"18",
		X"27",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"0A",X"16",X"0F",X"1E",X"1E",
		X"0F",X"9C",X"27",X"17",X"19",X"20",X"0F",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"27",X"0A",X"1E",
		X"19",X"0A",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"2A",X"0D",
		X"2B",X"0A",X"01",X"09",X"08",X"02",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",
		X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",
		X"0A",X"0A",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"1E",X"12",X"13",X"1D",X"0A",
		X"13",X"1D",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"1D",X"AE",X"0E",X"0F",X"1D",X"13",X"11",
		X"18",X"0F",X"0E",X"0A",X"0C",X"23",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",
		X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",
		X"0B",X"16",X"16",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"1D",X"0A",X"1C",X"0F",X"1D",X"0F",X"1C",
		X"20",X"0F",X"8E",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"81",X"1A",X"16",X"0B",X"23",X"0F",
		X"1C",X"0A",X"82",X"0D",X"16",X"0F",X"0B",X"18",X"0A",X"1F",X"1A",X"0A",X"19",X"18",X"0A",X"1E",
		X"12",X"0F",X"1D",X"0F",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"9D",X"0E",X"19",X"18",X"2C",X"1E",
		X"0A",X"1E",X"19",X"1F",X"0D",X"12",X"0A",X"1E",X"12",X"0F",X"1D",X"0F",X"0A",X"0F",X"18",X"0F",
		X"17",X"13",X"0F",X"9D",X"0D",X"1C",X"1F",X"17",X"0A",X"26",X"0A",X"01",X"00",X"80",X"11",X"1C",
		X"0F",X"0B",X"1D",X"13",X"0F",X"0A",X"26",X"0A",X"02",X"00",X"80",X"0B",X"18",X"1E",X"0A",X"26",
		X"0A",X"01",X"05",X"80",X"1D",X"1A",X"19",X"18",X"11",X"8F",X"0C",X"1C",X"1F",X"1D",X"92",X"26",
		X"0A",X"05",X"00",X"00",X"0A",X"1A",X"16",X"1F",X"1D",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"9D",
		X"0D",X"16",X"0F",X"0B",X"18",X"13",X"18",X"11",X"0A",X"16",X"0B",X"0E",X"A3",X"02",X"A2",X"0C",
		X"19",X"18",X"1F",X"1D",X"0A",X"17",X"1F",X"16",X"1E",X"13",X"1A",X"16",X"13",X"0F",X"9C",X"0C",
		X"0F",X"0A",X"0D",X"0B",X"1C",X"0F",X"10",X"1F",X"96",X"0B",X"1C",X"19",X"1F",X"18",X"0E",X"0A",
		X"1E",X"12",X"0F",X"0A",X"0E",X"1C",X"0B",X"13",X"98",X"1F",X"18",X"16",X"0F",X"1D",X"1D",X"0A",
		X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"0A",X"12",X"0B",X"1D",X"0A",X"17",X"19",X"1F",X"1E",X"92",
		X"0C",X"0F",X"21",X"0B",X"1C",X"0F",X"29",X"0A",X"1E",X"19",X"0A",X"15",X"13",X"16",X"16",X"0A",
		X"1C",X"19",X"0B",X"0D",X"92",X"1E",X"19",X"1F",X"0D",X"12",X"0A",X"21",X"13",X"1E",X"12",X"0A",
		X"0C",X"1C",X"19",X"19",X"17",X"8A",X"0E",X"13",X"20",X"0F",X"0A",X"0B",X"12",X"0F",X"0B",X"0E",
		X"0A",X"19",X"18",X"0F",X"0A",X"1D",X"13",X"18",X"15",X"0A",X"0B",X"18",X"8E",X"0D",X"19",X"16",
		X"16",X"0F",X"0D",X"1E",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"21",X"12",X"0F",X"18",X"0A",
		X"0E",X"1C",X"0B",X"13",X"98",X"10",X"16",X"0B",X"1D",X"12",X"0F",X"1D",X"0A",X"11",X"1C",X"0F",
		X"0F",X"98",X"1C",X"0B",X"24",X"19",X"1C",X"0A",X"0C",X"16",X"0B",X"0E",X"0F",X"1D",X"0A",X"0D",
		X"0B",X"98",X"0B",X"16",X"21",X"0B",X"23",X"1D",X"0A",X"12",X"1F",X"1C",X"1E",X"0A",X"23",X"19",
		X"9F",X"1D",X"13",X"18",X"95",X"0F",X"18",X"0E",X"0A",X"1D",X"13",X"18",X"15",X"0A",X"0C",X"19",
		X"18",X"1F",X"1D",X"0A",X"0A",X"0A",X"22",X"0A",X"02",X"05",X"80",X"0E",X"13",X"20",X"0F",X"0A",
		X"0B",X"12",X"0F",X"0B",X"0E",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0A",X"0A",X"22",X"0A",
		X"01",X"00",X"00",X"80",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",
		X"0A",X"0F",X"20",X"0F",X"1C",X"23",X"0A",X"0A",X"0A",X"00",X"00",X"00",X"0A",X"1A",X"19",X"13",
		X"18",X"1E",X"9D",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"0A",X"11",X"1C",X"19",X"21",X"1D",X"0A",
		X"0B",X"1D",X"0A",X"23",X"19",X"9F",X"27",X"17",X"19",X"20",X"0F",X"0A",X"16",X"0F",X"10",X"1E",
		X"27",X"0A",X"1E",X"19",X"0A",X"0F",X"1C",X"0B",X"1D",X"0F",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",
		X"9C",X"19",X"19",X"1A",X"1D",X"29",X"0A",X"0C",X"1F",X"0C",X"0C",X"16",X"0F",X"0A",X"1E",X"19",
		X"19",X"0A",X"1D",X"17",X"0B",X"16",X"96",X"02",X"22",X"0A",X"20",X"0B",X"16",X"1F",X"0F",X"0A",
		X"0B",X"1C",X"19",X"1F",X"18",X"0E",X"0A",X"0E",X"1C",X"0B",X"13",X"98",X"17",X"19",X"20",X"0F",
		X"0A",X"1F",X"1A",X"0A",X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",
		X"1C",X"0F",X"9D",X"8D",X"E7",X"8D",X"F3",X"8D",X"FB",X"8E",X"03",X"8E",X"07",X"8E",X"17",X"8E",
		X"1F",X"8E",X"23",X"8E",X"27",X"8E",X"2B",X"8E",X"3B",X"8E",X"3F",X"8E",X"53",X"8E",X"57",X"8E",
		X"5F",X"8E",X"63",X"8E",X"6B",X"8E",X"6F",X"8E",X"7F",X"8E",X"83",X"8E",X"87",X"8E",X"93",X"8E",
		X"97",X"8E",X"9B",X"8E",X"9F",X"8E",X"A3",X"8E",X"A7",X"8E",X"AB",X"8E",X"AB",X"8E",X"B3",X"8E",
		X"BB",X"8E",X"BF",X"8E",X"C7",X"8E",X"CF",X"8E",X"DB",X"8E",X"DF",X"8E",X"E3",X"8E",X"E7",X"8E",
		X"73",X"8E",X"EB",X"8E",X"EF",X"8E",X"F7",X"8F",X"03",X"8F",X"07",X"8F",X"13",X"8F",X"13",X"8F",
		X"1B",X"8F",X"23",X"8F",X"27",X"8F",X"2B",X"3E",X"50",X"99",X"09",X"36",X"90",X"33",X"0A",X"2E",
		X"A0",X"33",X"8B",X"2A",X"80",X"99",X"0D",X"30",X"80",X"99",X"8C",X"21",X"80",X"99",X"0E",X"37",
		X"80",X"99",X"8C",X"36",X"80",X"22",X"8F",X"36",X"80",X"22",X"0F",X"28",X"90",X"22",X"12",X"17",
		X"A0",X"99",X"10",X"17",X"A8",X"99",X"91",X"3A",X"80",X"33",X"13",X"24",X"B0",X"33",X"94",X"3A",
		X"20",X"88",X"95",X"2F",X"10",X"99",X"A3",X"2F",X"10",X"99",X"AF",X"23",X"D7",X"BB",X"42",X"4C",
		X"D7",X"BB",X"45",X"25",X"DF",X"44",X"43",X"34",X"E7",X"11",X"8B",X"28",X"16",X"BB",X"C0",X"30",
		X"80",X"22",X"45",X"4F",X"80",X"22",X"48",X"27",X"A0",X"22",X"3C",X"19",X"B0",X"22",X"4A",X"23",
		X"C0",X"22",X"CB",X"21",X"80",X"99",X"C9",X"24",X"60",X"33",X"23",X"59",X"60",X"33",X"CC",X"2A",
		X"40",X"88",X"CD",X"2D",X"1D",X"00",X"4E",X"35",X"63",X"AA",X"CF",X"28",X"16",X"BB",X"C1",X"33",
		X"46",X"11",X"D3",X"12",X"DC",X"AA",X"5B",X"5E",X"DC",X"AA",X"55",X"28",X"E4",X"AA",X"D4",X"3E",
		X"47",X"AA",X"DE",X"3E",X"47",X"AA",X"DF",X"14",X"54",X"22",X"60",X"0F",X"5C",X"22",X"61",X"0F",
		X"9C",X"22",X"FE",X"56",X"54",X"44",X"F7",X"11",X"68",X"11",X"E2",X"11",X"90",X"11",X"E4",X"11",
		X"7C",X"11",X"E3",X"6C",X"7F",X"99",X"E6",X"6C",X"6C",X"99",X"E5",X"11",X"B6",X"11",X"67",X"11",
		X"BD",X"11",X"E8",X"40",X"A4",X"44",X"6B",X"3A",X"AB",X"44",X"EC",X"5A",X"5C",X"44",X"F8",X"62",
		X"90",X"99",X"74",X"64",X"97",X"99",X"F5",X"58",X"B6",X"99",X"6F",X"5B",X"BD",X"99",X"F0",X"30",
		X"C7",X"33",X"71",X"23",X"CF",X"33",X"72",X"32",X"DC",X"AA",X"FF",X"58",X"CF",X"FF",X"F3",X"3C",
		X"58",X"11",X"DC",X"23",X"51",X"88",X"EE",X"20",X"51",X"88",X"FB",X"2C",X"13",X"11",X"D0",X"2E",
		X"DC",X"AA",X"79",X"32",X"E4",X"AA",X"C7",X"28",X"CA",X"AA",X"5A",X"2D",X"D4",X"AA",X"7A",X"2D",
		X"E0",X"AA",X"FC",X"28",X"42",X"AA",X"FD",X"12",X"C0",X"AA",X"5A",X"20",X"D0",X"AA",X"7A",X"20",
		X"E0",X"AA",X"FC",X"32",X"DC",X"AA",X"7F",X"2F",X"E4",X"AA",X"C7",X"11",X"B6",X"11",X"03",X"11",
		X"BD",X"11",X"84",X"2D",X"1D",X"AA",X"CE",X"2F",X"C7",X"33",X"81",X"17",X"CF",X"33",X"02",X"51",
		X"CF",X"33",X"F8",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
