-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "F50003F00FC00FC0FFFF0000005F0FC000030003C000C00001F41FBD00000000";
    attribute INIT_01 of inst : label is "5FC0000003F003F05555000003F5000000030003C000C00003E0000000000000";
    attribute INIT_02 of inst : label is "00000000C0000000FFFFFFFF03FC03C0000103FF000000000000000000000000";
    attribute INIT_03 of inst : label is "C003D55700030000FFFFFFFF3FC003C04000FFC0000000000000000000000000";
    attribute INIT_04 of inst : label is "01800000000000000000000000000000000000000000000003F0004000000000";
    attribute INIT_05 of inst : label is "00000000000003C00000000000000000F800C000002F00030000000000000000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0000000000F400E009D818C907C002C0F82FC003014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC6832558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "00001555C000C000FFFFEAABC003C00300030003201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "C050FA9401A405ABFA400C00006B0030CC00FA800424010BC000C64000000040";
    attribute INIT_0D of inst : label is "00C0000000C00000C000C000F6C9AAAA0000000000000000FA40180001AB000A";
    attribute INIT_0E of inst : label is "6A6798332A510000093E014E007F03FFFD00FFC00C60B38045A80000D929C90E";
    attribute INIT_0F of inst : label is "00C7000F104C00BE00610000318F00FFF906FF60BD00000014403780E600F000";
    attribute INIT_10 of inst : label is "FF000000FFFF0000FFFF000000FF00005FC0FF00FFD5FFFF57FFFFFF03F500FF";
    attribute INIT_11 of inst : label is "010000C00040030030903060060C090CFC0000000FFF000001E00A0000000000";
    attribute INIT_12 of inst : label is "AEA802C02ABA038040008000000100025E805E805E805E8030E420831B0CC208";
    attribute INIT_13 of inst : label is "0000FF000000003FAAAE550C2EAA0C150000005500001540CC00CCCC000C0CCC";
    attribute INIT_14 of inst : label is "0000C0F000000FFCD0003FD000010FFFFC00A000000F0002FFC0FF0000FF003F";
    attribute INIT_15 of inst : label is "3000FE00001E0002D4001500030A00690000000000000078735000000D0F0000";
    attribute INIT_16 of inst : label is "CE00800000400003FFFF0000000A00022A00640000C001E20000AA800000000E";
    attribute INIT_17 of inst : label is "000000000003000000000000000000000D00800001C4000B0000000000000000";
    attribute INIT_18 of inst : label is "84007800007A0085C000000000FF0000F000F800007F001F0180800009000009";
    attribute INIT_19 of inst : label is "D1D0000001F30000C0000000000000005000E4C0000100C6F040000000C10000";
    attribute INIT_1A of inst : label is "E2F88E103FF332B70000555000040557FFFC08BC3FFF1EE8800055500001055D";
    attribute INIT_1B of inst : label is "DF03FFD7C3DFD7FF68030CA7C009C009DF03FFD7C3DFD7FF00030003DF40C001";
    attribute INIT_1C of inst : label is "7F55FAAE05551FFF000095803F003F0C0098009C000000003F003F00004000C4";
    attribute INIT_1D of inst : label is "00009580000000000034024303240034FFF8A800FD79AAAA2FFF002AFFD0BFF4";
    attribute INIT_1E of inst : label is "000000000000000000000000000000005555000055FD00005555000000000074";
    attribute INIT_1F of inst : label is "000000000FFC0FC057F000007D7F0BC017F5030A000000000000000000000000";
    attribute INIT_20 of inst : label is "3F5F000000010000F5F507007F500F8000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "000F2F4700170000FC00747EF50000001F5F000000010000F57D07007F503E00";
    attribute INIT_22 of inst : label is "000003BB000900000000FBB058000000000000FB000900000000FBC058000000";
    attribute INIT_23 of inst : label is "0011002B010900335150FA00581073700000002B010900000000FA0058100000";
    attribute INIT_24 of inst : label is "0151002B010901735150FA00581073700151002B010903535150FA0058107370";
    attribute INIT_25 of inst : label is "0151002B010901735150FA00581073700111002B010900335150FA0058107370";
    attribute INIT_26 of inst : label is "0151002B010900335150FA00581073700151002B010903735150FA0058107370";
    attribute INIT_27 of inst : label is "0151002B010900335150FA00581073700151002B010903735150FA0058107370";
    attribute INIT_28 of inst : label is "282F007D025F0007FE0ADF40FD6080000454002B01090CDC5454FA005810DCDC";
    attribute INIT_29 of inst : label is "00A200070025001EFE28DDD0FFD680000282000700250007FF8ADDF4FFD68000";
    attribute INIT_2A of inst : label is "000F2F7D025F00007C00DF7EFD60BD80002F147D025F0000FE00DF45FD60B400";
    attribute INIT_2B of inst : label is "000100000000001FD0702E800000FA900038000A0000001F0B00E8000000BD00";
    attribute INIT_2C of inst : label is "000100000000001FD0706B800000FAD0000100000000017FD0702B800000AAD0";
    attribute INIT_2D of inst : label is "0BB400100000001E0720C1000000AD00003400100000000A0700C1000000E800";
    attribute INIT_2E of inst : label is "0035000300000009D700F000000058000038010A0000003A0B74E8000000BD00";
    attribute INIT_2F of inst : label is "0BBD000F0000000B5F20FC000000F800000D0030000000001C00C3000000C000";
    attribute INIT_30 of inst : label is "0282000700010007FF8ADDF4D5508000282F007D001D0007FE0ADF4055008000";
    attribute INIT_31 of inst : label is "002F147D00150000FE00DF455D00B40000A200070001001EFE28DDD0D5508000";
    attribute INIT_32 of inst : label is "00000008004000000000020040400000000F2F7D001500007C00DF7E5D00BD80";
    attribute INIT_33 of inst : label is "0000000300030000000082C00CC000000000000E0290000000000B0030C00000";
    attribute INIT_34 of inst : label is "00000080004C0000000020001000000000000000000000000000802011810000";
    attribute INIT_35 of inst : label is "0000002000320000000008000C00000000000020003000000000080086000000";
    attribute INIT_36 of inst : label is "000000380033000000002C000C000000001400C0000000001400C60000000000";
    attribute INIT_37 of inst : label is "282F007D00000007FE0ADF40800080000C340000000000550400000000000A00";
    attribute INIT_38 of inst : label is "00A200070000001EFE28DDD0080080000282000700000007FF8ADDF408008000";
    attribute INIT_39 of inst : label is "000F2F7D000000007C00DF7E8000BD80002F147D00000000FE00DF458000B400";
    attribute INIT_3A of inst : label is "BBE00030000000732FD01800000040087BC000300000001C0FBC30000000D000";
    attribute INIT_3B of inst : label is "2BC04090000000070FB4300000003400BBC00030000000280FAB30000000A000";
    attribute INIT_3C of inst : label is "FBC000300000001C0FB830380000D0007BF00030000000703FAC300000003400";
    attribute INIT_3D of inst : label is "2BD0F030000000A01FA0301300002800AB80DC300000001C0BAD30050000D000";
    attribute INIT_3E of inst : label is "303AD0E0002C0000E8002BBC140100007BC00035000000180FBC700000009000";
    attribute INIT_3F of inst : label is "C300C30FC955955509C390C35503555F0000FF553CD5000000000AA8C03C0000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0000AFC00FC00FC00000AAAA000003FA00030003C000C00000000EEC00000000";
    attribute INIT_01 of inst : label is "03F0FA0003F003F00000FFFF0FC000AFFFFF0003FFFFC00033F30A00FFFF0000";
    attribute INIT_02 of inst : label is "AAAAAAAAEAAAAAAAD555D55503FE03EA000000070000000000000000FFFC0000";
    attribute INIT_03 of inst : label is "EAABC003AAABAAAA55575557BFC0ABC00000D00000000000000000003FFF0000";
    attribute INIT_04 of inst : label is "004000000000000000000000000000000000000000000000004000C000000000";
    attribute INIT_05 of inst : label is "000000000000000000000AA800000000FF00E00000FF000B0000000000000000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0000000000402AFE10412BFA00402FEAFFFFE00B0000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C943";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "000000004000C0004001FFFF4001C00300010003155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "C000E60800000006E6A40C9005A60318C300E41800C00296C000C00000000000";
    attribute INIT_0D of inst : label is "0900000000180000FFFFC000F831F75D0AA0000000A80000E480093006260C18";
    attribute INIT_0E of inst : label is "FFFF030FFFFF000900110549003F00FFFC00FF004410B210FFFF6000FFFFE490";
    attribute INIT_0F of inst : label is "09C30033020D094D00060018FFFF093FFFFFFC98D00008008030F018D260D800";
    attribute INIT_10 of inst : label is "FF00AA00FFFFAAAAFFFFAAAA00FF00AA0040FF805400FFFF0015FFFF010002FF";
    attribute INIT_11 of inst : label is "20805740020801D5B5003030005E0C0CFC00FC00057F0FFF005007C000000000";
    attribute INIT_12 of inst : label is "00000B00000000E00000F0000000000F0AD6805E8AD4805EB54030C9015E630C";
    attribute INIT_13 of inst : label is "0000FC000000000FFFFF000C3FFF0C00CCCC00000CCC0000C000CCC0000000CC";
    attribute INIT_14 of inst : label is "FFF040300FFF0FDCF8000140000B0000FC00F000000F0003FFC0FF0000FF003F";
    attribute INIT_15 of inst : label is "C8007500038000010000400001BD02410000FD00000000070000F3F000000FFF";
    attribute INIT_16 of inst : label is "4000CC00000101CF00000FF00010000155408000006B00260000550000000000";
    attribute INIT_17 of inst : label is "0000000000030002FFC000000FFF00000000CF30000000CF0000000000000000";
    attribute INIT_18 of inst : label is "8000A800000A0057000000000015002A80001400000A00A80018180010000090";
    attribute INIT_19 of inst : label is "C00082E0004102C0C200C000002000000000C2E0000002E04000A3F0000002F0";
    attribute INIT_1A of inst : label is "FBD0E3E007FB3BD00000000000810210FFD09FFC07FF3FF80000200000100080";
    attribute INIT_1B of inst : label is "C50BF7C3C00EC37DAAAB2503EAFEC009C503FFC3C00FC3FFAAAB0003EAAAEF80";
    attribute INIT_1C of inst : label is "2F00FFFF002207FF000000183F003F0103030070000000003F003F00000C0030";
    attribute INIT_1D of inst : label is "000000180000000000CC018C0010009C3FFC7FE0F72EF7DF3FFF0BFFFFC0FFD0";
    attribute INIT_1E of inst : label is "000000000000000000000000000000000000AAAA03FFAAAA0000AAAA00000000";
    attribute INIT_1F of inst : label is "000000000FFE0FEA000002A007C107F800C007FD000000000000000000000000";
    attribute INIT_20 of inst : label is "0001000000002A005340EB400C00BF4000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0282140D0000003EE0A0DC05C000AF000001000000002A0252D0EB400C00FD00";
    attribute INIT_22 of inst : label is "0000005700000000C000F540000000000380001700000000C0B0F50000000000";
    attribute INIT_23 of inst : label is "000002F700000033C000F7E000003330000002F700000000C000F7E000000000";
    attribute INIT_24 of inst : label is "000002F700000173C000F7E000003330000002F700000173C000F7E000003330";
    attribute INIT_25 of inst : label is "000002F700000353C000F7E000003330000002F700000373C000F7E000003330";
    attribute INIT_26 of inst : label is "000002F700000033C000F7E000003330000002F700000353C000F7E000003330";
    attribute INIT_27 of inst : label is "000002F700000373C000F7E000003330000002F700000373C000F7E000003330";
    attribute INIT_28 of inst : label is "1FB6001E0007000367BDED007400F000000002F700000CCCC000F7E00000CCCC";
    attribute INIT_29 of inst : label is "007B000100000001D7B4EEC07740F800017B000100000000DAEDEED07740F800";
    attribute INIT_2A of inst : label is "02BE3D1E000700032FA0ED1F7400F0003EBF001E000700033FAFED007400F000";
    attribute INIT_2B of inst : label is "00000000000000035D7005000000FFC0003500010000002DD700500000005E00";
    attribute INIT_2C of inst : label is "0000000000000003D75005000000FFC00000000000000007D75005000000FFC0";
    attribute INIT_2D of inst : label is "013E00070000000FAF74F4000000FC00003E00070000002FAF00F4000000FE00";
    attribute INIT_2E of inst : label is "000A000000000038E800C00000000B000BB500010000000DD700500000005E20";
    attribute INIT_2F of inst : label is "0138002D000000200B745E000000C200003E000700000003AF00F4000000F000";
    attribute INIT_30 of inst : label is "017B000100290000DAEDEED00000F8001FB6001E0290000367BDED000000F000";
    attribute INIT_31 of inst : label is "3EBF001E000000033FAFED0001A0F000007B000100290001D7B4EEC00000F800";
    attribute INIT_32 of inst : label is "000E0024000000000B0030C00000000002BE3D1E000000032FA0ED1F01A0F000";
    attribute INIT_33 of inst : label is "0000000200000000000000800400000000000008000000000000020041000000";
    attribute INIT_34 of inst : label is "00E000CC00000000B0003000000000000000000000000000E0B0C30600000000";
    attribute INIT_35 of inst : label is "00000014001300000000140024000000000000140040000000001400C0400000";
    attribute INIT_36 of inst : label is "0000002000000000000008004000000000320041000000200C00010000000800";
    attribute INIT_37 of inst : label is "1FB6001E0000000367BDED000000F00000000000000002500000000000002860";
    attribute INIT_38 of inst : label is "007B000100000001D7B4EEC00000F800017B000100000000DAEDEED00000F800";
    attribute INIT_39 of inst : label is "02BE3D1E000000032FA0ED1F0000F0003EBF001E000000033FAFED000000F000";
    attribute INIT_3A of inst : label is "507F0004000022D5F400000000005E34007A00100000B2D5B400100000005E30";
    attribute INIT_3B of inst : label is "F07A0000000002FFB40040000000FE38507F0010000002FFF41410000000FE00";
    attribute INIT_3C of inst : label is "CC7A00400000C2D5B4350C0000005E00007A00300000D2F5B400300000007E38";
    attribute INIT_3D of inst : label is "B07A4000000002FDB43700000000FE00C07A4004000002D5B40C400000005E02";
    attribute INIT_3E of inst : label is "BAD5001D00000170570A70070000240005E00010000030AE2D4010000000E830";
    attribute INIT_3F of inst : label is "C309C390FAAAC0AAF0C300C3AAA9AA93FFFF28EABE3A0000FF55CC3CC2BE0000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFF03FFFFC0FFC0FFFF0000FFFFFFC000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "5FFFFFFF03FF03FF5555FFFFFFF5FFFF00000000000000000000000000000000";
    attribute INIT_02 of inst : label is "FFFFFFFF3FFFFFFFC000C0000003003F01FE00000007001F0003000300030003";
    attribute INIT_03 of inst : label is "C003D557FFFCFFFF00030003C000FC00BF400000D000F400C000C000C000C000";
    attribute INIT_04 of inst : label is "018000000000FFF5FFF5FFFFFFFFFFFF5FFFFFFF00005FFF03F0004000000000";
    attribute INIT_05 of inst : label is "FD00FFFD000003C000000000007F7FFF00000000000000000000000000000000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0000000000F400E009D818C907C002C000000000014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC0032558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "00001555C000C000C003C003C003C00300030003201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "0050FA9401A405ABFA400C00006B00300C00FA800424010B0000064000000040";
    attribute INIT_0D of inst : label is "00C0000000C00000C000C000F936AAAA0000000000000000FA40180001AB000A";
    attribute INIT_0E of inst : label is "6A6498302A51000001DF01F6000000000000000017409F8045A800001929090E";
    attribute INIT_0F of inst : label is "00C4000C10B4025000FF000F31800000090600606600F00074C00B0026003000";
    attribute INIT_10 of inst : label is "AAC000C0AA2A0000A8AA000003AA0300FFC0FFFDBFFFFFFFFFFEFFFF03FF7FFF";
    attribute INIT_11 of inst : label is "ABA000C00AEA030030903060060C090CC30000C000FF0C0001F85FC000001F55";
    attribute INIT_12 of inst : label is "AEA802C02ABA0380FF00FFC000FF03FFA17FA17FA17FA17F0000155000000554";
    attribute INIT_13 of inst : label is "5400BFC0000500FF557FAAFF3F553FEAFFFFFFFF3FFF3FFF0000000000000000";
    attribute INIT_14 of inst : label is "AAEC38CC3AAA3FC0D00C33DC30013555FF00FC00003F000F3FF0FFC003FF00FF";
    attribute INIT_15 of inst : label is "30000000001E0000FE001500030A00690000FE000000007F471CAAAC310F3AAA";
    attribute INIT_16 of inst : label is "30C030C00C300C31FFFF300C000A00002A00640000C001E20000FF800000000F";
    attribute INIT_17 of inst : label is "0000FC00000000FFE800000000AF000330C030C00D700C319400C300005B030C";
    attribute INIT_18 of inst : label is "8B007F0003FA0345FB00030003FF03008B005F0003FA03410000000000000000";
    attribute INIT_19 of inst : label is "9140C0C0013000C00000F40000000007D0C0000000C100009040C0C000C100C0";
    attribute INIT_1A of inst : label is "9FF461F033DC1948001A08000004000223CCF7242DB01C17801A080000010008";
    attribute INIT_1B of inst : label is "FFFCAAA83FFF2AAA97FCF3583FF63FF7FFFCAAA83FFF2AAAFFFCFFFC20BF3FFF";
    attribute INIT_1C of inst : label is "FF55FAA2057F1FFF000200003F003F0000001400000000083F003F0000000000";
    attribute INIT_1D of inst : label is "000000000010000200001400000000003FF8A80DF206AAAA2FFF702A5550BFF4";
    attribute INIT_1E of inst : label is "FFF0FFF0FFF8FFE001F000D00F400700555503D055550000555507C000300020";
    attribute INIT_1F of inst : label is "FFA0FFFE0003003F17F000004500002B000002FFFFFFFFFFFFFF002A2AFF0000";
    attribute INIT_20 of inst : label is "3F5087FFB50000030145FA000000A00000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "2FC0303B0000009C00FE7B0300000D00BF507FFF0000000E0151FA0000008000";
    attribute INIT_22 of inst : label is "000003BB000900000000FBB058000000000000FB000900000000FBC058000000";
    attribute INIT_23 of inst : label is "0000002B010900000000FA00581000000000002B010900000000FA0058100000";
    attribute INIT_24 of inst : label is "0000002B010900000000FA00581000000000002B010900000000FA0058100000";
    attribute INIT_25 of inst : label is "0000002B010900000000FA00581000000000002B010900000000FA0058100000";
    attribute INIT_26 of inst : label is "0000002B010900000000FA00581000000000002B010900000000FA0058100000";
    attribute INIT_27 of inst : label is "0000002B010900000000FA00581000000000002B010900000000FA0058100000";
    attribute INIT_28 of inst : label is "00000000025F000000000000FD6000000000002B010900000000FA0058100000";
    attribute INIT_29 of inst : label is "000000000025000000000000FFD60000000000000025000000000000FFD60000";
    attribute INIT_2A of inst : label is "00000000025F000000000000FD60000000000000025F000000000000FD600000";
    attribute INIT_2B of inst : label is "000100000000001FD2707FC00000FA900038000F0000001F8B00FC000000BD00";
    attribute INIT_2C of inst : label is "000100000000001FD2707FD00000FAD0000100000000017FD8703FD00000AAD0";
    attribute INIT_2D of inst : label is "0BB4001E0000001E4720ED000000AD000034001E0000000A0700ED000000E800";
    attribute INIT_2E of inst : label is "003D000300000009DF00F0000000D8000038010F0000003A0B74FC000000BD00";
    attribute INIT_2F of inst : label is "0BBD000F0000000B5F20FC000000F800000D003D00000000DC00DF000000C000";
    attribute INIT_30 of inst : label is "000000000001000000000000FFD0000000000000001F000000000000FD000000";
    attribute INIT_31 of inst : label is "00000000001F000000000000FD000000000000000001000000000000FFD00000";
    attribute INIT_32 of inst : label is "000B0009004007AFAE00F6004040E00000000000001F000000000000FD000000";
    attribute INIT_33 of inst : label is "0ABF000000030000D7003C000CC0000000030000029007A05C00F00030C00000";
    attribute INIT_34 of inst : label is "00BA009F004C000AE78060001000800002B4000000000002BAE09F601181FE00";
    attribute INIT_35 of inst : label is "022F001700330000FDD0D4004C00D0000BAF001700310007F880D400C6000000";
    attribute INIT_36 of inst : label is "032D00030033000078C0C0000C00C000002B00C70003000BE800D6000000E000";
    attribute INIT_37 of inst : label is "00000000005F000000000000FD4000000C030BBE00000057E800B0105F808A00";
    attribute INIT_38 of inst : label is "000000000005000000000000FFD40000000000000005000000000000FFD40000";
    attribute INIT_39 of inst : label is "00000000005F000000000000FD40000000000000005F000000000000FD400000";
    attribute INIT_3A of inst : label is "B80C0030003B007340D01800150040087808003000EC001C40BC3000EC00D000";
    attribute INIT_3B of inst : label is "280840900153000740B43000B0003400B808003000EC002840AB3000EC00A000";
    attribute INIT_3C of inst : label is "F808003003B0001C40B830383700D0007808003000DC007040AC3000DC003400";
    attribute INIT_3D of inst : label is "280CF030005400A080A0301354002800A808DC30003B001C40AD3005B000D000";
    attribute INIT_3E of inst : label is "3010D014002CDC00400040BC140102A0780C002000EC001800BC2000EC009000";
    attribute INIT_3F of inst : label is "C360C306C055F55500C3F0C3556355565454FF550000D4C0545500000000DC57";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFAFFFFFC0FFC0FFFFAAAAFFFFFFFA00000000000000000000000000000000";
    attribute INIT_01 of inst : label is "03FFFFFF03FF03FF0000FFFFFFC0FFFF00000000000000000000000000000000";
    attribute INIT_02 of inst : label is "FFFFFFFF3FFFFFFFEAAAEAAA0003003F003F0FF80003000F0003000300030003";
    attribute INIT_03 of inst : label is "EAABC003FFFCFFFFAAABAAABC000FC00FC002FF0C000F000C000C000C000C000";
    attribute INIT_04 of inst : label is "004000000000F500F500FFFFFFFFFFFF005FFFFF0000005F004000C000000000";
    attribute INIT_05 of inst : label is "D000FFD00000000000000AA8000707FF00000000000000000000000000000000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0000000000402AFE10412BFA00402FEA000000000000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C003";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "000000004000C0004001C0034001C00300010003155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "0000F60800000007F6A40C9005A703180300F41800C002970000000000000000";
    attribute INIT_0D of inst : label is "09000000001800000000C000F60EF5F50AA0000000A80000F480093006270C18";
    attribute INIT_0E of inst : label is "0000030C00000009006103F800000000000000000010AF000000600000002490";
    attribute INIT_0F of inst : label is "09C000300241093B03FF003F00000900000000986FC0F40010204E0812601800";
    attribute INIT_10 of inst : label is "FFC800C0FF3F0000FCFF000023FF030005F03F80FD407FFC017F3FFD0F5002FC";
    attribute INIT_11 of inst : label is "75D05740075D01D5B5003030005E0C0C038003002A800000005C07F000000000";
    attribute INIT_12 of inst : label is "F7C00B0003DF00E0D400FFC0001703FFF52B7FA1F52B7FA10000000000000000";
    attribute INIT_13 of inst : label is "0000FF000000003F55FFFFFF3FD53FFF0000FFFF00003FFF0000000000000000";
    attribute INIT_14 of inst : label is "C00C078C30003EC0F800ABEC000B3AAAFF00FC00003F000F2BF03FC003FA00FF";
    attribute INIT_15 of inst : label is "C800200003800000D400400001BF02410000FD0000000007AAACCF3C3AAA330F";
    attribute INIT_16 of inst : label is "30C030C00C300DB00000300C00100000FFC08000006B00260000550000000000";
    attribute INIT_17 of inst : label is "0000500000000015000000000000000330C030C00C300C300000490000010186";
    attribute INIT_18 of inst : label is "5500030001550300FB00FF0003FF03FF55000300015503000000000000000000";
    attribute INIT_19 of inst : label is "C0004240004102400000000000000000C0C082E000C002E04000633000000230";
    attribute INIT_1A of inst : label is "FFD01C9C07F706EF00000180008102103BD0639C07FB33870000218000100080";
    attribute INIT_1B of inst : label is "FFF4F7FC3FFE3F7D5554DAFC15013FF6FFFCF7FC3FFE3F7D5554FFFC1555107F";
    attribute INIT_1C of inst : label is "7F00FFFF825507FF001000003F003F0000000000001000003F003F0000000000";
    attribute INIT_1D of inst : label is "000400000000000000000000000000003FFC7FF4F001F5753FFF1FFF0000FFD0";
    attribute INIT_1E of inst : label is "FFC0FFFEFFFAFFFC00F003C00F0003C00000AFEA0000AAAA0000ABFA001000FC";
    attribute INIT_1F of inst : label is "FFF8FFF4000B00BFA80A02A0003E0000000007FD5555FFFF5555AFFFFFFF0002";
    attribute INIT_20 of inst : label is "7FA05FF400002A00AC00FF400000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "3D2D140D00000BC01E5FDC05000000F81FE8BF5000002A00AD00FF4000000000";
    attribute INIT_22 of inst : label is "0000005500000000C000D540000000000380001500000000C0B0D50000000000";
    attribute INIT_23 of inst : label is "000002F500000000C000D7E000000000000002F500000000C000D7E000000000";
    attribute INIT_24 of inst : label is "000002F500000000C000D7E000000000000002F500000000C000D7E000000000";
    attribute INIT_25 of inst : label is "000002F500000000C000D7E000000000000002F500000000C000D7E000000000";
    attribute INIT_26 of inst : label is "000002F500000000C000D7E000000000000002F500000000C000D7E000000000";
    attribute INIT_27 of inst : label is "000002F500000000C000D7E000000000000002F500000000C000D7E000000000";
    attribute INIT_28 of inst : label is "00000000000700000000000074000000000002F500000000C000D7E000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000007740000000000000000000000000000077400000";
    attribute INIT_2A of inst : label is "0000000000070000000000007400000000000000000700000000000074000000";
    attribute INIT_2B of inst : label is "0000000000000003DDF005000000FFC0003D00010000002DDF00500000005E00";
    attribute INIT_2C of inst : label is "0000000000000003F77005000000FFC00000000000000007F77005000000FFC0";
    attribute INIT_2D of inst : label is "013E00070000000FAF74F4000000FC00003E00070000002FEF00F4000000FE00";
    attribute INIT_2E of inst : label is "000F000000000038FC00C00000000B000BBD00010000000DDF0050000000DE20";
    attribute INIT_2F of inst : label is "0138002D0000002E8B745E000000EE00003E000700000003AF00F4000000F000";
    attribute INIT_30 of inst : label is "0000000000290000000000007F400000000000000297000000000000F4000000";
    attribute INIT_31 of inst : label is "000000000007000000000000F5A000000000000000290000000000007F400000";
    attribute INIT_32 of inst : label is "0000002400000053F00030C000005C00000000000007000000000000F5A00000";
    attribute INIT_33 of inst : label is "0002000200000002EB807D800400A800000B00090000005FAE00F6004100E000";
    attribute INIT_34 of inst : label is "000F00CC00000035004030000000FE00000000000000002F0F00C306000075C0";
    attribute INIT_35 of inst : label is "075C000B001300033000E0002400E080011C000B0040000B35D0E000C040C000";
    attribute INIT_36 of inst : label is "017E00270000020BBD40D8004000E080003F004300000017FC00C1000000D400";
    attribute INIT_37 of inst : label is "00000000000F000000000000FC000000001D01030000027F7FB8F8000000D060";
    attribute INIT_38 of inst : label is "000000000000000000000000FFC00000000000000000000000000000FFC00000";
    attribute INIT_39 of inst : label is "00000000000F000000000000FC00000000000000000F000000000000FC000000";
    attribute INIT_3A of inst : label is "5000002E000020000000370000008034000400B80000B0000000B80000008030";
    attribute INIT_3B of inst : label is "F0040372000000000000E00000000038500000B8000000000014B80000000000";
    attribute INIT_3C of inst : label is "CC0402E00000C00000350C0015008000000400300054D0000000300054008038";
    attribute INIT_3D of inst : label is "B00040DC000000004037DC0000000000C004402E00000000000CE00000008002";
    attribute INIT_3E of inst : label is "BA00000800005570800A2007000027B0040000B800003004C040B80000004030";
    attribute INIT_3F of inst : label is "C30FC3006AAAC6AA60C306C3AAAFAA03FFFF00000000D4DCFF5500000000CCD5";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
