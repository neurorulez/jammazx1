-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_7L is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_7L is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_7L_0 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"3571080A5A00A00003FF080A5000A0000078000003E02A0003D700AAD5C0BF80",
		INIT_02 => x"0355002ACD56A02000A5002A4D5CA0200005002AFFC0A0209573080A5FC0A800",
		INIT_03 => x"002A00FCA8000FF00002003CA0000F00000000FC000000F00000003C00000F00",
		INIT_04 => x"002A00FCA80000F00002003CA0000000000000FC000000F00000003C00000000",
		INIT_05 => x"002A00FCA8000AF00002003CA0000A00000000FC000000F00000003C00000A00",
		INIT_06 => x"000000070000FE000A0202C202800E00000000BF0000F840000000BF0000F800",
		INIT_07 => x"000000BF0000D000000000170000FE00000000170000FE00000000070000FE00",
		INIT_08 => x"288200FF0A28FC00000000BF0000D400000000BF0000D400000000BF0000D000",
		INIT_09 => x"000007FFAA08F8402A8006FF8000A00020AA012F0000FFD0000002D700005E00",
		INIT_0A => x"00000D0F0000E8FB00000D800020029B00000D0000032BF80002000B02A8BF90",
		INIT_0B => x"0000009E0000A03C0000380C00000F080000200C00000F020000000C00000F00",
		INIT_0C => x"000000BF0000F8400000003F0000E000000000BF0000F80000003C0A0000B600",
		INIT_0D => x"20000A8100084BFC00002FE80000001C04002FE810D02D5C00002FE800002D5C",
		INIT_0E => x"029500B4420001400295009048800180029505BC422000C0029500BC488800C0",
		INIT_0F => x"00000C2C0000B030000000000000000000000543000093F00000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000F000080000000CF570000A00F000003C000003D57000000000000003C",
		INIT_12 => x"BFBF0155BFB8550000003FFF0000FFF0028002EB0A00AE00000000BF0000F840",
		INIT_13 => x"0000000000000000000A3FFFA000003C00000000000000000000007F0000F400",
		INIT_14 => x"000E07E880000350000B03E880000300000A17E8C0000340002A57E8A0000354",
		INIT_15 => x"000A1FFAA0008FF4000A1FFFA000A8F4000A1FFFA000FA84000A0FFFA000FFA0",
		INIT_16 => x"000A0FFFA000FFA0000A08FFA000FFF0000A1A8FA000FFF4000A1FA8A000FFF4",
		INIT_17 => x"000A3FC0A000083C000A3FF0A000303C000A3FF8A000103C000A3FFEA000403C",
		INIT_18 => x"00001FFD0000557400001FFD0000557400001FFF0000557400001FFD00005574",
		INIT_19 => x"000A3FF8A000243C000000000000000000001FFD000055F400001FF5000057F4",
		INIT_1A => x"00003FF40000183C00003AFF000001AC000A003FA0000C00000A357FA000025C",
		INIT_1B => x"000A3F00A000C03C00023D07A000003C00003D7FA000040000023FF8A0000C0C",
		INIT_1C => x"000000FE0000FFFF0000007F0000FFFF0000007F0000FFFF0000003C0000FFFF",
		INIT_1D => x"00003CFF0000FFFF000000FF0000FFFF00003CFF0000FFFF000000FE0000FFFF",
		INIT_1E => x"0000FFFF0000FFFF00007FFF0000FFFF00007FFF0000FFFF00003C7F0000FFFF",
		INIT_1F => x"000044FE00000000000044FD000000000000447F000000000000447F00000000",
		INIT_20 => x"00000000000000C000550009054F00030000030000000000F150C00055006000",
		INIT_21 => x"0000000000026181150500004000010380000249000000000000C04054540000",
		INIT_22 => x"20005000800300005450000900000000C0030000000800140000000005156000",
		INIT_23 => x"20005000800300005400000000000000C0030000000800140000000000150000",
		INIT_24 => x"00000000000003AF00000000038100000000FEB0000000001080000000000000",
		INIT_25 => x"00000000000003AF0000000002EA00000000FEB0000000002AE0000000000000",
		INIT_26 => x"00000000000007F500000000000000000000D7F4000000000000000000000000",
		INIT_27 => x"00000000000007F500000000000000000000D7F4000000000000000000000000",
		INIT_28 => x"C3FFC3FFFF1F3FEAC000C0000000ABFFFFE38000FFFF00000000FFFF00ABFFFF",
		INIT_29 => x"C3FFC000FFFF0001C000C3FFFFFFE000FFFF557FFFFFFFFFFFFF0002FFFF0000",
		INIT_2A => x"FD0000000000000052BFFFFFD080FFFF0000000000007FFF00171300F00B0000",
		INIT_2B => x"FFFFFFFFFFFFFFFFA000000000000000FFEAFFFF0000FFFF00070000F0000A02",
		INIT_2C => x"00002D5E000002E000000B5F00003C0F00003D540000F2F400003C0F00003D54",
		INIT_2D => x"000BF0BDFFFF0000F0F07E070000E000FFFF0000E0007E0F0000000B0F0FD0BD",
		INIT_2E => x"00FF00FF00FF00FF00FF00FF00FFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_2F => x"0000000000000000FFFFFFFFFFFFFFFFFF00FF00FF00FF00FF00FFFFFF00FF00",
		INIT_30 => x"000000FF0000000000FF00FF00FF00FF00000000000000000000000000000000",
		INIT_31 => x"00000000000000000000000000000000000000000000FF00FF00FF00FF00FF00",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"00ABD000EFD0BFFFF000BFFFB00FFFFD0003402A42D00000FE00002F3FD0FFFF",
		INIT_35 => x"005FFFFFCF80EA00E003AFE0FEA8FFFF07F85FFF0FC0F87F000000000000AB00",
		INIT_36 => x"B330000F70A100003F0300FF5003FFC0FFFFFF01F800FFFFFFFF07FFF001FFFE",
		INIT_37 => x"20FC8F4334002D2C04C54B2214AA0A001420030A1C80F000FFF0AAAA1554BFFF",
		INIT_38 => x"15FFFFF8FFFF0000FFFF0001FFFFFFFFFFFF0015FFFFFFFFFF80FFFF0000FFFF",
		INIT_39 => x"02CF0000FFF000AA0000FFFA0800AAA0100001FD00000FFF0000000000000000",
		INIT_3A => x"FFFFFFFFFFFFFFFF0000A00015FF0000FFFFFFFFFFC3FFC3FFFF0000FFC30003",
		INIT_3B => x"0000FC7F002AFE000000000080000000FFFF1FFFFFC3FFC3000000007FC30003",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"000000070000FEFF00020000FFFFB400000CBFD000000290FFFE3C1F0000E000",
		INIT_3E => x"0000000000000004100100000402204080000080000020000800081002000000",
		INIT_3F => x"0000040100000004040000080000000008000010000000008001001000100000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7L_1 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"1AAE3FB0AA00300003EB3FB0AA0030002FE502574F9CD7C002B10303C280C3C0",
		INIT_02 => x"00EB0003FEAF0EFC00AA0003BAA40EFC00AA0003EBC00EFCFABF3FB0EB003000",
		INIT_03 => x"02FD02FD7F807ED000030014F000040000280055000052D00000001500005400",
		INIT_04 => x"02FD02FD7F807FD000030014F000050000280055000052D00000001500005500",
		INIT_05 => x"02FD02FD7F807ED000030004F000040000280055000052D00000000500005400",
		INIT_06 => x"3E01002FD000F54004050FEB4040AFC0AB4100D706F85C002F41009707F05800",
		INIT_07 => x"0007015F40BCF8000BF4002F0000F5400B80002F0000F5402F50002F0000F540",
		INIT_08 => x"3F0002C303F40E000000015F1FE0F8000000015F02E0F8000000015F05F8F800",
		INIT_09 => x"00000D7F00BFF000D5402FC310005800FE00002F0000FD7000AA2FC3A8000FE0",
		INIT_0A => x"000054FF0380FFB4000054FF0038F950000056FE000C55540004002501D7C3F8",
		INIT_0B => x"000005570020FD5400001EAF00005FA400001EAF20005FAD0000000730005F00",
		INIT_0C => x"AB4100C206F80C0000050275403CFE002F4100D707F05C000800157F0000D550",
		INIT_0D => x"27A01FFE0A98958402D00FFF0780800002D00FFF07C0C00002D00FFF0780C000",
		INIT_0E => x"002A000F8000D030002A005D81006070002A00558440A050002A004B8190E060",
		INIT_0F => x"00950600560002900000000000000000000F0002F000A1C00000000000000000",
		INIT_10 => x"0000000F0000C0000000CF000000F00F000003C000003C03000000020000D550",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"1FFF0000FFD40000002ABFFFA000FFF8BF410FFF07F8FFC0AB4100D706F85C00",
		INIT_13 => x"000000000000000000550FFFFF80C0300000000000000000BD0002C301F40E00",
		INIT_14 => x"083F0157F780000008BF01FFFB800000087F01FFF3800000083F01F5F3800080",
		INIT_15 => x"02FF07FFFF80FFD002FF07FFFF80FFD002FF07FFFF80FFD002FF07FFFF80FFD0",
		INIT_16 => x"02FF07FFFF80FFD002FF07FFFF80FFD002FF07FFFF80FFD002FF07FFFF80FFD0",
		INIT_17 => x"00550FFAFF80803000550FFFFF80C03000550FFFFF80803000550FFFFF80C030",
		INIT_18 => x"000006AB00008000000002AF00008000000002BE00008000000002FA00008000",
		INIT_19 => x"003505FFFC00C0500000000000000000000003EA00008080000007AA00008000",
		INIT_1A => x"00D40FF8BF80243000580FFD2F80603000700AFD1F80C1A00015002FFE00CC00",
		INIT_1B => x"001D0780F000C00000080400D000C80000000007D780C3000000001FF000D200",
		INIT_1C => x"0000005400005454000000540000545400000054000054540000005000005454",
		INIT_1D => x"0000505400005454000000540000545400005054000054540000005400005454",
		INIT_1E => x"0000545400005454000054540000545400005454000054540000505400005454",
		INIT_1F => x"0000005400000000000000400000000000000054000000000000005400000000",
		INIT_20 => x"000002A00200061300000090A48203030080C49000000A80821AC0C000000600",
		INIT_21 => x"06000542080384000000009020000801C0300012009085400008003000000600",
		INIT_22 => x"06000050400100000000000000000C0340000000009005000000C03000000000",
		INIT_23 => x"0600000040010000000000000000000040000000009000000000000000000000",
		INIT_24 => x"00000000000001F00000000002D500000000C3D00000000015F0000000000000",
		INIT_25 => x"00000000000001F00000000003400000000043D0000000000070000000000000",
		INIT_26 => x"000000000000007A00000000000000000000EB40000000000000000000000000",
		INIT_27 => x"000000000000007A00000000000000000000EB40000000000000000000000000",
		INIT_28 => x"C3FFC3FFFFCF0500C000E02F0000FFFFFFF000001FFF00000002FFFF954AFFFF",
		INIT_29 => x"C3FFC00AFFFFAA00C000C3FF3FFFF000FFFF0000FFFF0555FFFF0001FFFFC000",
		INIT_2A => x"50000000000002AFBFFDFFFF56FBFFFF0000400000023FD4B007E000FA00000B",
		INIT_2B => x"FFFF5FFFFFFFFFFFF400000000000000FFFFFFFFFA80FFFF00010000F8003F03",
		INIT_2C => x"00003C0F00002F7E00003CAF00003D5F00003EA00000F5E800003EEF00003EA0",
		INIT_2D => x"00BDF0F000000000F0F007E000007FFF000000007E000F0F0000FFFD0F0F0BD0",
		INIT_2E => x"00FF00FF00FF00FF00FF00FF00FFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_2F => x"0000000000000000FFFFFFFFFFFFFFFFFF00FF00FF00FF00FF00FFFFFF00FF00",
		INIT_30 => x"000000FF0000000000FF00FF00FF00FF00000000000000000000000000000000",
		INIT_31 => x"00000000000000000000000000000000000000000000FF00FF00FF00FF00FF00",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"AF7F0004F4007FF4000BFFFFFEAAFFF0A008081D2F4002FDA80000BFA140FFFF",
		INIT_35 => x"0001FFFF4FFEFFFAF803FFF8FFFC5500007C817F2FF0FF8707FF002FFAAA5B80",
		INIT_36 => x"53380F0F001C8040150A00FFBC00FFF01FFFFFE0FFE01FFFFFFF01FFFE00FFFF",
		INIT_37 => x"3C70E102B080D2FCA065030E5550604002FC01C500C040000000057F0000FFFF",
		INIT_38 => x"0005FFFF7FFFE8001FFFE000FFFF1FFFFFFF0000FFFF057FFFFEFFFF0000FFFF",
		INIT_39 => x"2FCF00A8FD507FFF0000FFFF0F80FFFF00000050000003FF0000FFFA0000AAA0",
		INIT_3A => x"FFFFFFFFFFFFFFFF0000FFA000050000FFFFFFFFFFC3FFC37FFF0000FFC3000B",
		INIT_3B => x"00AAFC15D07F55400000000020000000FFFF07FFFFC3FFC30000000007C30003",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"2800000000E07FFF02B500005FFFD000003CFFEA0000F400FF5F0C00E0007C00",
		INIT_3E => x"0000001000800801020800010000000002000000000000008004402000200000",
		INIT_3F => x"0000000000000000000000000100040800000000000004000100020100000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7L_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"0FAA1FED6800140003AA1FED6800100008240383303069C00C3C01EB30709440",
		INIT_02 => x"00290011AAC07BF400290011AAF07BF400290001AAC07BF403AA1FED68001400",
		INIT_03 => x"00FD007F5EF0FD00003C00000E00000000FD000050F02D00003D00005E000000",
		INIT_04 => x"00FD007F55F0FD00003C00000500000000FD000050F02D00003D000055000000",
		INIT_05 => x"00FD007F5EF0FD00002C00000E00000000FD000050F02D00002D00005E000000",
		INIT_06 => x"07EA00BFA800F8800055041F5400D0403FAA0BC3ABF40F8017AA0BC3AB500F80",
		INIT_07 => x"002A022FABD0FF0007D000FFAA00F88003EA00BFA800F8801F0200BFAA00F880",
		INIT_08 => x"0F550FEB57D0AFC000AA022F05D0FF00002A022FABC0FF0000AA022F80F4FF00",
		INIT_09 => x"005E0C3FABDDFC00C2AAFFEBA0000E0077EA00FFB500FC3000003FFF0000FFF8",
		INIT_0A => x"E000005501A05554E000007F00C6FFE8E00001FF0033FA80000A00B0AA83EBFF",
		INIT_0B => x"080002410080FFA00000055070000154000001507000015000001EB4700007AD",
		INIT_0C => x"3FAA0BC3ABF40F80002A0F30ABF4FFC0052A0BC3A1400F8002000AFF00204180",
		INIT_0D => x"01C207FF83E0EE40000101FF4BF8C00008EB01FFEBF8C00008EB01FFEBF8C000",
		INIT_0E => x"1A030000CC001F0830000000CC005D0C10030000C400558C10030000C8004B84",
		INIT_0F => x"09AF006AFA60A90000000000000000000387000FD000F0000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000A80F0000C00000000FAB0000D2AF0000ABEA000007AD000000010000EAB4",
		INIT_12 => x"011400004500000002C37DF70E00DDF441AA047FA904F4403FAA0BC3ABF40F80",
		INIT_13 => x"0000000000000000000001FF07F0F0000000000000000000742A0FEBA050AFC0",
		INIT_14 => x"0E5F0015DBC006000E1F0015DBC000000E1F0015DFC000000E3F0015FBC00010",
		INIT_15 => x"0FD5005F5FF0F5000FFD005F55F0F5000FFF005FD550F5000FFF005FFD50F500",
		INIT_16 => x"0FFF005FFD50F50005FF005FFFD0F500055F005FFFF0F5000D55005FFFF0F500",
		INIT_17 => x"000801FF87F0F000000001FF07F0F000000001FF07F0F000000001FF07F0F000",
		INIT_18 => x"2D00005F0000F000000B005F4000F0000000005F02D0F0002D00005F0000F000",
		INIT_19 => x"0A02000F8780FC000000000000000000000B005F4000F0000000005F02D0F000",
		INIT_1A => x"0030007F0C00B000058101F047500C00001801F427F01800002400FF1FF0F100",
		INIT_1B => x"0090007F0600F0000A90000B6000FC00069300030070F0400A96000B86A0F100",
		INIT_1C => x"002A00002A2A0000002A00002A2A0000002A00002A2A0000002A00002A2A0000",
		INIT_1D => x"2A2A00002A2A0000002A00002A2A00002A2A00002A2A0000002A00002A2A0000",
		INIT_1E => x"2A2A00002A2A00002A2A00002A2A00002A2A00002A2A00002A2A00002A2A0000",
		INIT_1F => x"222A0000000000002202000000000000222A000000000000222A000000000000",
		INIT_20 => x"00600000030358410150000009230100C0C0412509000000C860004005400000",
		INIT_21 => x"006000000C00100002A1090048000C0380100004090000000021C01042A00060",
		INIT_22 => x"000000000C03000000A0090000000002C030000000000000000080020A000060",
		INIT_23 => x"0000000000000000000009000000000200000000000000000000800200000060",
		INIT_24 => x"000000000000003A000000000FE000000000EB000000000082F8000000000000",
		INIT_25 => x"000000000000003A00000000080B00000000EB0000000000F800000000000000",
		INIT_26 => x"0000000000002F9F00000000000000000000FDBE000000000000000000000000",
		INIT_27 => x"0000000000002E1F00000000000000000000FD2E000000000000000000000000",
		INIT_28 => x"C3FFC100F5430000C000380500005555FFFC000001FF00000AAA5555AFFF5555",
		INIT_29 => x"C3FFC003FFFFFFFFC3FFC3FF0000FC00FFFFFAA8FFFF00000000000000004AAA",
		INIT_2A => x"500000020000B874FFFF5555EA8F5555000000020ABF8400F400000050000015",
		INIT_2B => x"FFFF0000FFFF00000000A00000000000FFFF0000FFFE003F00000000000C3FCB",
		INIT_2C => x"00003C0F00003C0F00001E0000001E2D00003C000000F03C00003F7F00003C00",
		INIT_2D => x"0BD0F0F0BFFF0000F0F0007E00000000FFFE000007E00F0F000000000F0FBD00",
		INIT_2E => x"00FF00FF00FF00FF00FF00000000000000000000000000000000000000000000",
		INIT_2F => x"00000000000000000000000000000000FF00FF00FF00FF0000000000FF000000",
		INIT_30 => x"00FF00FFFFFF00FF00FF00FF00FF00FFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_31 => x"FFFFFFFFFFFFFFFF0000000000000000FFFFFF00FF00FF00FF00FF00FF00FF00",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"FF3D0000002F1F4000BF5555FFFF5540F03C2C007D0C0BFCF0030055FFFF5555",
		INIT_35 => x"A000C0FF05FF555F000055000000000AE000FEA51FFCFFF8000080020AAAFF40",
		INIT_36 => x"011C0F0F0007C003C0FF0055FF00555081FFFFF8FFFF01FF3FFF0055FF805555",
		INIT_37 => x"0F305001D2E02FDA18753307555F8E0011FD0040017F0080FFFEF80101555FFF",
		INIT_38 => x"8000FFFF015FFFE801FF5000FFFF0155FFFF0000FFFF0001FFFF5555F8005555",
		INIT_39 => x"A1C5F81C40001FFF5554FFFF0000FFFF0000C00400AA015017FFFFFFF4BFFFFF",
		INIT_3A => x"FFFF5FFFFFFFFFFF0000555500000000FFFFFFFFFFC3FFC3015F0000FFC3002C",
		INIT_3B => x"FFFF0000800F0000FFE0FFFA001FAAA0FFFF007FFFC3FFC3FFF8000000030003",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"07A0057F00F8FFFF000000030FF7400000F0FFFF00004000FFE0000015A00780",
		INIT_3E => x"0000000100010000000000000010040400081010040040000200800000000000",
		INIT_3F => x"0000000441010040008100000800000004100404200000000204001000400000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7L_3 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"016A0154C0000000017A0154C000000001C2007FAE40C00001C20015AE004000",
		INIT_02 => x"00030000AD40154000030000A940154000030000AD401540017A0154C0000000",
		INIT_03 => x"00FE0000ADF00000003C00000D00000000FE0000A0F00000003E0000AD000000",
		INIT_04 => x"00FE0000A8F00000003C00000800000000FE0000A0F00000003E0000A8000000",
		INIT_05 => x"00FA0000ADF00000000800000D00000000FA0000A0F00000000A0000AD000000",
		INIT_06 => x"000000D70000FD0000FF0000FC0000000F000D7F03F0F5C000000D7F0000F5C0",
		INIT_07 => x"0000007F0000D70001E000D70000FD0000F800D72000FD00018000D72000FD00",
		INIT_08 => x"012A041FA100D0400000007F0A40D7000000007F2F00D7000000007F0240D700",
		INIT_09 => x"008A01FD84000400200041FF1400D70000120041A200FF4000BF1F7FF800F7D4",
		INIT_0A => x"380100005EE6000028010000556300002801005557C35555001400D70008FF41",
		INIT_0B => x"0180000055E05555200300003E000000000300003E000000000300403E000140",
		INIT_0C => x"0F000D7F03F0F5C000000D7F0140D04000000D7F0000F5C00B55555502400000",
		INIT_0D => x"0C7F007FD5FC540000000015007C000004170015C2FC000004170015C2FC0000",
		INIT_0E => x"050900000600005803C90000030000580A090000070000583C09000005000008",
		INIT_0F => x"0C1D00007030000000000000000000000FC1000042A000000000000000000000",
		INIT_10 => x"0005000000000000CF0B0000D00F000003C000003C03000000020000D5780000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"00000000000000000FEB0000AFC0000001020000010000000F000D7F03F0F5C0",
		INIT_13 => x"00000000000000002FA0000500FC40000000000000000000002A041FA000D040",
		INIT_14 => x"05EA0000FFE0004001FB0000BF00000025FE0000BFC00000A5FA0000BFE80000",
		INIT_15 => x"3FF000000FFC00003FFF000000FC00003FFF0000F00C00000FFF0000FF000000",
		INIT_16 => x"0FFF0000FF00000000FF0000FFF00000300F0000FFFC00003F000000FFFC0000",
		INIT_17 => x"2F80000518FC40002FA5000560FC40002FA1000580FC40002FA2000580FC4000",
		INIT_18 => x"FFC0000003FF0000FFC0000003FF0000FFC0000003FF0000FFC0000003FF0000",
		INIT_19 => x"2FA4000518FC40000000000000000000FFC0000003FF0000FFC0000003FF0000",
		INIT_1A => x"3AE20005818C4000001000000C00000025A10000405C00002FB8000424FC1000",
		INIT_1B => x"2F96000500FC50002FA0000506BC40002FA10005A2BC40002FA4000518FC4000",
		INIT_1C => x"007F0000FFFF0000007F0000FFFF000000FE0000FFFF0000007C0000FFFF0000",
		INIT_1D => x"7CFF0000FFFF000000FF0000FFFF00007CFF0000FFFF0000007F0000FFFF0000",
		INIT_1E => x"7FFF0000FFFF0000FEFF0000FFFF00007FFF0000FFFF00007CFE0000FFFF0000",
		INIT_1F => x"667F00000000000066BF000000000000667F00000000000066FE000000000000",
		INIT_20 => x"000600AA00030A8F0000000000C00000C000F2A09000AA000300000000000000",
		INIT_21 => x"00002A2A020300000000000092400001C08000020000A0A88186400000000000",
		INIT_22 => x"0006A8A000000000280010000000C0030000000090000A2A0000C001000A0004",
		INIT_23 => x"0000A80000000000280010000000C003000000000000002A0000C001000A0004",
		INIT_24 => x"000000000002001D0000000001500000A000DD00000000004154000000000000",
		INIT_25 => x"000000000002001F0000000005150000A000FD00000000001450000000000000",
		INIT_26 => x"000000000000050A000000000000000000006814000000000000000000000000",
		INIT_27 => x"00000000000007EA00000000000000000000EAF4000000000000000000000000",
		INIT_28 => x"C3FFC00050010000C00005EA002AAAAA5FFE000004000000FFFFAAAAFFFFAAAA",
		INIT_29 => x"C3FFC001FFFFFFFFC3FFC3FFC000FE2AFFFFFFFFFFFFFA800000AFCA0000BFFF",
		INIT_2A => x"00002A4B00008780FFFFAAAAFFCAAAAA0008002FFFFFC0007544AAAA0000AAAA",
		INIT_2B => x"FFFF0000FFFF00000000FC0000000000FFFF002AFFFFA0140000000000001500",
		INIT_2C => x"0000055400001405000001550000015000001554000055500000140500001554",
		INIT_2D => x"BD0BF0F0D0000000F07E00070000FFFF00070000E07E0F0F0000FFFFBD0FD000",
		INIT_2E => x"00FF00FF00FF00FF00FF00000000000000000000000000000000000000000000",
		INIT_2F => x"00000000000000000000000000000000FF00FF00FF00FF0000000000FF000000",
		INIT_30 => x"00FF00FFFFFF00FF00FF00FF00FF00FFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_31 => x"FFFFFFFFFFFFFFFF0000000000000000FFFFFF00FF00FF00FF00FF00FF00FF00",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"FC00200002FF04020BFFAAAAFFFFAAAAF010FC00103E2FF0400FAAAAFFFFAAAA",
		INIT_35 => x"FFA8803500150000000000000AAA0AFF55030C0081FF001500FF40075502F4A0",
		INIT_36 => x"000E3F030001F00700FFAAAAFF80AAAAF81FFFFFFFFF801F0FFFAAAAFFF0AAAA",
		INIT_37 => x"0F121CE6CB40F7BD6305033157AAE1000050000000377FF00005FFE82AA00017",
		INIT_38 => x"FE00FFFF0000FFFF001FAAAAFFFFAAAA57FFE000FFFF0000FFFFAAAAFFE0AAAA",
		INIT_39 => x"C100FFF4000005500000FFFF0000FFFF00AA0000CFFF00000015FFFF4055FFFF",
		INIT_3A => x"FFFF0057FFFFFFFF0000AAAA0000AAAAFFFFFFFFFFC3FFC30000AAAA57C3AB50",
		INIT_3B => x"FDFF0000F80100005550FFFF0005FFFFFFFF0007FFC3FFC35555FFFA0003AA83",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"007F000080FE5FFF000000003F4000000BF0FFF400000000F1FE000000000040",
		INIT_3E => x"0010004004000010004200000100000002001080000080408000000011000000",
		INIT_3F => x"0000000002002008000000000004000000000000000004008000400000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
