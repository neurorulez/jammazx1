-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D7AA183889EAAB2B0B8A02200A0946094690B3FFFFFE00A0C1FEA7A3D3F3EDB5";
    attribute INIT_01 of inst : label is "D973DA258046ED4C4322AEB3DFC9B54D4135AF7841AD814A2F549FA3CAFA0298";
    attribute INIT_02 of inst : label is "87E6CF07E79C96FD405406EDE5DAC8E6111E30028E1A003099FB0CCDB3B6007A";
    attribute INIT_03 of inst : label is "77CF921AE98012490000DD2B57F8747EE11FC54D2E9FC87CF72D3EE807D75DF7";
    attribute INIT_04 of inst : label is "299A9E0882A237FFD57F70C5549C679E89DBA312E20375533E87D85ACFC55CDF";
    attribute INIT_05 of inst : label is "7599DA40024800C0006934AEF8A2F081D28F35605B86B0000055EE638E1A70A4";
    attribute INIT_06 of inst : label is "ECE0004C00018001300006000CD25A5DF718A9938A605056AE03AF15D78AE3C4";
    attribute INIT_07 of inst : label is "0A0904124AFFF679F65B7274DF25A3BD3294BF7A7F0CB517C7C40DA458614BFC";
    attribute INIT_08 of inst : label is "A695050470071A8D518B5B42D16891B03F22209208010061A3ABFBFB57DDF3EF";
    attribute INIT_09 of inst : label is "28D94FEA365A3FDC80BC78061800100007C01002000D9007C3F9164A0E3366F1";
    attribute INIT_0A of inst : label is "DE8C902366C4D9E7532EF532E00403093108B820B1845F5F89050DEB5305111A";
    attribute INIT_0B of inst : label is "9E53EF95859300008190220E124D29BD20AADEB572514509570074424DE9DEDE";
    attribute INIT_0C of inst : label is "288E0840F2C33FFEDB6DB6D87FFC6318C3FFFFFE186185E7B9A55CB392440775";
    attribute INIT_0D of inst : label is "C37ECAF174DE84D1117117A67A45A6D04814538C7BF84D1348052000026A300B";
    attribute INIT_0E of inst : label is "4903B29233434350369BD37C8942A8007B5A346784AA97E908B5D725068812C9";
    attribute INIT_0F of inst : label is "3FFF6DB6DB6C3FFE318C61FFFFFF0C30C2F3C000000000000400154015122464";
    attribute INIT_10 of inst : label is "CFAEB48A908A53F3E534822905DE2D4140E1A2457326157C150B0593C750B059";
    attribute INIT_11 of inst : label is "90D113192740470C3084C755161108326EB3BB4B2FFFEDCFFE2A0200F082F20B";
    attribute INIT_12 of inst : label is "777B12EEED9BE589BE59484EA1674375571CB91898E93A8166A3B4375541CB91";
    attribute INIT_13 of inst : label is "3CC504034925F0348438BF05AB82807C8A274B3022677F3CDF0F0FCFBFBFBF88";
    attribute INIT_14 of inst : label is "5385F88724A041111F148D0220980C80D3052D984526E90624AA35705B2D8110";
    attribute INIT_15 of inst : label is "74954404A284209392E2A04B255599EECF8FE53A8B2BFCC7E95826B626B728FA";
    attribute INIT_16 of inst : label is "04909F7CB12201AA90805691E667979FACC64CF7709DCB9B964D453B8411C218";
    attribute INIT_17 of inst : label is "17450AAA3DD89DF435233A8A8E3968BFC7438F74265E3A76F01C2C1580B03002";
    attribute INIT_18 of inst : label is "8B55DA228262DA59227C79B100446339C81D110836A87BB84D10354541A6C451";
    attribute INIT_19 of inst : label is "5240662C98CD18C90C26508C220046E884A04801C70693A5324BC51493102558";
    attribute INIT_1A of inst : label is "D55FD5D23CF309B88A0A189A004460A649E86A933A8876E207870488C479D282";
    attribute INIT_1B of inst : label is "21EEC44D76B54949EF313FFB16FED33593B24CDF68E5A135722722A3F37FDF7F";
    attribute INIT_1C of inst : label is "1311276CA93B6504C1860048168F73DDDDBBBBBAEDF73BBBB8F7777DC6ECF762";
    attribute INIT_1D of inst : label is "3DDD67F8DE3DDD67FECD75634B5AADBC7972C89ED47BA6DFAB0C449DB2A4ED94";
    attribute INIT_1E of inst : label is "EECF3775D5575DCDB3BAEADE3DDD67F8DE3DDD67F8CEB9FC6FBACEB9FC6FBADE";
    attribute INIT_1F of inst : label is "A8D4681009AD88136E65FC9600E004164111B22AB0BF259F8F651CFBD4D9AABA";
    attribute INIT_20 of inst : label is "000000033CFAC8F3CFAC8EC96F1273CB8D8D8D8D8D8D868686868686E3636351";
    attribute INIT_21 of inst : label is "5E509B6DB036E65FF2E817E4A93E74A5D199AC92FC9E52FC0000000000000000";
    attribute INIT_22 of inst : label is "000000000000000000000000000000000000018F298E492164CC8B9BEC4F25BC";
    attribute INIT_23 of inst : label is "7BE9F9B89F33AA352CD6C97E4F297E0000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "71880182C0D881D34EAC0D33851739A2E41D7113A6FD5A800820299932209729";
    attribute INIT_25 of inst : label is "E01054604ED5CED40A8006829313FFA483296001A8D400C0B660549880F22201";
    attribute INIT_26 of inst : label is "B2BA4A8BC0D7B4E39878881BE6E2EC95EEC982ED7789B402D26A4983A001AC09";
    attribute INIT_27 of inst : label is "E9F423AAD4A19A83996664B996EAA22509AD3B649FBD9A779E5E5CD3923A7337";
    attribute INIT_28 of inst : label is "02A3DCB026AC53674B5294B5AD4A5294A5105B4D0167D44552C0A820220EA04B";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE9C3";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "E039483018CF3CB71F6D2B044364CF40EBC401FFFFF8592DCAFBCD6603E38D93";
    attribute INIT_01 of inst : label is "5B6376800C8C16048CBB3B4D65524C0159149507589D373770FFBFFE970964FD";
    attribute INIT_02 of inst : label is "2FD0A77414ED60818018022A1C5407AC96BF7CD330FC69C12B086CCEB3393669";
    attribute INIT_03 of inst : label is "460736880A20800000000544753F7E22C7AB348FFA364CF13468702AA1593411";
    attribute INIT_04 of inst : label is "492D83D7DDD7C2A88082808A31882FFE5BFB195C6B993FE7A434126223EF2140";
    attribute INIT_05 of inst : label is "B28039480150034001E21A1EF9034382E16819E03D8B5000000DDE4B905682E2";
    attribute INIT_06 of inst : label is "57E0002C00078003B0007E000AC46D3DB8199D3407601015E8259406DA036D00";
    attribute INIT_07 of inst : label is "D325B24001800081015C04596F4CD8C46E242CABFF2DEFBFCE76D28CC76C99BD";
    attribute INIT_08 of inst : label is "48075617017040975A19292B9DEE5377AC2FB920711B221AB01401092583679E";
    attribute INIT_09 of inst : label is "42A41400A00015F5FDCE8707E002077FF827E7FC380E07F8003A005BA17E3127";
    attribute INIT_0A of inst : label is "FE27FC8A033302015D9815D99911FEA0EBD6671607EB33E66C91BA4065767443";
    attribute INIT_0B of inst : label is "6878192D7B69000024C67FA1E5004010B7FE2406556468A67841387FF246BAFE";
    attribute INIT_0C of inst : label is "23712919CA6AFFFEDB6DB6D87FFC6318C3FFCF3C104104E38219F36CF82D104D";
    attribute INIT_0D of inst : label is "D0941F3680095C16A9EA9F1AACC80A0EB138E529480221A4332EC615E71E865C";
    attribute INIT_0E of inst : label is "C22E4B2592EAEAF58001002634EE43DB7F28858F91EEF985B806A55610D3345C";
    attribute INIT_0F of inst : label is "8000000000000000000000000000000000000000000000000480460102F0D5A5";
    attribute INIT_10 of inst : label is "5EBAA3115B4BFA17ADE0BC45BF2401D58BE8308BA172CB1F62097B69F22097B6";
    attribute INIT_11 of inst : label is "3516B6AF849AD54591AE08DA24BBAD77092D60109921946701CB67DA36181C20";
    attribute INIT_12 of inst : label is "0168A4021A208D6012A81A2477D8D448A4920225B57C2457D85A4D448A592022";
    attribute INIT_13 of inst : label is "902CABF02CCC66E7D17DC5B03E5F5D28A0A57AD68F4BB4894BABABDAD6D6D6D3";
    attribute INIT_14 of inst : label is "C8181651F7D531ECC84354BDC30B4476FAEF91E8F3902BA221D62A1A8090A5EC";
    attribute INIT_15 of inst : label is "7E526E1190AB72725EE690E773E165C087B7FDAA42C2045730C0DADA49C42423";
    attribute INIT_16 of inst : label is "05C7AD20725523B25AD898EA808164ACDB54021084415662ACF135C037DA7736";
    attribute INIT_17 of inst : label is "AE3AE67CA04C47DBB24A8331107785405C0EA8191146F8A7F59D40A01402C961";
    attribute INIT_18 of inst : label is "E4697554372736E00482FD4DD977B5228B622293DB7D480221A83D35E1F823AE";
    attribute INIT_19 of inst : label is "D4CD5000C2818122A910FED4184D6D01A2349801F801B687A9FD4FDEFADADACF";
    attribute INIT_1A of inst : label is "08D7F7BCAB43D3D2D0D0D9505B59109A538F547A4C133AC6FA248E329695A418";
    attribute INIT_1B of inst : label is "7B143AF01DEFEE9221064B180B3B66D924A49B6DB542D64208408C455D770222";
    attribute INIT_1C of inst : label is "2C59CAB6CAD5960B12C934B51935877D5F30414011A83AFBE98A8282AC518A1D";
    attribute INIT_1D of inst : label is "6B5EB52D4E7B9EB471201084F037EA7A83753109889C44268541372E59AB7248";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAADEFFFFBD6F5EEFBF9D6B4E7BDEB42D4C7B9AB5214E";
    attribute INIT_1F of inst : label is "05028133E0B96D689211320CB24B2CC421CCA66E66268324E748A84FB9680000";
    attribute INIT_20 of inst : label is "00000001746B1E1746B1E9B0DA64E5961010101010104848484848482424240A";
    attribute INIT_21 of inst : label is "A4E3410019892113689CC4D0140D096E22A601289A04A8980000000000000000";
    attribute INIT_22 of inst : label is "00000000000000000000000000000000000000D65B9A0A296AC71EB3FB2AC369";
    attribute INIT_23 of inst : label is "0B0ABAB70694445B7300844D02544C0000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "E92C5BC40063720406035002B8C02B181F13A6BC004C0053FEF77C3785A97640";
    attribute INIT_25 of inst : label is "570F771B2B0D0B0D99132E6AE28892BDB27B84CBC508F7BDC44CDE034BDEF7BA";
    attribute INIT_26 of inst : label is "9C0575F7E63FCF77D0FB961190D803E0101456B402601BAE800CA022C4CBCAB8";
    attribute INIT_27 of inst : label is "00D02FCF2DE89DAB43CD0F1438ECE5A34412142DA0E93094A1D2B00C06A18E69";
    attribute INIT_28 of inst : label is "16500233030E81D1DDF7BDFFFFDEFFB9CE7FB7DAAB8E4CDCF74E556856D0FC3D";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6127";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "E1B8403980A99427070B080A02484740085401BFFFF811D543F94D7719E99B81";
    attribute INIT_01 of inst : label is "03424A1008888A04203332150552C8C25000A21A508112214175C228550047ED";
    attribute INIT_02 of inst : label is "2FE4857482F5EA978060024EBC9D468090352093A6524D91AECB688922A63349";
    attribute INIT_03 of inst : label is "4450248288A400000000110B3042120A2480A5419834C9F535425A83E8044144";
    attribute INIT_04 of inst : label is "908B9AF75DFD57FFD7FF7782010C2B401BE0A85A2B690AA7ECB45A61FFFB0451";
    attribute INIT_05 of inst : label is "A180B2C0004002C0024CAB2833A84981F25EA8603515100000B0E843C93E49FC";
    attribute INIT_06 of inst : label is "CED000CA001B40046800C50010996450649CBB724ED0100389050C8286414320";
    attribute INIT_07 of inst : label is "0008241000FF969D977D5535DF7C71506C742D23FE2DE597CFA22E0DD77988B6";
    attribute INIT_08 of inst : label is "6E8150D3ED3EDA82500A49481C0E11CB8CA91C3239BFFE03300429E151CD6186";
    attribute INIT_09 of inst : label is "0A805402A00FC2008A04671F9802177FFC0217FE38F217FFC0021294A0373881";
    attribute INIT_0A of inst : label is "4547F42A03B43EF7FDA1FFDA1FE0854855FE820876FF43E676E1290801705840";
    attribute INIT_0B of inst : label is "05C3F7F35EB30000388023002140C81924A810801708002850FE32F7E1080101";
    attribute INIT_0C of inst : label is "4201BE11FDC280000000000000000000000000000000000003A14FD6B847E045";
    attribute INIT_0D of inst : label is "D0440F51C528069049E49FBC96DC9E10F92CB4A529720547400F07951483001E";
    attribute INIT_0E of inst : label is "63429201218989AD02819037252280485A0C940790EBF9892E80E170D0021458";
    attribute INIT_0F of inst : label is "20000000000000000000000000000000000000000000000000D0587F04E02435";
    attribute INIT_10 of inst : label is "5CF3F3C2524A5B173F72AF092511A05410E800E10362812A822B1EB2A220B1EB";
    attribute INIT_11 of inst : label is "6C141C8B950295451968215084150A440820B6DBF7DE7D46526A0210346A19E8";
    attribute INIT_12 of inst : label is "2219B4427B352D0A528892049124B05135548780E45CA8B1249A8B1513554878";
    attribute INIT_13 of inst : label is "04824904404F6786BA986BD429FFDD5FFDDB46948A507FF6D62626B64242425A";
    attribute INIT_14 of inst : label is "026B7C5086837F8682840408BC4EA404114AA12C558482E8E184EAD486A03787";
    attribute INIT_15 of inst : label is "09506F9D45EB7C719EA2AE8070694794C7BFFD229288DAD6118CFEFE6F55A977";
    attribute INIT_16 of inst : label is "7D063BE83429218A9488CEBA53A1B6F66FD204526409DBB3B7D9552AA451EB7F";
    attribute INIT_17 of inst : label is "4D7B06F690F50E6D26291199985AE56DD2C92437421FA1E4BDF540A09612F17D";
    attribute INIT_18 of inst : label is "2A41C2803487A6F5A6E16178C937D21A4A3337FB6EA929320543F9555F9006B0";
    attribute INIT_19 of inst : label is "D44D2BC68AE523A72502F087504F478520218F81FFE12496A1481954D290C05D";
    attribute INIT_1A of inst : label is "227DD7F691295342A0A0E42083419D9BC3EE705202737EB4FA3C6810841EE612";
    attribute INIT_1B of inst : label is "2DFE8057EF3AAFFBBDF7EAD75DADF36FF6FECDB6FD2767E337667776160002A8";
    attribute INIT_1C of inst : label is "7E79FFDFEFFEDF5F9AE9B5FD4F9FBAA80AFFFEABFFD5755156FFFD5FF7AAFF40";
    attribute INIT_1D of inst : label is "6749477CD25EC735839FE9C418BD5E0EA37C39F78CD664336641B7FBFD3FDF6D";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAAC463C84734824A4614AC1477496674D04EC315E416";
    attribute INIT_1F of inst : label is "01A044220D1D48B66E6CD9FEA2EA2D373489A286699B7FFE1AFF37B4EFB98000";
    attribute INIT_20 of inst : label is "BBBBBBB954DAD1154DAD181FF760E7DC1A081A081A080D04040D040D06820681";
    attribute INIT_21 of inst : label is "80F1B0410A66E6CDF6D5336FBB36E96F33B7FE366DFEF66FBBBBBBBBBBBBBBBB";
    attribute INIT_22 of inst : label is "777777777777777777777777777777777777769F72936BA92CAFD63BFF217FDD";
    attribute INIT_23 of inst : label is "2A21B2B19B77066B7BFF8B36FF7B377777777777777777777777777777777777";
    attribute INIT_24 of inst : label is "AD2C83F40C30FA14A642590AA850AB0A0BD101AC294C85535B777C53892B16A8";
    attribute INIT_25 of inst : label is "57DD069DEB14AB14A3E00C78F3AFEBEDAA738403F420FDBDC74046804BF6B6FA";
    attribute INIT_26 of inst : label is "188272EBE75FD7F5C0F9A7D0BCEA1DC43DF7AA3D0EA87D4250C8287AE403E10B";
    attribute INIT_27 of inst : label is "CA09AA2C00C3A80A4A012824A0A6CC334042360924C8A092B5CAC42E04A5CA2F";
    attribute INIT_28 of inst : label is "0410C600010081B39FE73BDE739CEF3DEF400390BF0848C9EFC4414004006E71";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4100";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "C9193018982050A381214A9204824B04185200BFFFFC11D7C8FE64D6F8F8F2A9";
    attribute INIT_01 of inst : label is "C4F767CEEEEE98379DBFFE116A9926604D8C37189C822AAC20C620A9918847A8";
    attribute INIT_02 of inst : label is "042F6845233182A0000004C7A18F4015571BB806C59C031499CB8C5FB9799CF6";
    attribute INIT_03 of inst : label is "0A400026300000000000810D8443088CCE28A5A0C410F371B4564CE02B2CF3CF";
    attribute INIT_04 of inst : label is "02288902AA2AA802A02A0842340B333E0858863D87BD233301ABCBD267E92539";
    attribute INIT_05 of inst : label is "E2B1BBC001C0015001640808F913EA83C0AB0AE07701D0000041C8BB05562AE0";
    attribute INIT_06 of inst : label is "B940013800250000A000540002C83C11E2909DF147407061BD0716838B41C5A0";
    attribute INIT_07 of inst : label is "4020825004A87270F23B75659F641D5D06C869C85F989D77A1AA5BA09C8A9981";
    attribute INIT_08 of inst : label is "2624474354357718088918203CE2528C8864587E9445DE02554429FF2CF9269A";
    attribute INIT_09 of inst : label is "88804402203FD5FDDFD4A000000000000000000000000000000004CC823623E5";
    attribute INIT_0A of inst : label is "9A8590A20280596BF502FF5036C0910A331C0803378E06C45A424FC250671012";
    attribute INIT_0B of inst : label is "7E9DA4FA24FFFFFF9084A3016140C81948A27C2506705120DFB022CEC7C09A12";
    attribute INIT_0C of inst : label is "96C4D4B7F5DC40000000000000000000000000000000000039836C9FB044C28A";
    attribute INIT_0D of inst : label is "41F40D76950814234B74B7EC72A54FE359ACF3DE73FC077312461F9A3A2A548C";
    attribute INIT_0E of inst : label is "C502910129DB535102819034042A8029B33D58F7CE87B10A4A25506744A00000";
    attribute INIT_0F of inst : label is "E000000000000000000000000000000000000000000000000090400210E038F5";
    attribute INIT_10 of inst : label is "D8E3E092646B56362D61B24A45FC8911C0A0A848420001E0AA2964FE08A2964F";
    attribute INIT_11 of inst : label is "9177132B01D600001CC449732C723B2211CFDBED24964BC412414A101030B082";
    attribute INIT_12 of inst : label is "2211B046D3B1222A1085AC061526451C21C6292899580E152610E441C2DC6292";
    attribute INIT_13 of inst : label is "04D6180D006523A0C50972616D8A8220A08B347D435C2DB6954F6D547E7C7E58";
    attribute INIT_14 of inst : label is "1A6D1404B0E1362A03012C625854681A0738001D5706A07AC286D71652021222";
    attribute INIT_15 of inst : label is "8562A748F50130EE2D47BD442A683305779C2882C6E8CFC01499FCFE6C512C70";
    attribute INIT_16 of inst : label is "788876DE53A9C296F69E6714E6E0B2B265A78467B80CD9B9B35B65AA8893CA23";
    attribute INIT_17 of inst : label is "0B4129273DB00825625358888CC8F064E67BCF6C02DA93FFBAF60018010070BE";
    attribute INIT_18 of inst : label is "404FC0400A11F23F6BC169EAAEAACED5C91116190CEE73FC0573DB65BEC03013";
    attribute INIT_19 of inst : label is "ACAC63FD074E24CB4E02D29B415BCCE8C126987E001C9124A02218C61C53CC4C";
    attribute INIT_1A of inst : label is "0A5777D73C78480270F0C060030CCF3D9156F11C6A1374B72AD8C55294CE62F7";
    attribute INIT_1B of inst : label is "7D542AFDAB1C8F7AC62374626DC4B5BC9F13D6F25EFB7B711223322356A0AAA2";
    attribute INIT_1C of inst : label is "B7332C5D9962CCEDC9A48EDBADAC9AA80AF000000380700402AAAAAAB556AA15";
    attribute INIT_1D of inst : label is "4852148521405005B0CDB044CA0C4444E1042893157AAD5D2BBC8CB174E58B23";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAA80485214852140500405080A4290A4290240802400";
    attribute INIT_1F of inst : label is "04A2C2FE5B4E291325257CF30B30A0932CEF44766CAF3CB2CE254C944CB48000";
    attribute INIT_20 of inst : label is "BC16BC1668D2DA268D2DA84F31304A4F4AD84AD84AD8A56C2C652C6552B6128B";
    attribute INIT_21 of inst : label is "D63090C701325257D25095E7C91E40235595B772BCF232BEBC16BC16BC16BC16";
    attribute INIT_22 of inst : label is "29D7C829D7C828829D7C829D7C829D7C829D7D293B5C3957A74C8CF04CB43CC4";
    attribute INIT_23 of inst : label is "F9C55D588F324AA11ADB395E79195E829D7C829D7C829D7C829D7DD7C829D7C8";
    attribute INIT_24 of inst : label is "200E9150529A4C1014004C5008850110B084448828480A4991330A5949136CE2";
    attribute INIT_25 of inst : label is "F7C866A6C297C295B4AA46E56FA24D5410314691514A491CAE09522A60AA7039";
    attribute INIT_26 of inst : label is "142EDEBBF3D7F594100339866F30AEA16EC32A9854C2AE4BC56022906E91492D";
    attribute INIT_27 of inst : label is "2A02E454408DC81C3950E56395BD75B58091336E817430433C0CD461502C220F";
    attribute INIT_28 of inst : label is "951AD462929800BE96A52B4A5694A52D6B52429095447BBEA5F5620800882570";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8427";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "1A510001D0041090902D28060134AF0129E4103FFFF855A908F96C446DEDBB82";
    attribute INIT_01 of inst : label is "3218BF08498C80C694313A20A7F36E828800100208A033280106AA08050956EC";
    attribute INIT_02 of inst : label is "10263DC61BB582C7FFFFFBCE279C488066F4ED7F2976BFAF6B1E6AA3220CEA1D";
    attribute INIT_03 of inst : label is "1042A4820080000000004A278013B8034E0D28F64100073F47D252760D249249";
    attribute INIT_04 of inst : label is "D9DD008A2888888A0220221B5F12143480532DDF7B970AB70B72D80C20214411";
    attribute INIT_05 of inst : label is "05F802F80EF806F006E08212980A648091188060381A30000088D202D4B0A59C";
    attribute INIT_06 of inst : label is "887800DF001BE0037C002F801DC101253A4D038520FBB0961CA02E54172A0B94";
    attribute INIT_07 of inst : label is "524DB761412AB630B62136A9A0650517D7A0A18D00500658102A52FBDA1BBA80";
    attribute INIT_08 of inst : label is "4881C093A93A92120832495A5D22A79D89455C04D000228B14952CA020954514";
    attribute INIT_09 of inst : label is "12889444A2028AAA282880000000000000000000000000000000039584566502";
    attribute INIT_0A of inst : label is "0145B8CA22742685F2A11F2A192192102176800143BB42DCE4A0920813E02840";
    attribute INIT_0B of inst : label is "720E130C736D00002896C701A593502892C020813E0800A898CE27CEDA088901";
    attribute INIT_0C of inst : label is "DA412A354A88C000000000000000000000000000000000000222726CB39B2018";
    attribute INIT_0D of inst : label is "8084900248104A026B06B01656AF6D824DAEB0842FA8466443631E7C200506C6";
    attribute INIT_0E of inst : label is "CA6CD925050101024302A05494A40169426C70982B0FF3249481D3E0B0017048";
    attribute INIT_0F of inst : label is "C0000000000000000000000000000000000000000000000001901F80028060B8";
    attribute INIT_10 of inst : label is "59E7E741495166566F671D04962120701B4000A06D23021D555C336DD757C336";
    attribute INIT_11 of inst : label is "24226C8B318A9504040021A28B223300230E6936D349B24CD3416C50204A1368";
    attribute INIT_12 of inst : label is "A39B3041DBB1287023A7804052909018B186828364598C529050C9118B886828";
    attribute INIT_13 of inst : label is "531049206DC343A0FEF3C8944E22A808A2A278D4339A3FFF840404064240404C";
    attribute INIT_14 of inst : label is "00FB454730CD38A4A8A52D4AA57CBCA3764CA80D933277432A17368654A824AD";
    attribute INIT_15 of inst : label is "016682501A881D61BC0F120667A865343850098444D00900C2BAFCFC6C114478";
    attribute INIT_16 of inst : label is "80034932C64D063C671EED305EE5F7376F82045FD0899BB3371E28AAACA26DF6";
    attribute INIT_17 of inst : label is "2EA3376617E08E654AC1119999D8D66D82E105F022C467D1B1960EEB5F2A4FA1";
    attribute INIT_18 of inst : label is "28894800303BA0712FE9A2EAAA23D08171333A5D2CCC2FC846672A28F9421A32";
    attribute INIT_19 of inst : label is "01AC223C0A5C75DB8422431491698BB80546B800000124EAB003180618E2589D";
    attribute INIT_1A of inst : label is "885D7F661C2D671641C4E540DE19137A40F790184F0207610A64A057189CE7C3";
    attribute INIT_1B of inst : label is "87015503677A8E498C6B68C68D8CBB2D9632ECB65C3363637EEE7EEFC6822282";
    attribute INIT_1C of inst : label is "365A6CDEF366D78D92C928DF8D989E02A050000002805000038000001C0380AA";
    attribute INIT_1D of inst : label is "2308C2308C2308C3339B71F4BE3C4C4DE30D1FFF1DD6793306D929B379CD9B4E";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAAA5611846118461184611A5611846118461184611AD";
    attribute INIT_1F of inst : label is "440206AE698871366CEF31C72F72B0BF2CA90C774DE671B6DE6417F4CED38000";
    attribute INIT_20 of inst : label is "EBE94141421D80D423C8041C73F0CFDC4242C0C0404060602020616110103088";
    attribute INIT_21 of inst : label is "C05DA4414166CEF347D0BCCE5B7CE90777736F2799C7379BEBE941414143EBEB";
    attribute INIT_22 of inst : label is "81FD5FD4A80A81FD4A80A81FD5FD4A80A81FD4BFF24147041C7885A0092171CE";
    attribute INIT_23 of inst : label is "04B61181BE6F4EE8B9B783CCE3DBCCA81FD5FD4A80A81FD5FD4A81FD5FD4A80A";
    attribute INIT_24 of inst : label is "AD2E4864212176A054D3D14AC854AC0A895062A54089A50541E419632D9D78CA";
    attribute INIT_25 of inst : label is "5B2C6A892A582A58BC4B61F774ADA3E15A7326D865295410914D9EA14471F461";
    attribute INIT_26 of inst : label is "32A111240A20494501053252410A919511107C45482A416C148CAA2A06D869B2";
    attribute INIT_27 of inst : label is "1021C464090A213A40090004003755DE08528FC2140E011BB06EC4807DB00C69";
    attribute INIT_28 of inst : label is "D05422CB03B28890B4AD694A5295A5294A4924B2AA002EEEA5154588189106B0";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6E35";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "325B6021D984549494253936CDB6EB092974023FFFFAD5FB5BFE82664BEB9FAB";
    attribute INIT_01 of inst : label is "4A9488719BAC1018E6D77B003556C8180A699043CBC13AA90422A821DA3B57DC";
    attribute INIT_02 of inst : label is "9C3FA740D4AD041FE07E022AC45590D6C6600781AA43C4A9A1E17330CCC33299";
    attribute INIT_03 of inst : label is "6C9AB6B6DB80010402085247169350D2943128A909811D210053C32A00A28A28";
    attribute INIT_04 of inst : label is "001800228A0A0A080282829B712A5C74DC3AB85A3337B541BA3E10AAA82189B6";
    attribute INIT_05 of inst : label is "04F802F80E780670064000001000418080080020100010000000400200100080";
    attribute INIT_06 of inst : label is "A8C00058000B000160002C000580000020000300004390001820241012080904";
    attribute INIT_07 of inst : label is "492493701DF4969B96F49549204E0724462D30AA40F446C8386E5288F2CA9C50";
    attribute INIT_08 of inst : label is "6E9262D3ED3EB696C93B6D73BDD6C7B018477CE455DFFE4B72D4DA8B3714E79E";
    attribute INIT_09 of inst : label is "3A93D40EA4F2A0A82204C8000000000000000000000000000000025AC8722033";
    attribute INIT_0A of inst : label is "234C80E84E14BAEF50A5F50A4DE49138132A9165F3954A4436E6D869204239C9";
    attribute INIT_0B of inst : label is "214A09012805000039826724A5C07A04DA648692042924E9087E62424029ABAB";
    attribute INIT_0C of inst : label is "5649FE77224A40000000000000000000000000000000000003A42900908FE4CB";
    attribute INIT_0D of inst : label is "460C1AB36C064E526B86A841018108A20168A0000800986749272F9030C7224E";
    attribute INIT_0E of inst : label is "C626C965DA1010A22DA4740C14A64909422914883B469106DE920042D2496183";
    attribute INIT_0F of inst : label is "40000000000000000000000000000000000000000000000001605FFE02826CA0";
    attribute INIT_10 of inst : label is "48A2A1C96D513A1225211726D307A49889A313E4940C13C28009280420009280";
    attribute INIT_11 of inst : label is "74A23E990C8AD68A7050A4C29366631079E40482492006444959265259EA51A9";
    attribute INIT_12 of inst : label is "6D6A298A0A0241380E94A09C5348D2D8ADB29791F4C864534856CD2D8A8B2979";
    attribute INIT_13 of inst : label is "290B24926DC1EB92451940D485775F575DF7625109083EDB6840428D4143434C";
    attribute INIT_14 of inst : label is "0F89E50492453E96949496247CC8651A9128A40903182A06EC96E2621EA6369F";
    attribute INIT_15 of inst : label is "F1C3079A57843DEDAD871F0860252713187818B45858F78008CADDDD4C3645B0";
    attribute INIT_16 of inst : label is "7A31008452CD32944612EC340209A6A64D601D9001315AB2B55A28B924A3AEF2";
    attribute INIT_17 of inst : label is "28002104040030412A70611111D098492090C1080D6E07D804E38342684D7CBD";
    attribute INIT_18 of inst : label is "A90B4124A861272364A5F24000AA8844312222110AEC08009868FA28C7846002";
    attribute INIT_19 of inst : label is "389C0DE5B2E3605A404CE217D6CB1CA2098498000001B68B8624BCB24A42C8D8";
    attribute INIT_1A of inst : label is "750A0214000B460A8286FC864EC99D5BD9DEB24A4603A6A8017CE1921096A4C7";
    attribute INIT_1B of inst : label is "0155400255AD5E91294A4A94A928220904A08824120A4A4224444444B57D57FD";
    attribute INIT_1C of inst : label is "A4780817C0409EE91AE9AA90A914E2AAAA95555554AA955554AAAAAAA554AAA0";
    attribute INIT_1D of inst : label is "695A5695A5695A5699124C949456A869880C9524C8945122C4B9A0205D01026B";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAA84695A5695A5695A569584695A5695A5695A569584";
    attribute INIT_1F of inst : label is "72399CFA7B552124494811040B44F8A5A68B6445450241245241412E892D0000";
    attribute INIT_20 of inst : label is "AAAAAAA9575AA01575AA02105A2E04AC63736373E1F171F9B8B0B9B1B87C78E6";
    attribute INIT_21 of inst : label is "BEA146CB294494810494A0485224A572222249C409042408000000000002AAAA";
    attribute INIT_22 of inst : label is "015555555555540000000015555555555540009232A2AD6935E4E49014284168";
    attribute INIT_23 of inst : label is "C825D0711245244B1124F2048212055540000000000015555555540000000000";
    attribute INIT_24 of inst : label is "E5AED9749E315A702C49DF6B4B56B56ACDD892BCE03895D7597F583305FF286B";
    attribute INIT_25 of inst : label is "77C872CDAE0E2E0CB7636571F5B493E4CB6906D975A5D5DD896DDEB156F2237A";
    attribute INIT_26 of inst : label is "10B1316C1F684BE7998133DC998ADD859DFE82A36F2B716F170CAB7B86D96DBC";
    attribute INIT_27 of inst : label is "584E44ED8BDCC96E7039C0E703155493134AD310028D4734A6529932C686466F";
    attribute INIT_28 of inst : label is "555633DB04F6039D9CEF39CE73BCE779DE492FB6BF21CCCCE7464558159576B6";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C35";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "B11C9818C0711444C6108491349226B4001048FFFFFF23A9E5FF46E2C9F9C9B8";
    attribute INIT_01 of inst : label is "C473CA94B88C19B5A9911B136D480471A7C6438826CE932DF1BC8AABD50C8EA8";
    attribute INIT_02 of inst : label is "6800650132B592200000064F249E4000E97B159A4E8ACD381B388CCC3337147A";
    attribute INIT_03 of inst : label is "82638041048001200240E0920859110E084582600010E5F4F10E8E20031861C7";
    attribute INIT_04 of inst : label is "FFF7FF280AA00AA002A802E1908B386B2ABDC82A2D33ABA28A1358386421B609";
    attribute INIT_05 of inst : label is "FB07FF07F107F90FF93FFFFFEFFF3E7F7FE7FFDFCFFFEFFFFFFF3FF9FFCFFE7F";
    attribute INIT_06 of inst : label is "113FFFB7FFF6FFFEDFFFDBFFFB7FFFFFDFFFFEFFFFBC6FFFF7DFDBEFEDF7F6FB";
    attribute INIT_07 of inst : label is "24924911247FD650D6371125906609DC22406E48A0797CE01DC709844420CD19";
    attribute INIT_08 of inst : label is "0149090B10B1014C24C58D8C0E472910C8123A130330030019C3F8A390CB4104";
    attribute INIT_09 of inst : label is "88A4452229180A00828E50000000000000000000000000000000064893122088";
    attribute INIT_0A of inst : label is "02A49620DA0A4101505215052012CB88B9114CD10B88A6440012415481098424";
    attribute INIT_0B of inst : label is "84A16DB28DB30000848D928210460A824991114810949214B781224241140202";
    attribute INIT_0C of inst : label is "0124090262E50000000000000000000000000000000000003852C5B790E01220";
    attribute INIT_0D of inst : label is "AC54423954412129C49C480CB3660F08DFEEBDEF79B826D0A6CA96598FB09D94";
    attribute INIT_0E of inst : label is "41D9A4D089CBCB50928C15044211046CE7980A607E7291124148810909249A6E";
    attribute INIT_0F of inst : label is "2000000000000000000000000000000000000000000000000080007E1811026A";
    attribute INIT_10 of inst : label is "C8A2A0242404CA32252040924C9052427656C81227BA4862A82B8DB22280B8DB";
    attribute INIT_11 of inst : label is "C209804902600924CB8E522948DDD6EF041092D92D92DBC42404D90823053014";
    attribute INIT_12 of inst : label is "331BB3664B38A68882CC18230866083603094C4C024813086701A083602094C4";
    attribute INIT_13 of inst : label is "8DE49A4D924542CB911C320A58A2A008A0AB85300EA4BFFFC72F2D4616161619";
    attribute INIT_14 of inst : label is "198970484BB0B040474A4691024924421B9050188910201A3042265860518040";
    attribute INIT_15 of inst : label is "0F190A81B29850E60CF040E120B29108E0741E4125283CC3B449BCBC2CD91270";
    attribute INIT_16 of inst : label is "01E1965D2938A9412D4A6612F221B6366D963673704D9B3B3798826C86085836";
    attribute INIT_17 of inst : label is "81A99457BCB06964032BD8888CDAC564964B2F2C1A4433E6879374A41483C963";
    attribute INIT_18 of inst : label is "14A4C410072DDAB802D328600022C232C4111A9D4FBB79B826D82882410D2A99";
    attribute INIT_19 of inst : label is "027F7A20416700C32C12594C8DFDB5E18252C8000004018089910A0D7529662C";
    attribute INIT_1A of inst : label is "2AA02837B37909213DB8C339B034443E62861975320D2EA606861F594A5CE360";
    attribute INIT_1B of inst : label is "0155400B673E8EDCC621746205CCBB2D9732ECB6597171719233222216802800";
    attribute INIT_1C of inst : label is "17152E5CA972C405C184005C058C72AA003000000180300554AAAAAAA554AAA0";
    attribute INIT_1D of inst : label is "695A5695A5695A5650CB68460D1D4D0C111608B60472371B620C04B97025CB00";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAA84695A5695A5695A569584695A5695A5695A569584";
    attribute INIT_1F of inst : label is "85C26037241E94132426CC96A77A7E160000130010D925B709672DB4CDB08000";
    attribute INIT_20 of inst : label is "55555556EA5A9E2EA5A9E189736442DF1C0C1C0C1E0E8E06474F464E67A3A709";
    attribute INIT_21 of inst : label is "94389820CC32426C92C61B24899250AB11116C136496B367FFFFFFFD5557FFFD";
    attribute INIT_22 of inst : label is "ABFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAAAAAAB0BFF5D0B086C659E915C0225CD";
    attribute INIT_23 of inst : label is "796319E8C9228225D8B689B24B59B3FFFFFFFFFFFFFFEAAAAAAAAAAAAAAAAAAA";
    attribute INIT_24 of inst : label is "221F22C25E8C011114240094842948852026280222084A2F0F00888910118314";
    attribute INIT_25 of inst : label is "BF298BA01221D222C18488E060C2CEADE4051722C253C0F28292254C3E568BA4";
    attribute INIT_26 of inst : label is "114CBC700EC873412180CC216465208A42298108909484D0E87214C43722D341";
    attribute INIT_27 of inst : label is "E890D31644E110811F847E11F8C4465004A1970C8D343872B84AC443C0087121";
    attribute INIT_28 of inst : label is "47008649129208C6E6398C6318C6318C73A490C8409E000031A22360060FAC39";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA611";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "312218190061160404800000B000461094B000FFFFFEA30091FE0391C8F8C091";
    attribute INIT_01 of inst : label is "C4218A52B9981804A1911310080804D38540861842CF0225A8A08A2BD0028C88";
    attribute INIT_02 of inst : label is "6BC0E000B210821000000644A4894084A53F3498469A4C18123884441117142A";
    attribute INIT_03 of inst : label is "455380208A8008001000D04314D9009E0C258060890D8DF4F10A0E2001104145";
    attribute INIT_04 of inst : label is "001000AAA0000AAAA80002D050041C4A832AA82A0D13A100AE15483844018501";
    attribute INIT_05 of inst : label is "0100028000800080008000000000800000100000000020000000800400200100";
    attribute INIT_06 of inst : label is "1180001000020000400008000100000000000200008000000000080004000200";
    attribute INIT_07 of inst : label is "0000003400FFD2515247152CB026015C12440058C06150901882098244408C8B";
    attribute INIT_08 of inst : label is "0101010A10A1018840AD4C4A0944A44008001016033A20242183F8AB10C81041";
    attribute INIT_09 of inst : label is "1892C40600080800A80D50000000000000000000000000000000064802B22081";
    attribute INIT_0A of inst : label is "9A94846002A94101544A1504A00AA55855012A090A8096440008091001011200";
    attribute INIT_0B of inst : label is "05D12DB7049300008280200000D01A0000211100101200128780A24351529A9A";
    attribute INIT_0C of inst : label is "028400A022D6000000000000000000000000000000000000384A0C9390560A41";
    attribute INIT_0D of inst : label is "C04408311C00843106906804372F25804FA799CE7998161090181C5D0A2A5030";
    attribute INIT_0E of inst : label is "4102804089C3C3500384340400020068A5180C50704291000900810100005848";
    attribute INIT_0F of inst : label is "2000000000000000000000000000000000000000000000000000000050300468";
    attribute INIT_10 of inst : label is "C8A2A20000001A32252008000190404040E08000032205280021049282021049";
    attribute INIT_11 of inst : label is "80015809044005141A8440610B0010AA082096596DB649C40008022030043410";
    attribute INIT_12 of inst : label is "231111464110A31801040816016E00540511080AC04822016E02A00540011080";
    attribute INIT_13 of inst : label is "4CD241210001222A141A720841A80020AA034E380884ADB6C70F0D4515151508";
    attribute INIT_14 of inst : label is "198160402A28A020272926488140A022055048188110200200A2040440498020";
    attribute INIT_15 of inst : label is "04411880B000C0C208400043298311007860102014383D8C9649F4F464550170";
    attribute INIT_16 of inst : label is "008196CC0120B000210A6610F220931324860573702C89191388000A80004224";
    attribute INIT_17 of inst : label is "03AB14533CB00B2C222318888CCA452486430F2403423092470B44A014038943";
    attribute INIT_18 of inst : label is "1084C0000224F0980240682000224610C0111ACD64027998161800000000AAB1";
    attribute INIT_19 of inst : label is "182A6220A9A431890C0A41080178816081428800000401820400001146214468";
    attribute INIT_1A of inst : label is "802A801332780901B1B18030004444340604014622811A4202801451084843A1";
    attribute INIT_1B of inst : label is "0155555922140C4CE72336720CE59964B3966592C86323319233222212AAAAAA";
    attribute INIT_1C of inst : label is "331064CC8326440CC18400C80C8A7200001554000080155554AAAAA005548000";
    attribute INIT_1D of inst : label is "6118461184611846D0C9284C0808060610E008928472301962140193300C9900";
    attribute INIT_1E of inst : label is "0000000000020888A2AAAA846118461184611846118461184611846118461184";
    attribute INIT_1F of inst : label is "0D86C0620017101324265CB2E62A28128200200000CB2C920B2D0C9064908000";
    attribute INIT_20 of inst : label is "55555556BE29082BE290808B214422571818181818188C0C0C0C0C0C4606061B";
    attribute INIT_21 of inst : label is "0418941008324265B2441965C9964009111124332CB2932FFFFFFFFFFFFD5555";
    attribute INIT_22 of inst : label is "54000000000000000000000000000000000001095DCF022908A1090E94062C85";
    attribute INIT_23 of inst : label is "3B619818CB220220489219965949975555555555555555555555555555555555";
    attribute INIT_24 of inst : label is "215C0600408800301400005280252904A014000060080A8E02220A1900210012";
    attribute INIT_25 of inst : label is "9A2D48200A94CA96A18018C04026DC0B22215C0601438028864015283F84A090";
    attribute INIT_26 of inst : label is "1528A8400C481210518428132C24A0A9420B82885092840A64E812823406082B";
    attribute INIT_27 of inst : label is "F848809962D19C430D0C3430D044445302818D0401F4107214485423C0046201";
    attribute INIT_28 of inst : label is "0600868000A000C2C631CC6318C631CE63000AC46B15444431E23150454E1824";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAA81";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
