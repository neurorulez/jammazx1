-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FDFFBBF35CA77DEBADEC4E12AF333241819818A23D8D49BCAF6DA9064D3E5503";
    attribute INIT_01 of inst : label is "051589350B90D1A2B057002003D1DF471ABCF6E90E7B7210CD2B80FF6D9B3BAE";
    attribute INIT_02 of inst : label is "DAECCD6476BBB5F97A30187838D04A3D0E91428F41EFCFF691AC1349B1492280";
    attribute INIT_03 of inst : label is "BB3FC3EF0BC8508A235A8BE9D02217D4224F053E243723A00A22E48326333591";
    attribute INIT_04 of inst : label is "D02099BF641E413E08447AB19A7E27D6CC89D8F3D9F2809401FEDEB13E408EC7";
    attribute INIT_05 of inst : label is "EF97CFA1EF7EF3FCFCF68555EAEC444D3D6B2847FD14D0B2C4EC84FF87C3F57F";
    attribute INIT_06 of inst : label is "34CBF109682A948202760DBEDB7170C160C83319A51D96000089F39912BF5755";
    attribute INIT_07 of inst : label is "D9F9CF1DB99F39E3B2D9BE78FD924FB79EF3E57F3BFC1C1C093FD11C294049A9";
    attribute INIT_08 of inst : label is "96EB77B05CD4CF75FBBD26497BB3C9BB3D4CF178ECFCE78EF339C6CF9E3BBDB5";
    attribute INIT_09 of inst : label is "86688DFA67FAAB47E8B44CF5FE79B4887F5D757DB40081015ED1EF8AA527D4F6";
    attribute INIT_0A of inst : label is "2B48624896036A8609C08101B0D7A28A6648D1A5D9A5DAEA2B42BA71138899A2";
    attribute INIT_0B of inst : label is "8C89704038526001C9934A6164D2D849901364A059C826C83B4C22C83A4C2248";
    attribute INIT_0C of inst : label is "69269A49A69A49269BF3245A8B304030112D402D0914B4520AD3088043103525";
    attribute INIT_0D of inst : label is "A69369269269269B69A6DA59269A59269A4DB69A69A6924B6D92596592492492";
    attribute INIT_0E of inst : label is "10C104B04B28A10638C06144200204228B24F24B24934F00200E38C069A59659";
    attribute INIT_0F of inst : label is "49279A68208228A28208228A29308308308348308308309A49249249249001E0";
    attribute INIT_10 of inst : label is "25291096C8AE6574E2751665AD4A5908172634E026603624926B4D0410451456";
    attribute INIT_11 of inst : label is "5EEA1115A0215EEA1115A0214997186EAFED0FB1C87E0D630034A3498D02C479";
    attribute INIT_12 of inst : label is "D576B9EFB13A4656385C22ADBFACB807EA40DD66B35D2DB659A1FA3FFC13521F";
    attribute INIT_13 of inst : label is "B9AFFB6CFECC1DF59A3BDD9B972D96793F58CB9691CE73ACC72003D5272D5255";
    attribute INIT_14 of inst : label is "3D4E97B89C439F4BAF3FD66444444445D64DB2C927C33BEAE7ACBD06E358C635";
    attribute INIT_15 of inst : label is "724CC065B6FFD0C016416B01923212E66AC1660D6073FDB6DB2EB6493E163BFD";
    attribute INIT_16 of inst : label is "8CC1981CFF6DB6FBB59FC58245FA3851BA2BCA2D23492C51B4AC94EEE5BF4ADF";
    attribute INIT_17 of inst : label is "F6360E2416DBA5D6E96493F43F8EBA91A4961CDA564A7772DFA3EF6502566658";
    attribute INIT_18 of inst : label is "315853148541D7535653292AE380139A93328691E41FA4B27B316ED018B1CD14";
    attribute INIT_19 of inst : label is "E93680019FC3424AA9A860602664283A39031A44737DBFF907041FB965039F55";
    attribute INIT_1A of inst : label is "9C8C2A733A7F2CE2C0725A5FE7DC0BB8E55E215010D12F0404C59645D6D973A9";
    attribute INIT_1B of inst : label is "96B9B9FB8CCEFE25CDCB044388D0DC6C6EE2AFFE969C2B77152AFFA4C0B7DFB0";
    attribute INIT_1C of inst : label is "650E8475F3B87AEF8EEFF39CE7203DC1FE438E8688BAB677BFFFF73567759AFD";
    attribute INIT_1D of inst : label is "D9698EC225A04AD96F69DE00044A54454068D8DBE6C6CB6CC31C30F567666AAB";
    attribute INIT_1E of inst : label is "499057FA23FCFE3EA597503EF65C6D7F1E38C45A921E22EDCFBFF744C9FDB13B";
    attribute INIT_1F of inst : label is "60415056FA2E1C8813A00DECAC9A997CD390134C1301051765A34D933C109380";
    attribute INIT_20 of inst : label is "FB4BC68086E01BF02C27E39D24C4B4F3AE8B001719EFFDDB213EC01AF02F4ACF";
    attribute INIT_21 of inst : label is "4D0BDC7C76B2BDD9FF373FDA3DF28514EF265BEA205D68B3D6E058001B5FB764";
    attribute INIT_22 of inst : label is "2804A1428140250A147AAC52630B6B9EE5B9DEF93EB60803E61536FE67AEF791";
    attribute INIT_23 of inst : label is "0000000008000000000000004002AFF004000008080008000010101010004020";
    attribute INIT_24 of inst : label is "0101010100010A140050A810A140050A0121A0B0000000004040404000200000";
    attribute INIT_25 of inst : label is "2012000000000808080808000050A80285028540142B80BB8000004000000001";
    attribute INIT_26 of inst : label is "00161F7A00000008048000000002020202020000142800A140A140050A400440";
    attribute INIT_27 of inst : label is "B04150916439D1BF5FFF00400004024000000001010101010001000000040000";
    attribute INIT_28 of inst : label is "86CE77185E7F3C40779E67BAE618767CC3AE871F0F1E31B0D66F0011400EDD49";
    attribute INIT_29 of inst : label is "B9B5D58EA5F26D14DDA6D64E6727F4376E9F3CF9FCF101C24C673B8E78D47984";
    attribute INIT_2A of inst : label is "6523B2285E986CFBD344AAAAA79159DD2001D94D8DA693F6E7CF99939E9ED25C";
    attribute INIT_2B of inst : label is "669F2CCD6A006088001408CF93A58B0F19DF67D2BF28677F72D468A02D6DA15F";
    attribute INIT_2C of inst : label is "FBFEDD5557FD57F9F3269E6BE853CEB3F3E7F87F38B41A2D3177C00A8A0AD24B";
    attribute INIT_2D of inst : label is "677FDFFE5D6C5A913DF9E4E6C7D7B8DD9136DBDD86FEBFBE653D6FE366EFE97F";
    attribute INIT_2E of inst : label is "64B26FA34D6952151142B629A20AD2250D34FFD42EFF1E913BB96FF55C855CE7";
    attribute INIT_2F of inst : label is "A345ACE8E5F66AA16211752BADAAD62CA41EB8270ECDD150D114800812A40809";
    attribute INIT_30 of inst : label is "007FB74827DCA275CED255E68224EBE7134EB14CC8DA54B3533E35306765CE57";
    attribute INIT_31 of inst : label is "60282E604C0802401FC0FF2AA505FC490000100496990D4100040F209B7F8000";
    attribute INIT_32 of inst : label is "04096CC96E000081798565FC0017A71105180020569189B4C0000AAA0029A7F8";
    attribute INIT_33 of inst : label is "50663C1F0000AABC6944600027A48E0EE35000280FFBCD3F000017F848E38B00";
    attribute INIT_34 of inst : label is "054118D1F8001555E1A020014AF00348C00005550011BC0040EBE000C7780002";
    attribute INIT_35 of inst : label is "444444427800800007C0DA600005051897930400222159A00003FFC0CF6DC420";
    attribute INIT_36 of inst : label is "314463FFF7339C6FDFAA6EED77719B85D886E4973319BB5C8A66ED501DAAB5C4";
    attribute INIT_37 of inst : label is "12999166809FAE993207474A285E7A53322DC93FBFBEE1A72834BF7EEFD438E9";
    attribute INIT_38 of inst : label is "042E15001991566885B28951B5609594282A5145432596E9F6D8832C13D2A933";
    attribute INIT_39 of inst : label is "85279CE41667E8288877C815A308F8B6AC88540340022ACD7089555910886833";
    attribute INIT_3A of inst : label is "FAD4948D2548DA564A7772DEAF93BE1C6E6FEAABAF5EB97AF4567F4BE7FE7399";
    attribute INIT_3B of inst : label is "E06A1C6CDF44AE1F1C902AD60E13F3EFFB32C0DE01693C42E755F37DB6597EB9";
    attribute INIT_3C of inst : label is "840A080C0282181CAAE49CFF0DBFB7EDDBD7BF5F7875299CF955B12B657CC9C5";
    attribute INIT_3D of inst : label is "D683087A2B0ACACF8823E06A2462E08CE4CF3CF3CC97DC214D058888A9308602";
    attribute INIT_3E of inst : label is "55494866D486A7D412F543EDDDDDCDC517980256B9A6019B200A19AC22D2ACAA";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "57C1494126EF3FDF70255EE2E3FFFC17FFFDB49A453F62DBB07E6C260566CB27";
    attribute INIT_01 of inst : label is "719D94069F4D2E13B25809242513B029D9C01AE6F10C7DE0DE2D1185B4B08812";
    attribute INIT_02 of inst : label is "6830140A1A0CD3268DC13C8A6AF32A6730582A998677D78BD31C86DFE86DB3FE";
    attribute INIT_03 of inst : label is "0061A7DE9409C949A601C03616656812652008465670AC8312E58A1302105020";
    attribute INIT_04 of inst : label is "2656D60600D284BD39D98B94B852C09A27314000A085E72F3B025AD608CD9CCC";
    attribute INIT_05 of inst : label is "026121C0D4004842B82DF6782C80501AC485ADD8177FFD2960034D82312530D3";
    attribute INIT_06 of inst : label is "00D1032EB3D4200A79B80820164A4A0A4E13701D43980C8888000BE45B43CF31";
    attribute INIT_07 of inst : label is "0B28C38720B51870E60B0A1C0092CFBCBF77D7EC8208C8C8C040089D0CAD0000";
    attribute INIT_08 of inst : label is "261E0FF185B85C9FAEEE88D81C151DC15385F5C5859461C3E718085A870E041E";
    attribute INIT_09 of inst : label is "331BBBA82E0147F2446485CF8AF69264802888816577F954A7F7D03B3743B9C0";
    attribute INIT_0A of inst : label is "3F2C8689D20869C211689D04B44AB4CB829A5B225F821B34338892B919333300";
    attribute INIT_0B of inst : label is "A4C83040311922000DB75BE74D96B1C31001642051E086C83B0882C83A08C2C8";
    attribute INIT_0C of inst : label is "49A49249259269A5967A040C07004602430D0430CB55ACC208CB30804340E521";
    attribute INIT_0D of inst : label is "64926DA69A69A69B69A6DA592592592592492496492492492492492492492492";
    attribute INIT_0E of inst : label is "B2CB2CB28A24F24C147A4104B2CB2490C10430000000432C82C10C1249649249";
    attribute INIT_0F of inst : label is "41051040000400010820C208300C71C30C71870C31C70C1220820820820F7860";
    attribute INIT_10 of inst : label is "4B932144C5291E50983D224E6719C63BDCD06F325820864000100028828A20A4";
    attribute INIT_11 of inst : label is "608D3B7EF2FB608D3B7EF2FB54B4D70518777CEFB7EFFF3F005AE5741300881A";
    attribute INIT_12 of inst : label is "E67C57A433AF15CDE1BD57F526B79C952912A65A2904C165A6DC986E16BDF888";
    attribute INIT_13 of inst : label is "E50A10585884D1110BA204C0810005A69310A78423FEF588A340013202CC3477";
    attribute INIT_14 of inst : label is "E7B0DC03D002500FAF5F932444444444600060B0D20C8A7F03ECFF07EB18C6B5";
    attribute INIT_15 of inst : label is "C9AEC90205861962EDF21B5308CEB4DAD9B0764EE4C58205948B45B687246116";
    attribute INIT_16 of inst : label is "0EC9D93160816522D168691D0E1870D07F13E40561C3D22115FCBC2CB37E4448";
    attribute INIT_17 of inst : label is "FE7E6F4170B20144B058693E5FD610B0E1E92C8AFE5E1659BF25A4929F8D8F76";
    attribute INIT_18 of inst : label is "13F8F2BD0F01EBF1FEF2FA78F400040FC2210F88D03F2C5124B20041731B6DB6";
    attribute INIT_19 of inst : label is "164B2C99ADDB312EB8FC97EA4C40847EF4B941B0EC90A000343D80825C64EDAF";
    attribute INIT_1A of inst : label is "EF3993129593969ED4EE852839E059C069FD607D992DB6A6F2C9493325A69CD2";
    attribute INIT_1B of inst : label is "A724CBFD451C506B02E028E6117BE0C23F076153292BD2D8689188C91F2DA24B";
    attribute INIT_1C of inst : label is "6D204F93B3B9FDCFDC1EFFFFFF33FDCF6D2FD9BDFC7DDAECBC0FD97AB3683F65";
    attribute INIT_1D of inst : label is "1AA8F8997E3F8E65A156A8DE263EACCDDE7CE4C7E7667DAD1996BBA62626C791";
    attribute INIT_1E of inst : label is "F3B7DD29DFC86BBD4D1D0ED28387D4B17EFBDED43EA75196BE9E98EEDAB4A312";
    attribute INIT_1F of inst : label is "CC237725687BCE908BD3DB7B75C76BA20CE6328D31912E3C69466A3B61B931B7";
    attribute INIT_20 of inst : label is "F46E585DA7C3B507C23EA52A65AD3969627647BC71DA357252C9B97343F49994";
    attribute INIT_21 of inst : label is "2E4435FF9BFA3B68814A7BB8FE0A4A8B5F56D5A679680444FB05DB789B90BF91";
    attribute INIT_22 of inst : label is "0800204091204489136AAFA93F9C7B18D2B1A1A0505AFE7C2A87D1A7FE1310CD";
    attribute INIT_23 of inst : label is "0A142850AC58B162C58B162C6A6ADC1403060000060C04000008000808080422";
    attribute INIT_24 of inst : label is "0002000080008204281021489122C48916949410000000400000800020314285";
    attribute INIT_25 of inst : label is "021200000008000010000400041020008122448112242A157800204000000100";
    attribute INIT_26 of inst : label is "103D557DC0010100848000000200000400010001040800204891204489FAFAA4";
    attribute INIT_27 of inst : label is "5B0A6B96F63F6F4D76D0E0408080424000000100000200008001800000060408";
    attribute INIT_28 of inst : label is "F097A486838D7DB72059D8CF15A6B74730FE1B7E75E9DB8F7ACAB3B237740000";
    attribute INIT_29 of inst : label is "CAF97FDE1DCFBB3E22F121F794CFFFC41840430E35F6D814B34BD2438F2B162B";
    attribute INIT_2A of inst : label is "B7A56AEFE3DEA5D23F3F7FFFF937EB0F66760482DFEDBFEDF211076721C1EFB6";
    attribute INIT_2B of inst : label is "034041050FB5F65E794D65AB6A9C40C4C2445A47CBC116B0501BA913D612ED80";
    attribute INIT_2C of inst : label is "FF2911998002AAA0CECDC01C2BEA2F404488211CC05C6637120C000780A9F835";
    attribute INIT_2D of inst : label is "10A0040116A6AF34DE10985A5E64885736164B26D4015419DB838835910210ED";
    attribute INIT_2E of inst : label is "3E56DAAEEA9BB67ED9DDEDFB7BFFBF7F6583404185015E6EC680B005521289BE";
    attribute INIT_2F of inst : label is "4C673A243B898D56B259A717C03548D6F48802BF825A2EF5F9291FFDEF59FEFF";
    attribute INIT_30 of inst : label is "000028082DF5D78AA3689AAAA468668154BA4F911DEC3E446D7E47BDC81203AC";
    attribute INIT_31 of inst : label is "0428281BB3F0004017A50000040100368000141460C4A400041000332CBF8000";
    attribute INIT_32 of inst : label is "150082D48000062401BA8F78000501E047E8E10102206E4B400204440211BA60";
    attribute INIT_33 of inst : label is "D400196802AA00038EE5500101E34331BEA800280BC2321008A015C2546E8001";
    attribute INIT_34 of inst : label is "0AAAE02E000001542D5000074A988CB780000000FEEDC7F208015DE752A00000";
    attribute INIT_35 of inst : label is "EBEBEBEEF4008082A02725BF8040007CBA25F8004001E5500003FFC0D002B841";
    attribute INIT_36 of inst : label is "005A8000182955068004850B82894158A0A850F83C94178E0E8FA785490010EB";
    attribute INIT_37 of inst : label is "2A75FA08C6F83B5F88F0299864E94C4EBF0925B86082220E448378DDB420704E";
    attribute INIT_38 of inst : label is "3190C8B29CBDB70448B8CDF526B95DC24345682A6AD16CB48B635AD0E921FDF8";
    attribute INIT_39 of inst : label is "F89D5E98A018CD9EC4C8116ABD6F01453AD9B4B62CA7B6E486425A75B36B6533";
    attribute INIT_3A of inst : label is "3E0925870F808AFE5E1659BEBEA01C20DE1E05316BB5AAD6AA0E00B809FD7A7D";
    attribute INIT_3B of inst : label is "CCB599934C92ED7B792B198E7329D1B00805EF48F2A2F1A50687A59145A69F23";
    attribute INIT_3C of inst : label is "0C1A222200A8800600828084382FBFE1DFBE2CE6245230BD0C6848B0978040CF";
    attribute INIT_3D of inst : label is "43450D3880002027010788000200BA0277C18618624AACC00A001860030CC220";
    attribute INIT_3E of inst : label is "202BC424C808AFB0033D006DDDDCDDC4FFA800D5F25EA54D0C180081803A0200";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "000080102CECEA5CD94F6F4BA84446D63E232CCB2AB03090CF6B9512A519CC02";
    attribute INIT_01 of inst : label is "0B5505C4EF4F1FEEA1700830209D68C396F29A3DD94C1BBA7C380883692C0C60";
    attribute INIT_02 of inst : label is "4325018280C02C9923B11C0A2AF1233841022ACE6977D82509181492DCDA4882";
    attribute INIT_03 of inst : label is "551852214628804EB90954CA18018C18018C056819B03A2483013A895004864A";
    attribute INIT_04 of inst : label is "8D1928D48442C07B4331832961A313D8C9EECC20B48AC55628E21B189CA118E6";
    attribute INIT_05 of inst : label is "1D4EA79824F22B222A69E64A65A0541179E64C6029461A49922675F8C8ACBB30";
    attribute INIT_06 of inst : label is "1259ECCE59E6E873B3B50BA9D4F8FA30FA26704F291BA8A8A8A800A6747F3FF1";
    attribute INIT_07 of inst : label is "4BCD6DD406B9ADBA844B336E81201498AE746A923C0AEAEAE27C044F89634088";
    attribute INIT_08 of inst : label is "B7C865D1A5AA5E100880261250974C897AB5F50DA5E6B6EA05AD4A5CDBA820DB";
    attribute INIT_09 of inst : label is "088000012F004CB24644A5FA42F803877EA80280155D595FE6555799245381D0";
    attribute INIT_0A of inst : label is "41004088900046A6AA648802224BF008401AF8A05080508988B9810228000010";
    attribute INIT_0B of inst : label is "04481000080116D65C3400C00D007802121924B451EE04C8000000C800000008";
    attribute INIT_0C of inst : label is "2000000001001000040D449A90044810084D9AB95B701E22044000304A090224";
    attribute INIT_0D of inst : label is "4001124104104100000124000100000100000004000000024900104100000000";
    attribute INIT_0E of inst : label is "0000000042080001002018282002080002000043043000001242000000410410";
    attribute INIT_0F of inst : label is "000000014414510514414510530820861861C618608208082082082082048068";
    attribute INIT_10 of inst : label is "EDEB6B99F1C56F266BB7145425A84A1AD4AFA9C19E2014400410020000000000";
    attribute INIT_11 of inst : label is "2153CB8B5D12E153CB8B5D12E5389F8B3BE97D7FBBEEFDBF007863ED5B0326BB";
    attribute INIT_12 of inst : label is "F8FD372821FF1FC1843FC15458171C0A009150A150385D0A953BF9741CAAABCF";
    attribute INIT_13 of inst : label is "F0520F428170B692E36DE0754A970A857FFA8FBECBFEFF3D1B80007F9CDEC21F";
    attribute INIT_14 of inst : label is "DA7BA7746DA62C679F3E4664444444446A06E156AFAEA037EBE5FF03E779DEF3";
    attribute INIT_15 of inst : label is "0BC880E3742DF69DB7631FF18B7276D653AC542A403454742A946AB57EC93A09";
    attribute INIT_16 of inst : label is "8A85500D151D0AA51AADD24AF7F966F27B7FFF39ECD3AEFAE7FE9CE127F91F51";
    attribute INIT_17 of inst : label is "3E3E02431E85028542A957F6F7FCEAF669D77973FF4E7093FC8F28E187CD4635";
    attribute INIT_18 of inst : label is "C3FCFA3FCF43EAFCFFFA7FFBE240025FFAA20DF3263C8F9047A0E1C011000000";
    attribute INIT_19 of inst : label is "4D36D274E8CC999A6C5408FE13223BA3BCC619D456D94D55019D8C80FC4FFD7F";
    attribute INIT_1A of inst : label is "BB4CC286E6741983FC6DED3A47D209A472F26789E01F66C2624281216A95771E";
    attribute INIT_1B of inst : label is "D5043B5A4613846C09F0086944ACD2D4FE96EDC4E514D54A8CCC22388B541F3C";
    attribute INIT_1C of inst : label is "719C76E24A491F29F04118C631B1890C48CC0718D6C142F80232D2585470A54D";
    attribute INIT_1D of inst : label is "DC70CCB1FE378D05A58F6C9E3632CC8D9F50FCFC17B7B50E9082AB871514DBE6";
    attribute INIT_1E of inst : label is "E297E9A8602206013E5D3DE3121CB6A5A34D4CE63B29930F7A965AA8E8C7CA82";
    attribute INIT_1F of inst : label is "FD663221447F12E4B269B600D5B50BB4A0C6A2AEA0326E3E75544A2A3BAB20D7";
    attribute INIT_20 of inst : label is "FA975C5966E33537CA372D6AE4ABA9793C7865BF7C13B4E890C9F33B43F491F4";
    attribute INIT_21 of inst : label is "CB5625BF8AEBBE18017A7BEEFE004C87B04755A4F120256F2B4FDD7C92941119";
    attribute INIT_22 of inst : label is "24509102706281820615512FD78C5296A3AD313050DAFC7F3332513A263B0049";
    attribute INIT_23 of inst : label is "091024409C103040C103040EC0C100240B0200181400040010383830382914AE";
    attribute INIT_24 of inst : label is "0103010281018812244881182060C1820541C1D000000040C040C040A0310244";
    attribute INIT_25 of inst : label is "8A56000000080808080804001C48816204E0C10B040FC0EB9010004081020503";
    attribute INIT_26 of inst : label is "B154157681820520948000000206020602050203102450911820628182A0AAE4";
    attribute INIT_27 of inst : label is "66B09CDD99961DBCA4CF408102904A40000001030103010281008B142C522C50";
    attribute INIT_28 of inst : label is "F1D9CFE9BDFB5DE604022025F7C98DFBE0479D313B74ED73EAE2EE3C3CCDB1B6";
    attribute INIT_29 of inst : label is "2A96811EFDF9CA2AFED7E73BF7DBE4FBA7456497ED779C674CACE5EDF38E6ECC";
    attribute INIT_2A of inst : label is "D9BAEB82008385E2E59311104D3DABEE786D35B312592D4970882898D15E9849";
    attribute INIT_2B of inst : label is "1DC449400B352CD43340C51D3F0CF8F8C202EC47389C8D40ABA3CEE4D9FF477F";
    attribute INIT_2C of inst : label is "B0969E1E1555555411195B15CEB382C86EDF31DFB74FA7D3C6F3800B00012BDD";
    attribute INIT_2D of inst : label is "A55031E117A7EDD7DFD0E25A58C0801D9C9B4D8D18AAAA0222BEEE464CA76012";
    attribute INIT_2E of inst : label is "67BB6B3B3C79D221E7768EE3B37233744A1B3C15A9C15FFB3C30CCBAA089C1D7";
    attribute INIT_2F of inst : label is "3FD96B874D27F1F6CBB6593C24C79ED92740DBA610EDEFC4A1C5B9F1CC2DF2FC";
    attribute INIT_30 of inst : label is "FF81B77DF222A08288F39C5924E844C1985A3280D528EA436D76ED058ED3B4C9";
    attribute INIT_31 of inst : label is "00787E7DB001010000370000040103F6E6001806002FD40000C0000B64BF8007";
    attribute INIT_32 of inst : label is "002002AE2000200981997178010140CDF8098001028072D940000333FF965A00";
    attribute INIT_33 of inst : label is "FC19E3E0E0010000001BD0200DEC20B64AA00068199AB8D08002BDFCFF909440";
    attribute INIT_34 of inst : label is "1AA1C6E400A940004E4000034A8CECB682131001F76E3470004900342DE80010";
    attribute INIT_35 of inst : label is "BFEABFED84F0A08000F725BF80000029E96DF802400955400003FFC0C4978800";
    attribute INIT_36 of inst : label is "880340AA93D407F82FF94FF297F32BE455D9AA33C007E82BF1455280030004EA";
    attribute INIT_37 of inst : label is "CB082CDB33100382E3193877A75B5A6105D267400B4D218D7B59BE0DB3D10025";
    attribute INIT_38 of inst : label is "0F6EF3275389C4DC7327A757CC7371339CD9CCD98D0A8142255165435712084C";
    attribute INIT_39 of inst : label is "3CC205BC6D203264FA602C8810387644CB3A3440C9C1389F77AE6196644C1B2A";
    attribute INIT_3A of inst : label is "BD28F7B34E7D73FF4E7093FEBEFB7C12E8AA11B14EC53F14FDA739504A0016E0";
    attribute INIT_3B of inst : label is "BB4745B6B6E85760CDCECE8C1CCC0417801A334338A5CA71C68804E20A957C89";
    attribute INIT_3C of inst : label is "658C800C86AE90BF8B6577019502143D0A2902A244D934BEED8FE8EFD9B654E6";
    attribute INIT_3D of inst : label is "DE9B7A7BABEACAEFA8A3E0EAACE274BEFD5F7DF7DCDDDEB17FC5CBD8B97BB6CA";
    attribute INIT_3E of inst : label is "BD8FF982FEA33C2561F757EDDDCDDDC4F7680473954FE2E52B8B5DED63D6ACAE";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "5451854015E77F9F1404C2E96844476A02203D75C51FF0897001E910214A4500";
    attribute INIT_01 of inst : label is "0F4390D0EC3E75CE33BC019C04CFB4C30F8AB08A1559442E2497080648061820";
    attribute INIT_02 of inst : label is "0307018380C164C9333438C861C2BDCEF984A7739EE3C43F8C5C9000969A4802";
    attribute INIT_03 of inst : label is "19B47831E500C05557D704090E21CA0E21D285521D12153681E17488011C060E";
    attribute INIT_04 of inst : label is "AB995A0AC4060064CE2DC3AD2F61603AE944C21A2D4613B09D96394B0075173D";
    attribute INIT_05 of inst : label is "852281B13E22070A841C2BA2118500474AD7B7AC0C73C665F3536C05CC98B418";
    attribute INIT_06 of inst : label is "1A0C18A3D1C44429613A1C80422022203204F188090C815577550846A64303F3";
    attribute INIT_07 of inst : label is "E80569520E80AD2A40E8A14AA26D200B8403D4E34304D4D4E0020442882940C8";
    attribute INIT_08 of inst : label is "8175F865F46643880444B78365D0EA5D00F40283740694A90CAD7F4052A4A0AA";
    attribute INIT_09 of inst : label is "99999C0320807C3815D3E4083A1C4B6683FD55603C00050213272037AA32049A";
    attribute INIT_0A of inst : label is "15001089524409C2444895200440A40944885220468001911919191911999998";
    attribute INIT_0B of inst : label is "04C8204020112200099301624480108910C964824B0040895100548950001489";
    attribute INIT_0C of inst : label is "1000040041001001017A4D8079544A020264C010993014A2544015324A09C220";
    attribute INIT_0D of inst : label is "0000900100100100000124100000100000000004000000000000000000000000";
    attribute INIT_0E of inst : label is "00800000800800020020000820000800000820800820000C0080002000000000";
    attribute INIT_0F of inst : label is "0041001001000040001000040008208208208208208208001041041041000044";
    attribute INIT_10 of inst : label is "49C71800D9115E8101B6005200A40100422505E1962000400410020020800824";
    attribute INIT_11 of inst : label is "50D182A21B1510D182A21B1526682EB410657EFFF3F27D1F004C60C08300007A";
    attribute INIT_12 of inst : label is "C07E0B681314B2C1041FA04C301418869482C2603008040601691E2C2C262C08";
    attribute INIT_13 of inst : label is "B087190280D251B1A6A30073460F0601239947A643CEF50C03100238A92D0019";
    attribute INIT_14 of inst : label is "8AD73094DA9A5B619F1F2624444444456200E0C0244EA04D01ACFD07E358D6B5";
    attribute INIT_15 of inst : label is "8ACF4829101926D9236B1FE2EB752C091112EA7CA4104210180D060120ED8219";
    attribute INIT_16 of inst : label is "5D4FA9041084061349841B62619E26D2BF45F1012CCF8A8845B5946A71BC91D0";
    attribute INIT_17 of inst : label is "D47661104203118CD462123E53D4049667C52822DACA3538DE45686FE498B022";
    attribute INIT_18 of inst : label is "C3E8F53C4F03FEFCFAF578F9E140015FC5D80D80001E4C304313C78843734734";
    attribute INIT_19 of inst : label is "CD36D264454A95D46610887C7321B3154CFBF5B41BE9E7F5078C8A0824CC8E2F";
    attribute INIT_1A of inst : label is "33E2F58EF4685FA5F884EC3A76CA099460F0298BE8F648C57B898CA326B16794";
    attribute INIT_1B of inst : label is "F3AEF80A478199228D5E1C794D0DCAE01E5624E49D18D351CEEFB220AB3598EE";
    attribute INIT_1C of inst : label is "3BBE6E8E3C348BD0BEC01431087745AAE58CF3BDF9E87A1C006D392FD02984E2";
    attribute INIT_1D of inst : label is "2E63EE20213A75A2F13E78A9BA758AEEA93573501BCAC797155DD43DEEAAFBF3";
    attribute INIT_1E of inst : label is "79B24598280C6780EC2F9C820296DE71123ADDCCBEB919BE518870FC78F58518";
    attribute INIT_1F of inst : label is "6FBAAAB5C46FC25CD775F7289C39A8E0BDE75EF7759FBDB6BB7EBBDCB2547DE2";
    attribute INIT_20 of inst : label is "9DD3C81D257BA79261AB673A47891C37E91FD6B7980B66CA0A98D519E13C70DC";
    attribute INIT_21 of inst : label is "5CD6F440E9E48658FF1EC0E20304F8BF3F4BA73CF5235D600E148FA2E9C20CB8";
    attribute INIT_22 of inst : label is "244881027060C10206C5514113DE855A4E34C8BA38F04EA4A2B238B22F365BAE";
    attribute INIT_23 of inst : label is "8812244884183060818306095515241C0204080C040004080030181010180CA6";
    attribute INIT_24 of inst : label is "01010100810289122048910830608183048A0A30000000C0C040C040E0112244";
    attribute INIT_25 of inst : label is "0652000000180808080804080C48910204E0C182040C5550302040C081020701";
    attribute INIT_26 of inst : label is "3068A80180000303958102040E0202020201020710244881182060C10245415C";
    attribute INIT_27 of inst : label is "7CA28C2A298B18B24040C0000180CA40810207030103010280008910244A0C10";
    attribute INIT_28 of inst : label is "21E36E49B95304C9300228B91049AB82C8AA8E292B54A4F2CE28EFAA7DDDB7B6";
    attribute INIT_29 of inst : label is "385D800130114137D43EC229508024B32707B4C54C13206BEFF1B73959CCECCE";
    attribute INIT_2A of inst : label is "F89445C39042743824BA1110486F3886576F33B3C08240001BE1A8B0A0FA14D9";
    attribute INIT_2B of inst : label is "0D02A2822B75ADD617C85F25591458988308304C631706905CE2C76CDED9E692";
    attribute INIT_2C of inst : label is "00F707E00000000C114DFB9F27206928CB9464474F43A1D08EFFFFFC0002BED3";
    attribute INIT_2D of inst : label is "C008141150E099B186286C0E0FB1883EAF09C6BBE000010229F4A163EF456A1E";
    attribute INIT_2E of inst : label is "E7B361561BD8BC39B6358D635FB6717CD54B0277E92500954666F9AF5A888C98";
    attribute INIT_2F of inst : label is "FB9CC197783F713AF9661C5C6DC5A55F1298862A93EC09A768BD1A95FDFA964F";
    attribute INIT_30 of inst : label is "000022A2828202000DA9AB248FCD2AEB15D634D08DFCCA6239025884C4CB3789";
    attribute INIT_31 of inst : label is "00D0566004000080200400000C03308000000A0A0180047802200004003F8000";
    attribute INIT_32 of inst : label is "002A058020000466024001000000110000080081020018007F000888FE400200";
    attribute INIT_33 of inst : label is "AC184008000140001800480001E2204002508060100200100102A940F0009400";
    attribute INIT_34 of inst : label is "3AB5C00100003A80830008034A869000C00010000000040010081084002E0000";
    attribute INIT_35 of inst : label is "554000100400008150C4002002000055E00100020008AB000003FFC02000F000";
    attribute INIT_36 of inst : label is "00000000080030006000D001A807540CAA195532AA05540AA805500004444215";
    attribute INIT_37 of inst : label is "8D7C249B2F502CC2479CB24F06B2972FB49A56C83A0BA1257B591198800A0000";
    attribute INIT_38 of inst : label is "0F6D7F27CBD9F6FF7DB7B7A74FD53DBBEEB9CCCDCB598CD43F117B1312DEA566";
    attribute INIT_39 of inst : label is "A4DF43806DBA3E45F70A1D98103C0E6AE1E3207DC9FB3EDB6BC6BDC3C667D9DF";
    attribute INIT_3A of inst : label is "FD5C24B33E0422DACA3538DEAF899C0AC803115C50F143C507218668E0050E05";
    attribute INIT_3B of inst : label is "3B676FACFEE9B83E9DDCC42E5E885100410793C71CE3CE79347A31CB46316C49";
    attribute INIT_3C of inst : label is "AC58AA6208A0AA023087DF439201FA16FD08003EE78A9E87158B3ED2F86E8628";
    attribute INIT_3D of inst : label is "4110453890A404071413828042042A02002082082275D4460018582103044204";
    attribute INIT_3E of inst : label is "084BC188E2412D22657620EDDCDDDDC563380061BB47C5E515146082842A4240";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "1AB5107208EC0244D4B8B9806C45DD3E0AEC0C107F95446A35402CBA054239B7";
    attribute INIT_01 of inst : label is "08EC550A961D2C398A0A15045543BB2111907767003BB6074A85DDA091287E04";
    attribute INIT_02 of inst : label is "0103008380404110452CA291550B3842946C2410D3082E09C31AA4924864BD82";
    attribute INIT_03 of inst : label is "0882A75A9685ED630DF20A50C3752D437534EC1356ED0E09D875125D010C020E";
    attribute INIT_04 of inst : label is "26524224F2FED6CB9C019394DC1240DA2608420F9794DDA6EC4E9C532F4F144E";
    attribute INIT_05 of inst : label is "40100B804F0504012CA92B0814844492D284C75A800000A125425D291696B891";
    attribute INIT_06 of inst : label is "E341200297948CC0CA39082211505240564173D340880680BB3AADD88B57FF0D";
    attribute INIT_07 of inst : label is "8A921520DAA242A4158A04A908241009A402F6A0D2A4D4D4D1152EEC56B59512";
    attribute INIT_08 of inst : label is "11948DD9C545508AB41A0C942F169BF166D50239C5490A90754A1C512A411A02";
    attribute INIT_09 of inst : label is "080082D6A95554A054C3D508228362C5D60A82928A800EA20DB30CDB5A6A6DA0";
    attribute INIT_0A of inst : label is "0902105A920088820081A10042D4000800494020418000088088088800080009";
    attribute INIT_0B of inst : label is "045A02108403468D20344BA02D52E000B4492D806000001B0D02101B0C02105B";
    attribute INIT_0C of inst : label is "100000000000000004DB0D12E900D200040D12A00344B816C34084145408006A";
    attribute INIT_0D of inst : label is "4100924004004000014000000104000104024904104100024900104100000000";
    attribute INIT_0E of inst : label is "2002082002002000000410000082080002080002082000282080000210410410";
    attribute INIT_0F of inst : label is "0040001000040001000040001008208208208208208208200000000000041040";
    attribute INIT_10 of inst : label is "A08342CDC0603C3230302E653DCA7396E548E51A50E000410410820820820820";
    attribute INIT_11 of inst : label is "8C0D422B5450CC0D422B5450D334B289A9F28E01C8710E830003E4140B01A898";
    attribute INIT_12 of inst : label is "FF716032ABAC55D5A1C2AE0A07684AD14E0A170B8542E0702A4AB92CA3A6A042";
    attribute INIT_13 of inst : label is "A45AB01CA2293C7450786A468D18803A57023B8009C632813B400332340E2541";
    attribute INIT_14 of inst : label is "96905D29474F0533AF7E01A444444444E80660054A8E0DB283A13D00EF3BCE73";
    attribute INIT_15 of inst : label is "A420AD0381C05B76CCAF94AAC8CFBC1DD11B414256889301C2E0702A4F826CB2";
    attribute INIT_16 of inst : label is "682855A224C070B81C0AE0949C392064BC11C474A053442213A8A5A1C2380465";
    attribute INIT_17 of inst : label is "034377D4F0385C2E0702A5782B8A645029A21509D452D0E11C02B21AF799DE23";
    attribute INIT_18 of inst : label is "03D0F8BE0FC1C0F0F4F8FC7EF520152F88010E70D81C039090AB162DF1C20000";
    attribute INIT_19 of inst : label is "32C924DEAD1B316D3A02B6154CC58EF8E4BCE12A89994578BB2D8C6945550E8F";
    attribute INIT_1A of inst : label is "A938B123C15412832AC5802115E953D2FBFDB82ACD25BDAB60282A2BA02A5452";
    attribute INIT_1B of inst : label is "319A8A0901118803565B5D342202E9E28F4F40414B7DD0146CBB81539B01D34B";
    attribute INIT_1C of inst : label is "0A7859BA4E4E93193094252DAD316D5B698C9B9EF5F562994042FC52B41920F4";
    attribute INIT_1D of inst : label is "42B52260090A45B0F9923E4932652888C9044060120317E104012051C0842715";
    attribute INIT_1E of inst : label is "125269394D0489514E0FCACB41A2BF79A34C28E8E77852121BB6BC021484C229";
    attribute INIT_1F of inst : label is "47223333FDEA5036C2B6F751580DAAF877210441889588B50E2411A182A4A032";
    attribute INIT_20 of inst : label is "8432292C034587D2651A14A143002CA6C12C127414127B2509048411F9120282";
    attribute INIT_21 of inst : label is "0B084502AAE0062000188061820DD2E9101087DE3AA3CC8007848224C8C95DE1";
    attribute INIT_22 of inst : label is "244891223060C18304D4414103DC8210168501297D7E42241DCA7D219D57AF08";
    attribute INIT_23 of inst : label is "8912244894183060C183060C5555269C070204080C000C000030101818180CA6";
    attribute INIT_24 of inst : label is "0101010180018810244081382040C102060A2A30000000C04040404060512244";
    attribute INIT_25 of inst : label is "065200000018080808080C000C4891224460C18306091555502040C081020701";
    attribute INIT_26 of inst : label is "3060AA8A8000030194800000060202020203000310244891382060C18355015C";
    attribute INIT_27 of inst : label is "4E966BC793D0282C40F540000181CAC0000003010101010181028910244A0C10";
    attribute INIT_28 of inst : label is "280C9004908D46B991211540A824899139B84A7C51A147450C3EBB277670D01A";
    attribute INIT_29 of inst : label is "E1027FE1980CBAE92A492990BA201B4891600242351AE235BB0648108D6BB16B";
    attribute INIT_2A of inst : label is "138E80FCF3F600280C209110412630DA4DF6981A52C96549692084484D21EF27";
    attribute INIT_2B of inst : label is "090965C20D35B4D6534945294A1550908A6050544042345A540A011152124584";
    attribute INIT_2C of inst : label is "B562A0000000000208B0204043B4371540820002D341A0D029FFFFF000000491";
    attribute INIT_2D of inst : label is "000506AADCEC8140C359CCEEE94BB406273BDD3400000041144AD0B9BBB2A9AC";
    attribute INIT_2E of inst : label is "9A6C9E0D96B4214A9CC94A5290A529CA551D54E8D690002C884090AA0C52E41F";
    attribute INIT_2F of inst : label is "48371A851309055290CC87401214285271E50819FB128A210C6B148359488443";
    attribute INIT_30 of inst : label is "00005F7775DF75DDD04A024924ECC4A4EC9E66CA153F0A58314363EC09425128";
    attribute INIT_31 of inst : label is "1050500200000180278400000A0A78C000000802618000700008000C001F8000";
    attribute INIT_32 of inst : label is "0408110000800111842000180061582300000411080008003F00055500C00000";
    attribute INIT_33 of inst : label is "290060000001500F18000800497810C00024054011C400000022AD50F0002800";
    attribute INIT_34 of inst : label is "0000018000002AA90100000040033000000002AAF880000008A8020400070000";
    attribute INIT_35 of inst : label is "BBAEEEE00000008000040000000228FDE0000000144DF2000AA9554010007100";
    attribute INIT_36 of inst : label is "4888800000000000000000000000000200040008007000E001D003AAA71406BB";
    attribute INIT_37 of inst : label is "68E7610AE2D2AB761454A8A8E5CCE81CEC2945CD6B29CAED6DD24B1875608055";
    attribute INIT_38 of inst : label is "A89D4CE7C278E4A24C0464E202B30C2261A52B3E38542E050933481CA56DFFC1";
    attribute INIT_39 of inst : label is "64B96E82902144B56CE9132A14251143126CB29D39EF1C94EA480E24D961C702";
    attribute INIT_3A of inst : label is "3A2142814DB109D452D0E11EAEC05C29D292CD1744FD13F44E5E1B0DE7FBBB97";
    attribute INIT_3B of inst : label is "0D94E0814997B92B733BBB89516851AD1C05854452A254A588561180803A5F20";
    attribute INIT_3C of inst : label is "0448CC80E048C982200DFDA07553B734DB80500A448612012A2848B01303CA8E";
    attribute INIT_3D of inst : label is "40451038800020074043840408880042000000000055FD001000080201011220";
    attribute INIT_3E of inst : label is "A0273807C8281E1100B0146DCDDDDDC4E7C5F406125154750040408008000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "17C80440B5C56BD72858B19EFE66646327304FBEF0900A42B941063609513425";
    attribute INIT_01 of inst : label is "08C91522970DA51923CB096C25364A3131931AA8018D5002C36D991093B9AD01";
    attribute INIT_02 of inst : label is "340C1A060D020102042B24925322B6C214CCA5B0C3183C498658E6DB69259902";
    attribute INIT_03 of inst : label is "088084421479C95966460390F2652D7265348E02564D6ED19E65131B04206810";
    attribute INIT_04 of inst : label is "3652511D98C004F518CB97A1802642BA8E18E00994809984CC033AF2194C5D88";
    attribute INIT_05 of inst : label is "2984458646483016F86D2ACD4220501A4014ED0A550451052808484810C07015";
    attribute INIT_06 of inst : label is "06C2A76697B5B95A5AF0E9348A030619120BF7E0106931B319109A911B67FFFD";
    attribute INIT_07 of inst : label is "10F296AA730E52D547105CB544240202008F095CE490C0C0D8254CD864A5C038";
    attribute INIT_08 of inst : label is "11900F25885180E3C14FCCDCA02096820D180E9B08794B550452B8872D545F1F";
    attribute INIT_09 of inst : label is "000803BCC049474E85EB982DCC032A54E60800178C4003121242129D184C7825";
    attribute INIT_0A of inst : label is "0B000118324018A240158B2008C008880158456040C000080000880880088808";
    attribute INIT_0B of inst : label is "05181C2C8023060002B141108C100420B0490C80400001580B00411802000158";
    attribute INIT_0C of inst : label is "00410000010010410064AC504C08C10000AC544C2304011602C0004640022060";
    attribute INIT_0D of inst : label is "0100000100100100010124000004000004000000000000024900104100000000";
    attribute INIT_0E of inst : label is "2082000082002002080410082082080000080000082002080080002210010410";
    attribute INIT_0F of inst : label is "1040041040001000040001000200000000000000000000200000000000009048";
    attribute INIT_10 of inst : label is "10838420C2008C080430C1D08084234A92084412D53000000400020820020800";
    attribute INIT_11 of inst : label is "8AAD7734A6548AAD7734A6549D66965D66E07C0F83E07C1FFF80780223FC111C";
    attribute INIT_12 of inst : label is "FF70002A628490E2B0C16E5DA8402C9490529A4C26114884D00A38AD2E715411";
    attribute INIT_13 of inst : label is "A2029221BC9381112502C35214291450470403C105C73042030FFC30400C0881";
    attribute INIT_14 of inst : label is "0214D929569815A9EFDE082444444444608C4A8A08BFCBFEA1B23DF8F7BDEF7B";
    attribute INIT_15 of inst : label is "1CB9894D22149B7258AB1452A8CA75C4578C887844AA8CA21148844052B44A92";
    attribute INIT_16 of inst : label is "910F712AA328844229154D108938A1483C81E0823063810409A0C63008382054";
    attribute INIT_17 of inst : label is "8C4C6A20244221108844047903C1011831C08204D06318041C102A52CEAC44F1";
    attribute INIT_18 of inst : label is "0FC3F07C3F3DC0F0F0F07878F81FF80FC0047C0401DC101052E20C1925E69A69";
    attribute INIT_19 of inst : label is "12492DCD940D756F1B14B20A42200652F2B10578C0345FD6352898A006550C0F";
    attribute INIT_1A of inst : label is "0B32B648CB47524114E790A414C0E781E0F0322AC924BE99690D30AD74D0405B";
    attribute INIT_1B of inst : label is "6F01E0078B5E356CB0F6CF3111D1C0C10E0610494931DA6A6EBB0551BBA6954B";
    attribute INIT_1C of inst : label is "D8794BD3F9F877C77DBFC21463751F686E4F2718C8DE941FFF9F9BF6975F3A6B";
    attribute INIT_1D of inst : label is "B71370250B5AFE8BB692AC2AAFAE6ABBAACFA3A3ED1D09BBC040450A0D4C6715";
    attribute INIT_1E of inst : label is "B66AAA6E1FF879FD4AB996B94DE3F636AD5534A1AD30D6529EDD9BBBB7385660";
    attribute INIT_1F of inst : label is "A5ABAAA16974DC94D61046FE256A50B6517240DB44508BFBD868E3464E40447A";
    attribute INIT_20 of inst : label is "0E3529070B289DAAC1D994A35B38481EC9060C3AABF4B2AC0405402B65528542";
    attribute INIT_21 of inst : label is "5903184084C687D9FF78007282A1C6895F0DFDBF3C691C31D335B7AEFE85F304";
    attribute INIT_22 of inst : label is "2040810210408102056AEAFBEF9C94218A6303405B5957AE1DCF5B4DDBD3352B";
    attribute INIT_23 of inst : label is "8912244894183060C183060EAAAAC66C060408181C081C000010303030380CA2";
    attribute INIT_24 of inst : label is "010101018000881020408108204081020575D5F000000040C040C040E0512244";
    attribute INIT_25 of inst : label is "0E5600000008180818081C081448912244A0C183060EEABFB000004000000101";
    attribute INIT_26 of inst : label is "307D575781020701948102040A02020202030001122040810830408102BABBEC";
    attribute INIT_27 of inst : label is "4E5B6B32D7B9A0268599C0000181CAC0000001030103010381038910244E0C10";
    attribute INIT_28 of inst : label is "2303285377020099625CCCCA2A53720E18909876E4CB928E7ABA9972B6221242";
    attribute INIT_29 of inst : label is "21908021A0270483691B14E538441B83870E29BC0802609899C1963707298A39";
    attribute INIT_2A of inst : label is "16E7B641944A2831963919986473EAEAE56242427FEDBFEDC7431327376C0409";
    attribute INIT_2B of inst : label is "A1044108C75CBD7675CBDF609826C10306C000E41AECC8D9A81A9B0952005580";
    attribute INIT_2C of inst : label is "EF19E00000000000E6736CB69B5D2A1868D0044254221108C600000015544C11";
    attribute INIT_2D of inst : label is "0004852904B48F210252D84B4E2EDC22725F6F620000009CCED15498998490E3";
    attribute INIT_2E of inst : label is "1A6DB265B69D7A4A1D8BCE7395AF395E4A93E456AC1200846B0A975AA312D9F0";
    attribute INIT_2F of inst : label is "4A7632D596494D0A965DA6841B340152CCD5A859D8368A6B9B2958B1CB4AAD56";
    attribute INIT_30 of inst : label is "007E1F5F5FD5F57D785A56FBADE86500EC9BAD065BED1F58E6006696686A996A";
    attribute INIT_31 of inst : label is "00050664000000802FC800000AAAFC00181100A09000000080020F00001F8000";
    attribute INIT_32 of inst : label is "04016900011504447840001800282B1200030000541190000020200000800000";
    attribute INIT_33 of inst : label is "01660000000156BF8000040802228C000050005057E00000000002B820002804";
    attribute INIT_34 of inst : label is "0055F90000002A29E200058282A120007E00000501000180000A2FC800011100";
    attribute INIT_35 of inst : label is "BEAFAFA000F0008007C8001F800445244000FC002220A2000002AA8020000800";
    attribute INIT_36 of inst : label is "060A8C00000000000000000000000000000000000000000000000000000148BE";
    attribute INIT_37 of inst : label is "2A74A02C6A54824A005224A844EC6CCE9404B5CCDE9732836DF6F4A9AE488704";
    attribute INIT_38 of inst : label is "289D4C6B220BC8A44E6464D312954F2271A1282E3A31188E49374A3884480460";
    attribute INIT_39 of inst : label is "A29CD4E08241449564A5412952A4D14F1860BC9D1AC17914EA594E30C179C544";
    attribute INIT_3A of inst : label is "3C0208C18E0204D06318041D4E841FC0C102A5775E0D7835E00C6A080005520C";
    attribute INIT_3B of inst : label is "8D94C8804C97C2613929B12C412801448800056052A0D4A51253E3A404704C04";
    attribute INIT_3C of inst : label is "050A0000008000000005F7A87BFB81BFC0D7FF42D5F77103A6680A90160A410C";
    attribute INIT_3D of inst : label is "4045003800000007544380000000000000000000007DF40000000A0001400280";
    attribute INIT_3E of inst : label is "02130210C1104C088830886CDDDDDDC4B303F9081030A5431004008200000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "D6ED835020A7D65CD868C669044444F614213441358566C94F05ACD2201B6DD1";
    attribute INIT_01 of inst : label is "0E23C298426E31C478270E103088DF821CBE5A390F2D121A4693C47248042D60";
    attribute INIT_02 of inst : label is "62302110188D25CB761BD66323BC313C4F24244F49DC392C980F300496924402";
    attribute INIT_03 of inst : label is "99BED06343E6E404104104D9C9B087C9B09FB427091B13946930666918C08440";
    attribute INIT_04 of inst : label is "C9091C1AB34A52364221F3E3896F039F9CCDE839BCF201900DFB19381EE60467";
    attribute INIT_05 of inst : label is "EF0787F9666B636E6860821A4D2054C308471667DC400241D203647DC989BFDD";
    attribute INIT_06 of inst : label is "D268F896C1C04025253F0DC4E06464246024381FEF8DC5B33B33F884243FFFFD";
    attribute INIT_07 of inst : label is "48D94C9BD48B299371483664FD92CB66840FEEF37FF6C6C6E03FE2489B184688";
    attribute INIT_08 of inst : label is "92E2F551B46A4366D37BB3047292E6A92EA40EF0246CA64D93298A4599373BDB";
    attribute INIT_09 of inst : label is "80088ED521FC1CA58040A43A4A1DA3067CA2AABEBF9553E4BA5717D9E91268B0";
    attribute INIT_0A of inst : label is "0B48015ABE801A268011A34008D0089A015A4568014800800888080000888008";
    attribute INIT_0B of inst : label is "055A54BD802B5690023440008D100020B4DBADA4C000011A0348011A0248015A";
    attribute INIT_0C of inst : label is "100104004000004101FF8D144008D32400AD50002B54020680D20046D0022468";
    attribute INIT_0D of inst : label is "4000924004004000000000104100104100000000000000000004000000000000";
    attribute INIT_0E of inst : label is "0000080080082000000000000000002082082082080000080082002000400000";
    attribute INIT_0F of inst : label is "0041001041001040041001040200000000000000000000201041041041008048";
    attribute INIT_10 of inst : label is "EF7F7BDFFDFF7FF7FBFF3E5EF739C671882705E9075200010000800020800824";
    attribute INIT_11 of inst : label is "1EF0828B59031EF0828B5903200817801BFF8FF1FC7F8FE3007FE7FDDF03EEFB";
    attribute INIT_12 of inst : label is "C07FFFAF3C3206684A31715CBA10D666859CE0703C1C4E0711217F37FA02A08F";
    attribute INIT_13 of inst : label is "BDFBDB8226C185D9810BC621428647112FFBFBBEF9FEFFBDFFF003FFBFFFF77D";
    attribute INIT_14 of inst : label is "0847239C1E009F219F3FF7E2222020202605C0E025ED99EBE1ADFD06EB5AD6B5";
    attribute INIT_15 of inst : label is "72ECF671381BE489230308590B7010124124670CFB3AE5B81E4E07013A491BDB";
    attribute INIT_16 of inst : label is "8CE19ECEB96E078381C1D24261FF3E77BB7DDF7DAF5F7EFBF7BEB5AFF7BFDF5E";
    attribute INIT_17 of inst : label is "EB2BA2C8C70389E0F27112F6FBBEFED7AFBF7DFBDF5AD7FBDFEFAF6382092424";
    attribute INIT_18 of inst : label is "F3FCFFBFCFC1FFFFFFFFFFFEE7E007EFBFFB8FFBFE1FEFD07B3C64EEC073CF3C";
    attribute INIT_19 of inst : label is "EDB6D224C5879190CC56088B376231051CC711873668BD5CD1848FB266031FFF";
    attribute INIT_1A of inst : label is "3BC0C88434281D22164CEC3B62FF19FE7FFFA380A6B24C8C61F5C0397711278C";
    attribute INIT_1B of inst : label is "9106A80B24C2F064D9B07DBBC4ACFFFEEFFFEF658C860BCB80C4736403BC8D64";
    attribute INIT_1C of inst : label is "258464E00001152152F5108421B909886A7C077BD4974A0B43329A18C8A5856C";
    attribute INIT_1D of inst : label is "885C84212B22C4D8B6D86D0A623881888A781010109095A4C33C31E2666632C6";
    attribute INIT_1E of inst : label is "C392B5EC75380650638DB22DE23CB6B6F1E7C6B0B1B701184AD45B4C48CB7330";
    attribute INIT_1F of inst : label is "E4322221685F234A33619CD4D43D08B5DA9232C433100A2E25672B391E303382";
    attribute INIT_20 of inst : label is "9387C01894E36DA2C227631A04A438713819022E3C3BB5D80019C0BD617CC1CC";
    attribute INIT_21 of inst : label is "CD04A40052A18AF0812E00AE83F8480C30A20D84303504432B65892DCB875150";
    attribute INIT_22 of inst : label is "20408102304081020445011043ABD318C2319FB019D8582FE21A1ABA257B7488";
    attribute INIT_23 of inst : label is "081020408C1020408102040900011FFC060000080C000C000010101010180CA6";
    attribute INIT_24 of inst : label is "0103010381038912244891383060C18306202030204081C04040404060310204";
    attribute INIT_25 of inst : label is "0E5600000018180818081C081C48912244E0C183060D0015702040C081020703";
    attribute INIT_26 of inst : label is "204A00038000030194800000060202020203000310204081182040810210540C";
    attribute INIT_27 of inst : label is "71A2840908923191C25FC0810380CA4081020701010101018001881220460818";
    attribute INIT_28 of inst : label is "964AF22C8CFF046861C7376DE20C19B9E8ED974D9B366C79EA024428388D21A4";
    attribute INIT_29 of inst : label is "29978031EC78C5BC96E4E71AF380247EBD591653FC11A5E766657B0CFAC6FED6";
    attribute INIT_2A of inst : label is "481041221C421410E58F11104829A8285069A1A38080094059970CD8DF961879";
    attribute INIT_2B of inst : label is "AC070071382740998274018E03861E1C01D266603440403FF9E0C4641CC90632";
    attribute INIT_2C of inst : label is "A5F688002EEEEEED39A99679C4B1E23B62C7A0C5BB81C0E0000000003BBBB2C1";
    attribute INIT_2D of inst : label is "0EBFB5FF04340DD347F0B05B58DAD41DC81269CC015FF5A73726C7EF66E9E0BE";
    attribute INIT_2E of inst : label is "E112431228C685A322242148523884610F117FFCFEFB01BBBC30EDF5566858DD";
    attribute INIT_2F of inst : label is "6388C106682C7030E122180B24C0841D024E58264DC98184F08C12A56E60B858";
    attribute INIT_30 of inst : label is "00000288220882208CE5290414E84EC312CB1A84C02C6A72290238868683A681";
    attribute INIT_31 of inst : label is "002D298003F10485200000000A0A0000000015556800000000AAA0C0001F9550";
    attribute INIT_32 of inst : label is "055090000000111006000060A02028E000060000100E000000444111FC000060";
    attribute INIT_33 of inst : label is "2918000000015503800004040A28700000504050500000000000028700000000";
    attribute INIT_34 of inst : label is "0054E0000000282A10000022808F00003E404004F80003E000AA0FC000000004";
    attribute INIT_35 of inst : label is "40055000020024801800001FD01001660000FE002002A0000002AABF000000A8";
    attribute INIT_36 of inst : label is "00A2800000000000000000000000000000000000000000000000000000000015";
    attribute INIT_37 of inst : label is "850C26DB030FADC2670812C31612122184D2461FBF1F6C857239365807C00000";
    attribute INIT_38 of inst : label is "CE4061061B1086CD6337165748C061BB1C0A848183C1E0E02C80638A12B20444";
    attribute INIT_39 of inst : label is "20C2C5276DA37240523BCC8618337C20C3021346418210DE0324A18604247033";
    attribute INIT_3A of inst : label is "BBFDF6BD7DFDFBDF5AD7FBDEAEFBDC3FFEFBF013044C113045A53D8342031484";
    attribute INIT_3B of inst : label is "7263046C9669FF5F8CC444071E835027FA52106708311E10F4E8607307112FFB";
    attribute INIT_3C of inst : label is "05080000000000000080A07B94D3F328F9E9D3A624099484F18320C6486E4461";
    attribute INIT_3D of inst : label is "4000003800000007000380000000000000000000000A8C0000000A0001400280";
    attribute INIT_3E of inst : label is "FDEFFDEFFEEFBFF777FF77C2222020208BFC06F7D9C8B1A94000008000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "546C81503083541088480822A40000741C0110A2B58550498F05AC50040A2543";
    attribute INIT_01 of inst : label is "8406821000781180D04708282194DF1708BE5A0D0F2D0A1A0AAB80F64800AD20";
    attribute INIT_02 of inst : label is "22100100088525CB72390476122022902E8020A445983B6495043000000120C0";
    attribute INIT_03 of inst : label is "911EC26303EA4008204202C9D0A007D0A00F942E002B23902A20262880000400";
    attribute INIT_04 of inst : label is "A0000A1A3148400F0801F3A1882C031E8C88E8395C73011808FB1AA016820883";
    attribute INIT_05 of inst : label is "E50287816628202E4040024944A5004118C41B17CC4209210911407D8484B01D";
    attribute INIT_06 of inst : label is "0201F4544120201604300C84422020102002B000000C813BB3BBF802103F0301";
    attribute INIT_07 of inst : label is "00D31CB9820A6397300034E5FDB64B6E110CA4303BF28282903FC0444000C018";
    attribute INIT_08 of inst : label is "9886C0811001006C57318000420204202C100C7180698E5C9663900539733101";
    attribute INIT_09 of inst : label is "0880044081F81807C0811030480122047C00003C11155044BC0487D983084020";
    attribute INIT_0A of inst : label is "090001889A00148B001489000A400A0C010C4420408000888880080888008000";
    attribute INIT_0B of inst : label is "014818248029120002910820A442002010480480000001880090018800900148";
    attribute INIT_0C of inst : label is "00010400410410000593A442080A444000840208210080020060004040020020";
    attribute INIT_0D of inst : label is "0000024004004000004000104000104000000000000000024904104100000000";
    attribute INIT_0E of inst : label is "0000002002082002080400400000000080000080000000002000082000010410";
    attribute INIT_0F of inst : label is "1000040001040041001040041000000000000000000000201041041041040000";
    attribute INIT_10 of inst : label is "00030000C0000C000030004000000252962E2480872400000000000000000000";
    attribute INIT_11 of inst : label is "DE60010100015E6001010001403004800BE00C0180600C030000600003000018";
    attribute INIT_12 of inst : label is "C070002790104260012149549800052200B05028100A44029123F823CE2A0027";
    attribute INIT_13 of inst : label is "A003D902264184D08109C011020502917F00038001C6300003000030000C0001";
    attribute INIT_14 of inst : label is "084687980C088F279F1E0020220222002605C0522FED995CE3A03D00E318C631";
    attribute INIT_15 of inst : label is "76644220101BC040140340540802009201242204A112D5900A0502817C2439D9";
    attribute INIT_16 of inst : label is "84408844B564029140A18902C5F820403801C0002043000001A084200038004E";
    attribute INIT_17 of inst : label is "4808200012010884402817F00380001021800000D04210001C00277140192224";
    attribute INIT_18 of inst : label is "03C0F03C0F01C0F0F0F07878E000000F80000C00001C00103B90408210B1C71C";
    attribute INIT_19 of inst : label is "800009042D034101A055048AA222202E0C87314D36E0BD5C51000FB226031C0F";
    attribute INIT_1A of inst : label is "92888242827810A81508002007C0018060F03300829001044084A42052017208";
    attribute INIT_1B of inst : label is "0402E0A700C270C4DB2679A18080C0C00E06006CC44249030480373202901F20";
    attribute INIT_1C of inst : label is "400440700A09042842E108421031808C6278077BC082000203705A8048C58069";
    attribute INIT_1D of inst : label is "904D04211E07885936484D1E646841991E28B0B005858188E31C116262630202";
    attribute INIT_1E of inst : label is "81079DCC40380C002191966CE438263650A2879860E6808840C2DBC480CB3110";
    attribute INIT_1F of inst : label is "B42222206054218A51A28C85801020348B1A108811304A2A444262121E101107";
    attribute INIT_20 of inst : label is "0305B028D82559A781415AD3882610120829832A282BB088001562AE63CAE16A";
    attribute INIT_21 of inst : label is "470280824992C0D88025040381F8840420A4198830910823034F107991060048";
    attribute INIT_22 of inst : label is "20408102304081020480015017BB110846109FB01998F07BC4301BB8406B7489";
    attribute INIT_23 of inst : label is "081020408C1020408102040815155FDC060000080C000C000010101010180CA6";
    attribute INIT_24 of inst : label is "01010101800188102040811820408102042A2A90000000C04040404060310204";
    attribute INIT_25 of inst : label is "065204081038080808080C000C40810204608102040955543000004000000301";
    attribute INIT_26 of inst : label is "3060A8A381020703958102040E0602060207020712244891383060C18345450C";
    attribute INIT_27 of inst : label is "40800090048811B9421FC0810381CAC0810207030103010381038912244E0C18";
    attribute INIT_28 of inst : label is "16CA76208C62220161C40768E20019B880A8C20C081025208008221020408010";
    attribute INIT_29 of inst : label is "01008130AA204FBCB0658C0863400022855900118888058400653B0C62000A10";
    attribute INIT_2A of inst : label is "452002A00CC00010C005000001140020204410122000080028B700001F968008";
    attribute INIT_2B of inst : label is "A4070040A0042014004201450146080A01D025603004407F59D04A6010D90436";
    attribute INIT_2C of inst : label is "101088001414141D20259269C811E03B66CF806039008050000000000117B241";
    attribute INIT_2D of inst : label is "054F95FF0232000161E000131010C00014006000008223A4072C478C00E98002";
    attribute INIT_2E of inst : label is "C000092020474E91014021C8706884C125187FD42CFA20A0381081F556205843";
    attribute INIT_2F of inst : label is "2341A804056468308211110B6DA08410A44E78404D818300510437EF3A21E8F0";
    attribute INIT_30 of inst : label is "0000480A82A0A82A0D84310414D01EC222430005C10CC2764409358002020043";
    attribute INIT_31 of inst : label is "0005018400000080200800050B0E0080004440A169000280000200C8001F8000";
    attribute INIT_32 of inst : label is "0010910018000444064000608022A8E200000000040E100000808000FC8001F8";
    attribute INIT_33 of inst : label is "0018400420015540100001000222708000A800555004000A0002AA8720005010";
    attribute INIT_34 of inst : label is "005401007C0028AA1200000290DE200000001554F90003E0000A200800018444";
    attribute INIT_35 of inst : label is "5550000000800000080800000001115A40000000288B52000002AABF20000600";
    attribute INIT_36 of inst : label is "0000100000000000000000000000000000000000000000000000000000000015";
    attribute INIT_37 of inst : label is "468C0002828FADC002840A62B53636518009441FBF5E648120348E5987C00000";
    attribute INIT_38 of inst : label is "452053024900825D51129504A440509A88184243414884526440514117B20C02";
    attribute INIT_39 of inst : label is "00A2C025002368204863CA0210287A25A2801506C080104902A2D34500282811";
    attribute INIT_3A of inst : label is "380000810C0000D04210001C0E801C00C003E8220CC83320CC123D8B42030084";
    attribute INIT_3B of inst : label is "600044249600F91F0C00088288035087FA12004600311800F0B4606002917C00";
    attribute INIT_3C of inst : label is "56AD5555555555555550A0F90480E70D73C1830604512000FB432086452E0081";
    attribute INIT_3D of inst : label is "6AAAAABD55555557AAABD5555555555555555555550AA6AAAAAAAD5555AAAB55";
    attribute INIT_3E of inst : label is "00030000C0000C000030004022022200970000001948A885AAAAAAD555555555";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
