-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "000F00030010FFE80000000000FF000000FF03FF3FFC3FFC0FF00BE003C0C0C3";
    attribute INIT_01 of inst : label is "F000C0000000000304002BFF00000000000000050FFF03FF00FF00FF003F002F";
    attribute INIT_02 of inst : label is "FFFCFFFAFFFF00000000FFFF1000FFFD00000000FFF0FFC0FF00FF00FC00F800";
    attribute INIT_03 of inst : label is "3F808005FF50FFFF0AAA0000BFFF0000FFFF0000003F0040FF808000003F03FF";
    attribute INIT_04 of inst : label is "FFFE0AF0F400FFF40AFF0000F4000FF40000D555A8000AFF0F000A0000000000";
    attribute INIT_05 of inst : label is "0A000FFC003F007F0007000FAFFC00030000FFFF0001FFFF52FF0000003F07FF";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "2B0003F5FF80800003A0FF40F400FFE2FFFFFFFF03FF0FFF2D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00FF000F";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282AC000D5553C0F2800";
    attribute INIT_0B of inst : label is "FC00FD00D000F0003FFAC000FFA0C000034003C001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "3FFFAFFF0000C0003FFCFFFF0FF00FF00000FFC000000000FFC0FFF0FF00FFC0";
    attribute INIT_0D of inst : label is "02E017F4FFFF0AFF0001FFF000030000000000030000000000005000BFFF0FA0";
    attribute INIT_0E of inst : label is "001F1FF0FFFF0000C0000000FC00A00F003FF00A00801FF4C00502FF80FF000F";
    attribute INIT_0F of inst : label is "0000000000005557FF850000FC00FFD0FF0000000AAAFFA002001FF400047FFF";
    attribute INIT_10 of inst : label is "000055FF3FFFFFFFFF02F000557FFFFFF400FF000AFF00030B801FD403FC03FC";
    attribute INIT_11 of inst : label is "55550000FFFF0FFF00000000000000050000000000020000000003FF3FC02801";
    attribute INIT_12 of inst : label is "0000000100A03FF0540003C003C003C0BFFF002B5F80000000000000001F8BFF";
    attribute INIT_13 of inst : label is "0000000002FC5002000000033FC03FC0000000000000000000000000FC000100";
    attribute INIT_14 of inst : label is "02F50000001503C00AC001FF02FF000200000000000040000000000000000000";
    attribute INIT_15 of inst : label is "AAA0000000000000FD55FFFF4000FFFF0000FFFF0000FF55001F00FF00E85FC0";
    attribute INIT_16 of inst : label is "0002000000000000000000003FC03FC0FFFFFFFF5003FF803FC03FC0FFFE0000";
    attribute INIT_17 of inst : label is "FFFFBFFF00000000000000000000000002FF000F4000FD00BFF002FF2FFF03FF";
    attribute INIT_18 of inst : label is "00000000FEA00000FFFF00000000F5404330A2080ABF000000B088A800000000";
    attribute INIT_19 of inst : label is "008C88A8FF80F000CCC380A20FFEFF8000000000800000007373208200000000";
    attribute INIT_1A of inst : label is "FFFFFFFF0000000000000000FFFFFFFEFFF8FFC00001007FFFFEE8000000055F";
    attribute INIT_1B of inst : label is "05FFFFFF0000005FF0000000001888A0000000140FFEFF80007F0FFE0FFF3FFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFD00BFF0BFF002FF0000F5000000140000000000006C888800000000";
    attribute INIT_1D of inst : label is "FFFFFFFF0005FFFF00000000FFFFFFFFFFF0FFFC0000000006900000000F0000";
    attribute INIT_1E of inst : label is "000000570000FFFF157FEA800000D5000000FFFFFD5402AB0000FFFF40000FFF";
    attribute INIT_1F of inst : label is "000000000000C00003FC03FC03FC03FC03FC4028800000000000000000000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
    attribute INIT_22 of inst : label is "100E006E000F0828E410E400C000A08000DD003F0003003FDC00F0000000F000";
    attribute INIT_23 of inst : label is "0000040E001D00000000E040D0000000003F003F0003002FF000F0000000E000";
    attribute INIT_24 of inst : label is "00000000010E000000000000E1000000003F00390007000EF000B0004000C000";
    attribute INIT_25 of inst : label is "00000000002000000000000020000000000F00370007004DC00070004000C400";
    attribute INIT_26 of inst : label is "000000000002000039FC2FD5B4000200001E002F001F0099D000E000D0009800";
    attribute INIT_27 of inst : label is "E7D815F80037028000000000000000000003000200020000B36CFC00D000AB00";
    attribute INIT_28 of inst : label is "FFFFFFFF745FAAAAFD40FFF0FC000000E73B00FE001E03A80000000000000000";
    attribute INIT_29 of inst : label is "BFF07F7D0000000080000000000000000FFF000F00040002FFFFFFFF03D1A002";
    attribute INIT_2A of inst : label is "008001BF00000000A800FF500000000000020000000000000FF811FD00000000";
    attribute INIT_2B of inst : label is "0000000D002D0000000080009000000000020003003600000000200070000000";
    attribute INIT_2C of inst : label is "00000000000000027800306006EC0000000000000000000030000FC000700000";
    attribute INIT_2D of inst : label is "2200103C0006000000803C049000000096D50000000097807ED0000000002A80";
    attribute INIT_2E of inst : label is "0028000E000F0000A000C000C0000000001E000F000F0000D000C000C0000000";
    attribute INIT_2F of inst : label is "00000000000B0000000000008000000000000008000D000000008000C0000000";
    attribute INIT_30 of inst : label is "00000000000300002000E4008000000000030000000200003350F000D0000000";
    attribute INIT_31 of inst : label is "000000000003000000000000D000000000000002000200000000CC0040000000";
    attribute INIT_32 of inst : label is "0099001E202F00009800D000E088000000E4000E80370000EC00C00070800000";
    attribute INIT_33 of inst : label is "0000002202FA000000002000FE000000000000CC082D00000000CC00E9040000";
    attribute INIT_34 of inst : label is "15F00BFF000007000000800000000000000000000A2A0000000000008AA00000";
    attribute INIT_35 of inst : label is "00000000000000002800008000000000000000000000000003D5BFF800000034";
    attribute INIT_36 of inst : label is "000000000000002B000000000000A00000010000000000000000010000000000";
    attribute INIT_37 of inst : label is "001C0000000000A8400000000000A000000000000000008B000000000000A000";
    attribute INIT_38 of inst : label is "00030000000000008F04BFE8000002FA043C0AFF00002BE0B000800000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000036000000000000A70000000000000000000000";
    attribute INIT_3A of inst : label is "00000000000000000F04BFE8000002FA043C0AFF00002BE00000800000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000096000000000000A58000000000000000000000";
    attribute INIT_3C of inst : label is "000B414002DFB847B00D0F80F008FFF27F0A000037A0EFFDF93485042AE00005";
    attribute INIT_3D of inst : label is "01F80350160A0000F4007FC01DF60010AA0880301FF430000000440008208000";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "000F000B00035FFCFFFF00000BFF003F00FF00FFFFFF3FFC0FF00FF003C002C0";
    attribute INIT_01 of inst : label is "F000E000000A0000C0003FF500000000000300000FFF03FF03FF00FF00BF003F";
    attribute INIT_02 of inst : label is "05F0FFFDFFFFAABF00000000C000FF5000000000FFF0FFC0FFC0FF00FE00FC00";
    attribute INIT_03 of inst : label is "0FF8F800D400FFFDFFFF0000FFFF0002FFFFFEAA00FF002FFFF8F800000F00FF";
    attribute INIT_04 of inst : label is "FFF5FFFC4000FF40FFFF000A400A3F40EAAA000005FF54000000050000000000";
    attribute INIT_05 of inst : label is "BF800350001F003F0003000FFFD400200000055500007FFF01FFC00A000000FF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "FFC00000FFD1F8000FFC05004000FF4005FFFFFF03FF0FFF1EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF03FF003F";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF4C000C0003EAD3EA8";
    attribute INIT_0B of inst : label is "F400FC00C000F00017FF0800FFFE2000C30303C02ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "0F507FFFA00000003FFC3FFC07D00FF003FA170000000000FFC0FFF0FF00FF00";
    attribute INIT_0D of inst : label is "2FF80040FFFFFFFF00000003FFF000020000000000030000C00000005FFF3FFF";
    attribute INIT_0E of inst : label is "A00101FCD5402ABF0FFF8000F000FF01000F40FF2BF801D00000A1FFF005003F";
    attribute INIT_0F of inst : label is "00000000AAAB0000FF40A0030000FF00FFE0FC00FF5005552FE80740000305FF";
    attribute INIT_10 of inst : label is "000000000FFFFFFF500FFC000000FFFF0200FC00BFFF00082FF8010003FC03FC";
    attribute INIT_11 of inst : label is "0000AAAAFFFF3FFF000A0000000000000000000000AF0000AFC000D43FC03FC0";
    attribute INIT_12 of inst : label is "0000000002FF05C00000AF4003C003C0FFFF0AFF03C0A80000280000000101FF";
    attribute INIT_13 of inst : label is "000000002FF0002F0000000114023FC0AAFF00000002000000000000FF00F800";
    attribute INIT_14 of inst : label is "03C0002A000001FA3FF0005047FF002F00000000000000008000000000000000";
    attribute INIT_15 of inst : label is "FFFF0000FFAA00000000FFFF0000FFFD00005550000000000080003F03FF0000";
    attribute INIT_16 of inst : label is "0003000000000000000000003FC03FC0FFFFFFFF0000FF4A3FC03FC0FFFF8000";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFF00000000000000AB00000FFD00BF0000F000FF402FFD3FFF0FFF";
    attribute INIT_18 of inst : label is "EA000000FFFF0000055FFEA800000000515053B4FFFF00000010003000000000";
    attribute INIT_19 of inst : label is "001000607FF0FE005441E8D301FF7FF028000000FA000000511130C300000000";
    attribute INIT_1A of inst : label is "7FFFFFFF0000000000000000FFFFFFFFFFFCFFF00000000FFFFFFFA000000000";
    attribute INIT_1B of inst : label is "00177FFF00000001FE0080000050000C0000000001FF7FF0000F01FF03FF1FFF";
    attribute INIT_1C of inst : label is "FFFFFFFFF000FF40FF400FFD0000400000000000FA800000000400AC00000000";
    attribute INIT_1D of inst : label is "FFFFFFFF000005FF02AF0000FFFDFFFFFFC0FFF4000000000000096000BF0002";
    attribute INIT_1E of inst : label is "000000000000057F0000FFFF000000000000FD500000FFFF000000000000C000";
    attribute INIT_1F of inst : label is "0000000000004000801403FC03FC03FC03FC03FCC00000000000000000000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
    attribute INIT_22 of inst : label is "020E000E003F000CC200C000F000E40000FB000F000300FFBC00C0000000FC00";
    attribute INIT_23 of inst : label is "011C008E000F0000F100C800C00000000026001F0003003F6000D0000000F000";
    attribute INIT_24 of inst : label is "0000005C002E00000000F400E0000000003F003F0003002FF000F0000000E000";
    attribute INIT_25 of inst : label is "00000000000C000000000000D0000000003F003E0003001DF000F0000000D000";
    attribute INIT_26 of inst : label is "0000000000030000077BFF00400029B2000E0037000300E4C00070000000EC00";
    attribute INIT_27 of inst : label is "F9E000FF00071FE000000000000000000000000300030001FF50FC004000BCD8";
    attribute INIT_28 of inst : label is "FFFFFDFF0005FFFFFFBCFDD0F400EF0017FC00FF00079CF90000000000000000";
    attribute INIT_29 of inst : label is "FF8B054000000280400000000000000005FF003F00000001FFFFFFFF0140FFAF";
    attribute INIT_2A of inst : label is "017F000400000000FF2885400000000000000020000000007FFF004000000B80";
    attribute INIT_2B of inst : label is "000100B0000100020000D4000000000000020049003300030000E40020000000";
    attribute INIT_2C of inst : label is "0000000000000001678018380074800000000000000000003E0007F000148000";
    attribute INIT_2D of inst : label is "D0600037000300000A47DC00400000001500000000009577000000000000FEFA";
    attribute INIT_2E of inst : label is "000C000700030000C000C00000000000000E000700030020C00040000000A000";
    attribute INIT_2F of inst : label is "000000080002000000008000000000000000000E000300000000C00000000000";
    attribute INIT_30 of inst : label is "0001000200030000DB00C000400000000000000200030000F900F0004000A880";
    attribute INIT_31 of inst : label is "0000000000020000000078004000000000000000000300000000B00040000000";
    attribute INIT_32 of inst : label is "00E4000EAADF0000EC00C2007E2A0000001E002F2EFF0099D000E000FE819800";
    attribute INIT_33 of inst : label is "000000CC9EFD00000000CC00FBDE00000022007823FF00002000F400F7A20000";
    attribute INIT_34 of inst : label is "0EBC556000000B00000000000000000000000000FBFB000000000000FFFF0000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000FAC095500000038";
    attribute INIT_36 of inst : label is "000000000000005D0800000000004000000000000000000B0000000000008000";
    attribute INIT_37 of inst : label is "00000000000007FF000000000000F40000000000000001DF040000000000DC00";
    attribute INIT_38 of inst : label is "0001000000000000E6BD0A5700000BF51FA6F568000017F8D000000000000000";
    attribute INIT_39 of inst : label is "00000000000000000000000200C000000000A00000C000000000000000000000";
    attribute INIT_3A of inst : label is "001F000000000000E6BD0A5700000BF51FA6F568000017F8FD00000000000000";
    attribute INIT_3B of inst : label is "00000000000000000000000200C000000000A00000C000000000000000000000";
    attribute INIT_3C of inst : label is "2D0500F4007C0000FE0081000002554B5000080001DCFF70FEF80C0005402800";
    attribute INIT_3D of inst : label is "0450800B015600004000FFF8FBF8000C590CFEF91F5251000A000000016A0008";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "003F000F057EFFFFAAAA555503FF007A03FF0FFFFFFFFFFF3FFC2FF80FF0F3CF";
    attribute INIT_01 of inst : label is "FC00F0000000000FBD50FFFF000000000003C15F3FFF0FFF03FF03FF00FF00BF";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFF002A0000FFFFF500FFFF00000000FFFCFFF0FFC0FFC0FF00FE00";
    attribute INIT_03 of inst : label is "FFE0E05FFFF4FFFFAFFF0000FFFF0000FFFFA80000FFD5FAFFE0E00000FF0FFF";
    attribute INIT_04 of inst : label is "FFFFAFFCFD00FFFDAFFF0000FD003FFD8000FFFFFEAAAFFF0F000A0000000000";
    attribute INIT_05 of inst : label is "AF803FFF00FF01FF001F003FFFFF000F0000FFFF1557FFFFFFFFC00000FF1FFF";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "BFC00FFFFFE2E0000FFAFFD0FD00FFFBFFFFFFFF0FFF3FFF2D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A03FF003F";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282AC000D5553C0F2800";
    attribute INIT_0B of inst : label is "FF00FF40F400FC00FFFFF000FFF8F000C7D30FF001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "FFFFFFFF0000F000FFFFFFFF3FFC3FFC03A0FFF500005550FFF0FFFCFFC0FFF0";
    attribute INIT_0D of inst : label is "0BF87FFDFFFFAFFF0007FFFEAAAF55560000000F00030000C000F543FFFF3FFA";
    attribute INIT_0E of inst : label is "007F7FFCFFFF002AFAAA9555FF00FA3F00FFFCAF02E07FFDF05F0BFFEBFF003F";
    attribute INIT_0F of inst : label is "000005550002FFFFFFFF0003FF00FFF4FFC0AD00AAAAFFFA0BA07FFD005FFFFF";
    attribute INIT_10 of inst : label is "0000FFFFFFFFFFFFFFEBFC00FFFFFFFFFD02FFC02FFF000F2FE07FFD0FFF0FFF";
    attribute INIT_11 of inst : label is "55550000FFFF3FFF000000000000005FC0002400000B0A400AC05FFFFFF0BEAF";
    attribute INIT_12 of inst : label is "0000000702FAFFFC540003C003C003C0FFFF00BF5F80000000090000007FEFFF";
    attribute INIT_13 of inst : label is "000000000BFFF50B0C03300FFFF0FFF000AA00000002000000000016FF00AF57";
    attribute INIT_14 of inst : label is "02F50000001503C0AFF007FF8BFF000B000094000000D0008000000000000000";
    attribute INIT_15 of inst : label is "FFFA0000AA000000FFFFFFFFD554FFFF0000FFFF0000FFFF807F03FF03FEFFF0";
    attribute INIT_16 of inst : label is "240B090202400030000C0000FFF0FFF0FFFFFFFFF50FFFE0FFF0FFF0FFFF0000";
    attribute INIT_17 of inst : label is "FFFFFFFFAAAA5555A400000A000200000BFF003FD000FF40FFFC0BFFBFFF0FFF";
    attribute INIT_18 of inst : label is "80000000FFFA0000FFFFA8000000FFD54330A208AFFF000000B088A800000000";
    attribute INIT_19 of inst : label is "008C88A8FFE0FC00CCC380A23FFFFFE060000000E00001A073732082001AA000";
    attribute INIT_1A of inst : label is "FFFFFFFF0003001800C00300FFFFFFFFFFFEFFF0000701FFFFFFFE0000005FFF";
    attribute INIT_1B of inst : label is "1FFFFFFF600001FFFC008000001888A00000007D3FFFFFE001FF3FFF3FFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFF40FFFCFFFC0BFF0009FF4000007D00A0000000006C888801600001";
    attribute INIT_1D of inst : label is "FFFFFFFF005FFFFF000A0000FFFFFFFFFFFCFFFF0940400080029416003F0002";
    attribute INIT_1E of inst : label is "000005FF0015FFFF7FFFFFEA0000FF505400FFFFFFFDABFF0000FFFFD000BFFF";
    attribute INIT_1F of inst : label is "030000C0C030F00C0FFF0FFF0FFF0FFF0FFFFABEE018806001800C0030000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "0FFD00150000028BDBC0D000C0008A0000E20020000000302C00200000003000";
    attribute INIT_23 of inst : label is "000203FD000200000000DF00C00000000000000000000020200000000000E000";
    attribute INIT_24 of inst : label is "0000000200FD000000000000DC0000000030000600050001300040004000C000";
    attribute INIT_25 of inst : label is "00000000000200000000000000000000000C00180000007EC000B0000000F400";
    attribute INIT_26 of inst : label is "000000000002000036B726C044000200000D00240018003AC00060009000B000";
    attribute INIT_27 of inst : label is "5FE4107800280000000000000000000000000002000300004D98480000000B00";
    attribute INIT_28 of inst : label is "DF0FED3489A0555502BEBC0903508A8099C40086000303800000000000000000";
    attribute INIT_29 of inst : label is "400E8082052000000000C00000000000F00000F207FB002D3C03D2F17C2E5E89";
    attribute INIT_2A of inst : label is "0B7E3E4000FD008053C000AD014000000009000100100000F0076E0200000200";
    attribute INIT_2B of inst : label is "0008000200120002000040004000000000010060004200000000C0000C000000";
    attribute INIT_2C of inst : label is "000000000000000000000F800110000000000000000000044800303801B40000";
    attribute INIT_2D of inst : label is "08001024000300000028180440000000B95500000000A9006B90000000002A80";
    attribute INIT_2E of inst : label is "000A000D000800008000C00080000000000D000400080000C000400080000000";
    attribute INIT_2F of inst : label is "000000000008000000000000800000000000000E000E00000000C000C0000000";
    attribute INIT_30 of inst : label is "00000000000200008800F400400000000000000000030000CD80400000000000";
    attribute INIT_31 of inst : label is "0000000000020000000000000000000000000000000200000000F40080000000";
    attribute INIT_32 of inst : label is "003A000D00240000B000C00060800000009B000D80380000D800C000B0800000";
    attribute INIT_33 of inst : label is "0000002002C50000000020006600000000000037080E00000000F000C1040000";
    attribute INIT_34 of inst : label is "D5F0FFFF0000C7000000800001780000000000000A82000000000000A2A00000";
    attribute INIT_35 of inst : label is "00000000000000009600026000080000000000002D40000003D5BFFF00000034";
    attribute INIT_36 of inst : label is "0000000000000094000004000000580000040000000000004000064000100000";
    attribute INIT_37 of inst : label is "8161000000000A1690000000000018000041000000000B344800020000005A00";
    attribute INIT_38 of inst : label is "000300000B5000008F00BFFF000002FFC03CFFFF0000FFE0B000800001780000";
    attribute INIT_39 of inst : label is "0000000000000000000000000036000000000000A70000000000000000000000";
    attribute INIT_3A of inst : label is "000000000B5000000F00BFFF000002FFC03CFFFF0000FFE00000800001780000";
    attribute INIT_3B of inst : label is "0000000000000000000000000096000000000000A58000000000000000000000";
    attribute INIT_3C of inst : label is "0AF4BCB70D00B87841F0F0370948000C8035E94137A0100002C07AD01514F005";
    attribute INIT_3D of inst : label is "7C07000B16F500600182803FE209201000B37FCF600030098010AB6408205428";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "003F002F000FFFFFFFFF00002FFF00FF03FF03FFFFFFFFFF3FFC3FFC0FF0CBE3";
    attribute INIT_01 of inst : label is "FC00F800C2AF0003F000FFFF80000000000F00003FFF0FFF0FFF03FF02FF00FF";
    attribute INIT_02 of inst : label is "5FFCFFFFFFFFFFFFAAAA5555F000FFF400020000FFFCFFF0FFF0FFC0FF80FF00";
    attribute INIT_03 of inst : label is "3FFEFE00FD00FFFFFFFF0000FFFF2AABFFFFFFFF03FF40BFFFFEFE00003F03FF";
    attribute INIT_04 of inst : label is "FFFFFFFFD000FFD0FFFF00AFD0AFFFD0FFFF40005FFF55550000050000000000";
    attribute INIT_05 of inst : label is "BFE00FF5007F00FF000F003FFFFF0ABD00005FFF0000FFFF07FFF0AF00B503FF";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "FFFA0350FFF7FE003FFF5F40D000FFD15FFFFFFF0FFF3FFF1EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF0FFF00FF";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF4C000C0003EAD3EA8";
    attribute INIT_0B of inst : label is "FD00FF00F000FC00FFFF7EA0FFFFFA00F3CF0FF02ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "3FF5FFFFFA83C000FFFFFFFF1FF43FFC0FFF7FC0AAA00000FFF0FFFCFFC0FFC0";
    attribute INIT_0D of inst : label is "BFFE01D0FFFFFFFFAAA9555FFFFD000B00000003000F0000F0000000FFFFFFFF";
    attribute INIT_0E of inst : label is "FA0707FFFFD5BFFF7FFFE000FC00FFD7003FD7FFBFFE07F4C000FFFFFC5F00FF";
    attribute INIT_0F of inst : label is "0AAA0000FFFF0001FFD0FA0F5E00FFC0FFF8FF00FFF55FFFBFFE1FD0000F1FFF";
    attribute INIT_10 of inst : label is "000000553FFFFFFFF53FFF000015FFFF5FABFF00FFFF00AFBFFE07400FFF0FFF";
    attribute INIT_11 of inst : label is "0000AAAAFFFFFFFF00AF0000000000000000300002FF9000FFF003FDFFF0FFF0";
    attribute INIT_12 of inst : label is "000000010BFF5FF00000AF4003C003C0FFFF2FFF03C0A80000BE0000000747FF";
    attribute INIT_13 of inst : label is "00290000BFFC00BF060118077D5FFFF0FFFF0000000B000000000000FFC0FE01";
    attribute INIT_14 of inst : label is "03C0002A000001FAFFFC01F5DFFF00BF0000000000004000E000000068000000";
    attribute INIT_15 of inst : label is "FFFF0000FFFF00005400FFFF0000FFFF0000FFF500005500EAF500FFAFFF05C0";
    attribute INIT_16 of inst : label is "300F0C03030000C000240003FFF0FFF0FFFFFFFF0003FFFFFFF0FFF0FFFFEAA8";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFF0000000202900AFF00003FFF02FF4000FC00FFD0BFFFFFFF3FFF";
    attribute INIT_18 of inst : label is "FFA00000FFFFA8005FFFFFFE00005000515053B4FFFF002A0010003000000000";
    attribute INIT_19 of inst : label is "00100060FFFCFF805441E8D307FFFFFCBE000000FF800006511130C380000680";
    attribute INIT_1A of inst : label is "FFFFFFFF0000000C00300180FFFFFFFFFFFFFFFC0001003FFFFFFFF800000005";
    attribute INIT_1B of inst : label is "007FFFFF05800007FF80E0000050000C0000000607FFFFFC003F07FF0FFF7FFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFC00FFD0FFD03FFF0250D00000009000FFEA0000000400AC00055800";
    attribute INIT_1D of inst : label is "FFFFFFFF00005FFFABFF0000FFFFFFFFFFF0FFFD500000256829400102FF000B";
    attribute INIT_1E of inst : label is "0000000100005FFF0015FFFF000040000000FFF55400FFFFAAAA55556AAAF555";
    attribute INIT_1F of inst : label is "0C0002404090D024F57D0FFF0FFF0FFF0FFF0FFFF00CC03000C003001800C000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "01FD000100303FFFFD00C000B000DBF00084000E000000C04800C00000002C00";
    attribute INIT_23 of inst : label is "0AEF007D00000000CE80F400C00000000019001A000000309000900000003000";
    attribute INIT_24 of inst : label is "000002AF001500000000CA00D000000000000030000000282000B0000000E000";
    attribute INIT_25 of inst : label is "0000000000FF000000000000EC000000003000110000000A700030000000C000";
    attribute INIT_26 of inst : label is "000000000000000006ED430040002750000D00380000009BC000B0000000D800";
    attribute INIT_27 of inst : label is "87F000C300043E180000000000000000000000030001000280100C0040004FF0";
    attribute INIT_28 of inst : label is "0B2D0255141AA80AF843522C090010F0100800C300053FC60000000000000000";
    attribute INIT_29 of inst : label is "00743A9D00002D68B0000000000001807A000BC10000BFFEF5E355001EB02850";
    attribute INIT_2A of inst : label is "0E8001FB0000000200D77AB001000100001F008880000000800015BD0000246A";
    attribute INIT_2B of inst : label is "0002000F000100000000000000000000000100B2004300008000180010000000";
    attribute INIT_2C of inst : label is "0000000000000000180007C0000000000000000000000000C1A0180C00146000";
    attribute INIT_2D of inst : label is "01A0003F000100000340FC00400000000100000000003FDD0000000000004110";
    attribute INIT_2E of inst : label is "001F000C00000000D000C00000000000000D00080000001BC000800000009000";
    attribute INIT_2F of inst : label is "0000000A0001000000008000000000000000000F000100000000C00000000000";
    attribute INIT_30 of inst : label is "0001000200010000A60000004000000000000002000100008400000040000A80";
    attribute INIT_31 of inst : label is "0000000000010000000080004000000000000000000100000000600040000000";
    attribute INIT_32 of inst : label is "009B000D80300000D800C20090820000000D00240C10003AC00060001201B000";
    attribute INIT_33 of inst : label is "00000037312600000000F0004C2400000020004F880000002000C40049080000";
    attribute INIT_34 of inst : label is "EABC557F0000FF000000FA000003000000000000540400000000000000050000";
    attribute INIT_35 of inst : label is "00000000000000001400004000000000000000ABC00000000FAAFD550000003F";
    attribute INIT_36 of inst : label is "00000000000001A2260000800000900000000000000000240200000000006000";
    attribute INIT_37 of inst : label is "0008000000001800000000000000090000000000000022201900000000002200";
    attribute INIT_38 of inst : label is "0001002B30000000E6BFFF5700000BF5FFA6F57F0000D7F8D000FA0000030000";
    attribute INIT_39 of inst : label is "00000000000000000000000200EA00000000A000EAC000000000000000000000";
    attribute INIT_3A of inst : label is "001F002B30000000E6BFFF5700000BF5FFA6F57F0000D7F8FD00FA0000030000";
    attribute INIT_3B of inst : label is "00000000000000000000000200EA00000000A000EAC000000000000000000000";
    attribute INIT_3C of inst : label is "92FA120007820007000216C0B002AAB4A506080001DC000B010702800000C7F0";
    attribute INIT_3D of inst : label is "03AD803401699EA8AFA9000704000C08A6F3000600A9502E5008D690016AF0A4";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
