-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D344D8649830C93FF5146EAA98D309A49B2A3FC00000139308C1D34C35B9352A";
    attribute INIT_01 of inst : label is "A11BAD08ED3C7686C0485372219AC0723067D599C661DDFC749A829999B502C4";
    attribute INIT_02 of inst : label is "DCDC90242A79A31EF61FD5863DFFBA674446856CAC51D8F78A17FBBEE99D1111";
    attribute INIT_03 of inst : label is "582A05618D6154197555346EB022026856D7FFFE976296EDF29B3A10E6071149";
    attribute INIT_04 of inst : label is "F9BD1337EF63A07A58B43C3CB5381D34DBB4A7698998498A6398261998560A81";
    attribute INIT_05 of inst : label is "78DA279A6B0AC0624711E60BEBE02191CA40362468822A2D742877800D5F3BD6";
    attribute INIT_06 of inst : label is "A259AA39999DF1AEBACD0697D66F3473DA39CC2A2B6779C8C3D40C62D0F03016";
    attribute INIT_07 of inst : label is "C003CFA5CB25F34DA04924D2E21E1DC8AF67A8CA68695955746BF3AA9D5B5CE9";
    attribute INIT_08 of inst : label is "4ABA10658940DDAACEF39187A7144814DA7795E6457374F8398F55F73BB0ADD9";
    attribute INIT_09 of inst : label is "10B2B2E8FAA4E235A29C46B411CB128739D7AF637951CA9BECE8F5900506BEC7";
    attribute INIT_0A of inst : label is "7A03E8CFAB0F4758BEF8DEFE3DEFF0D9BF9428F4DEFF7BFE4FE56C696684053D";
    attribute INIT_0B of inst : label is "5D5FFFD7D5F7D5F7FFF7D5F7D5F5D57557D0D3CCFF71CAE2558E38F137E2CD21";
    attribute INIT_0C of inst : label is "DDD7B6DFE4546F9E731ED66D4042C258F5D4F13CF054C13710921CBACE37A4DA";
    attribute INIT_0D of inst : label is "5556228328A9BAFB2EAE2A2C8289ABACFAEFFFE1FF999801E00051111400075D";
    attribute INIT_0E of inst : label is "AE14DD0119542DCF4EAB7B72D68E15915F339C3A4DA55555DDDAAAAAAAAD5555";
    attribute INIT_0F of inst : label is "187C0BABAFABAB51500DAA94F8280FFCFF69D8F4410052801C52CB9FF1C30A6E";
    attribute INIT_10 of inst : label is "A228A04A20A088CCCAF6F6CCE70F9F614B3EDCE4D249B8678F0DA6B2EFD66563";
    attribute INIT_11 of inst : label is "01007FC0820A4180000000000000000000000000000008F8ED380000007E048A";
    attribute INIT_12 of inst : label is "7095659E744B3A2746EB35C5CFB0CBC9A87E2C3BBC9EF6CAB72E63BD96C00400";
    attribute INIT_13 of inst : label is "4EF39187B697439A3E257580083BBB16EACE3987E0C5DAAA409EB6E905E81A54";
    attribute INIT_14 of inst : label is "966660000555500005555CDD3319FD4E1B82D9C8FFBFCA0E7390F963690CDAB2";
    attribute INIT_15 of inst : label is "658A09162A245D1240800F3A63DECC9BF80FDAA6559AA7775555500000000999";
    attribute INIT_16 of inst : label is "5AAAF80282AAA90002FBEFF9C633F992477E1ED378CA2B275638DEB2A2A3ACE0";
    attribute INIT_17 of inst : label is "54759C0CB14122C5448BA262A208431EE7226FE01F6D18656CDAFFFC2EABD410";
    attribute INIT_18 of inst : label is "D7DA19ACF659A1EA37882A43BDF8B743E9FF81D229AF2AAAAA86562EA67EBA54";
    attribute INIT_19 of inst : label is "EE75C1C0E3F53C4E04A6F1166C0D986D7F6A9BA294D2E93877EDD38E74D5BAF3";
    attribute INIT_1A of inst : label is "C6090D75EB60039309C246A67BFCC13BFC545F22A2D55F6AAFB5F34475576999";
    attribute INIT_1B of inst : label is "E0004800C53799BDA0DEFADF2BD9D642724D09B61AE733ACB7BF8F7BFE1FEB3E";
    attribute INIT_1C of inst : label is "C396277B4DC01053667E8FAC99BAC5C579629B986D9D9899DBE531BF1402261C";
    attribute INIT_1D of inst : label is "CA5219CB0E736B8E8F63D0FE6E1CFF8FF5DCDF3C1B35950BFB7AF0570EFDB266";
    attribute INIT_1E of inst : label is "B9F487118080098675B683EB785784FC4364620108E8D7FDBCC4500BC5567D99";
    attribute INIT_1F of inst : label is "E79CF6FFFFFFA676EC7134BFA761F2061C77EA94DFBBAC53C60E3171EF95B3F6";
    attribute INIT_20 of inst : label is "F18B8C1BAFF4D24D2397E3E71BA5E992E073CEFFFFFF2691EB92FEB976C3A7F9";
    attribute INIT_21 of inst : label is "4ED4BFCD27F66BA470230FDC4EBBBD8FF7B1D8D14F4561B77915151515B8E608";
    attribute INIT_22 of inst : label is "AE86BFC36B9402539CC62234A5A16639884272125397069D1BDE769AAFFEEBC7";
    attribute INIT_23 of inst : label is "2A2A33333335866EED8F4A6D2B616B1B5227349ED6D76975AD749ED6BA5D6B81";
    attribute INIT_24 of inst : label is "EB2AA0428853DAFA78CEF24C7501B5A5086D69420AED0A096193358F33332A2A";
    attribute INIT_25 of inst : label is "35E7E672C7494A3D37FF310947E8D6FBB6DDC8BE2324D5AE45FE6434428425DA";
    attribute INIT_26 of inst : label is "5218581E9A501C19A8009BC52EFF9DF847FDCCC622801BAD2754DF4FF290C3D2";
    attribute INIT_27 of inst : label is "2D7AC01673B3331215D7779030030FD7FFEFADB52B7BB89A3E689A1A684A9CC0";
    attribute INIT_28 of inst : label is "718B8C1E8149640243F183D235E66629FFDC758802FF398C6C7A98B1B92520F1";
    attribute INIT_29 of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA07375A2A7FBD8181BA7F94F7F44A3FBB9A";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2B of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2D of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0088C2619A34600003E7482E0F7A41B00046400000000D528201BA0229B04A26";
    attribute INIT_01 of inst : label is "8846744224F19A3000C4921C7D560C9C69D80C55576533899B4CDBD55078B0CA";
    attribute INIT_02 of inst : label is "3A90B72D50249AF24DC6AD3C4467FD11998A73E7E9C2179235B19FFFF4466262";
    attribute INIT_03 of inst : label is "AA84128C0A759C18F00BD1D9A6591DA71E755502715E752A0E00898A8A757210";
    attribute INIT_04 of inst : label is "03F04A842922A3355754CCCD55541BA028AA995A80A80A8AA0A86A0A9128A144";
    attribute INIT_05 of inst : label is "7C1BC7C08025CF29373ED4004361607E37A68059A1E6CE83418C97653E1155B5";
    attribute INIT_06 of inst : label is "8ED19AE050D2AF99A885B804001693CC68E6135CDC03EDE45F46DA6676B9B2AC";
    attribute INIT_07 of inst : label is "0000A28112004484B7E713C89F7755BF02CDA490A2AF912F515AF5642B3778F8";
    attribute INIT_08 of inst : label is "0DF82AAFF2EE119607DBC8BE818DCD241B0841161E41760F97792C2CC08B7006";
    attribute INIT_09 of inst : label is "4449A0AB8096059134D0B2225A3DE5D8004020B8401D6F4220E0E5E9B28616C7";
    attribute INIT_0A of inst : label is "D665A3988E511C74C10194AED94AB447285AF11194AE52B007E3414092219C74";
    attribute INIT_0B of inst : label is "2AAAAA82AAA02A0000002A02AAA22A8000DEFA2AB25520C47A2AACFA842B1B6C";
    attribute INIT_0C of inst : label is "DF004920001E105C73BE314AEDD5CEB9B73CE681F3E824B9325450022B84CA19";
    attribute INIT_0D of inst : label is "55565C29AA29EDAE2BAE28AE2971AEA9AF3F555F54F1C3541555FC105F800017";
    attribute INIT_0E of inst : label is "7D79CCBD63F3648013FDC077F0746C5DA080018CA19555557D7AAAABBAAD5775";
    attribute INIT_0F of inst : label is "794F0BBFBBAEBBEFBFBE0451515BE2C0011B420A000070CC004304828626BCE6";
    attribute INIT_10 of inst : label is "310D320308319999C31207F948D21FFE82614212D822BAFA2869558DB2AA82AA";
    attribute INIT_11 of inst : label is "010000400200000060000000000000000000000000000FE005A8000000528123";
    attribute INIT_12 of inst : label is "3400DB6999A6CCDA88000BA124244CAE65BD66420050009E6F1E417B31800400";
    attribute INIT_13 of inst : label is "07DBC8BE80056F4155908334919BFFB87E685997E4CDDB1C5B1D102AA92ACAE0";
    attribute INIT_14 of inst : label is "55A5AFFFF5555FFFF55552966737FE824C94000165B0002B483B02A98A521900";
    attribute INIT_15 of inst : label is "CB97D02E5D40B826864E51EEA6C425C400E0FAA9556AAD7D5555500000000A5A";
    attribute INIT_16 of inst : label is "2AABA082802AAD555024027B8266C3D7CC1EBBF6EA9DC44C82AE117044447CF5";
    attribute INIT_17 of inst : label is "888F9EB9123A0448A81104464E51CD3624871005C3F4AF2A0A1955577FFEC405";
    attribute INIT_18 of inst : label is "EA1B515B286236A024FE7AD80F7C6AD35C7720E54D82489D67DCAD7502818408";
    attribute INIT_19 of inst : label is "000C3BBAA6DF39A0CBCF62DAF452430CB16DA00C6D349A80280B4DDFFD452F07";
    attribute INIT_1A of inst : label is "0D6D6C9255118A2844582F6958FC3A044338E219C7189B8C4DC200232B22A644";
    attribute INIT_1B of inst : label is "5FFF224308AE7570B6BDAB5F5D3644D4B695B2DA6E5A8061E52BB652AD882662";
    attribute INIT_1C of inst : label is "3A4015CBA1001200155DF56BC4260AB8B34F251B09304C44044A1C45293C4069";
    attribute INIT_1D of inst : label is "0694C200AB4864DCDD0741C0B2DFFFC4AE416008D4A2E26CB2512120A9362459";
    attribute INIT_1E of inst : label is "44083100919100780C2CDE5EF4FD6EFDAED09B6857E7C832CB5CA99C098A0240";
    attribute INIT_1F of inst : label is "C8557A0000209540234D20088A6DE6CF3B88B1670608AB9DCF577BA506D60814";
    attribute INIT_20 of inst : label is "BBDDDEA08807ACDE4A400015C229005C802A4A0000200F25025C8FFBAFF40204";
    attribute INIT_21 of inst : label is "F22D6FC35BF16F1379C696624E167231986F3346304CCC4CC42A2A6E6E073872";
    attribute INIT_22 of inst : label is "E0DF87DA6FA65A4318E634B6F5B7E7318E631EF12B5B4B2C2C02A13A6BFEBADE";
    attribute INIT_23 of inst : label is "6E6E66676660207FF820D01F42AAFD57EF6A2109F0D9021BE24109F12084F817";
    attribute INIT_24 of inst : label is "3A2CF6E4D3A5B034955284DF27B85D57BB5755EF55ED8618083AA82166676E6E";
    attribute INIT_25 of inst : label is "A90215458E4C1B780A368DBC8891276F38E5C2FEB30ADB6E11BE35B7D1DEED19";
    attribute INIT_26 of inst : label is "4A2088E6268146A1D0E6A2A8098031FD9EC96A946F4CA0889A8E90969CEAAA08";
    attribute INIT_27 of inst : label is "4E4010002A2AA8DB4B7E5A0D3DD3DD8520B64E394588201EA3491EA740FEA5D9";
    attribute INIT_28 of inst : label is "BBDDDEA7098BA844549D1A00B91555C011BFA92A170245294D40495C213065E6";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE02A11106242491B1C4B4674B6201616F53";
    attribute INIT_2A of inst : label is "6666666666666666666666666666666666666666666666666666666666666667";
    attribute INIT_2B of inst : label is "6666666666666666666666666666666666666666666666666666666666666666";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "6666666666666666666666666666666666666666666666666666666666666667";
    attribute INIT_2F of inst : label is "6666666666666666666666666666666666666666666666666666666666666666";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "80864321CF9C5C3051B12BEBCF68D52401423FC000003A8A301C35D0A1064402";
    attribute INIT_01 of inst : label is "2F62B9FFA147DCEC40F921462CCC04462878884CC5415AABFDB292CCCC440482";
    attribute INIT_02 of inst : label is "E254671952802DD627A8390004688B81DEECAE8F4800AEB12D7128822E0777BB";
    attribute INIT_03 of inst : label is "8F41C0102848D91542AA25972493A2CAD4F2AAA8B274A74FF66112824D520542";
    attribute INIT_04 of inst : label is "43DCF9555BF762219801777600E9C35D09382A7689681681A2681A068A035420";
    attribute INIT_05 of inst : label is "355273420245C21A6509729C1481541B0EC754412228ACA2544D0147134166E7";
    attribute INIT_06 of inst : label is "2C910AA8C8D6190B27C0AC8494130578C2BC477F6633A94A5D44934026A920A7";
    attribute INIT_07 of inst : label is "20017BB4A9B5D7D9959EF77AB95B54190B442886CAEBD94A4772B5A9BD5A4E58";
    attribute INIT_08 of inst : label is "E62730A31CA95504275294BA95858921520814111314540105E39DA68A2D98A9";
    attribute INIT_09 of inst : label is "5401202AB08614A534C294A21A24215148447EF55474EFAABA3A202CA2C00224";
    attribute INIT_0A of inst : label is "FC74CAF54B705864C4F9DEFECDEFF416A5520005DEFB7BEA2562418A00A55159";
    attribute INIT_0B of inst : label is "7FFFFFD7FFF5555555555557FFF7555554AB7AA65B74A3746B269E7A55EDD248";
    attribute INIT_0C of inst : label is "202B249248221C410D35A1262A14348DED281449F9AF472F33974825E7556C50";
    attribute INIT_0D of inst : label is "5555ABFC00020205FFFA80017EAEFFFF0080AAB55551D5554AAAAFEFEA8002A0";
    attribute INIT_0E of inst : label is "36E9C82540B3C4045D56C224512A4848B0145F56C505555557FAAAABEAA955F5";
    attribute INIT_0F of inst : label is "10570144055540100400145061A2AFFCFA6E17FE0104A2880453CB3C71F034E4";
    attribute INIT_10 of inst : label is "0B4106C03908880042020035AFC4400E15554C6892100E88A4257306DBAE72E9";
    attribute INIT_11 of inst : label is "01000000000000000000000000000000000000000000081204200000003EDDF0";
    attribute INIT_12 of inst : label is "060B0DEA9DCB666CCC48082160B42C01347F6208050212D6142840A1E2000400";
    attribute INIT_13 of inst : label is "275294BA94A82900630750201610116A94A811034281120C524F4E83A00280E0";
    attribute INIT_14 of inst : label is "555AA000055550000555524E55B8FAF677970A41B725236755CAFAFEEBD45000";
    attribute INIT_15 of inst : label is "8F1ED83C7B60F03CA4CCDF58B78205C4DCFFC55555555FD55555500000000AA5";
    attribute INIT_16 of inst : label is "4AAAEA2802AAAD5556041269837783D76E34ABECB2D97678C49554E06666D417";
    attribute INIT_17 of inst : label is "CCDA82F1831B060C6C180686EEDA95BC08071369FE9FB20B40505554FAAA8155";
    attribute INIT_18 of inst : label is "2FD24AADB2BF15C868E538B8D56F6C00A1DD2424F97D221FD278D0D08341020C";
    attribute INIT_19 of inst : label is "82082A2AB78A05128A6DE28EDE5B8EA82F49200C392412002A5D05D739107507";
    attribute INIT_1A of inst : label is "0A41481F50252B38D2D2202D2E00B8107AADB3D56D8CCCC666665159ED9EE02A";
    attribute INIT_1B of inst : label is "3941020150D94ECC15C63241501B169EE4A0AE6CBCA9114177BFB37BFD85E3D5";
    attribute INIT_1C of inst : label is "C90573F3D5481248732759CE72AC0E6EDA69B4CE85F0B52B0B7B4AB62F3667A5";
    attribute INIT_1D of inst : label is "55B78AA36555401A1BD6F5B5DA97D57B7BDFBE1D1E9FBB48DB77B1B725DB36ED";
    attribute INIT_1E of inst : label is "69EC6266E6A24500083856739CC1C2050EC2915AD68E861B6D9CB9160CCE7A88";
    attribute INIT_1F of inst : label is "374FAEAB62BFD3314A4934236449368C2EECE1B59F520DDE8A5A52EC9E546947";
    attribute INIT_20 of inst : label is "529694B52D723693E90547F3AAAD5AD6A0490EAB62BF49F49AD6A14AC956201B";
    attribute INIT_21 of inst : label is "84E93AD24EB049A64862834C08B3557CC33D53DF024078A7A8F7337FBB15AE7A";
    attribute INIT_22 of inst : label is "401904C04BA0072842309165BF219084211902BE488A152855BA67730EA8F3D6";
    attribute INIT_23 of inst : label is "22A233323333ABB333EA8292084892449448652520918A0A400525200292902E";
    attribute INIT_24 of inst : label is "922810E038B6E6C6D44E6C91408889008B02402340A90E18EACF73A2333222A2";
    attribute INIT_25 of inst : label is "AD489335D7D89A6D18DB38A6CCE1B7FDBEF0D6FEA91A964ABF2A2524910A8910";
    attribute INIT_26 of inst : label is "9807C13807C93800C89C0789090439AD136DE652458CB52C6CC65DE90EF26939";
    attribute INIT_27 of inst : label is "6F569400498992884FFBA49DA5DA5ED58CE7EFBDEEDFA95801E97881E09883E0";
    attribute INIT_28 of inst : label is "D29694B5C8EAEE4756D4A930AD5332E806C2CDAA820B5CA52120D17AAF6269B7";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE049A58A2B1BD9898EF487793B1504C7DCB";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1F";
    attribute INIT_2D of inst : label is "1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
    attribute INIT_2E of inst : label is "1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
    attribute INIT_2F of inst : label is "1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "80260512C180481051996A8E938C02B440035400000000053184708855205242";
    attribute INIT_01 of inst : label is "6980AB48A34445A440C0042601DE94A60160AD1DF63558A1549292D9D8440948";
    attribute INIT_02 of inst : label is "02D60080120069960708550004E046415665A75FA8208CB02D23844119055599";
    attribute INIT_03 of inst : label is "AB1500AB1541115045826DC4A491B65A55E2AAA9A639A3C6522556C8C5677750";
    attribute INIT_04 of inst : label is "A9A8831199A66447FF98EEEFFE404708931C7E3381381380E0380E0382285112";
    attribute INIT_05 of inst : label is "115B71128204C8A28FA33713BD142B11846A514C602657094195D04F28042263";
    attribute INIT_06 of inst : label is "6E52905DD8045097A240388090018F6286B160E22235A64E914028E6D2847223";
    attribute INIT_07 of inst : label is "A002EF2ECDADDA6FC628A4122461501E088A0C135BEC6C6B4DAA100CD061660C";
    attribute INIT_08 of inst : label is "424A12FAD28C449AAB4C9D2284FCA6A51B449400380476A9358A84972C6888C0";
    attribute INIT_09 of inst : label is "5001A1816032240110448022CAF6BD1F18DC10C119C99788EDCD6B8A38C6D5DF";
    attribute INIT_0A of inst : label is "6D245EC18B50DD2046A44A58D4A585372112000D4A5D296280334088C1A55BCB";
    attribute INIT_0B of inst : label is "2AAAAA82AAA0000000000002AAA200000254384EC931EE41230D322011754000";
    attribute INIT_0C of inst : label is "AA81249249EA1CC208B2D07F8E317C359E0B0CE4FC8D252622831CE60C116449";
    attribute INIT_0D of inst : label is "FFFC0002AA81FFFAAAFE02AA8001FAAAFFFEAAAAAAAE2AAAAAABFAAABF80000A";
    attribute INIT_0E of inst : label is "AACCC58C3830C4C0410443013038F42EB1305016449555555557FFFEAAA9555F";
    attribute INIT_0F of inst : label is "49500405544554554551445079C0CF7EFA63A6F9410430C10C30C3DF75D12662";
    attribute INIT_10 of inst : label is "FB7DF6CF39F8000108C61004AC850008118541035A008302CEEE66A6590C3ED3";
    attribute INIT_11 of inst : label is "010000000000000020000000000000000000000000000A026AA0000000071DFF";
    attribute INIT_12 of inst : label is "60042D8A95496224446A010157966AE316FD6088C522A6462408B125C2000400";
    attribute INIT_13 of inst : label is "6B4C9D2284800D08401803964D2ABC8004227E9DF5CD8B8F88C60CE120600842";
    attribute INIT_14 of inst : label is "5555500000000000000008FFD6B100D25313D8D093D54E2C11632A62D3044980";
    attribute INIT_15 of inst : label is "4C08D81023604014ABFDD9C9D6632B0212CF7555555555555555500000000555";
    attribute INIT_16 of inst : label is "2000100008000400033C61FBCD66D838AC1E5994966C32289F3046802223920C";
    attribute INIT_17 of inst : label is "44724189E1DB03876C0E0329DFDDA6B310BC0855921935DB1849000080004000";
    attribute INIT_18 of inst : label is "8C4B18F7FA3DC77A3F002A07FDFA954A37F5015AABD8A81F5F22578805088A04";
    attribute INIT_19 of inst : label is "C6A459499672C338AC25B3CC5E4B0824E22EA11435743A185D440459C50D19E2";
    attribute INIT_1A of inst : label is "390C24C69571A9380088904F2B0120113AA5B9D52DC444E2227AF0BA0EA0ED28";
    attribute INIT_1B of inst : label is "79410202A1BBD99D86631580E98B9392CCA0362E39E311A05296352962A17B07";
    attribute INIT_1C of inst : label is "E39D9655C4656DB9C76288C5208AA6C44D3599C4249D900999230092A5D723EC";
    attribute INIT_1D of inst : label is "C6E608CF8C1126BEAF6F9AFECE3D7FC918C4BB14CFB1190649389DB16F499325";
    attribute INIT_1E of inst : label is "7E2D0331F5A01D804D181C3188888C0334D5D07805DC490964EDB797044627DA";
    attribute INIT_1F of inst : label is "B4F98FA92AF5C7604A20D5012660D02A3447E3BBDF93F54FAF5E7AE3FE63334F";
    attribute INIT_20 of inst : label is "F3D79EB935437BCFBFDD48A608CC7866207F17A92AF557DFFA6630F4C006292D";
    attribute INIT_21 of inst : label is "55BD10554C14ECA8E56019069DF3142A413942B529086286281111555518C4B8";
    attribute INIT_22 of inst : label is "6A94A89C2D4309CEF39DE436A4B19DE77BDE40F0100E01B806C831B2A7FE691C";
    attribute INIT_23 of inst : label is "BBBBAAAAAAADE3AAADABD0BD42404A06DE28B405B4586849289401B45A124AA7";
    attribute INIT_24 of inst : label is "0A86104E18966242ED06332E00880D0081014020416DD2C968EAADAAAAAABBBB";
    attribute INIT_25 of inst : label is "CC4BE7654992EB35484D20B047D3B9DA9D7C80DE18825A6806C1309720C8C509";
    attribute INIT_26 of inst : label is "049938009939209E39849C6D4A2B9AF9C524CEC755CEB9346645C449C23AF7F4";
    attribute INIT_27 of inst : label is "671FB0007F03B2092695249D55870B5487D5E75EF7D688A09810801819201819";
    attribute INIT_28 of inst : label is "F7F7BFBCAC42E56217F5CFFDDC676FAA82604491652F8B9E78F3B3608E4BACD3";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F268A2108D7755A24C11D4D140475AF9";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "03AF61A069D0310A5B88220D7FFC0C185155554000000D5883C90C128E060E14";
    attribute INIT_01 of inst : label is "D8149EC4AE64CF384039B38CCCCC958CCBC4A94CA0047521DF684B0CC951B829";
    attribute INIT_02 of inst : label is "025724C98481DA36AC4A310003FFDC71DEEF7836080091B55EAFFDC771E777BB";
    attribute INIT_03 of inst : label is "901222485C6445549622990906D1B9B79B6AAAAB7E7367CE528DDDEA4D720181";
    attribute INIT_04 of inst : label is "9005D91514C4DE619867999800696F3ECF3BCE73A63A23A4E83A0E83A48600D8";
    attribute INIT_05 of inst : label is "A0119A048A6028438424C299EE105CE374CB10F8606024A244443947034276E7";
    attribute INIT_06 of inst : label is "C88518D7CB140414092035272476D9C4ADE2400EEE3EE0EFF35B6054002E0B2D";
    attribute INIT_07 of inst : label is "900016D11211648286BAE572A86A46F629080E143605C06A1900A88D04623B40";
    attribute INIT_08 of inst : label is "1640B2B2148C5410BDC1DFE6B57AC4A08120483C785202550712A80C48CBB8C6";
    attribute INIT_09 of inst : label is "E4100B23403294A41452948AC805291B3B2A42C156A4878A840409020821C098";
    attribute INIT_0A of inst : label is "5C35B7894D559920472518C4E18C6C66099A105918C063120D4004900731DE76";
    attribute INIT_0B of inst : label is "2A2AAA80A280A280AA80A280A282A20000A908245B60B514BB869342150492C8";
    attribute INIT_0C of inst : label is "0000DB6DB7C25A70B13000310C919C2102AB04A582EE7C4EEE370B4024152441";
    attribute INIT_0D of inst : label is "00020000000000000000000000000000000000000000000000000000007FF800";
    attribute INIT_0E of inst : label is "616D80B46EA05242841429A7AC026019B0F22012441000000008000000040000";
    attribute INIT_0F of inst : label is "C114AAAFFFFFFEFFFFFBFBAF860CF2830411C514FFFF3DF1EBED3C208A08F6C0";
    attribute INIT_10 of inst : label is "04820930C606AEAC60CE9945ACB66FF8F2265C600C8CCB0844A4632CDB0E76C1";
    attribute INIT_11 of inst : label is "010000000000040000000000000000000000000000001C126D400000000F2200";
    attribute INIT_12 of inst : label is "CC489B1B1DE68678CC503A0B71BC0014C73F28CA64721EF6E912034B53000400";
    attribute INIT_13 of inst : label is "3DC1DFE6B5080F1540500055055546FCB4A8431146AC115F1B6A127710B20CC2";
    attribute INIT_14 of inst : label is "00000FFFF0000FFFF0000064CE2006E3C7F739C9B605758451832858C3044111";
    attribute INIT_15 of inst : label is "CE5C5BB9716EE1B868665FDCC429791E91E7A000000000000000000000000000";
    attribute INIT_16 of inst : label is "00000000000000000089DAE980C4A0288835551832D67672681157477777D304";
    attribute INIT_17 of inst : label is "EEFA6099CB8B772E2DDC37A8645FBE2159E47A5BC29C31CB7841000300000000";
    attribute INIT_18 of inst : label is "6C510A926896072000004000020000100000800004000020000100000A000CEE";
    attribute INIT_19 of inst : label is "B6407979C42AC12BBF798F6D9BDB0820C2450264B820D03074531914A41045E6";
    attribute INIT_1A of inst : label is "5D6660B350F5BB3208CA9F6CA1FE82167A2EB3D1758CEEC6777DF7264F74E408";
    attribute INIT_1B of inst : label is "3DD34B200011488906F7B17C4B9937B2CDF03C2F32611101463138631B890626";
    attribute INIT_1C of inst : label is "E1698271C5695F4EB22699CD22A88C4EDB65B4E8B587B0AB7B6322B725166705";
    attribute INIT_1D of inst : label is "CC8608B584550412122088384991005B398C960D86933B64DB61B1B324D9B384";
    attribute INIT_1E of inst : label is "782C82207520857F91381C739B898BF125DFC07104240C596CFFB5564CCC7239";
    attribute INIT_1F of inst : label is "6D4DAF29A2A5D234D820882D6C110BB8E0ECB7B3863600E639D9CEE096C6675C";
    attribute INIT_20 of inst : label is "4E7673B36167B601292948A20A8D50C6A069A329A2A5409492C6A108CB47421B";
    attribute INIT_21 of inst : label is "F7216A8052A1073841CCB648022EA53D92E243976A19C6AD4877777777118C98";
    attribute INIT_22 of inst : label is "08F0245846834B8C6719C4220013B9C6338C484E23705A006820D2416EAACB9C";
    attribute INIT_23 of inst : label is "22A22223222002A2200A12804A0A9054854028100488102008281524141A9234";
    attribute INIT_24 of inst : label is "000C52045992E6C2550E6D91529A88129F4204A6D0A8CB2C00A2A843222322A2";
    attribute INIT_25 of inst : label is "8D41D230DBE3830203586292EC97B3F81C7641411D028872022A01A2B408E041";
    attribute INIT_26 of inst : label is "A09C05809C05A09D04249D124E700809986DA443D5BBB362EEE84CDB663A6121";
    attribute INIT_27 of inst : label is "6754B00469A9162B2DB06DBE26E26620B497E71CE7D0ACA49C04849C04A49C04";
    attribute INIT_28 of inst : label is "CE5672B5ACD2ED66961489219D5222701AFCEDD165CA4884202D0360A98E0C0F";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0696C5D4169B101026D9B1918B85743448";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "806EE974D9B2D119BBE00C2D495B033C03777A400000002047E2002100408016";
    attribute INIT_01 of inst : label is "4A0B9250F25C896880000020E44055A0E341B0C45895906C8920DB800141B929";
    attribute INIT_02 of inst : label is "0C1AB4AF0E085A1F141B21924C40A80D9AA968160C9250F8B4F10ABAA03662EE";
    attribute INIT_03 of inst : label is "0A014020239410100002492232D5B4969D67F5717151776EB316758C0FC133C0";
    attribute INIT_04 of inst : label is "0B55103625480667F9FFFFFFFF9690C129BA4B7C40C40C4310C4310C40220450";
    attribute INIT_05 of inst : label is "71B3171E016528C18CA21164A775EA3314D73248B9A66EA46CDCB7572B4A46F7";
    attribute INIT_06 of inst : label is "481E1E5440180014300A93A470080941B4A0C8444452936650EB7095A0EE4A31";
    attribute INIT_07 of inst : label is "00010241320309805238EC76E123DD50044A6598168C87286B13FA26012262CD";
    attribute INIT_08 of inst : label is "524292031CA4D8146526CCA1D3D399B933432C52B164C685650EC0041B491100";
    attribute INIT_09 of inst : label is "74023F394096D2B4B2DA56925B052149004A8AC36480051B0D0D0B000029E898";
    attribute INIT_0A of inst : label is "DD7216872FD2BBF1ED68FEFE7FEFF5A6B31A492BFEFFFBE6CFF472B86160CA42";
    attribute INIT_0B of inst : label is "802AAAAAA02A02AAAAAAA02A002A00AAA9EDAB801B7005D2A34102E136041B69";
    attribute INIT_0C of inst : label is "FFFE104105169B4C4024820924385719A7D6EC98008DE54622A3025240366CC1";
    attribute INIT_0D of inst : label is "0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FF";
    attribute INIT_0E of inst : label is "54D038B5694EE59CC2A91D74088B40BBBE912436CC1000000000000000040000";
    attribute INIT_0F of inst : label is "5560051545050041504040110000EFFFFE73C7FC0000C20E1412C3DD75C0281C";
    attribute INIT_10 of inst : label is "00000000000222EDD33357C84109D0081A1CECE59E01BA698001401092894AB0";
    attribute INIT_11 of inst : label is "010000000000000020000000000000000000000000000C82100000000030C000";
    attribute INIT_12 of inst : label is "D4100106D9900440889A050DE0B514288603301B0D86D2EF400002010EC00400";
    attribute INIT_13 of inst : label is "2526CCA1D382A58554000000441FF021CAED5359552B635E5B5C232A442A1AC7";
    attribute INIT_14 of inst : label is "00000FFFF0000FFFF0000414EF3200DC53134801A54B6480634970A29B0D81C8";
    attribute INIT_15 of inst : label is "2D3A7834E9E0D0303F555969E6A623033AD07000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000008345CD8266BA7CCC74713032CC66404900D924EE66AAEC";
    attribute INIT_17 of inst : label is "88855D85060E04183810043F5550C735208C0CA1A559391B04C1000300000000";
    attribute INIT_18 of inst : label is "0CC3020920805280000000000000000000000000000000000000000000241499";
    attribute INIT_19 of inst : label is "0200ADAD66B5BB26AB15AAC8594310E0860C30043186030800C0B39EF5B98A31";
    attribute INIT_1A of inst : label is "AB6F60B7532B4B3101DA602D730181707A4DA2D24D8CCCC4444440146C568C3B";
    attribute INIT_1B of inst : label is "194102000088444312843642C45036D0D6CA990C24203205FFBF9FFBFCB3021C";
    attribute INIT_1C of inst : label is "004880678D9E9F4080169DED09B0480ED96490586D94B01B4B6301B7A5D64480";
    attribute INIT_1D of inst : label is "001439240063052120681A0001A35552AD292409B402336CDB5137B2C099B309";
    attribute INIT_1E of inst : label is "6A6C0EA07520050000AD4B5AD98D8E0B2071C520088008186C2BBDF608CD4148";
    attribute INIT_1F of inst : label is "4A056977572B201690E3AC726E9A243CA8CC9B67302548B41858C2C4015269D0";
    attribute INIT_20 of inst : label is "061630B24AD20002404AD9C01B39875CC000E977572BA120075CCE18EDC6E152";
    attribute INIT_21 of inst : label is "5D218FD863F6CC18C50E309928320E902620E9327DD843F41F66662222218D50";
    attribute INIT_22 of inst : label is "8472174D0ED75E310C6203A73937C31886303AC000004000000000007EAADB4A";
    attribute INIT_23 of inst : label is "A222AAAAAAAB0E2223060A5429CB26D9308C6C2F6218D856C4CC2E4236052114";
    attribute INIT_24 of inst : label is "D364D62CDBB6F6F6DCAD6DA576BBE1E6B97879AE5E1182A8D382230EAAAAA222";
    attribute INIT_25 of inst : label is "B98900169ADAC16B1C9A62B0CCAB676D39A56841BBA21E67473F6C86F72A59E1";
    attribute INIT_26 of inst : label is "048000048000248001208003018FBBA49A6DC000D5BAB24AC8AE089244A6300A";
    attribute INIT_27 of inst : label is "CE61D00000B0062B0D3A49BA60A604B148BECE69CDAD30240000248000048000";
    attribute INIT_28 of inst : label is "861630B1BED6CDF6B7A4600EB9801058A4C0CD95641ABC2011092561B16B05A6";
    attribute INIT_29 of inst : label is "00000001FFFFFFFE00000001FFFFFE000495F629125656049025092BC54BA502";
    attribute INIT_2A of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_2B of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_2C of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_2D of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_2E of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_2F of inst : label is "00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE00000001FFFFFFFE";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "8822613048921C3FF93772D1CA5601C44C913FC000003FDFB81DFFDEFFBF7F70";
    attribute INIT_01 of inst : label is "33068918B12444CF7FFFFF930D9FA6130C248F1DC672492044B7B419DC2E48E0";
    attribute INIT_02 of inst : label is "8AE600823214232722681E61B568881046648D4DF30D99396215A88220411199";
    attribute INIT_03 of inst : label is "91B2364000001101FFF92667C9014248E0D2AAFC9270874FF329925AC517DD46";
    attribute INIT_04 of inst : label is "015F7B99B4CC419E61980067FE000000193E227000000000000000000364EC8D";
    attribute INIT_05 of inst : label is "221C722224C52064878136A0AF7A4181C0469D67363B945983077105D1B622E7";
    attribute INIT_06 of inst : label is "33E5C90CD82597C3C650C0A89101A426A213442223B2489242693870D32E3947";
    attribute INIT_07 of inst : label is "FFFEDB25DB2592D91869A0D12586245890A11042C8704885862CA850B28F8644";
    attribute INIT_08 of inst : label is "C33E185AD6B267CFA4912484C96782C61C87B47001987930309ABFF248208EFF";
    attribute INIT_09 of inst : label is "9148C964314B284B5965096B2CB4A56508CF9E499CCD97CCFCFCF980000457C7";
    attribute INIT_0A of inst : label is "70E84C4D110C66227DFCFFF4EDEF6613E92186C6FFF37BD325519268108E2109";
    attribute INIT_0B of inst : label is "002AAAAAA00002AAAAAAA00000020000038C0CCCDB6DE6482B2CB24499F24004";
    attribute INIT_0C of inst : label is "0000C14815181A830313F96DB184089892EA022886AC77271B93DE79EC996E7C";
    attribute INIT_0D of inst : label is "00000000000000000000000000000000000000000000000000000000007FF800";
    attribute INIT_0E of inst : label is "1628864298A02D874D5689204B065E08BF919C96E7C000000000000000000000";
    attribute INIT_0F of inst : label is "3C90AAEAAFFAABFEAAFAEEBF0008000000000000C000000000000000000D1443";
    attribute INIT_10 of inst : label is "F03CF00F00F04000CC137145AF16400983246210E2228806AE6E67E2DB2C22CB";
    attribute INIT_11 of inst : label is "010000000000040000000000000000000000000000000800000000000030C00F";
    attribute INIT_12 of inst : label is "404FE49A845B6224476881936EB0C7E19643306C261332D73FFFFDFC92000400";
    attribute INIT_13 of inst : label is "64912484C880314C155005551175590015333FC6B0E19CCAA4C8C6201061485A";
    attribute INIT_14 of inst : label is "000000000000000000000EDC031102C773D38840B63FE6EC996CF8EEE3267CC8";
    attribute INIT_15 of inst : label is "0C895A12A5E848164C445C846278E000FCD8B000000000000000000000000000";
    attribute INIT_16 of inst : label is "2000100008000000005B407FCEA2617EC5AAF8B630D6222E4CB275902222D600";
    attribute INIT_17 of inst : label is "445AC001912B4254BD09024C44590B13C78003E5BE1F3103027C000000004000";
    attribute INIT_18 of inst : label is "AFFCD96CB25B18D8000040000000000000000000040000000001000005BFC604";
    attribute INIT_19 of inst : label is "CA3E3333E27A808A0B39D24F9E4BC93E1FF3E1543F7CBE082BE51504A61E1D02";
    attribute INIT_1A of inst : label is "0E929E7FDD2F6B3E04E5A02F2F00069D6326BB1935C46CE23671519DCDCCF04C";
    attribute INIT_1B of inst : label is "795302200133D999D8C630C0049BB722E950CA2C95BB99F27FFD3B7BD9C9F934";
    attribute INIT_1C of inst : label is "9BCEF651E6554D1AE66689CD14EF86C45B6DBDC9258C9049C96B0496641632EF";
    attribute INIT_1D of inst : label is "41664CE66CD9F29697E5F96EDF9BAADB3885B30F07B11192DB68B1392E59B32D";
    attribute INIT_1E of inst : label is "28EC122075200518FF3862739961A6008212418023DBE7D96CCDB9B7C4443DC8";
    attribute INIT_1F of inst : label is "6FDDADFFFF9F5768D820B4276E71B29E2C4656FBCBB6AC66FB5BDADDD82939F1";
    attribute INIT_20 of inst : label is "DED6F6BB6FFA37FB7BCFE7F64CDE5A2F201BADFFFF9F5DBDD82F31FAC057A01B";
    attribute INIT_21 of inst : label is "E49E3AA78EA870C86430C92C0D89250E5B935081822024826811111111D8C45E";
    attribute INIT_22 of inst : label is "3B8CEC74F2CD314AD294BCFCF3ED34A52B5BCDBFFFFFBFFFFFFFFFFFBD57DB9C";
    attribute INIT_23 of inst : label is "AA2AAAAAAAAC9A2AAC9B75B9D666CBB65E7814659DE028CB3834619C0A30CEE3";
    attribute INIT_24 of inst : label is "2E138CB39EB6E6C6F70432189C6E971C6BC5C71A31CF2AA92682249AAAAAAA2A";
    attribute INIT_25 of inst : label is "5E417768F3C88C2D09DB60C04646FBF5DC7C6021C981E1230CEB02780D8B0F5C";
    attribute INIT_26 of inst : label is "20000020000000000000000510141056636D8CF7C598BB6E0460E45B5332CBB0";
    attribute INIT_27 of inst : label is "F79600001B4BB60C05AB6DBA30A306D09E57F71EFBF7C8200000200000200000";
    attribute INIT_28 of inst : label is "DED6F6BC9C4AE4E2565DBBB05E7776280EC045BF12F95DEF6F798164CB2230BD";
    attribute INIT_29 of inst : label is "0000000000000001FFFFFFFFFFFFFE01B6DC3013CB838362DA19A5B8441C359C";
    attribute INIT_2A of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_2B of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_2C of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_2D of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_2E of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_2F of inst : label is "0000000000000001FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFE";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "80020100C080581FF1166AE9C43000AD04423FC0000000000000000000000062";
    attribute INIT_01 of inst : label is "211089083104448D400000368DDEA5368A20AD5DC221482845B292DDD8652041";
    attribute INIT_02 of inst : label is "8AD6008016102117222A1D209568004846648FCDE90488B92015A00001211199";
    attribute INIT_03 of inst : label is "8811022000110000000364EFA08126C8D4D2AAFC92208245F3055258C55755C2";
    attribute INIT_04 of inst : label is "204F731194CC47F99867FF980000000019162220000000000000000000220440";
    attribute INIT_05 of inst : label is "110A3116005500200203375F5085BD51A0441155320A984B4109700441962242";
    attribute INIT_06 of inst : label is "27548A1CD805B687A64085803001A420A210442222B021420160182070881023";
    attribute INIT_07 of inst : label is "00024924D92496D91069A0D0250D140001C120824848490F443A10E097054608";
    attribute INIT_08 of inst : label is "461A304A52A0468EA0428402C0B30B250A479C70115424A81082801228208A80";
    attribute INIT_09 of inst : label is "3001AA68718C20496184092A30B5AD4508C79EC11C499688C8484080001494CB";
    attribute INIT_0A of inst : label is "20C048410B444F42BCF84A58A4A5C813A11082444A592962002352F800840109";
    attribute INIT_0B of inst : label is "002AAAAAA00002AAAAAAA00000020000030622EEC939E220290C32201106E010";
    attribute INIT_0C of inst : label is "0000DA04050A0AC3068AF16CA1961CD457C2042806A5550C8A869E39CC112468";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "1200242358082D87CC02090009065C189F919C12468000000008000000040000";
    attribute INIT_0F of inst : label is "285001155000005555045014FBC70000018C38000104F2CF18630CE186010012";
    attribute INIT_10 of inst : label is "F03CF00F00F0088168D37004A71540009114600056028002AE4F37A649242643";
    attribute INIT_11 of inst : label is "010000000000000020000000000000000000000000000800600000000000000F";
    attribute INIT_12 of inst : label is "80002C8284492224457A00886E9047E3B4C2300A050AB253000000048A000400";
    attribute INIT_13 of inst : label is "E0428402C18021080000000000201808010A3C8CA0408A8AD2C446200060084A";
    attribute INIT_14 of inst : label is "000000000000000000000EDC448DFA555656C840931FA24C1128F84A490468CC";
    attribute INIT_15 of inst : label is "44894812A5A048124C444DCC9158E102F8881000000000000000000000000000";
    attribute INIT_16 of inst : label is "200010000800000000002DFFCD11604D22AAE422185222264430449022228604";
    attribute INIT_17 of inst : label is "4450C08891290254B409024C44498C8AC7840BE51C8991090068000000004000";
    attribute INIT_18 of inst : label is "A5EA9B6DB6DB10C8000000000200000000008000040000000000000004BF8204";
    attribute INIT_19 of inst : label is "EA3C3A3A5150810A0B68A2E4885988341EABA1141D743A0001E4104109151800";
    attribute INIT_1A of inst : label is "08435465A52F69920084A087220002152406992034C466623331518CE4CE4008";
    attribute INIT_1B of inst : label is "7D5142000133D998D04212C0448993B64DD08A65B4B311E31296292973010904";
    attribute INIT_1C of inst : label is "93C6E65344554D1A77630886108E86C44A289DC0249C9009C92900922C12324E";
    attribute INIT_1D of inst : label is "413208E24C11A286864190664D8A2A891084930513B1110A493891190E4B1624";
    attribute INIT_1E of inst : label is "68E40220752005547D1042210F00C60102528100014947CB25CD99B3C4443DC8";
    attribute INIT_1F of inst : label is "27D885FFFF9F576048413C072630909E244647DEC992AC727949CA49C83139F1";
    attribute INIT_20 of inst : label is "CE5272992FFA136933C7EFE608F44A3A203B0DFFFF9F1499C83A31F24013E089";
    attribute INIT_21 of inst : label is "849D1057441428802068A96C0499040E4B91408142502082081111111158C44C";
    attribute INIT_22 of inst : label is "6A8DA810A804114AD6B5A4D476A514A52B5A46800000000000000000D5555110";
    attribute INIT_23 of inst : label is "2222222222258A22258BD4BB5222D996CA281C21B5503843683C21B41E10DAA3";
    attribute INIT_24 of inst : label is "3A2285A28A12424269043B089422BD34224F4D091345020B62AAAD8A22222222";
    attribute INIT_25 of inst : label is "744037605141000709C920804657DED4F4DC01018801512004C02454258A0548";
    attribute INIT_26 of inst : label is "001800001800001800001807009401544124EEE7C498992C0644E4490390C390";
    attribute INIT_27 of inst : label is "BD1200003B0BB20804A9249A10A102709E45BD37BF7788001800001800001800";
    attribute INIT_28 of inst : label is "4E52729C984264C21249B394747776384E4044A620F91DCE667881208904001F";
    attribute INIT_29 of inst : label is "00000000000000000000000000000003B2586213C94141224A1CAC90C01C14DE";
    attribute INIT_2A of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2B of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2C of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2D of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2E of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2F of inst : label is "00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
