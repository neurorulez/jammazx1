-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_7J is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_7J is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_7J_0 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"3A3A27F4A0000800020027F480000800026000A80180280002A0027CAA801600",
		INIT_02 => x"00AA0000003E1FD8000A0000ACAC1FD80002000000801FD8BC0327F4F4000000",
		INIT_03 => x"00280F0C00000F000000003C00000F00002A0F3CA8000F000000003C00000F00",
		INIT_04 => x"00280F0C00000F000000003C00000000002A0F3CA8000F000000003C00000000",
		INIT_05 => x"00280F0C00000F000000003C00000A00002A0F3CA8000F000000003C00000A00",
		INIT_06 => x"00AA005002A88A0000A80005A800400000780B6AB400A78000A8016AA800A500",
		INIT_07 => x"2A8000A2AA00050000020000A8008A00002A000002A88A1400020010A8008A00",
		INIT_08 => x"007C2FBFF400FBE0002A00A2800000002A8014A2A8000000002A00A280000400",
		INIT_09 => x"017E021E00B00500002A03AA02F8DFD00E000050BD40B480007C3D5FF400D5F0",
		INIT_0A => x"0000F330000000870000F32F0000FD070000F390000015802F8007F6A800EA40",
		INIT_0B => x"00003F5100085FD00000083F0000FC000000003F8000FC000000003FC000FC00",
		INIT_0C => x"00A80B6AA800A7800AA03C2A028095F000A8016AA800A500200007F5000045FC",
		INIT_0D => x"00803696000899BC000010170000F81C0300116904C0445C000011690000445C",
		INIT_0E => x"0280050B0A80F1800280056F0BA0F3C0028000030BE8F980028005030BE8FC80",
		INIT_0F => x"00000FFF0000FFF00000000000000000000005410000A1500000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000FFF000007F00000030A800005FF00000FC3F0000C2A8000000FF0000FFC3",
		INIT_12 => x"000014AA0000A85000BC0000F800000000780500B400014000780B6AB400A780",
		INIT_13 => x"0000000000000000000002A00000F8300000000000000000002A3FBFA000FBF0",
		INIT_14 => x"0004001700008340000100070000830000000017400083400020401720008350",
		INIT_15 => x"0000008500006000000000800000560000000080000005600000008000000054",
		INIT_16 => x"0000008000000054000016800000000400000560000000000000005600000000",
		INIT_17 => x"0000023F0000F4300000029F0000C830000002A700007830000002A100007830",
		INIT_18 => x"00000A020000A02000000A820000A02000000A800000A02000000A020000A020",
		INIT_19 => x"000002A70000FC30000000000000000000000A020000A0A000000A0A000082A0",
		INIT_1A => x"0000028B0000F830000A05A0A000F85000003FF00000F3FC00002FA00000B8A0",
		INIT_1B => x"000003FF0000F81000080BFE0000F290000202F80000F8B4000002BF0000F0B0",
		INIT_1C => x"000000D40000CCCC0000005C0000CCCC0000005C0000CCCC000000300000CCCC",
		INIT_1D => x"000030CC0000CCCC000000DC0000CCCC000030CC0000CCCC000000D40000CCCC",
		INIT_1E => x"0000D4CC0000CCCC00005CCC0000CCCC00005CCC0000CCCC0000305C0000CCCC",
		INIT_1F => x"000044D400000000000044CC000000000000445C000000000000445C00000000",
		INIT_20 => x"00000000000000C000550009054F00030000030000000000F150C00055006000",
		INIT_21 => x"0000000000026181150500004000010380000249000000000000C04054540000",
		INIT_22 => x"20005000800300005450000900000000C0030000000800140000000005156000",
		INIT_23 => x"20005000800300005400000000000000C0030000000800140000000000150000",
		INIT_24 => x"000000000000000000000000007E00100000000000000000EF40010000000000",
		INIT_25 => x"0000000000000000000000000515000000000000000000005514000000000000",
		INIT_26 => x"00000000000000000000000001FF00000000000000000000FFD0000000000000",
		INIT_27 => x"00000000000028000000000000BF00000000000A000000007F80000000000000",
		INIT_28 => x"C3FFC3FFFF1F3FEAC3FFC3FFFE005400FFE38000FFFF00000000000000AB0000",
		INIT_29 => x"C3FFC3FCFFFF0001C3FCC000FFFF0000FFFF557FAA00FFFFFFFF0000FFFF0000",
		INIT_2A => x"FD030000E0003FAA5000000A0004FFFF0000380000007FFF00170388F00B1EAF",
		INIT_2B => x"0000FFFF0000FFFFA0000030000000000015FFFFFFFFAA0000070000F00C0A02",
		INIT_2C => x"00002D5E000002E000000B5F00003C0F00003D540000F2F400003C0F00003D54",
		INIT_2D => x"0009CC9255554000CCCC618600001AAA55550001600086330000AAA433339249",
		INIT_2E => x"0F0F0F0F0F0F0F0F0F0F0F0F0F0FFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_2F => x"0000000000000000FFFFFFFFFFFFFFFFF0F0F0F0F0F0F0F0F0F0FFFFF0F0F0F0",
		INIT_30 => x"00000F0F000000000F0F0F0F0F0F0F0F00000000000000000000000000000000",
		INIT_31 => x"00000000000000000000000000000000000000000000F0F0F0F0F0F0F0F0F0F0",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"00ABD000EFD0BFFFF2BF4000400FFFFF0033402A42D00000FE28FFD03FD003FF",
		INIT_35 => x"FFFF0000CF8015FFE003AFE0FEA8FFFF07F8FFF8083F07FC000000000000AB00",
		INIT_36 => x"B330000F70BE00003F03FF0052FCFFFF005FFFFEFFFF000100FFF800FFFE7FFF",
		INIT_37 => x"E0FC7C8334002D2C04C54B2214AA0A001420030A1C80F003FFF000001554BFFF",
		INIT_38 => x"EA00FFFF0000FFFF0000FFFE1FFF00000055FFEAFFFF0000FFFF01FFFFFFFFFF",
		INIT_39 => x"02CF8000FFF000AA0000FFFF0000FFFF200B01FD00000FFF0000FFFF0000FFFF",
		INIT_3A => x"FFFF0000FFFF0000FFFFFFFFEA00FFFFFFFF0055FFC3FFC30000FFFF0003FFC3",
		INIT_3B => x"0000FC7F002FFE000000FFFF0000FFFFFFFF1FF5FFC355430000FFFF0003FFC3",
		INIT_3C => x"00000000000000A500D10003F4049E000000E000000000001A00600000000000",
		INIT_3D => x"000000000000603C000000002B4B000000000B00000000008FA0000000000000",
		INIT_3E => x"0000000000000004100100000402204080000080000020000800081002000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7J_1 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"1F45284F5C00CC000B91284F0000CC00014E013CA0782900003F023CF0003C80",
		INIT_02 => x"0064003CBEDBF1280035003C51F4F1280000003C46E0F128E7AB284F5900CC00",
		INIT_03 => x"02D0050500007D00000000160000A40002FD07BD7F807F800000001500005400",
		INIT_04 => x"02D0050500007D00000000160000A50002FD07BD7F807F800000001500005500",
		INIT_05 => x"02D0050500007D00000000060000A40002FD07AD7F807F800000000500005400",
		INIT_06 => x"01FE00032FC0C7402BFA0000BFA0000000BE3D57F80055F000BE001DF800D000",
		INIT_07 => x"03F801D3BF40C000000B0003FBD4C740007E00032FC0C74000AF0003FBD4C740",
		INIT_08 => x"00FF1409FC00805017FF01D3E000C00003F801D3BD00C00017EF01D3FA00C000",
		INIT_09 => x"02FF0545FF4000002ABF000DEFF5D00001FF0000FF8051500057000054000000",
		INIT_0A => x"000041C001800000000041FF0008FD54000043FE000155405FFB0007FE2870C0",
		INIT_0B => x"0000102E0000F80000000E994000D008000218196000D0A4000200397000D600",
		INIT_0C => x"00BE3D57F80055F003FA00FDBFC0405000BE005FF800D4000000002F0000B804",
		INIT_0D => x"00B600940098232402F800E02F807E0003F000E008C03E0002F000E008803E00",
		INIT_0E => x"2E1F005ED5002B202E9F005ED7409F602E1F005ED7D0DF602E9F005ED7D59FF0",
		INIT_0F => x"0095071F5600F4D0000000000000000000AF00A80A00AA000000000000000000",
		INIT_10 => x"0000FFF000003F00000030FF00000FF00000FC3F0000C3FC000000FD00002AAF",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000007C0000F40003FA0000BF00000000BE0000F800000000BE3D57F80055F0",
		INIT_13 => x"0000000000000000005501FCE8003F30000000000000000002FF0001FE000000",
		INIT_14 => x"030800A80700F800038800000B00F800034800000300F8000308000A0300F880",
		INIT_15 => x"0000007800000000000000780000000000000078000000000000007800000000",
		INIT_16 => x"0000007800000000000000780000000000000078000000000000007800000000",
		INIT_17 => x"005501E5E800FF30005501F9E8007F30005501FCE8007F30005501FCE8003F30",
		INIT_18 => x"000007F400007F40000007F800007F00000007F900007E90000007E500007E50",
		INIT_19 => x"008507FCE2007DD00000000000000000000007FD00007FD0000007FD00007F50",
		INIT_1A => x"02D501E7E800FF30004701F6D800BF30005B05BEE0003E5002550FDC698033F0",
		INIT_1B => x"00A501FFDF8076D000B50DFF6F8037D000BD03FF68003CD000AF07FDCE007ED0",
		INIT_1C => x"0000005400005454000000540000545400000054000054540000005000005454",
		INIT_1D => x"0000505400005454000000540000545400005054000054540000005400005454",
		INIT_1E => x"0000545400005454000054540000545400005454000054540000505400005454",
		INIT_1F => x"0000005400000000000000400000000000000054000000000000005400000000",
		INIT_20 => x"000002A00200061300000090A48203030080C49000000A80821AC0C000000600",
		INIT_21 => x"06000542080384000000009020000801C0300012009085400008003000000600",
		INIT_22 => x"06000050400100000000000000000C0340000000009005000000C03000000000",
		INIT_23 => x"0600000040010000000000000000000040000000009000000000000000000000",
		INIT_24 => x"000000000000000000000000002A00000000000000000000AA00000000000000",
		INIT_25 => x"00000000000000000000000008BF00000000000000000000FF88000000000000",
		INIT_26 => x"0000000000003F800000000000150000000080BF000000005500000000000000",
		INIT_27 => x"0000000000001F800000000002F40000000080BD0000000007E0000000000000",
		INIT_28 => x"C3FFC3FFFFCF8500C3FFE050FF800000FFF000001FFF00000002000095400000",
		INIT_29 => x"C3FFC3CAFFFFAA00C3FEC0003FFF0000FFFF0000FFFF057FFFFF0000FFFF0000",
		INIT_2A => x"500000007800BD5000000AFF0000FFFF0000070000023FD40007E3EFFAAAEAF4",
		INIT_2B => x"AA00FFFF0000FFFFF4000038000000000000FFFF057FFFFF00010000F80C3F03",
		INIT_2C => x"00003C0F00002F7E00003CAF00003D5F00003EA00000F5E800003EEF00003EA0",
		INIT_2D => x"0092CCCC55550000CCCC061800006AAA55550000860033330000AAA933332490",
		INIT_2E => x"0F0F0F0F0F0F0F0F0F0F0F000F00000000000000000000000000000000000000",
		INIT_2F => x"00000000000000000000000000000000F0F0F0F0F0F0F0F000F00000F0F000F0",
		INIT_30 => x"0FFF0F0FFFFF0FFF0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF0000000000000000",
		INIT_31 => x"FFFFFFFFFFFFFFFF0000000000000000FFFFFFF0FFF0F0F0F0F0F0F0F0F0F0F0",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"AF7F000CF4007FF4ABF4000B00AAFFFFA030081D2F4002FDAABFFF4001400FFF",
		INIT_35 => x"FFFFAA00CFFE0005F803FFF8FFFC5500007C7FFF2F0FE07F07FF002FFAAA5B80",
		INIT_36 => x"53380F0F001F80401502FF00BFFFFFFFE0017FFFFFFFE000003FFE00FFFF0FFF",
		INIT_37 => x"FC701442B080D2FCA065830E5550604002FC010500C040000000FA8000000055",
		INIT_38 => x"FFFA1FFF8000FFFFE000FFFF01FFE0000000FFFF0055FA80FFFF001FFFFFFFFF",
		INIT_39 => x"2FCF40A8FD507FFF0000FFFF0000FFFF0E2F0050000003FF0000FFFF0000FFFF",
		INIT_3A => x"FFFF0000FFFF0000FFFFFFFFFFFAFFFFFFFF0000FFC300438000FFFF0003FD0B",
		INIT_3B => x"00AAFC15D07F55400000FFFF0000FFFFFFFF0000FFC300030000FFFF0003FFC3",
		INIT_3C => x"000000000002A264000B00005680506900009000000000002460C00000000000",
		INIT_3D => x"00000000000006F30000000003B400000000B700000000007C05000000000000",
		INIT_3E => x"0000001000800801020800010000000002000000000000008004402000200000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7J_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"06FF0F92BD00C0000EFF0F92BD00C0000FC30394FE203EC00F8300E8EE403D40",
		INIT_02 => x"007E0006FFB086F0007E0006FF9086F0007E0006FFB086F00EFF0F92BD00C000",
		INIT_03 => x"0F0D00005F000000003C00030E00F0000F3D007F5F00FD00003D00005E000000",
		INIT_04 => x"0F0D00005F000000003C00030500F0000F3D007F5F00FD00003D000055000000",
		INIT_05 => x"0F0D00005F000000002C00030E00F0000F2D007F5F00FD00002D00005E000000",
		INIT_06 => x"281500005D0001003FAB0000ABF000000057000C5400C0002857000454A04000",
		INIT_07 => x"0075004054280000002F000057400100001500005D00010000FD000057C00100",
		INIT_08 => x"00AB0004A800400001D50040FA000000007500405400000003D500407F000000",
		INIT_09 => x"2FE10300542000003D5500007F404000081500004BF800C000FF0000FC000000",
		INIT_0A => x"60000000006000006000007F0036FFE8600001FF000FFA8001FD0001557C0000",
		INIT_0B => x"280002FD0030FFA00003000070000100000301007000010000031A2470000600",
		INIT_0C => x"0057000C5400C000005D0044540000000AD700045E8040000C000AFF00287F80",
		INIT_0D => x"01F200788CC03E9002BD00145FF83D000A7B0014C6C83D000A7B0014C6C83D00",
		INIT_0E => x"006B000008005AEC2A9C000008005AF80A6B000008005A780A7B00002C005E78",
		INIT_0F => x"090A006A8060A9000000000000000000005700502D00F5000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"FFFF57F0FE003F00FFFFF054FFFF2D50FFFF5415FFFFF85200BF00FEFFFF154B",
		INIT_12 => x"02EB0054BA00540001050008410020003E57000056F000000057000C5400C000",
		INIT_13 => x"00000000000000000FF8001407800F0000000000000000000BD700045F804000",
		INIT_14 => x"01C500800B005000018500020B005000018502400F00580001A580002B005018",
		INIT_15 => x"0020000000000000000200000000000000000000200000000000000002000000",
		INIT_16 => x"0000000002000000000000000020000000000000000000000200000000000000",
		INIT_17 => x"0FF2001487800F000FF8001407800F000FF8001407800F000FF8001407800F00",
		INIT_18 => x"268B005EE2F805002F89005FA2F885002F8B005FE2680500268B005EE2F80500",
		INIT_19 => x"01B800448640010000000000000000002F89005FA2F8A4002F8B005FE2688500",
		INIT_1A => x"0FF8019503E00F400FF8000F45A0FF000FE7001BD380FF000FDB0116E7808E40",
		INIT_1B => x"0368001501F005000168019D1FF0010009680055FF800F000BFC005401400F00",
		INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"00600000030358410150000009230100C0C0412509000000C860004005400000",
		INIT_21 => x"006000000C00100002A1090048000C0380100004090000000021C01042A00060",
		INIT_22 => x"000000000C03000000A0090000000002C030000000000000000080020A000060",
		INIT_23 => x"0000000000000000000009000000000200000000000000000000800200000060",
		INIT_24 => x"0000000000003E2A00000000001F00000000EA2F000000007D00000000000000",
		INIT_25 => x"00000000000000AA0000000007F400000000EA800000000007F4000000000000",
		INIT_26 => x"000000000000007F00000000000000000000FF40000000000000000000000000",
		INIT_27 => x"00000000000001FF00000000054000000000FFD0000000000054000000000000",
		INIT_28 => x"C3FFC3FFF543E000C3FF3800FFFF0000FFFC000001FF0000E000000000000000",
		INIT_29 => x"C3FFC3C3FFFFFFFFC000C00000000000FFFFFAA8FFFF00000000000000000AAA",
		INIT_2A => x"50000000000040000000555500005555000000C00ABF0400000051557FFF5540",
		INIT_2B => x"FFFF57D4AA0000000000A00E00000000000000000001003F0000000000003FCB",
		INIT_2C => x"00003C0F00003C0F00001E0000001E2D00003C000000F03C00003F7F00003C00",
		INIT_2D => x"0924CCCC95550000CCCC00610000AAAA55560000186033330000AAAA33334900",
		INIT_2E => x"0F0F0F0F0F0F0F0F0F0F0FFF0FFFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_2F => x"0000000000000000FFFFFFFFFFFFFFFFF0F0F0F0F0F0F0F0FFF0FFFFF0F0FFF0",
		INIT_30 => x"0F000F0F00000F000F0F0F0F0F0F0F0F00000000000000000000000000000000",
		INIT_31 => x"00000000000000000000000000000000000000F000F0F0F0F0F0F0F0F0F0F0F0",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"FF3D002F002F1F40FF40000502FF5555F0002C007D0C0BFCFFFC550000FF0555",
		INIT_35 => x"5FFFC0FFC5FF0000000055000000000AE000015F3FC3FE87000080020AAAFF40",
		INIT_36 => x"011C0F0F0007C000FF035500FFFF5555FE000FFF17FFFE00C00F5500FFFF0155",
		INIT_37 => x"FC304001D2E02FDA18750307555F8E0201FD001001500080FFFEFFFE0155A000",
		INIT_38 => x"FFFF007FFEA0FFFFFE005555000754000000FFFF0000FFFEFFFF0000FFFF5555",
		INIT_39 => x"01C5F81C40001FFF55540055FFFAFFFF0FFFC00400AA015017FFFFFFF4BFFFFF",
		INIT_3A => x"0055A000FFFF0000FFFF5555FFFF5555FFFF0000FFC30003FEA055550003502C",
		INIT_3B => x"FFFF0000800F0000FFE0FFFF3E1FFFFFFFFF0000FFC30003FFF8FFFF03C3FFC3",
		INIT_3C => x"0000000200284181000C0000300100A900001E000000000041B0000000000000",
		INIT_3D => x"0000000000002F400000000003400000000043B4000000000600000000000000",
		INIT_3E => x"0000000100010000000000000010040400081010040040000200800000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7J_3 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"012D004140000000013D0041400000000197005CC7403C0001970004C7001400",
		INIT_02 => x"000000005C4041000001000078404100000100007C404100013D004140000000",
		INIT_03 => x"0F0E0000AF000000003C00000D0000000F3E0000AF000000003E0000AD000000",
		INIT_04 => x"0F0E0000AF000000003C0000080000000F3E0000AF000000003E0000A8000000",
		INIT_05 => x"0F0A0000AF000000000800000D0000000F0A0000AF000000000A0000AD000000",
		INIT_06 => x"1FFF0000FFFC0000076A0000A740000000FF0000FC0000001FFF0000FFD00000",
		INIT_07 => x"3FFF0000FFF40000001F0000FFF000000F070000DFF80000007F0000DF400000",
		INIT_08 => x"02D500005E0000000FFF0000F50000002FFF0000D0F0000001FF0000FD000000",
		INIT_09 => x"7F7500007BFC00001FFF0000EABC00003FED00005DFD00000B6A0000A7800000",
		INIT_0A => x"C80000000A1E0000D8000000001F0000D8080055023755553EAB0000FFF40000",
		INIT_0B => x"3F80005500185555002C0000F8000000002C0000F8000000002C0050F8000100",
		INIT_0C => x"00FF0000FC0000003FFF0000FEA000001FFF0000FFD000002400555502FC5500",
		INIT_0D => x"2D950000694CB4003FFF0000807C54003C680000362C54003C680000362C5400",
		INIT_0E => x"3AC600008F00004E3C060000A600004E35C60000D600004E03C600008600005E",
		INIT_0F => x"0CBF0000FE30000000000000000000000A81000012A000000000000000000000",
		INIT_10 => x"FFFAFFFFFF00FD0030F4FFFF2FF0FFFFFC3FFFFFC3FCFFFF00FD007F2A87FFFF",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"2FFF0000FFE00000000000FC0000FC003EDF0000DEF0000000FF0000FC000000",
		INIT_13 => x"0000000000000000105F0000E0E0100000000000000000001FD500005FD00000",
		INIT_14 => x"0A0A0100D2800020021B0003920000000A1E0400928001008A1A000094A00000",
		INIT_15 => x"000F0000C000000000000000FC000000000000000FC000000000000000FC0000",
		INIT_16 => x"0000000000FC00003C000000000C00000FC000000000000000FC000000000000",
		INIT_17 => x"10FF0000F8E01000107A0000E0E0100010570000E0E010001057000060E01000",
		INIT_18 => x"F03F000003F00000F03F000003F00000F03F000003F00000F03F000003F00000",
		INIT_19 => x"105B0000F8E010000000000000000000F03F000003F00000F03F000003F00000",
		INIT_1A => x"051F0000E07010003FCF0005E3FC50003FDE0005A2A0500010470001D0E04000",
		INIT_1B => x"10FF0000E0A4000010FF0000E1601000105E00005DE01000107F0000E0E01000",
		INIT_1C => x"005C0000DCDC0000005C0000DCDC000000D40000DCDC000000740000DCDC0000",
		INIT_1D => x"74DC0000DCDC000000DC0000DCDC000074DC0000DCDC0000005C0000DCDC0000",
		INIT_1E => x"5CDC0000DCDC0000D4DC0000DCDC00005CDC0000DCDC000074D40000DCDC0000",
		INIT_1F => x"645C00000000000064AC000000000000645C00000000000064D4000000000000",
		INIT_20 => x"000600AA00030A8F0000000000C00000C000F2A09000AA000300000000000000",
		INIT_21 => x"00002A2A020300000000000092400001C08000020000A0A88186400000000000",
		INIT_22 => x"0006A8A000000000280010000000C0030000000090000A2A0000C001000A0004",
		INIT_23 => x"0000A80000000000280010000000C003000000000000002A0000C001000A0004",
		INIT_24 => x"00000000000007E700000000002D0000000076F4000000001E00000000000000",
		INIT_25 => x"0000000000000BE50000000000000000000056FC000000000000000000000000",
		INIT_26 => x"00000000000002F50000000000000000000017E0000000000000000000000000",
		INIT_27 => x"0000000000000015000000000000000000009500000000000000000000000000",
		INIT_28 => x"C3FFC3FF5001F800C3FF05EAFFD5AAAA5FFE0000040000000000AAAA0000AAAA",
		INIT_29 => x"C3FFC3F1FFFFFFFFC000C0000000002AFFFFFFFFFFFFFA800000AFCA0000BFFF",
		INIT_2A => x"00002A40200000090000AAAA0BCAAAAA0010550BFFFFC0000006AAAA81FFAAAA",
		INIT_2B => x"FFFF0000FFFF00000000FC0500000000AA00002A0000A03C0000000000001500",
		INIT_2C => x"0000055400001405000001550000015000001554000055500000140500001554",
		INIT_2D => x"9249CCCC25550000CC6100068000AAAA55580000618633330002AAAA49339000",
		INIT_2E => x"0F0F0F0F0F0F0F0F0F0F00000000000000000000000000000000000000000000",
		INIT_2F => x"00000000000000000000000000000000F0F0F0F0F0F0F0F000000000F0F00000",
		INIT_30 => x"0F0F0F0FFFFF0F0F0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF0000000000000000",
		INIT_31 => x"FFFFFFFFFFFFFFFF0000000000000000FFFFF0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"FC00203F02FFC402F400AAAA2FFFAAAAF000FC00103E2FF0FFF0AAAA02FFAAAA",
		INIT_35 => x"00578035C0150000000000000AAA0AFF550000007FF0001000FF40075502F4A0",
		INIT_36 => x"020E3F030001F028FF01AAAAFFFFAAAAFFE003FF007FFFE0F001AAAAFFFFAAAA",
		INIT_37 => x"FC121CE6CB40F7BD6305033157AAE10B0C50000000007FF0000517FF2BFFFFE8",
		INIT_38 => x"FFFF0007FFFFFFFFFFE0AAAA0000AAAAA800FFFF0000FFFF7FFFAAAAFFFFAAAA",
		INIT_39 => x"0100FFF400000550FFFF0000FFFF005503FF0000CFFF0000FA15FFFF4855FFFF",
		INIT_3A => x"0000FFA800550000FFFFAAAAFFFFAAAAFFFF0000FFC30003FFFFAAAAA803AB50",
		INIT_3B => x"FDFF0000F80100005553FFFFFFC5FFFFFFFF0000FFC300035555FFFF3FC3FFC3",
		INIT_3C => x"0000002A00180A0200030000869200000000AD00000000000AD0000000000000",
		INIT_3D => x"00000000003001E00000000000000000008002C0000000000040000000000000",
		INIT_3E => x"0010004004000010004200000100000002001080000080408000000011000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
