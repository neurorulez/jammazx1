-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D352A0B57FEA2A4977BB18080082410493A17FFFFFCF408389FEA7A3D3F3EAB5";
    attribute INIT_01 of inst : label is "208B53050688596AA08094500A24F28449614EA8FBC4F2612971B05C07AC02D0";
    attribute INIT_02 of inst : label is "FC616582249E4F061E45A982F7BBCB31445F77C419F84F77D72089804FBC4109";
    attribute INIT_03 of inst : label is "89BE341034499CAFCD9900410F7AFFA7DC55555E004169FDC262E38A88145499";
    attribute INIT_04 of inst : label is "51A089270943A937ABA93780076A8522A211668422D64C1728AB834409386F50";
    attribute INIT_05 of inst : label is "F34F2110D2108910805499B883E2D415122286315425C47E8BC40155075D544E";
    attribute INIT_06 of inst : label is "4250545C518B4A32A60292DDFF9EDFA597F9AC96C9BD51493C0A4F0060B24174";
    attribute INIT_07 of inst : label is "829D5134F22CF4224501505499A48FD17E8F9C5A14936A1964B02AA294A2545C";
    attribute INIT_08 of inst : label is "830615531605408A9A97523A1128A7118145084A0E87140824D26D52CB94E216";
    attribute INIT_09 of inst : label is "54CA121CA721674943381D902702F8AD58C58A4236918946074DE28A00013802";
    attribute INIT_0A of inst : label is "ACBBF6EDA9D7DA3F7015FCD31CB1CFBB6A38922B18201AA08422A43896244542";
    attribute INIT_0B of inst : label is "68CF672559C9A3322214A2AD08D47BE33410CF0324290E1D3E24543A90024B93";
    attribute INIT_0C of inst : label is "47AD5FA461F7309C57CBCF2C8700FB027D0826FA40DF4201AF3CAC83D9C9D672";
    attribute INIT_0D of inst : label is "D3C00083105B997A27D13197E27D1310DD4BC23475AD632AB2B16B4FE4D7C941";
    attribute INIT_0E of inst : label is "8D1E02012248B31CD4451055AB35BA8DE47A949DA2A5540509DBECA80000CBEF";
    attribute INIT_0F of inst : label is "8E768A955138B13B60BEE6310AAB24C678060B64F974BFA4538B0FE8690B7AB0";
    attribute INIT_10 of inst : label is "9151B89941926A66A948F3DB6F1BEAAB25E89F31AAAC97E27CC43752DF69452B";
    attribute INIT_11 of inst : label is "3C6ED10BDC99F6BF6234BAEDC4F5F02D4D368DC6FAF1F2EA72C4358AE44FAE82";
    attribute INIT_12 of inst : label is "88A1244A20890402A8F7389A218CE801380DB474542106A1EEF1346189D2E623";
    attribute INIT_13 of inst : label is "41D6193070CF2CCB571C7CE4CA58B91C696BC8BFA0C1028A5488B55488163416";
    attribute INIT_14 of inst : label is "2A44048F49C04A094EEC8C871E72E4247A4CEEC649D496F442C9C6982A908A8D";
    attribute INIT_15 of inst : label is "145FFFFD54E4164C4244C5C442B13686B1942E85391133788DE6B805211A1231";
    attribute INIT_16 of inst : label is "FB26114604623029EAC6BAA5A2AA0B34686E83545483427964C34290111791C9";
    attribute INIT_17 of inst : label is "2A88551C7AA801570B00337378DF741A66D0AF7DBC646754A7661364651397DD";
    attribute INIT_18 of inst : label is "006845ADA168B448DC8AA48A4CCE8D70C5F2D812B88F7399A39CD38191D29609";
    attribute INIT_19 of inst : label is "22E7BFF822726DCCCE49B8C34294A3110D7DC0BC7E82692858267E886AC18A31";
    attribute INIT_1A of inst : label is "D51100284406842221250C068413619260C34CC01030D25967F30100000C02B0";
    attribute INIT_1B of inst : label is "9232032823232520204400104A798668B10FC11028CBAFEA0114670029ED2FE3";
    attribute INIT_1C of inst : label is "10A78EF5A24BC6E930D0D10402032C320EC4A2C458A8D5402EC19E9410080166";
    attribute INIT_1D of inst : label is "000000009C4060000B640080036401F003654204404AD120482E819CA729C842";
    attribute INIT_1E of inst : label is "4A5569652AAAACD345656565655559EA9EAD555575DD9E6EEBAAAEBB9B6775D5";
    attribute INIT_1F of inst : label is "0000000000000000000000000000958AC0D05A0B42680632A8755570AA74D6A1";
    attribute INIT_20 of inst : label is "7BF7A77B4826D648F836A54A89FFC719E08ED57CFD7CCAD63CABA0288D3AA281";
    attribute INIT_21 of inst : label is "A79D13B846540BEF34B279FD3EE806F3CFBE87E687CB7FC25F7BEBD43C25B01E";
    attribute INIT_22 of inst : label is "A9BA10480000BA7868A8F51DAB51EC9705ACFC5BE7E5F11A0C6537A49134B2CC";
    attribute INIT_23 of inst : label is "6A66D00456D515F731C70C385214CD4F11115FBBE8BA4E33CFA27551897431BA";
    attribute INIT_24 of inst : label is "E402467A0483107A24F19EA8A0800D040468000340011DAD15FB5997FE934AEF";
    attribute INIT_25 of inst : label is "0000000000000000000F266D02F9DAE7A7F0CB54D07B7C3E07C00951A8BE3E20";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A480EAC280DD640080263924B2C96C90016CC01FFF1B9533B9FBCD6603E36BD3";
    attribute INIT_01 of inst : label is "6400615610D5FA3944364C9B2D5143EAAE9FE14B6415A52B5A83597D393D67CB";
    attribute INIT_02 of inst : label is "4D17E8104A28E0228F0030ABDF2D9E420C065B0CCA63065B2F8402F90622A5BC";
    attribute INIT_03 of inst : label is "B2405B74058EE5E27ABFA001216C64CDF89FC6B81224A3F348000735662AF04E";
    attribute INIT_04 of inst : label is "862D9050B4EE2C0110AC013DB6644885AC7A8B16E01A855B41300868DB9A0050";
    attribute INIT_05 of inst : label is "27164A2D02D76622DDF04E00E8001D59845DF2BCF268AA84B405455500E38A46";
    attribute INIT_06 of inst : label is "D59785D26A004788D4B549A0406D14806DB6CA05D51B2A1C599832ED0607840D";
    attribute INIT_07 of inst : label is "BCF36A71645925D189B25DF04E05549680E63A814A0907F80E06E52FFD2C85D2";
    attribute INIT_08 of inst : label is "B7297DE5E74BA7BBC1983362683C97B8AB2146E1C8F734BB0E012039C02796AC";
    attribute INIT_09 of inst : label is "AA92C6EB2C7E0B90F0D2B6E47AD45F5AA8A07BF426FD0DB5EC1FEBF9E9EB8164";
    attribute INIT_0A of inst : label is "D948000005ECA27259523D6D2B5560002F855FA723523B26B6B542C70F12AA86";
    attribute INIT_0B of inst : label is "1C2000008000F08A5527DEBEE4E9409886B5DF47FBF7D1B07E47F3EA5ECEE70B";
    attribute INIT_0C of inst : label is "17EEF0794690444098B256773A112C941679422CAF459EF34959DB1A00002000";
    attribute INIT_0D of inst : label is "84996585F2E864004117AA4004117AA39BBC78A156108E8C54D75E9F0D393585";
    attribute INIT_0E of inst : label is "2855FB72BD21258D5B6DA2E28C92215A47EC7A444B77868E3D24A56D9965A2DA";
    attribute INIT_0F of inst : label is "31912DDE1B09C7A481CA18C2EC45520A80A85D1000A97F8BC65C9001C489935E";
    attribute INIT_10 of inst : label is "462244E02A45FC00C9A167F3F7684C455001042A3115400410AAE6EF71C4BCF4";
    attribute INIT_11 of inst : label is "5EF503E07D70200425F92D0509C4427116CAD13FFF647704099B421C1080F3E7";
    attribute INIT_12 of inst : label is "550B9EAF5FD4EB997290CC434529F77F89369188BA527B55219886B6C048305F";
    attribute INIT_13 of inst : label is "B2AC69AECB147DDCBC8290755EE52D8281D401E4B99DB6D3B17E469AB6E9C7A9";
    attribute INIT_14 of inst : label is "8F682FE28403D41A999B312A5100817F1C21991890093200DC5A1F52DB5AD542";
    attribute INIT_15 of inst : label is "DE82AA71AAB6B2F3BDFA521BBFFEFE3F189A90B7ADAAA13D585AD377B5AC9E94";
    attribute INIT_16 of inst : label is "C47E2AACC231C1DA4B0ED2CCBCDB5EFBDB94F53D59F8FF932F387B5B78EE939A";
    attribute INIT_17 of inst : label is "46127DE6B54B02F2111622CF3A39DC6F9927B114471B108ADBD9A78897672504";
    attribute INIT_18 of inst : label is "220C8C9495CEF7295C3CF3CCC919B9CC5A0524A48C359E64ECE36A5ED636329E";
    attribute INIT_19 of inst : label is "D0C3BFF3FD0CB26221B2CC186ADBCE6CB1F2CD86E143A20CE234E14E840D83BB";
    attribute INIT_1A of inst : label is "0DE315720857211C628E40572123098668D1EC45551F17EA8FE54AE4292845E7";
    attribute INIT_1B of inst : label is "006B2FBB044C04B6521E525B26FAA2E1AB444555118CFF3C233887A498B61A3E";
    attribute INIT_1C of inst : label is "7BD1B208FC9B8A1874345821EE4A5CA72BC944788F3929C9D2E583FF7F64B6E2";
    attribute INIT_1D of inst : label is "000000017901E7FC0181FF7E0381F80003802E56092E19EA7AB1C87BF7AD6DEF";
    attribute INIT_1E of inst : label is "6927D9BB89B337B6C9B9B9B9B55553553554CC00000000000000041111455555";
    attribute INIT_1F of inst : label is "000000000000000000000000000080C042B89702E25C000E1AB031B418B09B96";
    attribute INIT_20 of inst : label is "2E7FABFE6B29492BAA31158CB50011231AD81FB6081DCD2A8970964EDE2396BA";
    attribute INIT_21 of inst : label is "E8DF88B1E98E403D3FE8C4C8502AA11830012FD080030E85C72273FC807FC440";
    attribute INIT_22 of inst : label is "F3D81200000000162D751AB8104A093526333EF806221292E427080DB4010A12";
    attribute INIT_23 of inst : label is "B23F600E02BD03EF25C82A41712496C1D1404EEBF148C417FF16FDCCAE36FC9F";
    attribute INIT_24 of inst : label is "1AA958F849CCD9FD12C07FCEC0809E0000B0000782012E0408FC0D1D9621A1EF";
    attribute INIT_25 of inst : label is "00000000000000000002E08D6466008ABFF2DE20045D017E2819529B7DFE63B7";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B6D02A0085B16A09ECBA10000002090400A07FFFFF41052BA8F94D7719E90AA1";
    attribute INIT_01 of inst : label is "62680570D0025A10402486004930C06B44554158A6C4438230F5085D1E2F01C0";
    attribute INIT_02 of inst : label is "91016801061827128E3402B829D646800743AC87540D43AC870269BD41902128";
    attribute INIT_03 of inst : label is "8C6C1017A40B156051A2A0000834B00DB89D5408FBF683FA3A1A0004A7855407";
    attribute INIT_04 of inst : label is "81204C382523E90221E9020484400021A0518604BA0395C3444868000B1A2CAA";
    attribute INIT_05 of inst : label is "C10C3994C294A78090540703289A05400709E2F85028EBFA86C4195501249386";
    attribute INIT_06 of inst : label is "1314F514506867A0A701DBEFBFF6E97DB6C9759710820A00300A04081A813D10";
    attribute INIT_07 of inst : label is "A7945010C330C521E120505407057F50D8202A82D281C01D0270A9AB7BA8F514";
    attribute INIT_08 of inst : label is "550C050514382FF902D65AFA030801BD3A8BD6F1C4F5140AC810384AE83CA098";
    attribute INIT_09 of inst : label is "A05AA4A1AA4A87E4F14551FAE8E8522923A3A1534850D142881FE1DF51720047";
    attribute INIT_0A of inst : label is "6F61ADA8CDB7B21B716DB3B66D74E2A6CA105A03441218A2A42092824F00382F";
    attribute INIT_0B of inst : label is "544429178A45D11A09316113046D217A14047F6480200D207E52FE88DECC829B";
    attribute INIT_0C of inst : label is "17FEAAED2A52E408CCDB7B5DC9193FECDF7CCDBEBB37D719EDED6FC90A45E291";
    attribute INIT_0D of inst : label is "FED1458F02F6B33F66F7FF33F66E7FFB6EF70499377BED6766E6779F88BD85C0";
    attribute INIT_0E of inst : label is "264C91A320D9F5BFD15112F7E67371CB23B751B54584140BBFB6582891459F6E";
    attribute INIT_0F of inst : label is "5AD51610513967F6E3E59CF706F66DACFCBC56CCDF6F87FC315E9BBDA4C2DDE1";
    attribute INIT_10 of inst : label is "BBBB50B76F33DE7CE9D9BFFEFC3707F66CFD9BFF1FD9B3F66FFEDBBDE79CC0A3";
    attribute INIT_11 of inst : label is "E6D90AC27D117CEE6E2D52D90DA7C369FB6F5B97FFBF778666D4639E6ECCB2E7";
    attribute INIT_12 of inst : label is "A00A492FE125BC3B5A526C0A14A448A0098708CCC2FF6D84A4D81436D973A6E1";
    attribute INIT_13 of inst : label is "3714D214299F455EE28A00D5D2F7AB8A11E98560D3E1028014D2A402ACF42414";
    attribute INIT_14 of inst : label is "0840F946F88EBC9685FF99A9495147CA3FC45F4CD4CDF046B496369C0A108259";
    attribute INIT_15 of inst : label is "D1894F5B02A42491234EB54922B46EC5D551AAA42900A3C90D83F184210D1DAD";
    attribute INIT_16 of inst : label is "E238A4964B51AB520A56D2892A8290995154A3061E1043E24800429069A12A16";
    attribute INIT_17 of inst : label is "A31451403B0A048FAB22324B3A59C262504135D70110841296512A500542B7CD";
    attribute INIT_18 of inst : label is "FE040524A40E0708156AA2AC4808F58056011562C829064AAC324A86941454A6";
    attribute INIT_19 of inst : label is "94CF2AA2A123DB68645F6C11429A820C8472AD022071B8A47BB02066002551AF";
    attribute INIT_1A of inst : label is "C8106B76058F61820C6EC58F61190C873E711C02B70C168A4DF54B0F69A64CB2";
    attribute INIT_1B of inst : label is "8617A87A033300009002101242FBA140C74302B704E43F0C6112202008260105";
    attribute INIT_1C of inst : label is "3190A209559B86387D3C40002A475C7D1DC2645D8B980CC0FD338046120004E2";
    attribute INIT_1D of inst : label is "0000000002A1E7FC3E05FFFE3C05F9F03C044210084C80DA1284C018C42188C6";
    attribute INIT_1E of inst : label is "880639CB37BC3871C1C1C1C1CAAAA9E81E843C00000000000000041111455555";
    attribute INIT_1F of inst : label is "0000000000000000000000000000028140700E01C238013560A2C0A160A11C73";
    attribute INIT_20 of inst : label is "3EFFAAFE0A0B6D4AAB11A442A142D23AFA8C5D68433D382AA452047FDE3B8438";
    attribute INIT_21 of inst : label is "4104828920D1D42A0660C1F25A83E865C75C2FE4E902322D512053D4A875C650";
    attribute INIT_22 of inst : label is "53F4000000002A6E48D692AD22502DA536067FA83460E09288A30F0927152A86";
    attribute INIT_23 of inst : label is "603C40060A712C7421E49E24FE4845CD6AEFA44510408615A086F8142D168485";
    attribute INIT_24 of inst : label is "70A8507C50D1DA1A36C9AFF1800084000460002302000A1551B68ACC24CAB283";
    attribute INIT_25 of inst : label is "00000000000000000002639BEEEE5ABA3FE2DE74DC5D7D7E2B51A0D12CBE7510";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "924488E0854024AF3EF20822820820D4418C543FFF9B39A838FE64D6D8F889C1";
    attribute INIT_01 of inst : label is "28225067448048026804948001A280505444505B0FC20A0210940140252C200A";
    attribute INIT_02 of inst : label is "404920A0545101400211283320DE62041511BCD5084C11BCC10825A411512800";
    attribute INIT_03 of inst : label is "B0FE105308C95960C19284080331314484F5B8CEE9D241EE30A8A82601255529";
    attribute INIT_04 of inst : label is "014668A0042A6D0120ED01029F260441451D14202895419D0102A24020081C01";
    attribute INIT_05 of inst : label is "8828AD5686D201240055291B2088911D0241014040205000BFC4085F8430C282";
    attribute INIT_06 of inst : label is "1A1249E21AA2EB009C2FB6492492C92EB37DF6FA0811A820A12A10080C281042";
    attribute INIT_07 of inst : label is "92231A828BA2848848059855291A0017FC045A0852A4420C50542125482649E3";
    attribute INIT_08 of inst : label is "5F2295722A75221CAAD75ABEDF8E1C9E11EA0263A96E3DC9F454880A629118D0";
    attribute INIT_09 of inst : label is "28407241272CB76540C55D9AB06973AD3B49A87EF81D9866E60DF182713D5047";
    attribute INIT_0A of inst : label is "647BE4E0D7B3BEC93924D597846983827B1A53853498296C9DA63508D400546A";
    attribute INIT_0B of inst : label is "7046631618C5411EE1142631294E7BF014C64F3606216C583E2654D1219D56EF";
    attribute INIT_0C of inst : label is "17BBFAAE60E7B80E66595998F3EE9B564D2CE49A1993437C656665F398C58631";
    attribute INIT_0D of inst : label is "535544E62A331912226E13912227E130E4E7953A7D8E432322AFB1CF868C8451";
    attribute INIT_0E of inst : label is "4E9E95B10E4C913DA2093A31332D9ED77A131C998D9D94B370DECEC95954CDB7";
    attribute INIT_0F of inst : label is "8C66367652947E1BED6CC629223224C57E8E4664695CAB2499060CC861A2C8E5";
    attribute INIT_10 of inst : label is "991110B9B39A6627A54C980C5E932232244889938CC89122264E3939EBAB4A39";
    attribute INIT_11 of inst : label is "6098D580814B94B25245DB6D8DA1A340FDF53C9C099971E23246311624469A45";
    attribute INIT_12 of inst : label is "1005082C2504C4A41CE7300A718E48AD00DB004452C321B9CEE015F09B96CD24";
    attribute INIT_13 of inst : label is "26C4DF37208914CA0A8A84C4CA50AF9A90256AE055AF2ABC12C404E29164A9D0";
    attribute INIT_14 of inst : label is "5B4EA50658E84688242588831C70F5283AC6424449A590744EC89E74AAD3981C";
    attribute INIT_15 of inst : label is "8626D916D2B491552B58206D2880A75C4873029DAD34D985AA0991BDE5322C08";
    attribute INIT_16 of inst : label is "222A90C568C83A9819A7566424186A0D45413A162CD04A511440CA528F312148";
    attribute INIT_17 of inst : label is "3412DB3003090820B2566360810503644821D4D3118084E2549D685E1984DEF9";
    attribute INIT_18 of inst : label is "DE14C48C101E7129D00B30FC718812A826A1178B6074C60AA6304EF2D31038E2";
    attribute INIT_19 of inst : label is "C48FBFF0E77AD9806F7B30414A54E3099879A2890255F8F4D591024622528435";
    attribute INIT_1A of inst : label is "ACDA326828CA811B464D00CA8198144B0601D615A40C169385E308228CCDF6A3";
    attribute INIT_1B of inst : label is "2776AE6383FE400010129A800011020DB587952400D82F8A8A3023068D590307";
    attribute INIT_1C of inst : label is "10A61E1413086404A0205041220F8CF03C2A514B294D4A0D2632C8C690002092";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000010A9401145401003D6AB5ED7BD842";
    attribute INIT_1E of inst : label is "F77802003FBFC0082E0E0E0E000002002003FC00000000000000041111455555";
    attribute INIT_1F of inst : label is "00000000000000000000000000001A0D00300600C018050080E100E080E19FF7";
    attribute INIT_20 of inst : label is "2B67E4794124AD7352B1B9A91942D3B183B87182413D4022991A847B8C919210";
    attribute INIT_21 of inst : label is "51C22333885957F5831049C24CE029045145042F504404942A8F03D8C966A16A";
    attribute INIT_22 of inst : label is "998480000000CF4B915082193898E4AAAD2EFE982858BAC4EE12CDC4014D0C80";
    attribute INIT_23 of inst : label is "046C40046833106459828A147001044411044415584A05199F0214431ECE4E91";
    attribute INIT_24 of inst : label is "52A1CD7C1A997B13FD680FFD800004000020400100001AD08015980E6E40808B";
    attribute INIT_25 of inst : label is "0000000000000000000901F2F8E7129C85F989BE9F48675E88D5B0A3AABD0D52";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "2490381AA55504A6DB4A132CBA936DD8510E955FFF75B03838F96C444DED71EA";
    attribute INIT_01 of inst : label is "804813E09021701342125A2DA5451011414050412019146B5AA2452061B06419";
    attribute INIT_02 of inst : label is "690DC00908A28A0208A409F0080411811A40081AD40340080C404AAB4059AED8";
    attribute INIT_03 of inst : label is "1200D92480B10F2E44B6120001800F4C049190A31224D30E9A12001406876830";
    attribute INIT_04 of inst : label is "0385514594A4CE05004E0516910C4885061A28BB52074F82042A5811BD101644";
    attribute INIT_05 of inst : label is "14514AA5146206876968302F61D2070045058330724051011000183F81A68A84";
    attribute INIT_06 of inst : label is "9462B0C61848BC111B064DA69B4934906882412497C2241145B48C2812846D01";
    attribute INIT_07 of inst : label is "1507184515451885A2D609683028222203F101014B04093108E245442145A086";
    attribute INIT_08 of inst : label is "A4204A252058B5B0035E6B94C24D30082035103595E479B120208129886A34A3";
    attribute INIT_09 of inst : label is "019FC089F40891FF8707E41F403C8010AC80807E401B942C02981D0127600156";
    attribute INIT_0A of inst : label is "6D6FEDE5963734DB65ADF9938C608396D311534C625463CD18C45E217828A8B4";
    attribute INIT_0B of inst : label is "0055E72079C80154C53C655337CC2F0118A5509EA0CCD58860AA824D69EC026C";
    attribute INIT_0C of inst : label is "EC11050C305F50AAECFB9B59A167333CD9634DB2C53658766E6D6FA179C81E72";
    attribute INIT_0D of inst : label is "C7F7DEB623363376EFDA3B376EFDA3304CEA8C182B58C16EEE63F7D8D52E15FB";
    attribute INIT_0E of inst : label is "0608D5B384DBB125C20A2733E67934B79AB319B4A5A8E8A351D71A73FFDF9FFC";
    attribute INIT_0F of inst : label is "18D296A3A2746A3AD1F18C6B2E6EED9DD2AD56CDDB84D78CB552199823D6E083";
    attribute INIT_10 of inst : label is "BF77BF33AB34C6ED64DFB03C1A368F6EEDDBBF3339BBB76EFCEC13BAA69ACC33";
    attribute INIT_11 of inst : label is "67D9700101E83307966F7FFE898822627FB5398801B80986E7C3E376FDDCF35D";
    attribute INIT_12 of inst : label is "000818B467178CDD185FD0AC508547244FBB44CCCB4BA580BFA158B8904C3965";
    attribute INIT_13 of inst : label is "AF9BF260A99B76823092121B81114592146D396A55AA25112552888B1574E1A2";
    attribute INIT_14 of inst : label is "518B4015F2B40340956D99A108339A00A79556CCD78D95580340B8ED14631311";
    attribute INIT_15 of inst : label is "C601C0C18B18A400A53AB428A44300505523A318C6229F6C11A105A8C6254DAD";
    attribute INIT_16 of inst : label is "865B228973411C11114854494410408991D434528C806C1A40008C62EBA6E002";
    attribute INIT_17 of inst : label is "71539A2033111011BC64B28D0169126A59651104451BB5884E08A74A922669B6";
    attribute INIT_18 of inst : label is "22849924AD2E9153640E38D58311948066053606406016664CB32C72E2312CC2";
    attribute INIT_19 of inst : label is "4488000846FC49845FA930C58C50C42A948308028969C8A4AA908976002040A0";
    attribute INIT_1A of inst : label is "2E8BB1492EE49039770906C480BD8681A7408A759C8C16838E122B3EED8774CB";
    attribute INIT_1B of inst : label is "8560AE0B833A42DB501A5AEDB669833D3006751C9EFFC0F3022F6306D7B91AF7";
    attribute INIT_1C of inst : label is "F7DDFE5753982F0810300419A40C02C0B0094B686F01280D9A3947FED924B2D0";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000002C510144C6DDB70E6873DEE7BFDF";
    attribute INIT_1E of inst : label is "0040020B00400000000000000000000000000300000000000000041111455555";
    attribute INIT_1F of inst : label is "0000000000000000000000000000A8543EC7D8FB1E60048B120625051205E004";
    attribute INIT_20 of inst : label is "40C04400210DE021FF1410A4124480A085300182101ECAA2A052956EC1851330";
    attribute INIT_21 of inst : label is "59EE04D3828DC417D9040A0642720F0C30C3102655210094A0A4801BF30611F7";
    attribute INIT_22 of inst : label is "5BA400200041D59201328A8011096E2280CA8209227569484C5BAB6927048045";
    attribute INIT_23 of inst : label is "9051FB88A0C722E9056A7953CE6CFE80C0414111136F898A1A201516AFB3CB85";
    attribute INIT_24 of inst : label is "95A38B848F0A594324645F03F3819F9C0CFCC067E6033C4048D817119608212D";
    attribute INIT_25 of inst : label is "0000000000000000000726BB587A80E8D00501AB046381815A37B68273C08152";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B6D24C5A9B546640492911A69A4924DC0626FA5FFF41301818FE82666BAB618B";
    attribute INIT_01 of inst : label is "A4E92042F24B285145924E6DA5410144540144499021040EF2872D2320112509";
    attribute INIT_02 of inst : label is "012CA1172820802432F49021490490924F4A090F5CC54A090965EA254A0DA6D1";
    attribute INIT_03 of inst : label is "9900C93794AD0531245A00000126202025B894A9DBB6980ABA5A44944B933C08";
    attribute INIT_04 of inst : label is "3365104094A607409207489090856A9525CA081B7A4801090CA96925B068C144";
    attribute INIT_05 of inst : label is "041042210C424B936B3C0808B27A49889F2D0C412B614410900008AA80A68A8B";
    attribute INIT_06 of inst : label is "8402FCF7C969260633240492002492010482410414CAC050409E03293A943529";
    attribute INIT_07 of inst : label is "1752C94104410096E6D2CB3C08428012023348114B82837D282265C42144ECB6";
    attribute INIT_08 of inst : label is "ED6C4C252868A09611CE39B44A0C141D34AF0877A5683881F0B05229E9389420";
    attribute INIT_09 of inst : label is "0C68690E8690D244C0181092E3015118AB8D992ECA4FB32250C215423DBC2B57";
    attribute INIT_0A of inst : label is "4C41090196A7AC52572900248858060491614905225329471084F23BCC45FDEE";
    attribute INIT_0B of inst : label is "81D920484812076C452405102108080060A100D632ECD08100E22469001E082D";
    attribute INIT_0C of inst : label is "0150512808100132ECD35311A088301CD8494DB08D3612734D4C4D0048121204";
    attribute INIT_0D of inst : label is "90B7DC642FA4222444AA2222444BA22C28949D0A92509044445B5A803D001480";
    attribute INIT_0E of inst : label is "42A455926C9528A136DE3FA24458241A4A2149271511A0E2D10490F11554124A";
    attribute INIT_0F of inst : label is "109C544683AC5A20954908482444492882C9648892690020A444911204A48027";
    attribute INIT_10 of inst : label is "222211A2222404484C912014D2248544489112A2111122444A8B0A2524920E92";
    attribute INIT_11 of inst : label is "59D544182138242410432491A9296A4A4049510805290D0444A742744888515D";
    attribute INIT_12 of inst : label is "492820A4041480849010411050110C2DD82A00888A422110208220B85050A107";
    attribute INIT_13 of inst : label is "AA8D5612811240E6825A1B54E234CF5A1F46A3F155246E35350A90AA15726CA0";
    attribute INIT_14 of inst : label is "230A801E41280EA0D06D19A108141400F2090488942918950EE0D04CB8C23150";
    attribute INIT_15 of inst : label is "323FC7D11A30B619A76AF4C9A4C228495DE7A7118C26B8583B4555918C254EBD";
    attribute INIT_16 of inst : label is "0662A69D6ACA0A106168C84D8DB6C348D8D6940FAE492603619918C7440194A0";
    attribute INIT_17 of inst : label is "63728C636B2120C54078C24647368DE54925B28A22C994AA4C48A54A9AA52000";
    attribute INIT_18 of inst : label is "FE749DB6B9DEEB634E869044D9199DC5C6453526C48089266459285242292186";
    attribute INIT_19 of inst : label is "45092AA045001201A0024102084856AA96822A16816B8964BBF2816E44A4496F";
    attribute INIT_1A of inst : label is "0A0B6AE86D8E86216D5D0DAE86BBA5D366CB5CD6342C16822217C828C08264EA";
    attribute INIT_1B of inst : label is "9556E56922AB32DB564A7A6DB511056D558856B42120D096BAA08036DC204D34";
    attribute INIT_1C of inst : label is "0810C324A0C02D4522A2C934A6681281A129572AE5552AAD482B934ACBB69286";
    attribute INIT_1D of inst : label is "00000000000000000000000000000000000026724D5E8DF97E10E90042100001";
    attribute INIT_1E of inst : label is "0080040040000000100000000FFFF60060000000000000000000041111455555";
    attribute INIT_1F of inst : label is "000000000000000000000000000080403E07C0F81E0000000204040402070008";
    attribute INIT_20 of inst : label is "26886E84695B7129AADA158D955D0C44C039E8E9B4DCFFFD5EA7B57DC365B6A3";
    attribute INIT_21 of inst : label is "625438A50D0A5FE8A42A0C23E32A00C30C309C3FD51A674EFBD6900FF31251F4";
    attribute INIT_22 of inst : label is "A0EA00001201A526990A4A89924A082E0ABB821ECCA772125AAB3B2DB46D369F";
    attribute INIT_23 of inst : label is "00004380000100600100090040000C003EFBAEBEB378952E3AB70DDC2D133BDA";
    attribute INIT_24 of inst : label is "9CA90885DB5E5BC17FC00C018381841C0C20C06106030800003000000C000001";
    attribute INIT_25 of inst : label is "00000000000000000002299FEB466C1AA40F454A6D071300EFB792B63641DB73";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "002921387F4572996CB63C924924924448D23FDFFFCA00C0C9FF46E2C9B994B8";
    attribute INIT_01 of inst : label is "111481090924D10C31492124906180145111050CA24186210C194C818C419124";
    attribute INIT_02 of inst : label is "069344C48C30C18B6D0A408465B2D868B0A365F0AB5AA365F69013A2A322124C";
    attribute INIT_03 of inst : label is "C82736804A6F6434F2B2000003111804A6CF6B3700002116452530439048C44B";
    attribute INIT_04 of inst : label is "481198634210511040511046CF732650D0730C4905220426223484924DD58850";
    attribute INIT_05 of inst : label is "861863318129904924C44B98244524264090DA24D9041401C24002AA86186044";
    attribute INIT_06 of inst : label is "C62802082494A00D4890924B6C92DB6592C92D92CC900118636232840146028D";
    attribute INIT_07 of inst : label is "4028246186618A60124824C44B8280384E24304C2088E4928C19109084130208";
    attribute INIT_08 of inst : label is "A7972293871615B1CC638CD12171C629836530A3986782140E511C8494C14631";
    attribute INIT_09 of inst : label is "1AEAC718AC618BCC012002B204031CC61893C5C26D7098972D8A115E83639C8E";
    attribute INIT_0A of inst : label is "6D7124A18736311B616DA5B62D65928246DC2E729D0A94104A531044401A0220";
    attribute INIT_0B of inst : label is "4367210448410D91301930D1942F7920DA31D0CE49125CF420EABD18697DE34E";
    attribute INIT_0C of inst : label is "0040452F6EF3704E66DB1B589B11B29E595164B3AD9674766C6D6D9BC8411210";
    attribute INIT_0D of inst : label is "F2E3050797B3199232C2B399232C2B32CCC660F161CC4B22222373885D8DE054";
    attribute INIT_0E of inst : label is "3C5B01411248B499882087B12331B09362B2749C59CA1A1B1596CD86898D4B6C";
    attribute INIT_0F of inst : label is "8C716728681362B2E96CC621822224E459ECF6665BCDAD6617070CC97686D998";
    attribute INIT_10 of inst : label is "911141B9BB9677263448B41A9B12E3222648CB33888899232CCCB331924860E9";
    attribute INIT_11 of inst : label is "6558C330A06BBDF6C326B6DD8883E220DB6E5DA505BF2DE332D8313724678E0D";
    attribute INIT_12 of inst : label is "04078E1531C2A6515EF3306D2FEDD0B2493340446153A9CDE660DA6A4BF3E431";
    attribute INIT_13 of inst : label is "02E053B8E08B0DF7056836559FB818683073E0748132914C89C14A6140690231";
    attribute INIT_14 of inst : label is "94A61C36DEE3CA199C6D889BDC9070E1B6F5C6C44C859A70CA198B2745294C4E";
    attribute INIT_15 of inst : label is "08603FE5616A09E618910B46190C49657208584A5A985988C05A41CA52922C42";
    attribute INIT_16 of inst : label is "798E18606008C80894A1752250413C66060D46240D20D0C09E60A529041B8318";
    attribute INIT_17 of inst : label is "843C329C2DD440F87F80FB3A87D0F0F8B6D8DCF3DCB66B6331B718B66898B6CB";
    attribute INIT_18 of inst : label is "030662C6C6072394C6114B8306E6B2B84BB8C1B9783F72D99786C58BA9CCC317";
    attribute INIT_19 of inst : label is "502695533332DB83665B704DA52BB180CA08C1CCC607B4160418C61F3057A530";
    attribute INIT_1A of inst : label is "83690C192435908520A32415908984C122486A50D08C169A4407EE9425EE2302";
    attribute INIT_1B of inst : label is "4319119C8445464909A10924926CD0AC9803D0D0800590E6299004F245291061";
    attribute INIT_1C of inst : label is "6334AF7D5088E30C1212248211E352358D2605C0B81CC0E42C854E2134924871";
    attribute INIT_1D of inst : label is "00000000000000000000000000000000000191093C856401004B64635AD6B5AC";
    attribute INIT_1E of inst : label is "00000000400000001000000000000FFFFFF80000000000000000041111455555";
    attribute INIT_1F of inst : label is "00000000000000000000000000007FBFC1F83F07E1FFFFFFFDFBFBFBFDFA0000";
    attribute INIT_20 of inst : label is "24A87EC794E04D94A879CA104D724633E14A0F12C97CE222BC50C8EA8B31CA04";
    attribute INIT_21 of inst : label is "6D44438212E0A42A800449CE8E24031861C768002AF58E81A7A3D035F01D70FD";
    attribute INIT_22 of inst : label is "D164002012488D0C0425307A4CA4AD02038EC21D226CC42501036E2403824124";
    attribute INIT_23 of inst : label is "FFFFBC7FFFFCFFDFFCFFE6FF3FFFFBFF805405401C38459C35CAAE64551A89D5";
    attribute INIT_24 of inst : label is "C67CA700E4633C3C023FF8FF7C7E7BE3F3DF3F9EF9FCF7FFFFCFFFFFFBFFFFFE";
    attribute INIT_25 of inst : label is "0000000000000000000E62492CE992248A07971A181706207AC14C09E700EE38";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "802020307F04629B64B028000000000D00E07FFFFFCA908709FE0391C8F89091";
    attribute INIT_01 of inst : label is "2010010100001C08200004000061801051540558A64186000035080104010100";
    attribute INIT_02 of inst : label is "0C0070800C30C3020A88008024B6580004816CC4A84A816CC540134081680008";
    attribute INIT_03 of inst : label is "8A6692100C626032962000000335344322882C1E000000044424200204001C09";
    attribute INIT_04 of inst : label is "2021986100024308004308068A22044060430C00240204078010800109181A00";
    attribute INIT_05 of inst : label is "8618633180200400001C0958000404040000822010301014864000AA851440C6";
    attribute INIT_06 of inst : label is "C62104144090A6010B01B64B64B2DB25B2496CB24C904018600E02100106820D";
    attribute INIT_07 of inst : label is "08344061866188010000401C09420290CE2518080180500A0C30208084020414";
    attribute INIT_08 of inst : label is "02460612021415208A1142C003208260816001830842003004700A005081A631";
    attribute INIT_09 of inst : label is "086883088820988CC10016226001488C18010504254109020482015301411A8C";
    attribute INIT_0A of inst : label is "253924A0841210093144949225218A8240182820140B000008423228CC086C66";
    attribute INIT_0B of inst : label is "4057210448410150201D61DB14A679601831904420A8185001CAA61869694348";
    attribute INIT_0C of inst : label is "510104266CF3702E66498948B39996BE4BD36497A592D4F3262524B3C8411210";
    attribute INIT_0D of inst : label is "56410512029319923242999923242990C642403071CC4322222221004984A055";
    attribute INIT_0E of inst : label is "0C1E01012248969090400291233391B92296449C5C88380914B24CA2AB8D4926";
    attribute INIT_0F of inst : label is "8C717220E01122964124C623022224C458A452664964AA2C16020CC8769248B0";
    attribute INIT_10 of inst : label is "91110199B996132638489C08891263222648C9198888992324643190B2C8C489";
    attribute INIT_11 of inst : label is "2308C100A27195B2C60E924C1C45071109244CC1049584E33250311324668A04";
    attribute INIT_12 of inst : label is "000504156082AC514CF3702C29CDA1A0493900444159AC89E660584B4992C460";
    attribute INIT_13 of inst : label is "03446110C08919140C78163108A008781123E132014203081981084100400430";
    attribute INIT_14 of inst : label is "108634148AE14208182488939C90F1A0A45582444C8C9970420818290C21084C";
    attribute INIT_15 of inst : label is "10200004412809440001084400014981820040084A1069808840710842122842";
    attribute INIT_16 of inst : label is "28AE10446000C90010819422408228244401860008000240944084214511810C";
    attribute INIT_17 of inst : label is "861402150C5000FE7FFF036A865490C99248E4515412294210D508942008924B";
    attribute INIT_18 of inst : label is "200456A62504A252C0018A014AAA232818A848A9AA155248B692448AA1444214";
    attribute INIT_19 of inst : label is "58C4D55E0332498066493045842A230088084088C20510140620C2142056851A";
    attribute INIT_1A of inst : label is "81610C500431000C218A04310008040302012440400C1694021C7B14274E2222";
    attribute INIT_1B of inst : label is "0219219004454400058000000378C0E00B01C04000209024300004A00D090020";
    attribute INIT_1C of inst : label is "21342F750087420830104000034350350D020640C81041806C848A0000000043";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000010200288944010009802908421084";
    attribute INIT_1E of inst : label is "0000000040000000100000000000000000000000000000000000041111455555";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000020000";
    attribute INIT_20 of inst : label is "1588188558A0051800388D088CB2461161040836C97D2A281C0028C883122202";
    attribute INIT_21 of inst : label is "414027830A41D0028224339A1E200130C34D6BC080561E08CF039C04B110785C";
    attribute INIT_22 of inst : label is "8070000080009D18081010550AC2A7440384401C256CD21600A36E2400412294";
    attribute INIT_23 of inst : label is "0000B800000200000200100080000800550005554A18020E25A0C954150A89D0";
    attribute INIT_24 of inst : label is "C6788400D0533A70008003FC70000B80005C0002E00010000000001000000000";
    attribute INIT_25 of inst : label is "0000000000000000000C42402DE9B6258C06153A30070C00624104118480C410";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
