-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "C4D89B0DC30004D5135E810F42A001E01B223FFFFFFFCD2309F3A6F2D9FEC850";
    attribute INIT_01 of inst : label is "464CCDC3364B0E2C92AA34080ED98A4A3D55555D1D3657B6D9847331BB3A8B3C";
    attribute INIT_02 of inst : label is "79825310B88125F64043895275512F49D1459ABC5FC2A24DF12CCD719966EB99";
    attribute INIT_03 of inst : label is "9F865474D5AAF37B51FF677741683865B7FDC966504F0D6F180C527EB542C48A";
    attribute INIT_04 of inst : label is "966AD942C893EB79D30B768FB3A37EC96FBD97B996612573AABE65C30026CA4B";
    attribute INIT_05 of inst : label is "0A8B82BD92524D901DFA6A2CA2CBFED77D12D51646A2C8F5BAA592896A4F2D7A";
    attribute INIT_06 of inst : label is "A5D0934D24DA0000001F7C2A49A6926D0FAB25366652922EFF64C93A09A19D24";
    attribute INIT_07 of inst : label is "D94FDA9556EA2E6AC180584CC09999981352A94B356CAC95D75BAA592B2D749D";
    attribute INIT_08 of inst : label is "33170CE5CEC2E8F3146DCE4588745AC2E07598138B7599BD4B38611254DCCA6C";
    attribute INIT_09 of inst : label is "7D7DDC41688022C914EED0670EFAA75BDC669D3F3DA3B4668415ABDDCF7DEE67";
    attribute INIT_0A of inst : label is "4B85CA915C514DDB6CEA8B4FE4185D6666227432DA5BDC5B09D2E9162B1582C5";
    attribute INIT_0B of inst : label is "B9307357DF74EDFF8DF9AA7A64B8B2FFDED197FEF6D7DC37B9B63E60A44F8427";
    attribute INIT_0C of inst : label is "738F1BE5C65083D980B2D9CAE548041D28CE467CD3F9B6D6BE1E3BB00BF3BEE5";
    attribute INIT_0D of inst : label is "EB09BC9F5CECB6CF139A58481A0681A04812068007E741312B9C7B4EAA763A77";
    attribute INIT_0E of inst : label is "6955ED5803FBBDEF3B7FDB045FE9FECDBB198784F98D123448D123111B9D6E5B";
    attribute INIT_0F of inst : label is "6E34583C2BF21A000AD2F9B5A91F1D04040100545AC00020801813C001C557C1";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC25C45A938C55214C8E5";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "24A49248F2F869E6DF1BCD3ED19A7DA797FDA7E92524949247776A20CA6C8ACC";
    attribute INIT_19 of inst : label is "B56999EE5D254539317D965E1F69F7BCDA9A79A796F34A6DF5BEDBC32CA95249";
    attribute INIT_1A of inst : label is "96722EA9B12A75C416BAA5EA66435523329D1292999BB3B721593B8924DCA985";
    attribute INIT_1B of inst : label is "FFE60DCE2854D58E609D2A3CC1629729E8BAA66AB31263391588731B952AF319";
    attribute INIT_1C of inst : label is "5BCACF2FD00DDB8D12110B742ABA1311EF5E585227BDB366619CCF3199986716";
    attribute INIT_1D of inst : label is "4E8C298A5DA6BB5BD0F1BF9747200D4E639665545F98C553C414009895C3FD27";
    attribute INIT_1E of inst : label is "A13469EE0D3FB3EAE07FA6B47D4F4D36535D161A9895A5574F96454DD6DC0800";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00044422200013A329ACAA8AA7BF3178";
    attribute INIT_20 of inst : label is "FBFC8533328F7580FBA777A82338CF7273F753EFAEC8517FEA9358466F79842C";
    attribute INIT_21 of inst : label is "DF7FD0A6DF5DD0A2DF7FD0A6DF5DD0A2DF1FE6B6FAEC8516FBFC8536FAEC8516";
    attribute INIT_22 of inst : label is "05FB2B3B2B3B2BBBAB3B2BBB2FFC55555513593E454D0EFE3EDA10D2DF5DD0A2";
    attribute INIT_23 of inst : label is "A4E4A626A4E4A6E4A4955FFFFEED74F9958D110085F08F847C298683E16E31E1";
    attribute INIT_24 of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAA0AAAA0000038570888250582208410F00224A4E4";
    attribute INIT_25 of inst : label is "BB3BDF9FAECEF7E7DBB3BDF9FAECEF7E7EBB3BCEEEEED72AAAAAAAFAAAAAAAAA";
    attribute INIT_26 of inst : label is "095D26E45B0D6CB108BE006250042122F80921880554909B916C35B2ECEF7E7E";
    attribute INIT_27 of inst : label is "286190DB21212C22310890445EB25711DCD2B734BC462F8038B50118BE024863";
    attribute INIT_28 of inst : label is "285BBBBBBBBB92BFEF053EB3D58E7617A6924D99C893385C9A6ECF16DB2A2D68";
    attribute INIT_29 of inst : label is "6199B3C39AC922DB248B6CBD965116AD44D3E7132DD844B76112DD854356112D";
    attribute INIT_2A of inst : label is "C667EED329249092576492425242537B6D2E8393364DE624D30C66CF0C7B3678";
    attribute INIT_2B of inst : label is "14BB94046A12AC0EB1140A02303AC288DD619448908A8989B12FA9AC92445893";
    attribute INIT_2C of inst : label is "0028052AC2000B391DCA20A914525512016159C3201080400280422C202B8B8B";
    attribute INIT_2D of inst : label is "901010360404000101012040400010ECAD451522925512A5614005D95A030804";
    attribute INIT_2E of inst : label is "D4288AE9259E8B10483A6204557492CE4188251D350A22BA4967A2C4120EA282";
    attribute INIT_2F of inst : label is "F83E4029D33987BE9747CD9350A22BA496722C4120E9881155D24B3D06209474";
    attribute INIT_30 of inst : label is "53B8BA3F154F00000231B1384485E415F86A5281452883024A2E7F300C49EA91";
    attribute INIT_31 of inst : label is "F55B1EAEAD8EB63C6218C426CF66177CBD4E39EE471238BABA3C7154EE2E8FC5";
    attribute INIT_32 of inst : label is "402773ACD78CB9C2ABA76FB8CA921919490D242002000D4D9ECC2E615593B7DC";
    attribute INIT_33 of inst : label is "4234F2CBE4D53294FB3D49714C82080092002010480082092000010492492400";
    attribute INIT_34 of inst : label is "2C8B55655A8B22955956A2D405015B77466AD4A0A10A0A19A432CF9DA340A1AA";
    attribute INIT_35 of inst : label is "955946A2D405435A76964954A2C8B55655A8B22955956A2F50D435376974954A";
    attribute INIT_36 of inst : label is "CCD412C92994590EAACA7516432AB29D45890240B76974944A2C8355651A8B20";
    attribute INIT_37 of inst : label is "46639614C66A2ACCD5C36891BBBCBEB267240020056CDC3D37F67FCE2F30368C";
    attribute INIT_38 of inst : label is "D27A69A274D3443371F4C3323879576E5037FCE06D1EFF32E002009E14423C28";
    attribute INIT_39 of inst : label is "FFFFB4BA1D2E87107739DBB18146697422F0421D020219CE65D7BEDF11DF273D";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFE31E77899D5292FAD4D9996A334782022F45BC04A3300A86E786115";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "FA9752E1A7CA4C5E3178479FDCB633F4D286403FFFFF849340E22B1A1FFF4129";
    attribute INIT_01 of inst : label is "C2ADF07176DEADCA2DF356D6F5BBE3E3F6FBBF3D38293F7DE17FFC7FA1ECFFF3";
    attribute INIT_02 of inst : label is "B4BBA3363F3000600926E2C5EAC099B7AB0363C0A00CF8008469235C23491AD2";
    attribute INIT_03 of inst : label is "ECE38A3FB38797FEBC202AD2B76B3DFD3FFBE733E1FDBBDD755680357879CD40";
    attribute INIT_04 of inst : label is "44009411B5E8BEC6ADC2EDA38BE9127B762FFBEF6E3A4E9C6DD239AFF884072F";
    attribute INIT_05 of inst : label is "BFFF7D7EFFBEDFF93D9FF8400000406DA409AC0DAD81B5F120D10804D7A2FBBB";
    attribute INIT_06 of inst : label is "F9378E38F3C76BDAF6AE5DEF041049205002002011C226AF462BB691A51B0B6A";
    attribute INIT_07 of inst : label is "4E0A475AED508D4E1B41F4A0FC01441A84AFB5A2004A0A0104120D108288404A";
    attribute INIT_08 of inst : label is "7E894D491EEBD96A7D21F3F5E968B75104FBDFDFE12F4F6BA60E387E4C0E0040";
    attribute INIT_09 of inst : label is "CAC5AEA4DAD91EB5EB15ADC2AD5D06EA0A7F9BEE5FD09A972BDCAF0BFFE5857E";
    attribute INIT_0A of inst : label is "02A15BC9280051A931E0BC93E93E0B2C0FB0B91346EA0B43CAFC9B0F0783C9E4";
    attribute INIT_0B of inst : label is "64006A3CF90574FF6EF537AC002A36F0FA0CB2A7D233A5997BFD03F97700ED01";
    attribute INIT_0C of inst : label is "EAE3A8AE510EDD16EFDFDF19CC3F2F7BFED6A03915F0F14F98CAA96D0B3A95DB";
    attribute INIT_0D of inst : label is "5121186878D77FE60192521085210852308D2355502FD5559DC58ED8F0AAA9C3";
    attribute INIT_0E of inst : label is "538446502B5EE30053D034B088740096FFC613610C4081122408110506BF0CCF";
    attribute INIT_0F of inst : label is "F658011458642A024B69F0C4EC5E1955555555154C154887003B84E000919AA8";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC49F217340CCF1249000";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "9676CB2F863EE7CF38E3BE71CE5DE39F20E7882C96B2CE59782802289CE92E1F";
    attribute INIT_19 of inst : label is "40A917CB680ECC12BCC633EFB8E3DE31CE5CE39F3ACF3C778E3BEF3C618DCB2C";
    attribute INIT_1A of inst : label is "4A471E4AA2345920243EC55805A1A611155F25AB0888A3F803441801084489EA";
    attribute INIT_1B of inst : label is "FFEA044F94184296A1964CFD43780133C4792A5E50A2A140185CB5089AC17508";
    attribute INIT_1C of inst : label is "7C9492536ECA64922922269A71025C6644A8F31C400804C0004A0017C00012DF";
    attribute INIT_1D of inst : label is "152B4E3001040392209D5B21A5C45272D34A998A9131862B28A04CBF2707B1C9";
    attribute INIT_1E of inst : label is "397AA3B8D67627E788F63AFB929C70200201282541294E207325AE734DB094AC";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF002BE69C52B2054A4E13310C56226BA2";
    attribute INIT_20 of inst : label is "44001FE0229C45A461B277BE046603FB01257C044003FC800000E288E54FE149";
    attribute INIT_21 of inst : label is "488003FC488007F848A203F848A207FC48A0101244003FC245101FC245103FE2";
    attribute INIT_22 of inst : label is "D76DD5C5C5D5D5EDC55555C545B7FFFFFFACE67EBBE92D2A2BCD562048A207FC";
    attribute INIT_23 of inst : label is "07474767054547050DB00AAAABE391FAAFE92A92CB6ACB565ABBBFA6D5FFFF73";
    attribute INIT_24 of inst : label is "CCCCCCCCCCCCCCCCCCCCCCCC0CCCC444445562AE14B73CA452CCF7B96B674707";
    attribute INIT_25 of inst : label is "7400A8025C010A803F400A80254010E8005400A505053B43CCCCCCFCCCCCCCCC";
    attribute INIT_26 of inst : label is "DFFBBC8ABFAFFD723CFE8AE5FD48F5F3FA2279156FFEFAF22AFABF75C010A800";
    attribute INIT_27 of inst : label is "DE7CFC5496F2E8CF6CC3F9EE31A4A65343BD70AD548D3FA2A96FD234FE889E45";
    attribute INIT_28 of inst : label is "CDB0505050505025033B95C5772B5B845B3E96FFFA40EE17AD97FEC008E77C9F";
    attribute INIT_29 of inst : label is "C82000EE525FFBAE4B66914229E6EC539B295C6FCAE5FB9FD7FCEE5B3BBD5FE3";
    attribute INIT_2A of inst : label is "E26AC903CCB2CECB371ACB3B3B2B2FB327C9BF92AC3ADD1061AB8003B904001D";
    attribute INIT_2B of inst : label is "6FE57FFDAFED9C95B23FBDB67256CBD9AB6504851ADB9696ACCB1AAF2BCB567F";
    attribute INIT_2C of inst : label is "FBEF7297D3C92D7BB13D53569A2FB6A9CFE9ABF6F54D5A6DF6D539FD34BB9F9B";
    attribute INIT_2D of inst : label is "B5ADADFF6B6B7FDADADED6B6B7B5A97DD3EE7BF3FDF7B94BE9E496FBA7DCF7E7";
    attribute INIT_2E of inst : label is "2B52565309304CB76D1495A93B298499265BB78A4EDC9D94C24C912DDBC5A5BB";
    attribute INIT_2F of inst : label is "6593D984B7FDE103E4D08124EDC9D94C24C112DDBC5276E4ACA61260896EDA29";
    attribute INIT_30 of inst : label is "BE2447808AF8D2B7BC484E80917B0A9A21142AA5ACCD56D5B7F8FF17A0008EFB";
    attribute INIT_31 of inst : label is "5A24EBDB127449D695A569C0370A2BC11599207F623313244783C8AF8911E022";
    attribute INIT_32 of inst : label is "6827D6027AB21703305809FF946DF3F236F8DBF5EF7B53906E145701986C04FF";
    attribute INIT_33 of inst : label is "4B40489203679DFA860BF495E74928B61024B05B09125A2D80892D16C04DB289";
    attribute INIT_34 of inst : label is "E4F21B2690D934C7C9E63E1AD39DA5E9DB353BFEFEBDAF507BE25900159B553D";
    attribute INIT_35 of inst : label is "C7C9F63E3BDB9DA4E9A4D9E43E4F21B2690D934C7C9E63E1AD39DA5EBE4D9E43";
    attribute INIT_36 of inst : label is "9134B49B3E87C9F4364DA1B26D8F93EC7C57BFBD4EBE4D9F43E4FA1B26D0D936";
    attribute INIT_37 of inst : label is "3438FC6283C517DD5E7695BC025BC924014A2264B7291273A92CBFC052157D85";
    attribute INIT_38 of inst : label is "220D96EF9B2DCBFC8B4D32F0F287A58929FBFC2AFB01FF069154AA13A3F6E0C5";
    attribute INIT_39 of inst : label is "FFFDFF26A7C9A92365B2F2552DB7BE4D454084334B6B7D95966F5F60456055B5";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFF7147523BE67B4FCE7080BEA7BEB57BB96D004E9620DD23FEBF0A93E";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "A29240694A9286DA5B6A9AEF9EE4DDFF52A23FFFFFFF89B840E92E1C55FE0018";
    attribute INIT_01 of inst : label is "214AE000242D4A66D2A0342D0A1BCC0C0A1C4607A90486929F4A0A281A0B0238";
    attribute INIT_02 of inst : label is "045C3549270A01E010424D1A1D524168754920B82147A26DAAA8115155408A8B";
    attribute INIT_03 of inst : label is "BD00042DB1E9616129A900502268A350D553524D1EAF818F01529130D018C05A";
    attribute INIT_04 of inst : label is "50A29454924BEC8D528D17EC3AAB4005C6B1441497D36A21DA375552052520DB";
    attribute INIT_05 of inst : label is "2B028247484100021F090A492403401A6D2415249624928528942892092F3202";
    attribute INIT_06 of inst : label is "D96E28A28A247398C72A551B555555514008490484FFA57C50025FF3D1BC5568";
    attribute INIT_07 of inst : label is "544800540CA2FFEC0200602A340405478048A928514A2225445289428A891114";
    attribute INIT_08 of inst : label is "6BA028491FBAF9FF59554FAD4A513E740842102AB212942B8100002BED1B2249";
    attribute INIT_09 of inst : label is "D309411B2B7D42590D2A4A214A29A5215552D4A535FA896A07108915E7902A51";
    attribute INIT_0A of inst : label is "82E90A75C9943B4205E8A1B3E92B94151F3091994EA1552A946CB62C562B158A";
    attribute INIT_0B of inst : label is "F2A7FA0D1E15F3F8AB0127AD00252808B9850545CC254510B4820371DE664A91";
    attribute INIT_0C of inst : label is "BAE2A57974063F5B1000D162E8711AD094820E8557F5EE4558EF83EFB92B7FEB";
    attribute INIT_0D of inst : label is "2D56107B6A82C2EAA8F7D210A4615A5610A46111112D24A9254707F0128383AB";
    attribute INIT_0E of inst : label is "7FC545A03382B9C73C283CE6952C7E17AAD93563FD44A902840A110044B554AD";
    attribute INIT_0F of inst : label is "14A801183B596894D322817C787E3A000000000052D54820802727000ED9FEEC";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA38D14E724E5FE4848DB";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "0090104BA404C75D35A218E38D54D74C61430A4820A402805A200AA014EBAC0A";
    attribute INIT_19 of inst : label is "D38C291264DC44C5B5EA212131C748ABA551C70D20A695431AA9A69441084200";
    attribute INIT_1A of inst : label is "981368869DB5345563683C91B195A6D7530463B37BA8A086AB28835FC95C4DA7";
    attribute INIT_1B of inst : label is "FF9A01C6B59BCE31A02A4D334069473521A21A39C511A0355A8D8D139A070D01";
    attribute INIT_1C of inst : label is "28D6FF79BC6F731B46335BDC599B9EFBF7ECFE5F66B6DAA334D54516A8CD350A";
    attribute INIT_1D of inst : label is "9FA9EF1AED25DBD723D9FDF2E76A7F7A8A0CDCDFD99AA37A7C0057FD3247A5E7";
    attribute INIT_1E of inst : label is "0F7BB3B6F674F7EF28F4BE50DF9C790012ED473731BDEB3379F6EB7ADB6B24A8";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF889106CE92E727EAEF1B9B86E4B33AE0";
    attribute INIT_20 of inst : label is "20474A82A20C5420228101870260051006BC41E20476A8001540A20060523948";
    attribute INIT_21 of inst : label is "8408C9508408ED50842ACD54842AC950842AAB2421566AA420476A8420474AA4";
    attribute INIT_22 of inst : label is "14904040405050D0D0C0C0C0C24900000010A07E83E94A015020F6508408E954";
    attribute INIT_23 of inst : label is "1151539353131313124FF555545289FA5FE944929282A41504A4496825224354";
    attribute INIT_24 of inst : label is "0FFFFFF0FF0000FFF00FF0F00F00F0505041502824A8CB6892A229AA8A911111";
    attribute INIT_25 of inst : label is "6550228A19550822B6154A08850542CA2145502FFAAF2B620F000FFFFFFF0000";
    attribute INIT_26 of inst : label is "B8F8A6CC0B2FEDC450BE8A899C514542FA231D1CF3E2A29B302CBFB785428A21";
    attribute INIT_27 of inst : label is "05514AC008242ECAA212D154F82034158E3163CC51142FA2A2679450BE88C747";
    attribute INIT_28 of inst : label is "7081144114411480520EC14111485006020BB2B1D092001AE4958ED6D20AA180";
    attribute INIT_29 of inst : label is "1A10815AC5000000100000000000000000000000000000000000000080002004";
    attribute INIT_2A of inst : label is "5CC3E5BA80249200014E001A5A5A58BC224938FEA2B6494061E042056B4A102B";
    attribute INIT_2B of inst : label is "00B0D0161A02E96AA504680BA5AA94885549253890A1D151E20E914A8AE8B10A";
    attribute INIT_2C of inst : label is "002884C5720A29CB41F28C2055C21442E6B90E68CA20815042885ED720A50525";
    attribute INIT_2D of inst : label is "DB9C9CE4E7273939C9CE4E7273939A75A251840A80144262B90514EB44A30815";
    attribute INIT_2E of inst : label is "922506A5695D742948A949129352B4AEBA14A554A08149A95A575D0A52AA494A";
    attribute INIT_2F of inst : label is "F723DBCA563944AF65B6414A48941A95A575F0A522A5244A0D4AD2BAF8529152";
    attribute INIT_30 of inst : label is "2802454C68A0908553460356880C60D0190002A5150A05280808AB542E80B81F";
    attribute INIT_31 of inst : label is "1348428AA5229084A52948425FCF2F108C1800A201800E02454D468A00D1531A";
    attribute INIT_32 of inst : label is "2582A8202BA328003C2C0A88069081114A4521014A521094BF9E5EA01E160544";
    attribute INIT_33 of inst : label is "5294D25975B4280259045F690A9245124849068924248144961240A24B000053";
    attribute INIT_34 of inst : label is "08A8904544822A25111128A7B8E7205058809685A1685212002DA42B6D9C0568";
    attribute INIT_35 of inst : label is "25111128A7B8E72051249159208AC904564822B25111928B73CC6205365B1512";
    attribute INIT_36 of inst : label is "801524922A241151208A8904544A2222516F71CC451249151208A8904544822A";
    attribute INIT_37 of inst : label is "323F982A6381075B9A2D256C528D6DB62B5226A0954A14A5EC652AD091014916";
    attribute INIT_38 of inst : label is "058924A512494A4512512EBCA0A2A5385A52AC029202AB0AA0CC665961AED050";
    attribute INIT_39 of inst : label is "FFFCA924A2492833A5205A150585124949188431512A2905264D5F0621461527";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFF71C74D155408C0DC048015DD28243191501465AE08CB136957DBD18";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "3202405E6CDC742AD0AADA6FF53CDDFB40BB543FFFFFC59820F0259827FE2529";
    attribute INIT_01 of inst : label is "F0719000288C41F65810A9B58B1BE454800C0A8289248412BA090244722D24D9";
    attribute INIT_02 of inst : label is "14042E22221A0120349B456B0550002C1541202B216812692253568B129AB47B";
    attribute INIT_03 of inst : label is "9B00043FF169E8412920041CAB81051D480602F4D89385330B8410204008F05A";
    attribute INIT_04 of inst : label is "54821040924D84216EE44FF550EA402495D67570D45922EA83A6DC68D424004A";
    attribute INIT_05 of inst : label is "234A92530A08248692490A492002405BDD001504952092A42095208009369892";
    attribute INIT_06 of inst : label is "9548410410495A52B4B1418AE38E38E5000A4924A7BDC5553803CB608688576D";
    attribute INIT_07 of inst : label is "77480A6749BA63D444C00C460C6C48C4890A852A410828240542095208094117";
    attribute INIT_08 of inst : label is "2E08218F4992D19DE8107EA8611C33413A12E2A23692F63D2794002DA4560240";
    attribute INIT_09 of inst : label is "771A714929340A4E7D4B0BF063E91184169A86B5276B99EA978A645634529B9D";
    attribute INIT_0A of inst : label is "86830A5479B8FE4E90BF706E1822B6975B718CA74D041780F3CAA5C5A2D168B4";
    attribute INIT_0B of inst : label is "B6B7A24B0CA4AFFEFF87266D4061073C93C73DE49E3DE69A221211E5B4014A95";
    attribute INIT_0C of inst : label is "228A2973459296E9548086F0623DA983523BBE1C92FFBFD4DA762F93B565EE33";
    attribute INIT_0D of inst : label is "2056003728185280A16D96A788A26A8EA389A26BEFA0A4AD27949348168E2FF2";
    attribute INIT_0E of inst : label is "7C041004022A5290A9BCB48304896001C67DC04B0F130C0CB130C0BBBE836420";
    attribute INIT_0F of inst : label is "1C0C310009283B2041E09C9881313F0000000000693FFF580145D803F0D9E2EC";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8004086F1484F0010064";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "209082097160F58658672C30C27D71D71A75D488248002920DDFDD5FE2598541";
    attribute INIT_19 of inst : label is "560885A731CF65C8107088383D7184F2C279658753EBADF5C6F2C30D14494240";
    attribute INIT_1A of inst : label is "40820803881A120221A80453020333C1A08420A180D2589313016981CE8E2880";
    attribute INIT_1B of inst : label is "FFCE04E2098C1814E0834729C122439908200E1A0000E1188C08A709CD0C2709";
    attribute INIT_1C of inst : label is "A656595C9D5319D9333938C65EA8E71132784A67ABF7FFAA2897C70A7A8A25E9";
    attribute INIT_1D of inst : label is "19A073AAC4258CC93A5C64B2D3265D9E887744464889311F665B0B1C3970546B";
    attribute INIT_1E of inst : label is "573DF15A7C2A93E4AE0A8F4C49CE9D0492C432B3919E67D59CB2679FFBED04C2";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0940AE21308066873E888E23E9119C9";
    attribute INIT_20 of inst : label is "2155388319DC23562813049E03264288829F1902045188000007380D67422A93";
    attribute INIT_21 of inst : label is "0408A714042A8314042A83100408A310042AA020204538A0215538A020443880";
    attribute INIT_22 of inst : label is "5292524252524252C2D2C2D2C24811111143383E476023AB2AAB3058042AA714";
    attribute INIT_23 of inst : label is "4949094B0B4B0B4B09204444450CE0F92DA034D2429A64D32695184534ABCD02";
    attribute INIT_24 of inst : label is "F000000FF0FFFFFFFFF00FF000FFFFAAFFAD35A6869518461A44E6812B494909";
    attribute INIT_25 of inst : label is "055402AA014400A28055082AA4144202290150855550CE030000FF0FFFFFFFFF";
    attribute INIT_26 of inst : label is "B2C0924E251CA58022DE610129C0948B7998790ACB024A493894729604500A20";
    attribute INIT_27 of inst : label is "21192A9249003470E2404013C8452A620D29830A6008B798404A7022DE661E42";
    attribute INIT_28 of inst : label is "000AFBEFAEBAFAA58590867D2C231C2E900B49B145BE50BADB6D8B2DBE58D0E9";
    attribute INIT_29 of inst : label is "8C98102660000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "270F76D4E9009202505290080A4808006CAA566C8F81408410136040919B0204";
    attribute INIT_2B of inst : label is "30BFC617B8C2F4EB7319C30B532DCC39D6E400CAE63C52D2C2749193E9292135";
    attribute INIT_2C of inst : label is "863090F75049A6D239A2AC2546411848EFA836878AA0951823091FF5049C9C99";
    attribute INIT_2D of inst : label is "B7ADADEDEB6B7B7ADADEDEB6B7B7A9B1185584A8C318487BA834D36230AB0951";
    attribute INIT_2E of inst : label is "829906B1B63630D321AE414C9358DB1B186991D720A649AC6D8D8C34C8EB8199";
    attribute INIT_2F of inst : label is "3403FDDA762E7E82552B46320A641AC6D8D8C34C86B905320D636C6C61A6435C";
    attribute INIT_30 of inst : label is "884151442A22D69559465350894C7487550BD9B4D453A5284928011536A06917";
    attribute INIT_31 of inst : label is "024800912500940295A5297A8B6F051898C9085111788B40514542A210545102";
    attribute INIT_32 of inst : label is "041001A04E8B6C43C2AE2844249005264A01280D2B4AD2F516DE0AA1E1571422";
    attribute INIT_33 of inst : label is "08E497DDA799A6927F9D4BE06900000041000000208000001040000008200000";
    attribute INIT_34 of inst : label is "6A110350881A8441D4220EDA52B4A0DC689AD6358D4350C0A4B9B6841F892423";
    attribute INIT_35 of inst : label is "41D42A0ECAD695A0DC14042A06A150350A81A8541D42A0ECA56B4A0DE5524220";
    attribute INIT_36 of inst : label is "181082808440D42206A110350883A8441DB4A56B4DC14042A06A150350A81A85";
    attribute INIT_37 of inst : label is "BBA80E0B7AE105DF6AAD04081064659623C2D845F2C183964D50C0541D010212";
    attribute INIT_38 of inst : label is "38A004A5C0096B440BCCAED5531A89D1CF4C044204080103103C1E9571ACD417";
    attribute INIT_39 of inst : label is "FFFEA0A04CAA52AB21D350743599E55281B353D28BF1A698CB48027A247A11CA";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFC5145E33B44A42B9648050D48C60555D20AFE4EBF789D8E4C4C4128";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "BB41682C68D0789AE26876509093BA1AE894557FFFFFACED03EE4F2C16FE8919";
    attribute INIT_01 of inst : label is "08C90B80549DCB48D034E1858B6F4C2C2A595695228690C9452B4685008B4A50";
    attribute INIT_02 of inst : label is "8864A427619D12A22F342D1A41A8202D06A1A4E6A94A31A00641320832099044";
    attribute INIT_03 of inst : label is "4A40042DB60D098DAEA21CAC89912D5CC553538586B1D630AF662041C0AD6B54";
    attribute INIT_04 of inst : label is "60449890D3688C816AEC05A9026D041351252106495ACA44010259225CD04224";
    attribute INIT_05 of inst : label is "AF2C59526B6CB2D5E50D95045045440416821A869950D32930D811410DA23213";
    attribute INIT_06 of inst : label is "D96D04104100C631AD2A5704000000024110A282140004E9204A2251D31D17F9";
    attribute INIT_07 of inst : label is "16A0834268B4312C2AC2CEAB6186A56C306B0DB0224C408914930D81122A0456";
    attribute INIT_08 of inst : label is "6C54697D8013535B59556A992948A18A978852ECE298D6C0D044102E48284544";
    attribute INIT_09 of inst : label is "9201232492590C20692B6109C945248417591242D15A8909C910481796420B58";
    attribute INIT_0A of inst : label is "0A15134D2658D2B49C0E74180CEF1689E1529BF157041682D22492180C060301";
    attribute INIT_0B of inst : label is "0818426A7289C80452053427E8A7AD100405688020288004020006B53E446A9E";
    attribute INIT_0C of inst : label is "471C74840A0AD49476D216939A398B1296B4E150270A111A4C785405C0421002";
    attribute INIT_0D of inst : label is "21A920246A935B2AD0B6D6C3B1EC790E4791E43AEAA9B4EC942844045BC854C8";
    attribute INIT_0E of inst : label is "8004140402090C1AD01322A4D43F9E08ACA5F57DF212265C302060FAEAA754A5";
    attribute INIT_0F of inst : label is "5F2F86FBAFDEB96DE7F6CC00ADF0F58000000000400000000787E01C01260113";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8AEDC677AD97F1930BE7";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "B6564B65456290514554828A2AE10410570417C592924ADB6D7DDFFD801B2D61";
    attribute INIT_19 of inst : label is "FBDADFE3F2ED76F9776829B8A41455482AE4105057082A8015C0082ED14C9924";
    attribute INIT_1A of inst : label is "7DFBEDB3987B97CEFBFB26F5FFCF7FF9AAA5FAE79CD57CA7779E27B9FEBF3BB4";
    attribute INIT_1B of inst : label is "FF8E83F6EFFCEF78E85BFFF1D0EDFFF9B7B6CE9DABD4E8BBBDEFC747FD378745";
    attribute INIT_1C of inst : label is "ACC6DB199D4B33DB66BB7ACD599A563376FA1A5666926CCAA897176AE08A25AB";
    attribute INIT_1D of inst : label is "1DA06B1DE451CADB6AC96DB6566D5E5BBACCCCCCD9DB3B3CAF7DD88510B04966";
    attribute INIT_1E of inst : label is "F0C820761E69381446092D58DB845A86A8E526B73DB9613359B6E15A69A097F0";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAF5559065FAC07686B1999B66933B84D";
    attribute INIT_20 of inst : label is "4C44A0A09915322420121517096FCDD996BA1884C44A0A000000008190476823";
    attribute INIT_21 of inst : label is "09AAB0100988B01009AAB01009AA901009A220A04C44A0A04D55A0A04D54A0A0";
    attribute INIT_22 of inst : label is "52029292829212820212928280014141415402015A202900C082206209AAB010";
    attribute INIT_23 of inst : label is "0A484A08084A4A0A0005050505500805682026FA4A1A70D2A293780514BBC542";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFF00FFFFFF555000D39A5169378045A4CE2A1290A4A4A";
    attribute INIT_25 of inst : label is "0112008B004580224015280AB4055A02A501129444440013F0F0000FFFFFFFFF";
    attribute INIT_26 of inst : label is "D68396EFF450818222C1950529489C8B06525D195A0E4E5B3ED54286155802AC";
    attribute INIT_27 of inst : label is "B61D67410C92C860CEC14B33B105A0C21909864060C8B065414AD322C1949746";
    attribute INIT_28 of inst : label is "FDF4410410411506520ED0226463082CD96592B01ED2C0B16DB581F6D2C0C0CD";
    attribute INIT_29 of inst : label is "2009C0E3075FEBAC5B26914229C6E8531B295C6F8AE5FA9FD7F8EE5BABBD7FA7";
    attribute INIT_2A of inst : label is "780C9A4ACDB64AD93902D92B692928001A6D20928092491CB28127038409381C";
    attribute INIT_2B of inst : label is "264042C80859008B2308A164A22C8811564480B18215B3B38652134B39D98328";
    attribute INIT_2C of inst : label is "B6CBB2A558E9E5CE677194ECC39B65D9D6AC6E4CC643B30B6CBB3AD58F901410";
    attribute INIT_2D of inst : label is "6B3909C84A4656B3909C84A4656B397732329D985B65D952AC74F2EA64653B30";
    attribute INIT_2E of inst : label is "8A9514B6D06064CD21AD454A9A5B6030324691D6A2A54D2DB418193348EB4569";
    attribute INIT_2F of inst : label is "1722D98A7E0160192498086A2A5452DB4181933486B5152A296D80C0C91A435A";
    attribute INIT_30 of inst : label is "8A8C91599229BCECCD5EDB5BBB6D72820126CE7C89011C9B24B3AA14B3644702";
    attribute INIT_31 of inst : label is "8B253161939A4E69EE399B2788C5845410DBF9BB3249928D91589B22A364566C";
    attribute INIT_32 of inst : label is "0007FEC1A8122D7FFCEDEFDF164A62C327349CD3CCF7164F118B08BFFE76F7EF";
    attribute INIT_33 of inst : label is "0A4300221161ACDA0049A24C6B00000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "461C0230E01187018C380C331CE62498A9938A1284A1204836C4000260853CC3";
    attribute INIT_35 of inst : label is "018C300C3398E7249B65BC30046180230C01186018C300C3318E62499249C380";
    attribute INIT_36 of inst : label is "1120ECB786008C30046180230C0318601847318E49B65BC30046180230C01186";
    attribute INIT_37 of inst : label is "B92FE84B3285951B8A3DB52C50CC6DB623DBB846F38307878D71AA9050254B56";
    attribute INIT_38 of inst : label is "280492458924B9EC88081C45867A80E1EF5AA80B9683AA0C3BFC0021E3BE5094";
    attribute INIT_39 of inst : label is "FFFCDB2D82492163A086605C369192490526F7820FA1AC34A22D0068EC28D0C8";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFF0A28E152032B4B2D0A8866A5ACE8444411EAC6FFF5CDF3698842038";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B308611B6AD36DBBB6EF4A20C1B25411619678FFFFFFB68BACE9767CD6FE8909";
    attribute INIT_01 of inst : label is "D4D994126C9DFB83CA946CA48B765CDC891C4647AF804EC9C14906A4486B22D2";
    attribute INIT_02 of inst : label is "132CA9AC445B17A06D366CD908F84D2423E0146EB2CA95048ED932CC76C99664";
    attribute INIT_03 of inst : label is "CA24B2C9274D4DEDAFA05DDD81956C5FCFFBCB0484959395254B740949ADEB76";
    attribute INIT_04 of inst : label is "740E91D009688E9162FCC929064F09B3CD0521265C5F794D0B02DB2ACCF0096F";
    attribute INIT_05 of inst : label is "A7664B52292C92CDBF2D9F40F00F00841784CF804D7009AD22DD03C265A2BA53";
    attribute INIT_06 of inst : label is "F87D75D75D705695842E1D0EBAEBAEBB503A87A05C0C5CFCA00B2054C94CB6C8";
    attribute INIT_07 of inst : label is "D6E811562AB645AC8A40E4B2C25586584A29A5BA0748E81D06D22DD03A0F40F6";
    attribute INIT_08 of inst : label is "060AEB4A593B95FF5F4F20BB6948B04156CA526EF6DAD6E83EA2492FECB89F00";
    attribute INIT_09 of inst : label is "D261236D9F6D27A328AB6BD5D9856CB1B7D9B265365ED50954F23936DB58DB58";
    attribute INIT_0A of inst : label is "1583BB5D69FBFAEED01DF616112FB6CD2155D997E731B636D6FC3F6EB75BADD6";
    attribute INIT_0B of inst : label is "1757E12A7E56D8044A0EB67531576D2F8855696C43A96CE8F6DB2B4722CA39F2";
    attribute INIT_0C of inst : label is "228A0E23C1DA50847259D691F93109561296A5155B08515CE166059AB1A10C3B";
    attribute INIT_0D of inst : label is "B37F0085EFB15BA9B1F7C2298E6298F22C8F22854440BCEC9514EE4AD61A0436";
    attribute INIT_0E of inst : label is "FFF84050820FA900B1AB73AEB71CFE40A40514AFF009102448C1A2055102D7B4";
    attribute INIT_0F of inst : label is "A0D000045021469218093389617DF92800AA0000400000004A00000001FFFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF512398852680E6CF418";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "9256D9254483E9A69A0B4D34D05A69A68869A20DB6B6DA492A20A08AF807ACA9";
    attribute INIT_19 of inst : label is "0425201C0D128906888924A0FA69A034D11A69A68AD34469A034D340C924DB6D";
    attribute INIT_1A of inst : label is "8204124C678468310404D90A00308006555A0518632A83588861D8460140C44B";
    attribute INIT_1B of inst : label is "FFF104091003108710A4000E2112000648493162542B11444210388802C8788A";
    attribute INIT_1C of inst : label is "2CD6DA510C5A225825B02A8BD912D43376A4D2D44440040641360C0AC1B04DEB";
    attribute INIT_1D of inst : label is "5D244A571C70329B62CB4DA60605D250BAC8888891110A242A490B458A104144";
    attribute INIT_1E of inst : label is "160F1854E308280502082858DA835380781924B1258B4A2251A62A5024919482";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF05155FC4520097494A11111448222A89";
    attribute INIT_20 of inst : label is "2CCB75B8FF1DFEE6A6118DE7380C1331C72ECE22CCA75BBBBBBBCB88E50AB489";
    attribute INIT_21 of inst : label is "85996AB385996AB385BB6AB385BB6AB385AEC34C2DDB75BC2CCA75BC2CCA75BC";
    attribute INIT_22 of inst : label is "93B60E0E0E1E9E369E8E0E0E8EDBFEABFEABCE61E2A5290101867C5985996AB3";
    attribute INIT_23 of inst : label is "307270D2723030323B6AAFFAAFFF3187CA2522B24BA24D124C99DE0664EEF803";
    attribute INIT_24 of inst : label is "FFFFFF000000000FFFFFF00000000AAAAA912224149D9F04527778018BD03030";
    attribute INIT_25 of inst : label is "C760F3B271D93CECB4724739039C818E40E7206FAFAFF2630FFFFF0FFFFFFFFF";
    attribute INIT_26 of inst : label is "98A9948A0332E9E23AC107C5DE48ECEB04731D9E72B676522808CB271D83CEC1";
    attribute INIT_27 of inst : label is "92DB27C02592E1724EC94833A36CA8531A19E6C6708CB041E1679232C11CC767";
    attribute INIT_28 of inst : label is "000AFEAFEAFEBD815B83DF997D694898492FB623F1B6E263EDB11F8DB6F262C4";
    attribute INIT_29 of inst : label is "87C0844628000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "7B4CDB4EC4924ADB7722DB6B6B6B68002341A4FE9D5A0DB12496021110F81088";
    attribute INIT_2B of inst : label is "A27A924E5A49EACB4A88C9272B2D2C95D69414B3B6B937972EDB138B999B9778";
    attribute INIT_2C of inst : label is "926993EF9659657A32199C64D38934C963CB2BC66671934926992E7965985858";
    attribute INIT_2D of inst : label is "918C8CE4E7231DB9C9C766327391895D17338C9A4934C9E7CB2CB2BA2E661934";
    attribute INIT_2E of inst : label is "5A34B5B7937BE1D32BED2D1A4ADBC1BDF0C994F6968D256DE0DEF864CA7B8599";
    attribute INIT_2F of inst : label is "0D6495D96C7B6807E1F8136968D2D6DE0DEF864CAFB4B4696B6F26F7C3A657DA";
    attribute INIT_30 of inst : label is "5B8F0B71E16D3DC5DECE4A68992987F6890E592C9D6B34B9259DFF25F2C54C3F";
    attribute INIT_31 of inst : label is "0BA621C9D2134848CF718912070943660883826631E18F8E0B71DE16E3C2DC78";
    attribute INIT_32 of inst : label is "004F766952BB6C80006900AB176863D3B636D8DBDC7792240E1286C000348055";
    attribute INIT_33 of inst : label is "4AD249205264A44B86B0E20D2920120904924000824124820024124020120120";
    attribute INIT_34 of inst : label is "D4B9D6A5CEB52E74A973A53398E72D99CBB18C93A4C932411269A61BE0C49C69";
    attribute INIT_35 of inst : label is "74A973A53318E62D99A0D97BAD4BDD6A5EEB52F74A97BA5231CC62D9BE1F973A";
    attribute INIT_36 of inst : label is "B374B41B2F75A97BAD4BDD6A5EE952F74A47398E599A0D973AD4B9D6A5CEB52E";
    attribute INIT_37 of inst : label is "BDFFFC47BFC79FBBFB3DB7B4DACC4D34645A884593BB378728B5BFCA5047EDCC";
    attribute INIT_38 of inst : label is "2D4492658924C9548D0C1C5B833B94C9CE5BFC8EDB93FF2EB001FE51E2BED88A";
    attribute INIT_39 of inst : label is "FFFCED06D7C3F4EBB482764524B5BE1FA5465A820B612C14AE2F212C652C54C9";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFF450442972A6959AC8E013284ADACC000160156DC0AEDB6684D4ABBB";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "229052004C9B000A002A4200E002101040203FFFFFFFE48900F82EF865FE40BC";
    attribute INIT_01 of inst : label is "6800880400080064430600351249040432699A9D01848612366A6041968D4C89";
    attribute INIT_02 of inst : label is "124D0788254901A0000114286D1848A9B461261C1FC102CB2000000300000009";
    attribute INIT_03 of inst : label is "3B4000249460206109A01501000480945551504936A345A2882110001000420A";
    attribute INIT_04 of inst : label is "101210409243B4224CA51485B0A3002541964DB0919000299266104C90349003";
    attribute INIT_05 of inst : label is "4248921B420124001D412300300340325D84918491B09234200404C2490ED098";
    attribute INIT_06 of inst : label is "9049A61A61A95AF7B5FA142051051055100801803010812832005B3181180524";
    attribute INIT_07 of inst : label is "25600A25432A335462826A62400C8C4801024008090821040542004048090805";
    attribute INIT_08 of inst : label is "2A0492C108B8414A68904E0010941140A052A4802012A498935492AA41580309";
    attribute INIT_09 of inst : label is "0B4E5440240048584D320A680268012105120497E528C8020D02010596508293";
    attribute INIT_0A of inst : label is "02802002144914BA9484146208A204133410849069A10420A5C825A04028100A";
    attribute INIT_0B of inst : label is "0070400310ADDB0DC1680225200000B8818245D40C05D442B4921E5178075212";
    attribute INIT_0C of inst : label is "20820460400006CB0080E0C882A52A24D52F361CB70B77C00A5E23C589637F61";
    attribute INIT_0D of inst : label is "01290136222A001291924491204812449120480014A1020003045240001622E2";
    attribute INIT_0E of inst : label is "00001054022B9CCE6D3FF28001A48080CA920915099020448912040010852001";
    attribute INIT_0F of inst : label is "0000010000000000000000241F169400A0020000C00000006C07E00000000000";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "0000000079104104100A08208150410408C1002000000000002A0A0A74411510";
    attribute INIT_19 of inst : label is "00000000000000000010C90410410220801041040882014100A0820594400000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "FF80000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "A2D6DB5D98031909121904C4D8CC2711666458263364B72A2084D5021AA8A108";
    attribute INIT_1D of inst : label is "99C9738B7C30FCEB44C06DB6C720DB9E2484444659988910660044A542646673";
    attribute INIT_1E of inst : label is "594E9176522CB435348CCF44598A9D84987E1213909863199DB6639C924C02C8";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF545550220B2226727388889220B338E8";
    attribute INIT_20 of inst : label is "60442AA3990D32002B83231604208510F2B211E60442AA141417A0042D122010";
    attribute INIT_21 of inst : label is "CC2A8150CC2A8150CC088150CC088150CC02201660452AA660452AA660452AA6";
    attribute INIT_22 of inst : label is "54DB13131303031B03038303036D55540003A221CAEA12AB2A497C70CC2A8150";
    attribute INIT_23 of inst : label is "44040464040604040DB00555500E80872B6A105A80DAA6D536A628A9B5114754";
    attribute INIT_24 of inst : label is "000000FFFFFFFFF000000FFF0FFFF000002D55AA82A668AA0A99A7AA68644444";
    attribute INIT_25 of inst : label is "311408880C4402221B11008880444062201110055005EA12F00000F000000000";
    attribute INIT_26 of inst : label is "52B3A6CE09BBB5B44CA08F60795135328278D9095ADE9A9B3826EED6C4502228";
    attribute INIT_27 of inst : label is "041048C24120066420121544580006A0598DB62365112823C80E5444A09E3642";
    attribute INIT_28 of inst : label is "000500055500168186688745121294260000499180001098124C8C00000C18E8";
    attribute INIT_29 of inst : label is "0062A14210000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0C912CB0A000000011000000000007FFE482419206A4525041088A85000C5428";
    attribute INIT_2B of inst : label is "94876491EC923E12381512487848E32C6471285A0522D070402CD4722A782007";
    attribute INIT_2C of inst : label is "2492243540BAAB1B5DC2228924D249120AA05CCB889A2492492251D40BA7C3C3";
    attribute INIT_2D of inst : label is "6F3939494A4A5273939DBCE4A5252AC5A844D1249249121AA055558B5088A249";
    attribute INIT_2E of inst : label is "912920207005344D520A4894901038021A26A905244A480818014D035482606A";
    attribute INIT_2F of inst : label is "140241825A344C8E4126401244A48081C014D135482922524040C008681AA414";
    attribute INIT_30 of inst : label is "2A61454C08AA56B511400353800D65459D0B94F55252A12249072A510E42601B";
    attribute INIT_31 of inst : label is "4108081084061017B5AD78021ECF2E5B1C0890A213409A60454D008A98515302";
    attribute INIT_32 of inst : label is "804A83A16A8A0840020F428882141021080C202F79DAD0043D9E5CA00107A144";
    attribute INIT_33 of inst : label is "84AD96496DB84A105B4D19621204020804904800804904024024924120924920";
    attribute INIT_34 of inst : label is "85222429152148890A45485AD694A05428085324C9124C92A012D9A814080130";
    attribute INIT_35 of inst : label is "890A4D484A52B5A056400A45485222429152148890A45484A56B5A054000A454";
    attribute INIT_36 of inst : label is "0808000149A90A4C48526A429312149A90B4A52B456412A4D485262429352149";
    attribute INIT_37 of inst : label is "32386A8243A8A10408800201042D6DB6AB0132ABF44080704C586A9609080051";
    attribute INIT_38 of inst : label is "1229249552492A45115422A0F404A9106B46A95000A8AA410BFDFEB41402C500";
    attribute INIT_39 of inst : label is "FFFE12092C824A670975003A5689641240B0E73155AAA3AD434541128A528912";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFC1040C55020000391612441549008000E40124040208039DC0BF88A";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "E520A401CF9B24149052400000C2000024333FFFFFFFE48820F808C27CFEE428";
    attribute INIT_01 of inst : label is "330E9061A76B0E6CB1E78716369D0B0B16308D885B0931B6B72E3878B386C799";
    attribute INIT_02 of inst : label is "32CB0298154813292493DB362E7091B0B9C2478E1FE3E649710C88618864431B";
    attribute INIT_03 of inst : label is "BBC32C2499703B1B1B2923370104B8F4B00020DB12E74DE798A531163084E41E";
    attribute INIT_04 of inst : label is "3136B4C124C19862C5AB348493B61B6C3593C49DA5B006389C2631C7A2612690";
    attribute INIT_05 of inst : label is "1AD3A40BC4DB6DB480DB6E1261261216DF09270924E1249D690C4D849306618C";
    attribute INIT_06 of inst : label is "9049C71E79CB5AD6BDF00072E38F3CE7049893093031C3073230D92130130D27";
    attribute INIT_07 of inst : label is "6DC24C39836E061A63827A62004C0C4009C4FA189B5A634D4DD690C4DA9B1A0D";
    attribute INIT_08 of inst : label is "1A099EA30124C10030B1CE61DCF611413233BD1B81B3AD38A19C30B806712612";
    attribute INIT_09 of inst : label is "DB8FDC926C0292598E36CC330E7807630C769DBDBD08D80605160B0C20B186F3";
    attribute INIT_0A of inst : label is "06836C239C41451FB4402C41F0B80DB70011348362630C63AD8001CC663B1D8C";
    attribute INIT_0B of inst : label is "16302481C9A913018B7B4245004C39EC89C28F644E0F648B8DB61D114027C610";
    attribute INIT_0C of inst : label is "208208634121024BCD363CCC46AD2E7CDDE9C236A40142E48A5606F083616BB1";
    attribute INIT_0D of inst : label is "610082125AEE369681000531485314C5214C52000407639A4304D249003606BA";
    attribute INIT_0E of inst : label is "0000040002393DCE336FCA000DE40100F8B28B1803A1428102040800101C2C63";
    attribute INIT_0F of inst : label is "00000000000000000000003DDD3D0E02A80282A0C00000007000000000000000";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "490924903B1D71C71C238E38E01C71C708F1C2324849212482800AA040005B3E";
    attribute INIT_19 of inst : label is "00000000000000000016DB075C71C2B8E15C71C702E38171C0B8E385B6D26492";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "FF80000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "BA7249CCB809191B923B8E4448CF331122C00832336D9733A68C65038CC9230E";
    attribute INIT_1D of inst : label is "0CF1398E1C603E71C4612492427049CF470444644CCC491046246022027F8732";
    attribute INIT_1E of inst : label is "E04000830010941527F0E5744B00CF09301F923691B13119CC92D1CD925E42E9";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF002AA0230BA2433C3988889320999458";
    attribute INIT_20 of inst : label is "3A650043AA4D5412294966948C188404729061F3A6500415401200266D10089C";
    attribute INIT_21 of inst : label is "674C840C674C840C674C840C674C840C675320333A6500433A6500433A650043";
    attribute INIT_22 of inst : label is "784B23232323230B2323232321255555555600019A939EAB2A494C18674C840C";
    attribute INIT_23 of inst : label is "848484248484848484900555555808066A539C5F204F227913C330B09E198498";
    attribute INIT_24 of inst : label is "000000000000000000000FFF00000AAAAAA794F2C3C330B30F0CC24C3C248484";
    attribute INIT_25 of inst : label is "3D998ECCCF6663B30BD998ECCC76667B331D9985555081060F0FFF0000000000";
    attribute INIT_26 of inst : label is "52A2C26640A2189987808E303B66161E0268530B4A8B0B0999028862F6663B33";
    attribute INIT_27 of inst : label is "6C70D9849A49A44799A425884C320338498512214661E0238C0E5987809A14C2";
    attribute INIT_28 of inst : label is "000555500000178DB4683404C7DCE727249A499C40019C9E924CE200018798B3";
    attribute INIT_29 of inst : label is "4660A10020000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "C4E32593B2492124908124848484800060000300430000910018828408CC1420";
    attribute INIT_2B of inst : label is "99253925AF24961618623C92585861C46C324E4C19C278D87124D83E6C2C7885";
    attribute INIT_2C of inst : label is "493C493C433CB2149CC4471238649E241A2194B3910C48E493C491C433C6C6C6";
    attribute INIT_2D of inst : label is "273939C9CE4E76D2929494A4A5252C8248886247249E240A219659449910C48E";
    attribute INIT_2E of inst : label is "214A4069218F36059C1A90A5203490C79B02CE0D4852901A48638D816706302C";
    attribute INIT_2F of inst : label is "C01A4104DB89CC8C00024194852901A4C638D916706A429480D2631C6C8B3835";
    attribute INIT_30 of inst : label is "04392087241256B621E12196C48669599F11E476669CC344936F019A060470C0";
    attribute INIT_31 of inst : label is "61080C9C84061017BDEF6C12090525994A06908089044838208672410E4821C9";
    attribute INIT_32 of inst : label is "120003E241081B43FF074201C23439791A1C68652B4A5824120A4B21FF83A100";
    attribute INIT_33 of inst : label is "E724B2DB25BF5BA0598E597BD624904924124924920924904904904904024824";
    attribute INIT_34 of inst : label is "05C3382E1DC170EE0B86705AD6B5B2366C4E61C8F23C8724CDB259C81003621E";
    attribute INIT_35 of inst : label is "EE0B86704A52B5B236400B8E705C7382E3DC171EE0B8E705AD294B234000B867";
    attribute INIT_36 of inst : label is "CC9E000171CE0B8E705C7B82E3DC171CE0B5AD69636412B86705C3382E1DC170";
    attribute INIT_37 of inst : label is "221073304132C21414C24002272524933321BB12D8CC9858E64E406709120021";
    attribute INIT_38 of inst : label is "96B2493764926C0261244114D9064E1C6B740664004C0193CBFDFEAE1841A660";
    attribute INIT_39 of inst : label is "FFFF3209480012224E59933B96EF40009092B5A865ACBACA45809DD313930E33";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFC1040E5D3284269B3C24DC177B438000AC0108400210809775BD896";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
