-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0B92300C0C481F961DD41F96273C033012301F960B931DDD303835350F611A1C";
    attribute INIT_01 of inst : label is "55550000311D0000744C00001115300C5444300C755D300C0FC316340FC41796";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF0000000000FF00FF00FF00FF00FF00FF300C300C";
    attribute INIT_03 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FFE40B16940AA00AA00AA00000";
    attribute INIT_04 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_05 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_06 of inst : label is "123020081DD42A282BA92A280F78022031342A2813362AAA30302A2A0FC32028";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF1F9728281E9C2A28";
    attribute INIT_08 of inst : label is "0DD1222A1DD408801D1C2A2A0FC328A80CC022281FD62AA80FC30A8200000000";
    attribute INIT_09 of inst : label is "0FC32A283FDF0A823FFF0A820C0C2A2A3CE40AA203032A2830302A2A1FD70A82";
    attribute INIT_0A of inst : label is "3FD70A820FD720000FC32A28303020201D942A280FD30AA20FC3282A0FC30880";
    attribute INIT_0B of inst : label is "FFFF3EBC8D1E3450448D1410848DD710848D141032342AAA1B1E20203A3C0A82";
    attribute INIT_0C of inst : label is "98040200755F0000C003169402101004755D300C7FFD300CFFFF3EBCFFFF3EBC";
    attribute INIT_0D of inst : label is "9FF600006559300C4961300C82820C3042812008096000002418000010240480";
    attribute INIT_0E of inst : label is "9006955612842828396C0000300C1C340C301824C0031694341CC28355550000";
    attribute INIT_0F of inst : label is "3D7C2008341C0000C003955603C016940C301824141684408550011241411824";
    attribute INIT_10 of inst : label is "300C382C3C3C000012840AA00820C143CBE33FFCC2839FF6800287D27FFD382C";
    attribute INIT_11 of inst : label is "FFFFFFFF0000000000000000FCECC080CCC4FFFD000000009884033212268CC0";
    attribute INIT_12 of inst : label is "8BB02181B2CD1B878D141B26CDBBB26EDF8B015C2C17C2093B3F020313337FFF";
    attribute INIT_13 of inst : label is "60615598D650AF56E238D28AB246D862AA28A42383C2579814428A888E578520";
    attribute INIT_14 of inst : label is "861C5141DFB4F2C509704D38A2AC91BA18A2422908ECF091566241057981655A";
    attribute INIT_15 of inst : label is "D1C13492292AC977956635144E288B26CDA6549A49E58EFACB1C5F791C5D7122";
    attribute INIT_16 of inst : label is "5519AC9460E6CF5269E5811C13492393AC9779566051473CA0B8B27FD5249E38";
    attribute INIT_17 of inst : label is "2C9A7DCB269BCB2650B92814B2DC6D5B75DA482682B66F2CDA67CB25D6B45566";
    attribute INIT_18 of inst : label is "608ECB26082FF1C5248A1849E3BA083BFD7149A2861A796E82164B26CDB8E6F1";
    attribute INIT_19 of inst : label is "7DD24CCCEDEE9654171BFC7FE7B779526741462C9422BF09B7B1597695666514";
    attribute INIT_1A of inst : label is "3B08AA9946242E6E299EDEE47DD259F07505CA7D397D394D094D0951111DDEE4";
    attribute INIT_1B of inst : label is "BCE888E4D1BD09D27DCB5935415467CA822A518908E658B41A52E94785D505C2";
    attribute INIT_1C of inst : label is "124D1BD0AD64D50559C0995B0B9182655CE656C6242E57749F7412D64D505467";
    attribute INIT_1D of inst : label is "C5E4CCCEDEE96537FFF1BFFF08EE18AE0939F070D0735D27DDAB8988697B947E";
    attribute INIT_1E of inst : label is "8BFAFEC1CB2C97E5D92947D9267D55515D5951595149414941797179717951FF";
    attribute INIT_1F of inst : label is "A181A2C9B4420219443FC24EFF251BD242C9C3532C485D710EB1217DE72C988F";
    attribute INIT_20 of inst : label is "30300303000000000C0CC0C00000000095D40F0724B09C0BC72423ABD44BC327";
    attribute INIT_21 of inst : label is "0002000000000000A00800000000000032320202000000000000C4C400000000";
    attribute INIT_22 of inst : label is "0220000000000000088000000000000000200000000000000080000000000000";
    attribute INIT_23 of inst : label is "0000000100000000000040000000000000000103000000000000C04000000000";
    attribute INIT_24 of inst : label is "00000000000000000000032103120000000000000000000000001C8C2C4C0000";
    attribute INIT_25 of inst : label is "000023339CCC0000BFFD40400000002000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "000048C084C0000000000000000000000000000200000000C0C0E8C8CCC4C0C0";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000003234313800000000000020000000";
    attribute INIT_28 of inst : label is "35FF3F0013170000F5FFFC33DCD4000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "FF5F00FF17370000DF7F02EBDCD40000FF5F00FF17370000FD5F32FDDCD40000";
    attribute INIT_2A of inst : label is "17CB0921CE0CACE3DF0B015C2C17C209FF5F00FF17370000FD5F03FCDCD40000";
    attribute INIT_2B of inst : label is "1F42CCA38F1614D067010450A701C45CA7010450A6310450A63104508BF45C10";
    attribute INIT_2C of inst : label is "B1C89F4D1A101E7D1A101E7D014BDF692A3707B43B7FECC38174A1287F3702A1";
    attribute INIT_2D of inst : label is "68A66701549494107C060BE049346141813490644D2400A44D249C491341272D";
    attribute INIT_2E of inst : label is "A24F01C89969E7AD79D4A169159249559665969A75A79635E45205E456582555";
    attribute INIT_2F of inst : label is "66F093510D98164F8915D0684114A4797C6464795C64612ACA1791D6219A23AC";
    attribute INIT_30 of inst : label is "B95953565991C90969D5465CD6859565596B5114B857456655D16A153416D38D";
    attribute INIT_31 of inst : label is "5A85A7927B622C714D6569A54515A5B92C60665A547192D6589DC219566A5117";
    attribute INIT_32 of inst : label is "A83C2085B3C9294F8D14096EEE3793EAE5276ACC90EAC606675A59269E4BF61A";
    attribute INIT_33 of inst : label is "50A16654D4589D9EC2B8E24A91CAD8628AA884A3B00E665C1442AA089D1B8424";
    attribute INIT_34 of inst : label is "87185045ED7CF1C918344E34A3A8A276286242293B20E0D1546A410568C55696";
    attribute INIT_35 of inst : label is "F04524D20AA6D937956605D44E28892EED2666527925BE3ACB1C5E7D1F5140E6";
    attribute INIT_36 of inst : label is "4655AD9071A2DC1E79A58314124D209FAD9359D65091473CA2B093FBC5648E78";
    attribute INIT_37 of inst : label is "2E927EC7269BC92E62710990B3D85E9776D64922A13A4FACD96BC92DE5785566";
    attribute INIT_38 of inst : label is "6382C92E0B23F1C526821A41E2BE0A33DCF56826861A5BE6811A492EEE34F4B9";
    attribute INIT_39 of inst : label is "7CD67F00FFA69558065FDFF3E5BF58D6548D472884628ECDA4FD597695664594";
    attribute INIT_3A of inst : label is "0ACCAA9945281FAA2B96FD687CD6787445C5DB391BF51BC51B0518150355FD68";
    attribute INIT_3B of inst : label is "BEE0B920E37538167EC749755114768E822A624539226970185AD987B5153406";
    attribute INIT_3C of inst : label is "1349385C9DA4C54578449A57281D91297D62754A07A2557C9D7C315A5C145563";
    attribute INIT_3D of inst : label is "F524FF02FE6945B7FCFDBFFF3B222B620A35D0F0D0734D67EE67AA045AB79772";
    attribute INIT_3E of inst : label is "BA3EFCC9CB2CB56DCA65761D17B954555E55525552455205523552F552F57377";
    attribute INIT_3F of inst : label is "A085B28994C202194733D30ACDED385E7209D01F1E805C752C3913B5C7ACAB43";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1555302411142FE91554030311101FF5151523291514363C1010303010140FC3";
    attribute INIT_01 of inst : label is "00000000300C0000300C00000000300C0000300C300C300C15142B2B14143979";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF0000000000FF00FF00FF00FF00FF00FF300C300C";
    attribute INIT_03 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF2968D8070550055000000AA0";
    attribute INIT_04 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_05 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_06 of inst : label is "2FEB300C262C0FC32EE8074333342BBA2B3A07432F692C6C3034303025380F86";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF2F6903122D6823E3";
    attribute INIT_08 of inst : label is "262E0F872EEA0CC02E2E0C0C2DF80FD2272D0D852FE90FC3253C2FEB00000000";
    attribute INIT_09 of inst : label is "2F690FC30FC72FF30FD72FC30C0C0C0C0FD23DF8030307433A3A30300FC30FC3";
    attribute INIT_0A of inst : label is "0FC32FFF0FC33A3C0FC30FC33A3A30302D7807432FE93DF82F692FF22FE92EE8";
    attribute INIT_0B of inst : label is "3D7CFFFFAABF1145ACC40020ACC461A0ACC420A02BBB2C4C0F0F30300FD72F7D";
    attribute INIT_0C of inst : label is "004020190000A0082968C0032968300C300C300C341C3EBC3D7CFFFF3D7CFFFF";
    attribute INIT_0D of inst : label is "C143382C300C9AA6300C86920C30414124180690100418240000200801202408";
    attribute INIT_0E of inst : label is "6AA96009141421480000369C2C38300C24180C302968C00300006FF90000AAAA";
    attribute INIT_0F of inst : label is "10043EBC0000382C6AA9C003296803C024180C300221682848800AA124188282";
    attribute INIT_10 of inst : label is "341C300C00003C3C05502148C28304107FFDC7D36FF9C1434BE14001341CBFFE";
    attribute INIT_11 of inst : label is "FFFFFFFF0000000000000000FFFECCC8C040FCDC000000004CC0211903316448";
    attribute INIT_12 of inst : label is "844677B799160BEFC4516459164445B3234EE46044AB14CFBFFF23330103373F";
    attribute INIT_13 of inst : label is "3080544CE129CC54C348179AC596C564878D2634BB02544CE218D210D254DD30";
    attribute INIT_14 of inst : label is "9ABC461ACCC20B1608034179E6B165B15925E7498D2AC0915130804544CE2151";
    attribute INIT_15 of inst : label is "1BC010637B7B1654D553280542302C5916A6D59249249ECE3BBC430EBC430E36";
    attribute INIT_16 of inst : label is "1802316570238A5649248DBC000237B7B1654D55328054B16EC2C580A5649278";
    attribute INIT_17 of inst : label is "91646D6459146459509D7822A73351A479534E34824490916648EC5953469513";
    attribute INIT_18 of inst : label is "58DEEC5B8DA02D85648C8F49278C9F780B61592323D2492327D2AC591648B530";
    attribute INIT_19 of inst : label is "716362220D74534426480A40A4454D55318854B16E378C6858C58D54D5131805";
    attribute INIT_1A of inst : label is "498D21D7567563511DD9E996716373F42109960D0D0D0D1D1D1D1D1DD5512996";
    attribute INIT_1B of inst : label is "71250D21D58D59F6CB33CB2CD6CC5712A349D59D5835D420A7601D2FC40C5863";
    attribute INIT_1C of inst : label is "235D58D58F2CB35B1D81D75C58D5875D7035D71675635C7DB2E0ACF2CB35B055";
    attribute INIT_1D of inst : label is "49222220D7453455CCC59CCC592759275A23F22C82A01F6CB06665559D265671";
    attribute INIT_1E of inst : label is "4EF6BD9A2C11633C53100BF311BD2525212121252529292D2D393135353199CC";
    attribute INIT_1F of inst : label is "E6B68B16469ADA0967F3079AAA3768869B168690EECC430E03BB310C38B1682F";
    attribute INIT_20 of inst : label is "03300003000000000CC0C00000000000BCDC3A033810CC7AC53825CC78B6C31A";
    attribute INIT_21 of inst : label is "000100000000000000040000000000000101313100000000C8C8000000000000";
    attribute INIT_22 of inst : label is "0100000000000000004000000000000001100000000000000440000000000000";
    attribute INIT_23 of inst : label is "000200000000000080000000000000000203000000000000C080000000000000";
    attribute INIT_24 of inst : label is "00000000000000000000003000000000000000000000000000000CC000000000";
    attribute INIT_25 of inst : label is "0203393CCCC00000DCDC000000003B3E00000000000000000000000000000000";
    attribute INIT_26 of inst : label is "00000C000000000000000000000000000000000300000000C0C0DCCC0000C0C0";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000330000000000000000030000000";
    attribute INIT_28 of inst : label is "3F003AFF0000232BFC32FAEE0000ECE800000000000000000000000000000000";
    attribute INIT_29 of inst : label is "00FFFFAF00002B3B01EFEFBF0000ECE800FFFFAF00002B3B23DEEEAE0000ECE8";
    attribute INIT_2A of inst : label is "0140E5448602F4B9230EE46044AB14CF00FFFFAF00002B3B21DEFEAF0000ECE8";
    attribute INIT_2B of inst : label is "A05605E0ABBB1145BD800020BD8060A4BD8020A0BF804024BF900020A4116A69";
    attribute INIT_2C of inst : label is "BF2800023B08461A3B18441280FC22213B20687648FF31EAAA76E5BA7F885BE5";
    attribute INIT_2D of inst : label is "5B64BF8050648C81082B5B22C410E3A0D42188BD124008BF0200C25A82DCB823";
    attribute INIT_2E of inst : label is "6382028E524927B279E6B249659E49EE92692D9E59E79AC9259EE9669A6BA596";
    attribute INIT_2F of inst : label is "57864691625D1518D48986759570F9019477790186765109064BE60426C024F1";
    attribute INIT_30 of inst : label is "5C20115520C0618D764223051594CC09447599107C20145709817542215528D4";
    attribute INIT_31 of inst : label is "5E9524927B26F1499575744201D5424CC6385744429CD19523CC52BD40779511";
    attribute INIT_32 of inst : label is "950265FF89563B2FD4115691154864371549940266170649675269659A6B25DA";
    attribute INIT_33 of inst : label is "20C05740C2A5DD10D20C265EE516D524A70D05B888CE5740C298C058D158CC74";
    attribute INIT_34 of inst : label is "AB78461AFC02091E08035235E4B964B54965D68D8E26E0114074910177021095";
    attribute INIT_35 of inst : label is "384C10635AFF1558D457098140381E91256AE4564924BF4A2BFC430E9CC30D3A";
    attribute INIT_36 of inst : label is "084211E540E3991A4924AF34000225FF91E55D1520C864717C8AE40495A49278";
    attribute INIT_37 of inst : label is "91645DA449545691635148E284BF616458D74D389108A0515688DE91514E8457";
    attribute INIT_38 of inst : label is "7B52DE93AC242D8567809E0D278C9E7C182D4867309E4827349E9E91164884F4";
    attribute INIT_39 of inst : label is "50E740AA1D34514C1688180895815D1522C464714DBB9E2079419D14C4570941";
    attribute INIT_3A of inst : label is "6B0531975579509D3E55E99650E771FC028587490F050F150F550F55D4552996";
    attribute INIT_3B of inst : label is "41E50C25E7457976C83FCB2CF748445E928DE7554971C46094AC0F67C7005863";
    attribute INIT_3C of inst : label is "139D79518F2C92DF2C45D75C7951971D41F1C55E54E75F71B0E8BCB2C93D91D1";
    attribute INIT_3D of inst : label is "482600A8D54D15D1FD01BF4049674967486BC3E8A0281F6C91E255958D665479";
    attribute INIT_3E of inst : label is "7D3AAED60C9143BC405C383F237505A500A501A506A50BA50EB501F504F5BB44";
    attribute INIT_3F of inst : label is "E5BA891E661ACA4974BF261E89BB6982895EA418FF88430E223F03C428F14BA3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "1FD7300C191C0FC31DD40B833338177517350B831F961C9C303830301A340F49";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F9603211E9413D3";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF000000000000000000FF00FF00FF00FF00FF00FFFFFFFFFF";
    attribute INIT_03 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FFFFFFFFFF0FF00FF0BFFE7FFD";
    attribute INIT_04 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_05 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_06 of inst : label is "0761300C0C842F692EE82F691B3C033021302F6907632EEE30343A3A0F92252C";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0FC329380FC82B69";
    attribute INIT_08 of inst : label is "0C84272F0CC00CC00C0C2E2E0FD22DF80D85272D0FC32FE90F960FC300000000";
    attribute INIT_09 of inst : label is "0FC32F692FCF0FD32FFF0FC30C0C2E2E2DF01FF203032F6930303A3A0FC30FC3";
    attribute INIT_0A of inst : label is "2FC30FD70FC330140FC32F69303030300DD02F690FC31FF20FC32D7A0FC30CC0";
    attribute INIT_0B of inst : label is "7EBDBD7E3C6D229A184C4504584896445848450423312EEE0F0F30302F7D0FD7";
    attribute INIT_0C of inst : label is "77BFFDEEDFF5FFFF40018002FCBFEFFBFFFFFFFFDFF7FFFF400180025695A96A";
    attribute INIT_0D of inst : label is "341CEFFBCFF3CFF3E7DBDBE7796DB69EF96FDBE7E7DBEFFBDFF7FFFFFEDFFB7F";
    attribute INIT_0E of inst : label is "3FFC3FFCE96BD697D7D7EBEBDBE7E7DBF3CFF3CF7EBDBD7EDFF7382CFFFFFFFF";
    attribute INIT_0F of inst : label is "C7D3CBE3DFF7EFFB3FFC3FFCFC3FFC3FF3CFF3CFFFFC3FFF3FFFFFFCFBEFF7DF";
    attribute INIT_10 of inst : label is "CBE3C7D3D7D7EBEBF82FF41FB7DE7BED20089006382C341C3EBC3D7CC143C283";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFCFF3CFF3FFFFFFFFFFFFFFFFF7BFFDEF333FFCCCFCCC333F";
    attribute INIT_12 of inst : label is "4E607B7BE1A447DB48A68291A4E6A9289565666A555555A5FFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "3D05590FC264E87AA3BC6863292D06FB44CEF63BD2935A0F4164EF98EF68DE34";
    attribute INIT_14 of inst : label is "65640A68AC6A01A446C0868618CA4B41BED133BD8EF464CD6C3D0575A0F41560";
    attribute INIT_15 of inst : label is "66481443878EA468D683E054913F2292A479A86186186D850664014464004039";
    attribute INIT_16 of inst : label is "C05A0A449D1377A18E18C26480403878EA468D683F05483A7AA8292C7A18E1BC";
    attribute INIT_17 of inst : label is "3A469E8691AAEA916462A00A7AEF8A4281A33438D12829AA4BA82A91A3281643";
    attribute INIT_18 of inst : label is "A0E38A920E7B1E4A187C3F8E1B6C2FBEC792861F0FE3861B0BE38A92A4EB798E";
    attribute INIT_19 of inst : label is "8A03FBBB878033FC0E9A47A47AC68D643F054A0A4038E8944C691A68D683D054";
    attribute INIT_1A of inst : label is "AD0EB4FBAD3ED3E6262229358A43C2D82F03AE874F870F870F874FAA2E666935";
    attribute INIT_1B of inst : label is "0ABB8EB87BC7BC71C771C71EE8CC0CAB63AEEB4FB53E2F6C03ED4F9B4052A043";
    attribute INIT_1C of inst : label is "43C7BC7BC71C7BA30FB0F8A4B4FB53E2A03E292D3ED3E01C71EC0C71C7BA300E";
    attribute INIT_1D of inst : label is "A23BBBB878033E7BEEEBDEEEBE90BE90BCE6D06BB01F871C769AABBB8F64D58A";
    attribute INIT_1E of inst : label is "8C4B10E82A8A4A2ED61D13761235AAAAAAAAA6A6AEA2AAAAA68E82828A869622";
    attribute INIT_1F of inst : label is "3979DAA42825E75A5BC8936280499CDA3AA4FA0C19840040F166100511AA4734";
    attribute INIT_20 of inst : label is "21300203000000000C48C0800000000017BE340D6318F0FA69632DC1F0746241";
    attribute INIT_21 of inst : label is "3337333B00000000ACCCECCC0000000023231313000000004040808000000000";
    attribute INIT_22 of inst : label is "3327333B00000000D8CCECCC000000003137333B00000000D4CCECCC00000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000010002000000004000800000000000";
    attribute INIT_24 of inst : label is "33373F7FFFFF0313EFEBFEFCFFFFFFFFFFFE3333767CFFFF9C8CCCC8FDDDC4C0";
    attribute INIT_25 of inst : label is "3FBE00090323FFFF0103FFFFFFFFEECBFFFFFFFFFFFFFFFFFEFCECCCC8C0FFFF";
    attribute INIT_26 of inst : label is "C3F33FBCFFDC282350443D3CF7CDC4C000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "3CBF37CEFFD8CFF2DAF0E4CC4040A7FD32362333377F01119FFFCCCC0D9DCAF3";
    attribute INIT_28 of inst : label is "3FFF3FFF02020101FFFFFFFF888044403FB7033801237D78C000F0FBCF3EF8CE";
    attribute INIT_29 of inst : label is "FFFFFFFF02220111FFFFFFFF88804440FFFFFFFF02220111FFFFFFFF88804440";
    attribute INIT_2A of inst : label is "FF558F57E6BD56F7D5A5666A555555A5FFFFFFFF02220111FFFFFFFF88804440";
    attribute INIT_2B of inst : label is "0AF807640FB023CE0E0051450E00D14D0E0051450F00C10D0F0441050F7F6049";
    attribute INIT_2C of inst : label is "27408624706085147040851404E147076333C313F32ADFB0200C4CF0E6B3AF4C";
    attribute INIT_2D of inst : label is "E00D0F00C10D2D022883EA84D02207041801200E1041500E104006F400F89107";
    attribute INIT_2E of inst : label is "060310103CF34D0CE38E04D30E30E30338D38334D3CF38134D38230E30E04E38";
    attribute INIT_2F of inst : label is "0ECAC70FA039702C9CB0CAE30771BBB40C2FFBB40C2EC760D0C20EE12EEB2FFB";
    attribute INIT_30 of inst : label is "090A1AB00A98802DE3A0438BB0A49C9042E10352290A040EB085E02072700B9C";
    attribute INIT_31 of inst : label is "FC0F0C30F20CF7F00C2DE12061CB2039C8320E42442CD8300B98B20C4AE00B52";
    attribute INIT_32 of inst : label is "1C3C0FEFB0B4630F3C23B40CE0F38FE1C3E0386CCCE3D0D00CF4D38D38C2BEB3";
    attribute INIT_33 of inst : label is "08940E428428CFA6F2EC0CF24EF0272E270783BAB15E0E4A0434EBC8CBE89D2D";
    attribute INIT_34 of inst : label is "01F00E388EB670347058F00F2F030C09E88D32ACAC2C66C44AE10061E0A05070";
    attribute INIT_35 of inst : label is "12CC4106F20BC3F0A40E90C5C262348FC3F0CCF0C30C2DD04178051405C11760";
    attribute INIT_36 of inst : label is "82074C4DC80630B8CB0C813C84104FA08C8FDA30099C0F773BB84EE10F8CB2F0";
    attribute INIT_37 of inst : label is "0CCEE90FE233FC8C05E7C2823EFADD4FF03207B197712FB33B2D3C8CD3F8040E";
    attribute INIT_38 of inst : label is "F0F2BC0E0E2E4B1F0E203E8B0E2C3EBAB14BC20E283EC20E283EBC0FE3F23E92";
    attribute INIT_39 of inst : label is "CC0BFFAAE51C33EC3E0E30692C9BD83009980F5F0330BC845F340F3CA40E8005";
    attribute INIT_3A of inst : label is "CB83B2B2CFF3F12E41AA0CF4DC0BE74C08CFFDCB3D0F3D0F3D0F3E2E08AA0CF4";
    attribute INIT_3B of inst : label is "6E2FEF2C6DCFD8F1C42DC71EFAD03E7232AE8FCFC3F24EF8323C3F0F0112C087";
    attribute INIT_3C of inst : label is "310FDBF3871C78EF7C2CF8E5F3F3312F87B25BF03CCFC79472F41831E73E07D2";
    attribute INIT_3D of inst : label is "83AEFFA858C70FFFABFFAA7FE8CDE8CDE9F78332C292C71C62CEAAAADD3CF342";
    attribute INIT_3E of inst : label is "9A0332707F9F0F3FC74D013B0029FFAFFFAFF1AFF9AFFBAFF38FF40FFC0FC03F";
    attribute INIT_3F of inst : label is "0FA0B83C4CF092CB2F08D07EC301FB0638FC8E897810051484A7411063730128";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0110302404403FBC1554171605140BB01010373C0111377D1010353505411A96";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF05413E3E05443D3C";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF000000000000000000FF00FF00FF00FF00FF00FFFFFFFFFF";
    attribute INIT_03 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FFFFFFFFFF00000000782DBEBE";
    attribute INIT_04 of inst : label is "00FF00FF00FF00BF00FF00FF00BF00FF00FF00FF00BF00FF00FF00FF00FF00BB";
    attribute INIT_05 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_06 of inst : label is "3ABA2008377C0A822BA9020227702AAA3B3E02023B3C28283030202025690A82";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF3F3D02023C3C22A2";
    attribute INIT_08 of inst : label is "277B0A823FFE08803F3E08082DE90A82266808803FFC0A8225692AAA00000000";
    attribute INIT_09 of inst : label is "2F690A821FD72AA21FD72A820C0C08081EC628A8030302023A3A20201FD70A82";
    attribute INIT_0A of inst : label is "1FD72AAA0FD72A280FC30A823A3A20203D3C02022FF928A82F692AA22FE92AA8";
    attribute INIT_0B of inst : label is "87D24BE104BC11042C0051472C0071C72C0051473ABE28081B1E20201A962A28";
    attribute INIT_0C of inst : label is "EFFBDFF7AAAA5FF782824281D7C7CFF3FFFFFFFFEBEBDFF78282414183C243C1";
    attribute INIT_0D of inst : label is "6AA9D7D79AA665599EB66D79F7DFFBEF9FF6FD7FFEBFF7DFFBEFDFF7EFDBDBF7";
    attribute INIT_0E of inst : label is "C553CAA3EFFBDFF7EEBBDD77C7D3CBE3DBE7E7DB97D66BE9EBEB9556AAAA5555";
    attribute INIT_0F of inst : label is "EAABD557EBEBD7D795566AA9D697E96BDBE7E7DBE9CBD397F22FF44F9EB66D79";
    attribute INIT_10 of inst : label is "CFF3CFF3EBEBD7D7EFFBDFF77D7DBEBE9416682995566AA9F55FFAAF8AA24551";
    attribute INIT_11 of inst : label is "FFFFFFFFAAAA5555CFF3CFF3FFFFFFFFFFFFFFFF7FFBDFFEE77BDEE7EDDBDBB7";
    attribute INIT_12 of inst : label is "0FF0370701D8432F04410F62D8BBB62FC000151451101500FFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "03103C008400C70C73603618F6180D860D0D803611D43C008510D80CD80C0F47";
    attribute INIT_14 of inst : label is "18B4061887B2C1D870F0C361862D8603618303600D807520F0031883C00850F0";
    attribute INIT_15 of inst : label is "3B4041046063D81C0F003141D0000763D83CF41041041C9C72B4071CB4071C46";
    attribute INIT_16 of inst : label is "0103DD81E10000D0410403B4041046062D81C0F003141D1D887C760B0D041070";
    attribute INIT_17 of inst : label is "1D80C307603BC760370760009672FD4F60700C371CF72C1D83CF876070F40F00";
    attribute INIT_18 of inst : label is "D0D807600D82C31D04000C4107000C70B0C741000310410003100763D8BC0ED0";
    attribute INIT_19 of inst : label is "CC01CCCCC734B1CC0F6030C30C31C0F0001C1F1D80360760C7F60F1C0F000181";
    attribute INIT_1A of inst : label is "400D0072D41D41C440843D12CC41F7043303D4C787C787C787C787C000003D12";
    attribute INIT_1B of inst : label is "CD01CD0C75075071C701C71CD0F21CD00340B507521CFC3001F007EF003C4303";
    attribute INIT_1C of inst : label is "81C75075071C7343C7C873CB507521CF2E1CF2D41D41CF1C71F00071C7343E1C";
    attribute INIT_1D of inst : label is "010CCCCC734B1F3D33351333510351035337003CC030C71C73222222C7F472CC";
    attribute INIT_1E of inst : label is "8049125847DD8D37570700170003CFCFCFCFCBC7C3CFCBC7C3CFCFCBC7C3CB33";
    attribute INIT_1F of inst : label is "860601D8F41818CB2C0CF3D8C00F61C611D88601CAD0071C072B401C701D8004";
    attribute INIT_20 of inst : label is "12300103000000000C84C040000000006BBC38191204E934541212CA25F44243";
    attribute INIT_21 of inst : label is "33393337011102224CC4DCCC4440888010102020000000008888444400000000";
    attribute INIT_22 of inst : label is "311B333701110222E44CDCCC44408880322B333701110222E88CDCCC44408880";
    attribute INIT_23 of inst : label is "0002000100000000800040000000000002020101000000008080404000000000";
    attribute INIT_24 of inst : label is "333B1515FFFF0101FFFF757DFFFE5555FFFF3135B9995555ECCCDCC4EEEE4040";
    attribute INIT_25 of inst : label is "282812060202FFFF2222BFBFAAAAD5D5AAAAFFFFAAAAFFFFA8A8DCCC8080FFFF";
    attribute INIT_26 of inst : label is "C9F97C5CBFCC5415E0881454FBDE404000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "2C7E3BCDBBE4DBEDE5F0D8C8C0C05BFF333B13373BBB0101AAAFDCCC466E4555";
    attribute INIT_28 of inst : label is "3FFF3FFF1115222AFFFFFFFF5454A8A83D6B12370211BEA4E0085AB78F79F5C5";
    attribute INIT_29 of inst : label is "FFFFFFFF15152A2AFFFFFFFF5454A8A8FFFFFFFF15152A2AFFFFFFFF5454A8A8";
    attribute INIT_2A of inst : label is "101400564B2BA45E8000151451101500FFFFFFFF15152A2AFFFFFFFF5454A8A8";
    attribute INIT_2B of inst : label is "C78D20973761001019C0450658C035C258C045065BC005025BC0050240001455";
    attribute INIT_2C of inst : label is "6A345218658C5208658C5208C094825A573202D12695A8561C59915B95623591";
    attribute INIT_2D of inst : label is "11001BC0050248C0484306D38101963945000C1900058C590005138CC38570D2";
    attribute INIT_2E of inst : label is "D50350040830821C30821830C20830850810850010000C404104408100114100";
    attribute INIT_2F of inst : label is "4985921650246458494185921234442B0159842B015B9A469D02818E11CE12EC";
    attribute INIT_30 of inst : label is "140574240541011F93100740E44C4951C5931E3534065C496193935025A40549";
    attribute INIT_31 of inst : label is "89481041361184A3015B911017521004407149C11004F4640545012DC5901E34";
    attribute INIT_32 of inst : label is "7C2850DF6304563F4100083BBF2282AE9E00A898008C9D2152891491450678E7";
    attribute INIT_33 of inst : label is "054D49C5D100D21801BC5289838D3C135F00C473605149C1D104CE14DE044D5A";
    attribute INIT_34 of inst : label is "7D241208B42AA30474A085289268D00F34D3017D3D1055A1C5933D1793103464";
    attribute INIT_35 of inst : label is "5C88144105A69E004C4951908155003A9E31908104106F0535A8130CC4824813";
    attribute INIT_36 of inst : label is "5012B90084D56445041071281000105A7980B424054D4A10CA60038E48504134";
    attribute INIT_37 of inst : label is "3940854A02E6C039548A0080D16B9A8200A50C7268660A84E20E803920A41C49";
    attribute INIT_38 of inst : label is "B20100383C13964811500D44114C0D34E4960511140D0411100D003ABE21694C";
    attribute INIT_39 of inst : label is "8801EA55842CB3D40C3865865960B52407454A08C0324138F42B1A484C497150";
    attribute INIT_3A of inst : label is "0704147387147144240009979801D098048FA503E50FA50FA50FE40C15004997";
    attribute INIT_3B of inst : label is "88118E1051C71471D41DC71CF1222C01410CD187075C9DA43125663F5230100B";
    attribute INIT_3C of inst : label is "F1071471471C40CFA61C63CA147172C60B98A18D1C51CB1871E41431C43C0BC8";
    attribute INIT_3D of inst : label is "0211AA5442CB1E7954A9556A04520452156A52618171871C44FA00BFB52C66CC";
    attribute INIT_3E of inst : label is "960112482208C922455B11560153AA0AAA0AAD0AA60AA80AA70AAA0AA10A8C6A";
    attribute INIT_3F of inst : label is "905F634083817E165AC4B2CC920334D22340C148A94C1208536E034102C4C514";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
