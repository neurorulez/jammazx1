-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "54292AA049326940A502940A502940A502940A502940A5007E132429B203E993";
    attribute INIT_01 of inst : label is "089B026254A2AE108B0803128C0B5C8AA71389C4E271383A674CE99D33A674ED";
    attribute INIT_02 of inst : label is "9679A953D064EC6F8A80FDCADF32815B0B003001139C89625DEF667791EA3010";
    attribute INIT_03 of inst : label is "C72AEC03953CABE54F22F913C8BE55F22F913C8BE44F227D3A959F33CD4F679A";
    attribute INIT_04 of inst : label is "307C14072AEC72A6C72AEC72A6C4018CE338CE3272A6C72AEC72A6C72AEC72A6";
    attribute INIT_05 of inst : label is "6AA1766CA36423F423642564256456AC6B03B06185CCBF0DFF1E79F3F43E51E1";
    attribute INIT_06 of inst : label is "92A3BC2CB84296C31658B210B2694BB34A7B0C7D0C7D43E915365FE15E02FF01";
    attribute INIT_07 of inst : label is "E54F2E7957CA9665F8E5FB82955E061251424BB3DE432EC7790CBB7DE4F2ED77";
    attribute INIT_08 of inst : label is "B926CAE5F393B72760E4ED5C9D85E89F4FDE8F83D7F4B97BCB9E5DF2EF953CBB";
    attribute INIT_09 of inst : label is "89F4EC3E84C04AC8002118F468002F3014114B533652B54AB3D048B0E69A69A4";
    attribute INIT_0A of inst : label is "D964109F7A76A012B6649B2C96FD6FD026D9F6CB1CB4025440810AC5E893D1BC";
    attribute INIT_0B of inst : label is "24B92592C5064EBDFC8206B2CB93E6FAF5268A9C9B16591527DE8DB6044F7264";
    attribute INIT_0C of inst : label is "FCAABA6E75CF37DCB9A2607175DE7AB68292039320499405D99024DA0692B42D";
    attribute INIT_0D of inst : label is "680AD71CF9D79EB800D10AC64C9B3F385005A22A16EAFCDCF38F5F5B1B1D57EA";
    attribute INIT_0E of inst : label is "BAAAE9B7FD7F0A4215CCCDF3F1109D6E4B5C3AF3D85D150BEAEA22FE7E4EBCEB";
    attribute INIT_0F of inst : label is "11096805A78AF35C899D28FD251FB2431CE9927BD1BD2F9B9BBBBFFFFFBBBBDF";
    attribute INIT_10 of inst : label is "79E5ED16BCFE5FFA3FCC65D6280C8328B86210C4231780C6431FF181DCA20160";
    attribute INIT_11 of inst : label is "56CA6B563581EE1FFF0C0A18843108C5F20319C0C7FC6D2F3BB579E79E79E79E";
    attribute INIT_12 of inst : label is "5FF2ECE6A6AF5D237CF813C1BE44F2651C8D152793B258927E2761BED995B692";
    attribute INIT_13 of inst : label is "F515403E6D6D2185AC77CF7CF7CF7CF7CB4559FCBF5C2BDCABF5CF2EFD53CABF";
    attribute INIT_14 of inst : label is "3D27FFFFD80C79C1CBFCB9525CB95024907F52DCA9502C15CE7E59A6BF5B016F";
    attribute INIT_15 of inst : label is "186C4438B11DE7BCCE7301625EB5C0AD2782AD00B001D9E08920FF1050FB30FB";
    attribute INIT_16 of inst : label is "F3A1C3B079D0E1F83CE870ED1EF4387E8F7A1C3B47BD0E1FC6344018457A4FCF";
    attribute INIT_17 of inst : label is "9FB57FABD8DEAFF7BBDF0152FAB6FDC68399BBFFD9FFEED1EF470ED1EF4387E0";
    attribute INIT_18 of inst : label is "1A3956CA8C76D94758E19D4725D1C7B7E5627F5B7927FFAFEBFEA94BF59DE9F5";
    attribute INIT_19 of inst : label is "8DD0178976C641CD4BB4EA0752ECA2248B12E772D9173AD0A239CAF57ABC73C7";
    attribute INIT_1A of inst : label is "00380003A000380403A040380403A040398EC659DBE105182D50066E235C073A";
    attribute INIT_1B of inst : label is "BA12BA59090A420CF05444442AAAAAA9555555AA98EC65880003A020380203A0";
    attribute INIT_1C of inst : label is "000C0000B4828500885045DD77E6BBF75DFDAEFFD772264898202925901247D4";
    attribute INIT_1D of inst : label is "0010011F2E59C99E723F917CA9E4CA06CBB20000101001001044090028805502";
    attribute INIT_1E of inst : label is "98B122742154C01E4CF3977EAFE54F2650116BC6308421042126305E00005801";
    attribute INIT_1F of inst : label is "A92D58C078136EC048098713C1A60C60A02E029685AF1F3CD9330F24DAAB5BB8";
    attribute INIT_20 of inst : label is "57E0A88FC0F0A45F82A27940F13F13B13B13F1E301E04F5EB01EA4DBB0D58C07";
    attribute INIT_21 of inst : label is "C0917C1A89EF145050F00622883828881888A2031146036AFC113D05A2FC0A38";
    attribute INIT_22 of inst : label is "BC516143C01A8A2070A2206A20880C45182DABF844F4168BE028605F02A03B02";
    attribute INIT_23 of inst : label is "9C7799CE38A94A5294A5A3E20BEBD495090DD3DA8A27B6E2A8E29C35215005B5";
    attribute INIT_24 of inst : label is "55119A244669EBA8F154466D369B4DA74900D37E6F8D01400101F9B3C259C779";
    attribute INIT_25 of inst : label is "13A212C49D109A7A623C55109A044269E988F114427833E233C59F119A7AEA3C";
    attribute INIT_26 of inst : label is "0002AE002024242020000024A4A0A0DF9CAFF5F8000F2B793B63636362440758";
    attribute INIT_27 of inst : label is "BE2169001591455AC5FCAD1A27FAB07449EAC1AB6EFAA13AA5BEAC8E96E09C00";
    attribute INIT_28 of inst : label is "21174B472F2EA04845D3D9CBCBA8121176B632F2CA04845D1D2CDF1358005410";
    attribute INIT_29 of inst : label is "BCBAA129176B632F2CA80845D9DACBCBAA021176B43372EA80845D3D9CBCBAA0";
    attribute INIT_2A of inst : label is "563581FCBA8029574B632F2EA04855D3D1CDCBAA021576B672F2EA84A45DBD1C";
    attribute INIT_2B of inst : label is "581E88BFB457E7ED38793939392C6C453AED386D386D38446EF86D2D386D386B";
    attribute INIT_2C of inst : label is "0C9C9C9C9A044446EEEEC4445178421242BC40255A56D7ACF697DFD68CDFCF45";
    attribute INIT_2D of inst : label is "54840C9C9C9C94840C9C9C9C94840C9C9C9C94840C9C9C9C94840C9C9C9C9484";
    attribute INIT_2E of inst : label is "88CF3C0283590592097392822412ACB899601C399C00C82A620B0C82A4984AA5";
    attribute INIT_2F of inst : label is "004483A6524CC00D8641AE49C94004483E49E65600644941AA6350468300AA49";
    attribute INIT_30 of inst : label is "2416CB654020064B244E1D05CF339001700F3C018724F6497CCE00741AE49C94";
    attribute INIT_31 of inst : label is "D37C9BF4DF99C4C212BB1209405C9622420B4B1B424C04A40504B4812A18AC48";
    attribute INIT_32 of inst : label is "C010BF7A010217EFC4A96E93F1AD6358D6318C635AD631AC7FE72EF972807A3F";
    attribute INIT_33 of inst : label is "E318D6B1AC6358D6B1F8102FDC83060103D76186197AF000102FDC830681EBB0";
    attribute INIT_34 of inst : label is "C71C73CDC0BDCB817B99579A134641E22F33FE0010108A865099404039AC48FF";
    attribute INIT_35 of inst : label is "A27BF982D2E0ADA44FF301FEF4AD694A33DF1CF3C73CF3CF1C71CF1C73CF3C73";
    attribute INIT_36 of inst : label is "40F503D40D50334DCED704CA2AA80AA07A80AA07A80AA07A80AA06A81AA07B13";
    attribute INIT_37 of inst : label is "6505D075407507D41F507D41D5075405503D407501D4075015405503540F503D";
    attribute INIT_38 of inst : label is "0D503503503503503D40D40D503503D40D40D501501D40D405501D40CF4CE2AA";
    attribute INIT_39 of inst : label is "0D648575844825B79291454A00880000088008095015407503503503503503D4";
    attribute INIT_3A of inst : label is "99A26082E9380749815A24A6880BA5C5444007499966882E972B0B41F55AB1AC";
    attribute INIT_3B of inst : label is "5BF69777C3E24EC9ABCD8F6F6F8C378F6BDC1656EBD904D14EC4239D12C2F640";
    attribute INIT_3C of inst : label is "6B5E1BFD57ACFF86CE9E74F3920DF37679BAEFC7A697E55FCF5C3EC3374D5F9F";
    attribute INIT_3D of inst : label is "F893332FC242F912EFF60F5C8A0F00000000000000003AA738E72739CE73A78F";
    attribute INIT_3E of inst : label is "2C0E5CF7FD4AC231854E9C0530A9C391D02FEBB0F61C7196250A5D6A414F9431";
    attribute INIT_3F of inst : label is "DE0F0634000602489B44F7B5979B39AD0DC59D0875B5135DAB2F444E29B4ADBB";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "03F2E01E8666A5D997665D997665D997665D997665D99764C0034CB1865F9187";
    attribute INIT_01 of inst : label is "64732666DA46F64D9D2B3727FCD862EEEC7E3B1F8EC7E3284D08A1342284D09C";
    attribute INIT_02 of inst : label is "077D905D1A61BC80178276150086AA333822F2CD9EB19AD68779CECE7B067639";
    attribute INIT_03 of inst : label is "D85C0D982E41700B805C82E41700B905C82E41700B805C86E43800BBEC8477D9";
    attribute INIT_04 of inst : label is "11AB2E585C8D85C8D85C0D85C0DD97C0701C070085C8D85C0D85C0D85C8D85C8";
    attribute INIT_05 of inst : label is "23E583400A008A908A008E008E00E6205324B2ED8FF89D40E820820C089B74F3";
    attribute INIT_06 of inst : label is "6C0A4080296624088484244424B0025ED8B22236223611B02F463FE9809C0F46";
    attribute INIT_07 of inst : label is "4E0274138095009C2C1C241DA3C1595E9B50B4D86890413886E34DA689041288";
    attribute INIT_08 of inst : label is "22CB2E2C246C00DC2C1B04C370921701B80360B06812C2843500A905402A09C2";
    attribute INIT_09 of inst : label is "440A90F1D69BD1A5F6C5991A01BAB184BC48DA39A035AFD78D7AD5831B25B383";
    attribute INIT_0A of inst : label is "884967A5854036B5A48B2CBFB23622459200BCD82426DE8F2D162EC815006843";
    attribute INIT_0B of inst : label is "6B0B5BB50E60DA634B259D76B5B49C0502E84D816C821259E9614016CED744B6";
    attribute INIT_0C of inst : label is "692AEF9013D71D61501685F2DC2585404BB527A44B22DF27D22D93679135AE1C";
    attribute INIT_0D of inst : label is "EEAC8E296B24005B970A2D2C31E1880972FA14776BBC692C40B66662222002BC";
    attribute INIT_0E of inst : label is "8CABBE45FCFF2F2F26C48525AFAA67871238E48028A338942D194714B4192005";
    attribute INIT_0F of inst : label is "C8DAC1120793F4391A9162243C46D6ABBFF8B69CA61A5664464642020202020F";
    attribute INIT_10 of inst : label is "94594AEE8B60A82D402127F339201819A1EC53DC8F71C3DFEB7FF6E70033664C";
    attribute INIT_11 of inst : label is "0406B3102992A64858AE3C7B14F723DC070F7E1ADFFDB040780F945945945945";
    attribute INIT_12 of inst : label is "A805484B41C700495113A09404E02741A3529A686A5682049E465C4E844105B5";
    attribute INIT_13 of inst : label is "0871ECC4F2259397BCA8A2CB28A2CB28A2BB04C150719E23700E805506803521";
    attribute INIT_14 of inst : label is "0A43FFFF051CFE929BFAD3695AD36995C8FF695AC36995481089D2C020882C40";
    attribute INIT_15 of inst : label is "60A48AC11226EC5D08620B037AF6D9BD93064D85809782111C91FF4962700270";
    attribute INIT_16 of inst : label is "64854A07B242A503D9215290EC10A948760854A03B042A500F3C893CCF0AE080";
    attribute INIT_17 of inst : label is "4196AD15517CD5AAAFAA5543BE9F46F91A5025BFF25FEB1EC915291EC90A948F";
    attribute INIT_18 of inst : label is "9805844CCC0F8980B4D6060085E02DEAFF850006D40C05F5C0F7E295403F12B6";
    attribute INIT_19 of inst : label is "01E01204D3854612A69CF12785A1250248234D32890ABC4803402C86C3600920";
    attribute INIT_1A of inst : label is "203A00038000380603A0403A060380403B0C670C79C0020074A0054D001A41B6";
    attribute INIT_1B of inst : label is "73370036F6A3EFB9803AFAFA866666666666663320C670D202038020380003A0";
    attribute INIT_1C of inst : label is "3F9DF792355FDF5E3FF1EFB600D300698032C019600760C1884647836F6FE30F";
    attribute INIT_1D of inst : label is "9E69A7C180A2962485C06C49724B9530604492493A79E69A79AAFEF15CE9F73F";
    attribute INIT_1E of inst : label is "4862C4A0B7FD4934B1242C03724B925CA939C61FF18C633CB747F370DB6DE9A7";
    attribute INIT_1F of inst : label is "7A5FBF4BD5A4EECD2DEF786C37FDFDEAEAD0545B9DFFBBF300BC15589F01F909";
    attribute INIT_20 of inst : label is "E51E577C7F1FD2947B5EE7BD1F71F77F77F71A3D6F5C91A3D6F5493BB3EBD4BD";
    attribute INIT_21 of inst : label is "FD5A52E57B9C4B96BD2BEA5C55CB5457AB72DCF56E28F405C4AB4BFA14A3C5DF";
    attribute INIT_22 of inst : label is "712E5AA4BFAB7355ED735EADC973D5B9A3F01712B92BE8D29717BF94BF5EF7FD";
    attribute INIT_23 of inst : label is "2B1AC2B08F77C6318C635684DF60A33F3A7CAF50A5CE94295FC55EB6B5F3EF02";
    attribute INIT_24 of inst : label is "8AAE77DAB9C254F12E6AB9C080402010C61208091938258B122424629682B1AC";
    attribute INIT_25 of inst : label is "FF75FFFBFBAFF297FD4A8AAFF7FABFCA5FF52A2ABFCF4F15CE7E78AE70953C4B";
    attribute INIT_26 of inst : label is "0020DC8014101014140000141410103921700B11249ADC96E5EBEBEBEA266BBF";
    attribute INIT_27 of inst : label is "E8CFC492E15BAA210ABBF5AA4AEFC6B8959F4A8D9DC3124316DBF757BB753800";
    attribute INIT_28 of inst : label is "F68195B0D0405EBFA06467341017BF681B198D0405EBFA0656F30066E0002E6F";
    attribute INIT_29 of inst : label is "41017AF6819198D0405EBDA06567341017AF681B5BCC0405EBDA06C6D341017A";
    attribute INIT_2A of inst : label is "10299281017AF681B59CD0405EFDA06C6D301017BFE81B5B0D0405EBDA0646F3";
    attribute INIT_2B of inst : label is "BC7FCD688701003B913B913B913AC53B912F906EC47AC52F907B912F906F9073";
    attribute INIT_2C of inst : label is "08B8B8B8B7AFAFA8505005050FC5EB2BCC09FFDFF739AD01000035AD922AFFE6";
    attribute INIT_2D of inst : label is "609008B8B8B8B09008B8B8B8B09008B8B8B8B09008B8B8B8B09008B8B8B8B090";
    attribute INIT_2E of inst : label is "6044B5B4403ACBC920B8C99E92417BE6410DA718833C0489E124C0489E782CC6";
    attribute INIT_2F of inst : label is "F3D248DFCB2D7BE66124173C64CF3D248D75E20CFBD09A65338B7BF6CA69172C";
    attribute INIT_30 of inst : label is "493FFDB6DB492FFDB7C18491AF10E7DE3696BCB0614D4BBEB4419E124173C64C";
    attribute INIT_31 of inst : label is "2C09524A8046FD2D3B57B7E5E5AF59CFAFE6E6BE97D7D67ECAFB4F5BF4AF77DB";
    attribute INIT_32 of inst : label is "7E7EFF85FFFFFFF27FFFEFEC00200840008000080200802000485C87C4F687C0";
    attribute INIT_33 of inst : label is "00400000200000108007DFFFE3FDF9FFFFD8BEFBEFFB0FFFDFFFE3FDF9FFEC5F";
    attribute INIT_34 of inst : label is "0D30D3401DF7B03BAD6AAA457AA0AAB5508400DB7DFB559CB87AC1E60050F400";
    attribute INIT_35 of inst : label is "71325E5281F93C4B22E6706420080200A99D30C30C34D34D30C34C30C30D30D3";
    attribute INIT_36 of inst : label is "AE0EB83AE2EB8A12F680CE4D1475C5D7075C5D7075C4D7075D0D7035C0D71952";
    attribute INIT_37 of inst : label is "5EB8EBABAE0EBA3AE8EBA3AEAEBABAE2EB83AE0EB83AE0EB8BAE2EB8BAE0EB83";
    attribute INIT_38 of inst : label is "E2EB86B8EB8EB86BA3AEBAEA6B86B83AE3AE26BA6B83AE3AE26B81AEA6E491C3";
    attribute INIT_39 of inst : label is "97540638E78F3976DA1964D80808000008080000EB83AE8EB8EB8EB8EB8EB89A";
    attribute INIT_3A of inst : label is "60739B011F2008FD83070B6BC60C7F84B45818FF9210B011FE024000BB98814C";
    attribute INIT_3B of inst : label is "FC7ED646ED87D4B8AA665FCD24BD7FD285B1C83260BCAA1E09452311E2A6FB51";
    attribute INIT_3C of inst : label is "04348007991C96205DBAEDD7780B8F8F49A34DBFACFA7648CDFBA2097ACDED55";
    attribute INIT_3D of inst : label is "4E045ADAE76FEFEBFBBE3F88A2AF00000000000000001FED75AEF16B5AD76E9B";
    attribute INIT_3E of inst : label is "4034AB0A1234248530AD56C0E7178EED743DC67BD394669A8C09C8316301AD2B";
    attribute INIT_3F of inst : label is "8822A5CC870E2A1C6135C8F8390A43E752CC873E99F93D2136361C64822890AE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "55E6CAAE3745B376CDDB376CDDB376CDDB376CDDB376CDD87C090CE4A6729C86";
    attribute INIT_01 of inst : label is "932A05409324A8614A9B821508568AF135D2E976BB5D2E5BA3746EADD5BA3751";
    attribute INIT_02 of inst : label is "C451384B0321E8628501B7F40EF4381A1699A7BB773D56F58A50A8B5A2FA68D3";
    attribute INIT_03 of inst : label is "B7D0AB33EA1F40FA87D0BEA5F42EA87D4BE85F52FA17503AA4A80EA289E24513";
    attribute INIT_04 of inst : label is "001D0A77D0AB7D0AB7D0AB7D0AB11C1C0701C070FD02B7D02B7D02B7D0AB7D0A";
    attribute INIT_05 of inst : label is "5462275B2A002A902A002A902E0025C142F220AD26FA0AE1A30EBF76ED9A7051";
    attribute INIT_06 of inst : label is "DB2AD821018AA482A915481500C454092A000AA40EA454070AD4D54A50A68ADB";
    attribute INIT_07 of inst : label is "BA25D52E89756E8B7D8B748B61B060658210C920DA45B6D24926DB4936924936";
    attribute INIT_08 of inst : label is "FD249BCB7FE857D0A4FA949F529DD52FA85F4093E8133EA1F50EA87D03EA5744";
    attribute INIT_09 of inst : label is "40EA91AE9874B6BA332650EA84C4CEF42AF7561BADAD6AB56B28B561E6D3497E";
    attribute INIT_0A of inst : label is "5849DD6EFD03842D6BF4926A5692692646A4A816019DA5B5D3B93085D40BAA1D";
    attribute INIT_0B of inst : label is "5ADAD6ADC7C035D2DDA60A45A8ADDA75405BC13E923600775BBF40E5A8B0BA4C";
    attribute INIT_0C of inst : label is "D9803EDA2828EBBF50E5A728CB3EF543CEAD307BA239327C3DD11C913C2D68B4";
    attribute INIT_0D of inst : label is "D331F3DE9592EAF419F7C7E03873A2C9931FEF9D7D96D9DE116333377777FD16";
    attribute INIT_0E of inst : label is "9000FB6FAB6AD3D3C1C2007A4ABF72ED1FCF325D71FECF3FC7F6F9EF482C974F";
    attribute INIT_0F of inst : label is "A616A4C1BD3407825624AA9215524583AE742596D41D5733311331133113315A";
    attribute INIT_10 of inst : label is "9A620CD4282FA15753BD21234C664915635A56B09AC406B782DAA74831EE983B";
    attribute INIT_11 of inst : label is "51A592E0A179084B5BA226D615AC26B1545ADF50B6A9D5DD4AAE9A61869A6186";
    attribute INIT_12 of inst : label is "A17D40EB536C110B05AEE9774BBB5D903D50025BA805BAECE0415831A014692C";
    attribute INIT_13 of inst : label is "CD8B333EC344CD494A34D30C30C34D34D435425F409A4B3D42EA97543E81F42F";
    attribute INIT_14 of inst : label is "00419249950A21F155533B9CAB3B9CCA60AA9CAB2B9CCA615A9DB311EAD1311B";
    attribute INIT_15 of inst : label is "508E62A13981EA3DA94B02C6DBACF4EB43132B01624DBBD12F29AA7180D480D0";
    attribute INIT_16 of inst : label is "F5A4D9D1FAD26CC8FD6936757E349B32BF1A4D995F8D26CEA41C211C0AC0F005";
    attribute INIT_17 of inst : label is "36E7B3BDBBA6767B74EC1003AB92BEADA94B7EEA9F754D97E3536657E349B3A3";
    attribute INIT_18 of inst : label is "3A49D3AE9C9275C92A55A1A90C52467B1A86D8DB1908F6561B1952D98DA09BC7";
    attribute INIT_19 of inst : label is "1051E4472B0584DD39582A714D57E1FC639FA486773B0A0A9B5A4EB75B8C9129";
    attribute INIT_1A of inst : label is "403C0603C0403E0403C0403C0603C0603D9963AE7460010839C00585040A0814";
    attribute INIT_1B of inst : label is "3B97CAB4D360AED16005005541E1E1E07878783C09963AC60603E0403E0603C0";
    attribute INIT_1C of inst : label is "736CEE1C20195D699C9B99F599FACCF9667EB33E5994D2A540E4EE2B6DB4C3CD";
    attribute INIT_1D of inst : label is "69A69B0EAAB77E6AF5C3AE57F6BF1482AAE5EDB6DDA69A69B6D8EF4D90B09512";
    attribute INIT_1E of inst : label is "E53970D0266B0EDBF357EE1F72BFB5F8A4D8B52724A5299026C52929249266DA";
    attribute INIT_1F of inst : label is "E360C1DA7C36AAA4298A6772B8431083031FBF8D9E9AB46EB5D0DA2EEE75B9B4";
    attribute INIT_20 of inst : label is "73461C5A118466CD1872D4A5896896896896870729F2D870729F2DAAA81C3DA7";
    attribute INIT_21 of inst : label is "138B3569CB5A1E6CE1F88EF2D9867ADA3BC87246386E4EB3B33C7F273668C702";
    attribute INIT_22 of inst : label is "6879B3D7E239C96619C968EF23C918E0B91ACECCF5F89C59AB1C49CD58706846";
    attribute INIT_23 of inst : label is "F5FD7F5FFECEA5294A52C5065695F6763230F6C3878DB0E1E5A5D6858D230A59";
    attribute INIT_24 of inst : label is "1E382518E0ABF03DF838E0964B2592C8A53D64B5BAB6070E183AD6E955BF5FD7";
    attribute INIT_25 of inst : label is "C68714263438A8FE0E7E1E382518E0A3F839F878E084C68714223438AAFC0F7E";
    attribute INIT_26 of inst : label is "A8347A800080908090800014849080B6BD70FB16DB6DFDAFC490909090722FC4";
    attribute INIT_27 of inst : label is "D99ABB6DB562DCF3CFDFF8B8FF7FE2F1F9FF9BA6DBA1B7E1B37DFCDC8DCDB6AA";
    attribute INIT_28 of inst : label is "C60E96F5BAB74F3383ACB76EADD3DCE0EB2D9BAB74F7183ADB66E8CDD820B676";
    attribute INIT_29 of inst : label is "EADD3DC60EB2D9BAB74F7183A5B66EADD3DC60EB6DDBAB74F7183A5BD6EADD3D";
    attribute INIT_2A of inst : label is "E0A17982DD3CCE0EB6DDBAB74F7383ADB56EADD3DC60E96F5BAB74F7183A4BF6";
    attribute INIT_2B of inst : label is "E06561DA375743D1110444451045104510504511110444504505105045104512";
    attribute INIT_2C of inst : label is "0909090906C550005500055009B68E8A86EE9369B5A96A219088D24F3DD912B0";
    attribute INIT_2D of inst : label is "9120090909090120090909090120090909090120090909090120090909090120";
    attribute INIT_2E of inst : label is "044550005814D300440E00E7008815500A00075083CF211EBA48F211EAAE2F37";
    attribute INIT_2F of inst : label is "3CE010A271C634D0780801C70073CE010A38820734E2400081C014C001240155";
    attribute INIT_30 of inst : label is "000A492580001A4925C1E023441079E782451126782071C71841E780801C7007";
    attribute INIT_31 of inst : label is "F815E4BF277E585A0AC8686828649249696020680D058414865AC230AC6B0080";
    attribute INIT_32 of inst : label is "3F7FFDFFFFFFFFFFFFFFD93C00000800100000004010840000AF703F80B4F703";
    attribute INIT_33 of inst : label is "00000000000842008007FFFFFFFDFFFFFFDFBC71E7FBFFFFFFFFFFFDFFFFEFDF";
    attribute INIT_34 of inst : label is "68A68A25D66B7BACD6EA657C72C1777B9EF401249E671648C9AB26A7EEE27B08";
    attribute INIT_35 of inst : label is "E0ED23E8529B7EFC1CD128998D6B58D60648A69A69A28A28A69A29A69A68A68A";
    attribute INIT_36 of inst : label is "7C15F057C15F0559BC564DC3116F82BE0AF92BE0AF83BE0AF97BE5EF97BE1FF0";
    attribute INIT_37 of inst : label is "F5F25F057C15F057C15F057C15F057C15F057C15F057C15F057C15F057C95F05";
    attribute INIT_38 of inst : label is "C9DF0DF25F05F0DF257C97C9DF2DF257C17C9DF2DF057C97C1DF077C1CFC3197";
    attribute INIT_39 of inst : label is "CC52084542012491060820860088000008800808DF2F7C95F25F25F05F05F077";
    attribute INIT_3A of inst : label is "59237200DC0C06E2069AA79EAE0B71428B5416E28CA0A82DC41CB1460C97050B";
    attribute INIT_3B of inst : label is "0C7A24103910D0163918A871C964BDDCBC5401408699A40E64B2D8E060215050";
    attribute INIT_3C of inst : label is "12808C12B445A4A3663331912816F0B2A002303950080CA0B40A0032D8A6E07C";
    attribute INIT_3D of inst : label is "9375B25FD04603104C55A7F0B16000000000000000000CCD99A251236CD98CDE";
    attribute INIT_3E of inst : label is "2A29D5C5D5C343830815A4B120108083C90612C8AB2CDC30120184809EBC4C92";
    attribute INIT_3F of inst : label is "D841423271E5C78B348CE63DBFDCD8522FCE470473A3C583CFC7886608AAB10A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "BC5325E299DC64C993264C9976EDDBB76EDDBB3264C99324F80B28B594586D93";
    attribute INIT_01 of inst : label is "264E20C40A70694A1A352A3828A13DE65A2D169B4DA6D3502A0542A8550AA154";
    attribute INIT_02 of inst : label is "10820150CB6488A597B3FC0480A6A33E31766E64CA0331484802108866062225";
    attribute INIT_03 of inst : label is "181291980B404A025016809404A02401680B404A02D0160095A810A4900B4920";
    attribute INIT_04 of inst : label is "11012D581291812918129181291D562A8AA288A2012998129981299812998129";
    attribute INIT_05 of inst : label is "8944FF00E804E84CE84CEA04EA04883E008883DC1B33E447A324D3AF4D9AFF23";
    attribute INIT_06 of inst : label is "27EA04E0352780CE84F402750293D2EDBE013A133A01D40C2E2D755DAFDD7A66";
    attribute INIT_07 of inst : label is "43C21E10F08784A885288610138A4A4C4B53124D6D9A5975966965F259EDB7C9";
    attribute INIT_08 of inst : label is "42492F1884094012960252C05A560580240048580B0A40B004A02C0160090878";
    attribute INIT_09 of inst : label is "4802C6A0921B89849A54F102D29090A4815DA13F8042100D10810B120B2CB751";
    attribute INIT_0A of inst : label is "3805771081601462190924BB7E13E135BE13A9312106DC4C24D2A78804800B40";
    attribute INIT_0B of inst : label is "846420420A65D50C6134908852E21181214445B124AE015DC420580C7988C496";
    attribute INIT_0C of inst : label is "455524105230C0204A0C75A628A081202BE3AC6C4AB25AB63625592559E212C4";
    attribute INIT_0D of inst : label is "44248A2DB5B69A11D28A2484D42782252A4914502AE9455C4292222222228069";
    attribute INIT_0E of inst : label is "25549040A8AA252535D69C36C540A5145228B6D32892289244914526DCEDB4C0";
    attribute INIT_0F of inst : label is "DDB11BB25D1BF569B198FA131F426C673DEB6056103D0E6666666644444466AA";
    attribute INIT_10 of inst : label is "9249888668102C2168293E4218A8BA2610C5618AC62EB9899E2AAF66993B760E";
    attribute INIT_11 of inst : label is "309C441F00443A68582560315862B18B8EE626378AABD2407878124924924924";
    attribute INIT_12 of inst : label is "2501625C0494E30F0910908484242120A05A0AC40B4C53A65E670A4E980C2722";
    attribute INIT_13 of inst : label is "5A6C2EE5C69AB53401A08208208208208321C2205A6DB9204802401280B004A0";
    attribute INIT_14 of inst : label is "280249250599A48211FAD36B8AD76AB85CFF6B8AD76AB85830810A4C30A7AF0D";
    attribute INIT_15 of inst : label is "06F99A0DE66DC638000A8A293242CB90BB6CD0C515B312191495AAC923D023D0";
    attribute INIT_16 of inst : label is "0348202281A4103140D20808A069040C50348206281A41011CC89F24CA2ACD9D";
    attribute INIT_17 of inst : label is "254AC506107418AC2EB114114172D0A9000034EA9A754D0A0680808A069040C5";
    attribute INIT_18 of inst : label is "000000000000000000000000200008AC4D4494921309A8A892E2B690293F1212";
    attribute INIT_19 of inst : label is "8001E00000600000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "4002040020400204002040020400204000000000007DFFFF8000002020404080";
    attribute INIT_1B of inst : label is "5D6D9E072CAA4362140000000000000000000000000000020400204002040020";
    attribute INIT_1C of inst : label is "AD9BBB52A4BA8637537D768C324639231C938E49C721C49931DDFCE072492532";
    attribute INIT_1D of inst : label is "B6DB6DC4E018848181600B485842C131382212DB76596DB6DB748DB8EEDB666F";
    attribute INIT_1E of inst : label is "00000001B4C0A934240C09004A42C216093E08CCA94AD669B42CA2064B6DD165";
    attribute INIT_1F of inst : label is "9338B12CD932B108B1321248641054A2626A4647DB9AA74B0000000000000000";
    attribute INIT_20 of inst : label is "A927918385614AE49C4718C5C30C30E30E30C284B364CC284B364CAC438B12CD";
    attribute INIT_21 of inst : label is "052B93791C5228CC89B22B475C644558A5194614A2AC14073B226C8AD724D460";
    attribute INIT_22 of inst : label is "48A32226C8AD1D71D11562946518528AB0501CE889B22B5C9B51C2A4DE470C15";
    attribute INIT_23 of inst : label is "21485210A41E8C6339CC20F5B4F4EBF2BABCCCA65259C9949925B6C8E73A7A03";
    attribute INIT_24 of inst : label is "AB23245C8CA36611B2AC8C80B0582C1688F60981DC6195AB57AE075C10521485";
    attribute INIT_25 of inst : label is "70E4758B8723A8D9C46CAB23A45C8EA36711B2AC8EA160C4750B0623A8D9846C";
    attribute INIT_26 of inst : label is "00007280151919191900001D191D0D24605802C16DBA1690B531313130AAACF1";
    attribute INIT_27 of inst : label is "8CCD44926ACA7631ABCF5EB34F3D6AE6D4F5EB14D3075147514F5C5ECD65A400";
    attribute INIT_28 of inst : label is "9499F91AD4DBB4A52E5F47B536AD294B9D91ED4DAB4A5265747B716530101E5B";
    attribute INIT_29 of inst : label is "536AD29499F91ED4DAB4A52E5747B536AD294B9FD1ADCDAB4A5265E47B536ED2";
    attribute INIT_2A of inst : label is "1F0044036AD294B9FD1AD4DAB4A5265E47B736ED29499F91AD4DBB4A5265F47B";
    attribute INIT_2B of inst : label is "91FEE126FBFC2054141414001555401540001541415540014140155414014144";
    attribute INIT_2C of inst : label is "000080808360000000000000030B6B6BDD516DB38C6339E14DA47CDF57671F70";
    attribute INIT_2D of inst : label is "1000000080000100018101810100000181000100010101810100008000808100";
    attribute INIT_2E of inst : label is "05DC14020110410804080882100810404020110BB104201828044201820AC020";
    attribute INIT_2F of inst : label is "10420182C105104221008104044104201820AEC4104201008101104201008104";
    attribute INIT_30 of inst : label is "5B2B65B2B2592B2592D8840305762082100C14022100C10415D8821008104044";
    attribute INIT_31 of inst : label is "0F086A43405229696B4DADA4A4A25B4DA4ADA4A49492B6D6DA694AD295AD16B6";
    attribute INIT_32 of inst : label is "00000000000000000000000000000000000000000000000000181E80D4D681E0";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "6DA4DA6491084922108DD873CB250A1850A400DB694AD3BC7651D9573FB1EF80";
    attribute INIT_35 of inst : label is "042090378C0D04000000024001080200012936DB4DA4934D36936DA69B6DA492";
    attribute INIT_36 of inst : label is "2080820208082230278C40000004001040410104040010404101040400104104";
    attribute INIT_37 of inst : label is "0082080020808002000800200080020808202080820208082020808202000820";
    attribute INIT_38 of inst : label is "0008208008208208202002080800800208200082082020020808002004200001";
    attribute INIT_39 of inst : label is "2000008000410208020000008800088008808080082020808008008208208202";
    attribute INIT_3A of inst : label is "86040181022C0815F84F1019C6040BF83A0C0815605690102AC0FF382620F802";
    attribute INIT_3B of inst : label is "C1092CAA105009420148A4304120000012C1942852C0AAD7EFE7D3E9F6BD9A51";
    attribute INIT_3C of inst : label is "1ADE907D26459BA4668A2451160042049251B21AC968C5B1B6425D5005B6100E";
    attribute INIT_3D of inst : label is "8001000008084400501117B0FCBA0000000000000000132111A22D685A19A299";
    attribute INIT_3E of inst : label is "00014040000000002040840100081080404502028000400448D0824480000040";
    attribute INIT_3F of inst : label is "30D04110081010200813401248220204001004210012100820243001A6820020";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "80583C034014AD5AB122448956AD5AB122448956AD5AB122960D1896AC4876C1";
    attribute INIT_01 of inst : label is "6EC0BC57AAED485932716AB402C250E890080412090080A0540A83506A054097";
    attribute INIT_02 of inst : label is "04101018EBB0028AD7EBB58738E724AAB232C6EDDC7012D08240018840CC266F";
    attribute INIT_03 of inst : label is "9E18C99B4C7A73D31E9CF4E7A63D31E9C74C3A61D38E9870E32888A080830001";
    attribute INIT_04 of inst : label is "9D51AC5E1849E1849E1841E1841D172A4A02A0A0E18C9E18C9E18C1E18C1E18C";
    attribute INIT_05 of inst : label is "B3154B044AB2C86AC8B2CA22CA22807D1C548374099AE942ACA49224591A774A";
    attribute INIT_06 of inst : label is "0B4A22C0C165032DA2251165111A93CC948CB288B2889444AE453554694F4A2F";
    attribute INIT_07 of inst : label is "939C9CE4E3271CA1472147582A125A58AB980416080880110432084092C10502";
    attribute INIT_08 of inst : label is "42492D21470E6E18C5C318F87313A63C39B863170E62F0C7A73D38E9874E3273";
    attribute INIT_09 of inst : label is "73D38A8C1689132DAAE5C5C39AB4B8E6A8DD92BD82052A102804102B892DB2D9";
    attribute INIT_0A of inst : label is "A8693228E18E57042D0924B32A1AA085BA082812A82248996D572EABA73F0E78";
    attribute INIT_0B of inst : label is "4A625085A800CB081164D010900510698C0A75E1248A084C8A387384C0128496";
    attribute INIT_0C of inst : label is "01D5305E24A28A3A73808486A948E1CE09042D4C4E725A36A6273925190429D2";
    attribute INIT_0D of inst : label is "0524DB6DBDB68A21929B763A1BB58C09326D36DA2017098C3123B33333B02A97";
    attribute INIT_0E of inst : label is "0554C16DA9EA64646AC94736E4153AF09B6DB6D134C26DD806136D86DA2DB442";
    attribute INIT_0F of inst : label is "5DC203BCD858096C42C25208DA4350B629480082E75E47000000220002220060";
    attribute INIT_10 of inst : label is "618512CB88EC38C386392E84B6701C112DCE6B9CCE776398F26AAB5640197646";
    attribute INIT_11 of inst : label is "A0C0803E8E2A2C6C5C7871739AE73399C58E631C9AAAD6644E08238E38E38E38";
    attribute INIT_12 of inst : label is "38E9C7CC0031360D15E4E72F3938C9C6B861EB4B0E30B33000688A80D0683005";
    attribute INIT_13 of inst : label is "2E7A2EDCFBA5BC3D41C71C71C71C71C71AB283D87341B4BA61C30E1874E3A71C";
    attribute INIT_14 of inst : label is "01019248A351EF2B9952B34BCAB34DBCDAAA4BCAB34DBC5F18D1146A29EC2E0B";
    attribute INIT_15 of inst : label is "CCC0C9998322E8DD91C4E84B62C6D9319BE441F42496331D1191AA996B510B51";
    attribute INIT_16 of inst : label is "CDD4E11AE6EA70AD73753856B9BA9C2B5CDD4E11AE6EA70898429EA2EA4C8040";
    attribute INIT_17 of inst : label is "3663A18D18A6343A34E8BAAAABCD3724C14C36EA9B754DAB9B93846B9BA9C235";
    attribute INIT_18 of inst : label is "B3941C20592D841296024A32AB24AC3A2A86D8DBDE4E54545B11524F0DAAC983";
    attribute INIT_19 of inst : label is "A5201802C8E8D2089644915484204C9A0C1CC38486A5A4420004A00281612812";
    attribute INIT_1A of inst : label is "40020400204002040020400204002040020100200CFDFFFF8CB008E029405382";
    attribute INIT_1B of inst : label is "9E618C1A65ADB0242005555500001FFFFF800000201002020400204002040020";
    attribute INIT_1C of inst : label is "249199924FAD60139121338011C028E0147202390113C1932ECCCDC1A6DB0320";
    attribute INIT_1D of inst : label is "B6D964EDC055241DE9CF4C327193093B703112D926596DB64939CC9A664B2264";
    attribute INIT_1E of inst : label is "8D4982619589492920EF4E7861938C9849200089294AD631945507044B64A165";
    attribute INIT_1F of inst : label is "B322C58C9B32881E292A9E4E279E70824248D6E7CA1AA50A802E0D3061644A9D";
    attribute INIT_20 of inst : label is "B41A9912A5A962D0686414A58208248248208B16326CC8B16326CCA2062C58C9";
    attribute INIT_21 of inst : label is "A58B41A192438CA0C9B72C645E42645CB9946797332F964B28326DCB16834644";
    attribute INIT_22 of inst : label is "0E321326DCB19179019172E6519E5CCCBE592C84C9B72C5A0D1912D068650A96";
    attribute INIT_23 of inst : label is "79DE7799EE3E1421294058849494F9433332DCC692E951A4B425D4A0A4226A25";
    attribute INIT_24 of inst : label is "CD32A454CA936C59B734CA8924924120141290194B60448997246505B0B79DE7";
    attribute INIT_25 of inst : label is "4086440A243224DB166DCD32A454CA936C59B734CA814486540A0432A4DB166D";
    attribute INIT_26 of inst : label is "FFCC62801404000C08000010141C08077873C3896C941C60C294909491332CC1";
    attribute INIT_27 of inst : label is "0222A492785232B59B4EDCB56D3B72D2DEED8B56C2275967596EDA5A2DB5A7FF";
    attribute INIT_28 of inst : label is "B504381CA24915AD49070D2892056B5041C30A24915AD49070C2AA1209020EC9";
    attribute INIT_29 of inst : label is "892056B5043C30A24915AD49070C2892056B5041C30AA4915AD490F0F2892056";
    attribute INIT_2A of inst : label is "3E8E2A012057B5041C30A24915AD490F0F2A92056B504383CA24915AD4907052";
    attribute INIT_2B of inst : label is "CFE47D891B01C611111111111111111111111111111111111111111111111100";
    attribute INIT_2C of inst : label is "0B8B0B0B8020000000000000021129699F292496842129496922603F3768723E";
    attribute INIT_2D of inst : label is "03000B0B8B8B02000A8A8A8A83000A0B8B8A02000A0A8A8A03000B0B8B8B0200";
    attribute INIT_2E of inst : label is "04CC14020110610844080882108810404020118991042118A8446211820A7018";
    attribute INIT_2F of inst : label is "1042118AC105104231088104044104211820A644104211088101104211088104";
    attribute INIT_30 of inst : label is "D96B2592B65B2964B2C8C42305322082108C54223108C10414C8821088104044";
    attribute INIT_31 of inst : label is "4E3263930C762B29694CACACACA2494DADA4A4ACB592B652CA6B4A5695A536B2";
    attribute INIT_32 of inst : label is "BECE0085FCF9E0103B16002FF1AC6318C6B18D6B1AC635AC7EDE9CF4E653E987";
    attribute INIT_33 of inst : label is "E358C6318C6B18C631FFCF80227EF9FCF828DD75F6050FFFCF80227EF87C146F";
    attribute INIT_34 of inst : label is "492693479BB58F376B00CE7152419F9CF8E400D92B5A7039024C29072C01A207";
    attribute INIT_35 of inst : label is "000094344124040000000240000002100109A6D349B4D36DA4934934DA49A6D3";
    attribute INIT_36 of inst : label is "20808202080821136044E0100004101000400100041010004101040400104124";
    attribute INIT_37 of inst : label is "0080080020008002000800200080020008202000800200080020008202000820";
    attribute INIT_38 of inst : label is "0008208208208208002002000800820208208082082020020808202000210001";
    attribute INIT_39 of inst : label is "568040209C6981143A000000848408088C0C0088080020808208008208208202";
    attribute INIT_3A of inst : label is "085C210000040006844D88A3600003063E0C000490FC90000C166E002201F471";
    attribute INIT_3B of inst : label is "98284402014008320300E03041200000041090285200BB976FF7F26D18D31E51";
    attribute INIT_3C of inst : label is "DAE18002A77B44E01930C986400050A32692820988402521A41E00300880740C";
    attribute INIT_3D of inst : label is "674EDA80A4ADE2E8414D131C051F00000000000000000DECEC1D80D836CECC56";
    attribute INIT_3E of inst : label is "52B4EB0B16BD2D65B1A342CCF33E5C7DFBE287A148B1EE9ABCDD61B7E5A7E3F3";
    attribute INIT_3F of inst : label is "19555E55441E2E3859E39C5E70E087105800DCB3CA5ABEA0D995BB50B24957A4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "556402AA216F1EAD5EFDEAD5EFDEAD5EFDEAD5EFDEAD5EFC57181ADD2D688C0A";
    attribute INIT_01 of inst : label is "FBDF2AE7C3BE2A7DEAD5EF33BC8C90F175FADD7CB65F2D5FEBED7F8FB1FE3ED0";
    attribute INIT_02 of inst : label is "8EEAC8E70302A4FA8621F44607B610113C9BB7BF7B5BBC6B0948CD6371783CE9";
    attribute INIT_03 of inst : label is "F91837F48E447223111808E047033011888C44722391988CC08806F75662EEAC";
    attribute INIT_04 of inst : label is "184D0E7918BF918B7918BF918B715F8C2318C230918BF918B7918BF918379183";
    attribute INIT_05 of inst : label is "7606465B220022902200229022003718AAA3DE47DD5CB84120138A142B74E581";
    attribute INIT_06 of inst : label is "9822902969EA850220190011004654C10A860C80088044010F839FE61864CFBA";
    attribute INIT_07 of inst : label is "7393981CE4E606EE35EE3486C1667F7F03006D36DB49268B6996D329345B4C36";
    attribute INIT_08 of inst : label is "99249A4E348C591CA52314A4729A662331667294CE53CCE046033911C88C0E72";
    attribute INIT_09 of inst : label is "602394E7DE65661F0BD7993304FAF6B43477CC1B2D98CDE6C63CE5C064D269E7";
    attribute INIT_0A of inst : label is "52019BC699C08759C2649268140040064436E70C18992B30F85EBC4A6604CC04";
    attribute INIT_0B of inst : label is "71998FF845C37FB18D46866F3E78D6118330A15CB2948066F1A670277E6672CE";
    attribute INIT_0C of inst : label is "B1FF985E3B1C79A4703306E826369980CDB93733267B367F99933D933DB9CF2B";
    attribute INIT_0D of inst : label is "3FBE79E49493EA2F5FF3C7761E3B01C1E3CFE79D5564B19A71F93939393F7564";
    attribute INIT_0E of inst : label is "D7FE6177FFBFF8F8ED87C3925BFFB48B19E7927D3CECCF1DC76679C24E249F43";
    attribute INIT_0F of inst : label is "66BC64D33A9582AB7CF22800C5000F14A30E7B37921514DDDDFFDFDDFDFFDF95";
    attribute INIT_10 of inst : label is "9A6A2C963963303949ED4A83EA64591FC6377C6EF1A5AC6AD5AFF25AB4CD9B33";
    attribute INIT_11 of inst : label is "D1371B8C5551EF71B14EF38DDB1ABC6D36B1AAD76BFC995B41AE5A69A6186186";
    attribute INIT_12 of inst : label is "3011C26A604B2102011CA0E507293B40267043F0CE171BCC017F4C6F24B44D98";
    attribute INIT_13 of inst : label is "89F13BC68277F4F69FB4D34D34D30C30C42550C660CB69266223919888C44702";
    attribute INIT_14 of inst : label is "1E2224930A878240F00B9AEE839AEBE9FAC1EE838AEBE97ED6AD6119C69CBD10";
    attribute INIT_15 of inst : label is "14EEA629BA95A5344A52439FD51BB4C6CEB576A1CECD5AF5ABADFF3DF0901090";
    attribute INIT_16 of inst : label is "916983D4C8B4C1CA645A60E4322D307A191698390C8B4C1CF2F0F028FF9852C3";
    attribute INIT_17 of inst : label is "933B808C0CA230181460AFAD102B0865EB9F967FCB3FE5D32AE60E532AD30729";
    attribute INIT_18 of inst : label is "0851810C84A2218A6070284A0442801844A24B698D405090AD024F7C16952F01";
    attribute INIT_19 of inst : label is "1440014C07071094603822210115234040030E52210E08995A128C241208A06A";
    attribute INIT_1A of inst : label is "201802018020180201802018000180001998E35D3200000030100707050E0A1C";
    attribute INIT_1B of inst : label is "4AE1EA209E2825E8E0055500001FE01F807F80C0098E35C00201802018020180";
    attribute INIT_1C of inst : label is "3648CD5A68AC4B7DD7D9DFE39DF1EEF8E77E7BBF39D6B176C57FD7A20965C3ED";
    attribute INIT_1D of inst : label is "EB2EB383A0A4E62791C0CC4E72731420E84569A699E59E59F59CFECB32A8B632";
    attribute INIT_1E of inst : label is "60004204277E0D97313C8E0672739398A1DBF7351729CAF027833BB9A69A76B2";
    attribute INIT_1F of inst : label is "D128D1AE4F135D6AADAB6975BA6DA853D3DDA7850A57CC5DC092C0088C13B320";
    attribute INIT_20 of inst : label is "3ECADF3619867AFB297E3295895891A95A918306B93C48306B93C4D57A8D1AE4";
    attribute INIT_21 of inst : label is "99EBEDADF8F78FA2F89EDC7D5BC17F5B79FC7F6E3EAD67F369BE26B3D7D977C3";
    attribute INIT_22 of inst : label is "DE3E8BE27B71F56F45FD6DE7F1FDB8FAB59FCDA6F89ECF5F6DDF4CFB697CDA66";
    attribute INIT_23 of inst : label is "AD6B5AD6B5E5E398E6399B86F9EA650EB1326DC2B34B70ACD075D882B5BB4DF9";
    attribute INIT_24 of inst : label is "8DFE3B17F8F13C189E37F8FE6F279BC9E3BBE42DA1AEC6CD1A34B684DB1AD6B5";
    attribute INIT_25 of inst : label is "5DAFC6A2CD7E3C4D46278DFEBB17FAF135189E37FAC44D8FD6224C7EBC4F0627";
    attribute INIT_26 of inst : label is "FFF2360024202030300000243430206DE6602314D34B9C9CC41A1A1E1FAAACD4";
    attribute INIT_27 of inst : label is "B1BC93CF276B9B9CBB069AB76C126ACADE69EB56F773517351669B5B6DB5CFFF";
    attribute INIT_28 of inst : label is "CE0B337133F76E7182CDD64CFDDB8C60B137933F76E3182C4DF4ECDFE024666C";
    attribute INIT_29 of inst : label is "CFDDB9CE0B135933F76E7382C4DF4CFDDB9CE0B337D3BF76E7382C4DC4CFDDB9";
    attribute INIT_2A of inst : label is "8C5551FFDDB8CE0B137D33F76E7382CCDC4EFDDB9CE0B337133F76E7382CDDE4";
    attribute INIT_2B of inst : label is "C2626198AF57018444504504445045044444445045051050450444451050451B";
    attribute INIT_2C of inst : label is "0E0E8E0E8CD000050000500019748A0A84E5DA4DE739EF20DA89968BF9BA1130";
    attribute INIT_2D of inst : label is "E5840E8E0E8E04840F0F8F0F85840E8E8E0E05840E0E8E0E85840E8E0E8E0484";
    attribute INIT_2E of inst : label is "204779B4DA34D34160BAC1E782C135D21B4DA34083CF058A6120F058A7980FC7";
    attribute INIT_2F of inst : label is "3CD058AE575C3CF0782C135D20D3CD058AEB820D3CD0582C17583CF0582C13CF";
    attribute INIT_30 of inst : label is "1218080584825A0101C1E4B1DF1069A682C57092782C534D3041E782C135D20D";
    attribute INIT_31 of inst : label is "8A0C426203DB58181AE16161617000E9696060610C2580B4175AC631AC6BA5A4";
    attribute INIT_32 of inst : label is "4131FF7A03061FEFC4E9FFD3F18C6B1AC6B18C6318C6B18C7F791088A0B49108";
    attribute INIT_33 of inst : label is "E358C6B58C631AD6B1F8307FDD81060307D7228A09FAF000307FDD810783EB90";
    attribute INIT_34 of inst : label is "49369948576FE0AFD7DA6B4C72C272F3B7B7FFA68CE39E6BD7C75F36E87F7877";
    attribute INIT_35 of inst : label is "20DF7A8B808F84001B8088F62000000107D1B4196D941961B49A6126D0650691";
    attribute INIT_36 of inst : label is "24009002400906088B8230000184901240480124049012404801240480120100";
    attribute INIT_37 of inst : label is "0090092024009202480920248092024009002400900240090024009002400900";
    attribute INIT_38 of inst : label is "400900900900900900240240090090024024009009002402400920241B200099";
    attribute INIT_39 of inst : label is "88014041010420C1068001000000000000000001092024009009209009009002";
    attribute INIT_3A of inst : label is "D92771835E281AF50295001F44057B81C0680AF5045C5815EF00CE001EDC62AA";
    attribute INIT_3B of inst : label is "9827B24443D92C9B41DE8618789780681717A5B363E79F910F05038146FFFF01";
    attribute INIT_3C of inst : label is "73DE8B6CE5E3BB22959DACED4A0445A2DFE6DF1F7C9242D97F49EB168E5B580B";
    attribute INIT_3D of inst : label is "BCA220734DD311511D051744BDC0000000000000000035A6D4DA96E9BA656759";
    attribute INIT_3E of inst : label is "00804000A04080AA091024AC2060900103C310C007818471325283061C521900";
    attribute INIT_3F of inst : label is "134C288628910346867E6E3704FA51528A0F0F0691930343260245A1202A904A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "543622A1B0673B76EDDBB76E993264C993264C993264C9923E3986CCC363DCC1";
    attribute INIT_01 of inst : label is "91138372E1130461C18187869E5C80F13399CCF67B3D9EF77EEFDFFBFF7FEFDC";
    attribute INIT_02 of inst : label is "C6798C13A1301E6FC3ACB4C0623A06838C89031221099C270739CCE733301891";
    attribute INIT_03 of inst : label is "F3058F3180CC06603305982CC1660A301980CC0660B305182CCA4233CC666798";
    attribute INIT_04 of inst : label is "166C8473058F3058F3058F3058F01D8C6318C6303058F3058F3058F3058F3058";
    attribute INIT_05 of inst : label is "4472065220DB20DB20DB2293329377C1FF77B5FD83BEA985A7D24D9325A4754C";
    attribute INIT_06 of inst : label is "9122932201908832091049984874441B6230C836C83661B187878AAE14E48572";
    attribute INIT_07 of inst : label is "60B305982CC1671E319E31E2C8616167210C6DB09261248B4D06DB2DA6124824";
    attribute INIT_08 of inst : label is "9924986E3182C3058460B08C0618C046020C04118283182CC14602301980CC16";
    attribute INIT_09 of inst : label is "146020B2D864E43233065E6034C2C23B3C731C932938C563C258E1CC749B4825";
    attribute INIT_0A of inst : label is "589289C63059C039C2649266C636636A4624349CCC992321911830F0C14180CC";
    attribute INIT_0B of inst : label is "70B385B873806CFB8C276F271B38CE3011F1901C921624A2318C16770EE1724C";
    attribute INIT_0C of inst : label is "A1AAB65A3859658C06770638BE363011CC3830B72029302C5B9014901439C66C";
    attribute INIT_0D of inst : label is "B1B2F3CDB1B6CC6C1873C6E41C3B0691830CE79A8274A9F251EB3B3B3B380074";
    attribute INIT_0E of inst : label is "12AAD9775755D1D1D70684B6D000BECA1BCF36D9B8D9CF1B26CE79B6DC0DB666";
    attribute INIT_0F of inst : label is "221CE44922DC839A5C218C363186C702094CBF37F30701BBBB9B9BB9B9B9B995";
    attribute INIT_10 of inst : label is "8E3A2C122B260330508E6B00402709C9CA7274E4F19224E593955F09A4C48931";
    attribute INIT_11 of inst : label is "51A73BE0FFBBE173A320029C9D393C64B09396C4E557C91B89A04E38E38E38E3";
    attribute INIT_12 of inst : label is "0A301A24034A3D030ED82CC1660B305A0C16207182C71CEC61614131B09468F8";
    attribute INIT_13 of inst : label is "F9C1B9B24E50E3E7BF186186186186186404464C06D3620C046033019828C146";
    attribute INIT_14 of inst : label is "DB1B2492856F16CC47518DC63989C0E3752AC63989C0E374C66C61D1E7903918";
    attribute INIT_15 of inst : label is "1CCF7639BDDF27E4DAD6B7948D19244E4C130E5BCA48DC4AC64155E59CD6DCD6";
    attribute INIT_16 of inst : label is "BD65BB9CDEB2DDEE6F596EF737ACB7739BD65BB9CDEB2DDCF66F73D65F981B87";
    attribute INIT_17 of inst : label is "B621C99E59A6793CB4F315415432886DBBDBB6D55B6AADF37AF6EF737ACB7739";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFDFFFF13CC6E2DEDB1903F9D99B0740DA6D8ADB21";
    attribute INIT_19 of inst : label is "7FFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "BFFDFBFFDFBFFDFBFFDFBFFDFBFFDFBFFFFFFFFFFF8200007FFFFFDFDFBFBF7F";
    attribute INIT_1B of inst : label is "19DDCA229208A499EC0AAAAA0FFFFFFFFFFFFF003FFFFFFDFBFFDFBFFDFBFFDF";
    attribute INIT_1C of inst : label is "3240C418849949481C8188619930EC98764E3B271D9470F1E04C4622292480E9";
    attribute INIT_1D of inst : label is "69A69A5223A0C363305182CC0660B6D488CC49B6C9249A69A6829E4133249990";
    attribute INIT_1E of inst : label is "FFFFFFFE4A3E0C861B1980CC04603305B68BE7A2F4A5ADCE4B86F8FD26DB0C92";
    attribute INIT_1F of inst : label is "C16CD98F1C174CE425C7C1A1904319CB0B27978EBC55EDDEBFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "32DECC36519462CB7B30B6B5BCDBCDBCDBCDB3663C705B3663C705D338CD98F1";
    attribute INIT_21 of inst : label is "D18B2DECC2F7061260B88C305D1B305A30C83046182E477365982E23165BC30A";
    attribute INIT_22 of inst : label is "DC18D982E230C17464C168C320C11860B91DCDB260B88C596F0C28CB7930DB46";
    attribute INIT_23 of inst : label is "8461184230C16318E73BD726198AE51A3034E1B6670B2D99C7759D12B5B3ADB9";
    attribute INIT_24 of inst : label is "0498FB8263E17198B81263EE673399CD61BCE424209C060C193890864F184611";
    attribute INIT_25 of inst : label is "1DB31EF0ED98F85C662E0498FB8263E17198B81263DE1DB30EF0ED98785C662E";
    attribute INIT_26 of inst : label is "00022600040808080800000C0C0C1C6CCC046034DB63011828CECECECE222EDE";
    attribute INIT_27 of inst : label is "7312B249246789188B2F58B22CBD72C858F58B22F7731373136F595B65B5EC00";
    attribute INIT_28 of inst : label is "4226A2C1A324421081A8B168C9108420602C5A32542108180B16AF8B99A4E564";
    attribute INIT_29 of inst : label is "8C9108420622C5A32542108980B168C9508422622C1AB2442108988B068C9508";
    attribute INIT_2A of inst : label is "E0FFBB7C9508420622C1A32442108188B06AC95084206A2C1A324421081A8B16";
    attribute INIT_2B of inst : label is "E0E461DB335778FFEAABEBEBEBEBEBEBEBFFEABFEAAABFFFEABFEABFEABFEABB";
    attribute INIT_2C of inst : label is "008000880C80000000002AAABC749484A4849248E739EF20DA8DCB7D1CD99230";
    attribute INIT_2D of inst : label is "1900008000888900000000888900018000898900008000888900000000888900";
    attribute INIT_2E of inst : label is "04CC1402011041080408088210081040402011099104201828044201820A4020";
    attribute INIT_2F of inst : label is "10420182C105104221008104044104201820A644104201008101104201008104";
    attribute INIT_30 of inst : label is "B6C49B6C4926C4926C48840305322082100C14022100C10414C8821008104044";
    attribute INIT_31 of inst : label is "80CC0660311984C4C632121B1B19B43A1A1A1A1242486D8DB1C4218C6210CC49";
    attribute INIT_32 of inst : label is "0000000000000000000000000E739CE739CE739CE739CE7381330198098C3019";
    attribute INIT_33 of inst : label is "1CA7294A539CE739CE0000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "4DB4DA6C645AC8C8B59A210C269A6043023BFFB6C4210C6881220486DACF5170";
    attribute INIT_35 of inst : label is "0049A7D803F604000800029001000010224926DB69B6D26D26D369269B6D36D2";
    attribute INIT_36 of inst : label is "200080020008000FD80380000004101040410104041010404101040400100100";
    attribute INIT_37 of inst : label is "0082080020808002000800200080020808002080820208082020808002000800";
    attribute INIT_38 of inst : label is "0008008008008008002082000800800200200082082020020808202088200401";
    attribute INIT_39 of inst : label is "D80F1CF1C73D71CF7E0000000404800084048800082020808008008008008002";
    attribute INIT_3A of inst : label is "F9FBF880FC0007E2879A8FEEA203F047C00407E09F82080FC53F1007D9DF07FD";
    attribute INIT_3B of inst : label is "90080418094008120040201043210000049104284280944AA040800428103000";
    attribute INIT_3C of inst : label is "EC740E96DA359283C49E24F12E0022A52691A21A8822040480D2852009A41004";
    attribute INIT_3D of inst : label is "73F0E3F8F4EB0500514503445410000000000000000039A710E25F69DA712789";
    attribute INIT_3E of inst : label is "FEBC7F8FF3E7EFA6BD7AFEF5D7AF4FDF7D79FD387F1F79E3A75C7D3A71F9FD3C";
    attribute INIT_3F of inst : label is "D34F35D334E9EBD3C79D67F1C73CFA63F78FD7AE99EBEBF9D7D7D61EBA79F7E4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "FC1027E000228000000000000000000000000000000000007E1802AC01534C03";
    attribute INIT_01 of inst : label is "48B90720C0862450A9414503940A48C89148A44221108812A25448891122244C";
    attribute INIT_02 of inst : label is "863888528100B42F82A534C1223200111A44A28911088A228F7BC6C631291541";
    attribute INIT_03 of inst : label is "53008511804C026013049824C126013049824C126013009801880231C4426388";
    attribute INIT_04 of inst : label is "1264045300853008530085300856158C6318C630300853008530085300853008";
    attribute INIT_05 of inst : label is "D2492E00600160496001620162010000000137998A2640C72753499325A47215";
    attribute INIT_06 of inst : label is "0062016021438096003000B00052C2492E1258125812C09107424AA93091A548";
    attribute INIT_07 of inst : label is "6083041820C10615109511A3A1D1515681002490492092482090002000400080";
    attribute INIT_08 of inst : label is "90000A45118003000460008C0014C026000C001182029820C126093049824C10";
    attribute INIT_09 of inst : label is "106080925452D2292285086080A2A2313C510A170035AFD7A2F850A452400165";
    attribute INIT_0A of inst : label is "700045A230408015A240002A5C12C1212C129D8A4C94969149142844C129820C";
    attribute INIT_0B of inst : label is "28914794514095E344252D629B944C3001A8C008001C0011688C1022A6532004";
    attribute INIT_0C of inst : label is "A0AA94CA3449248C023285149D3230088A14299200201024C90010001015AE38";
    attribute INIT_0D of inst : label is "A0A2410490928D2810C112E40C1F0611020582080861A0D05189999999980061";
    attribute INIT_0E of inst : label is "02AA5336541501011506849255559C5A890412519A5B044B72D820B24C049472";
    attribute INIT_0F of inst : label is "910AC22B62DA83490A90B8121702428082121AA5110101BBBBB99BBB99BB99B5";
    attribute INIT_10 of inst : label is "08212C1669060030408C642A286C0B18A96A52D4AB52025101455D2494A24528";
    attribute INIT_11 of inst : label is "7096800000006153A320225A94B52AD4B00944C051574B0B09E0482082082082";
    attribute INIT_12 of inst : label is "01300A600A1A9F060CD820C1060830400C100029820299A461412170909C25D4";
    attribute INIT_13 of inst : label is "F349A8B60CC0A6A295145145145145145205C20C0049290C126083041804C026";
    attribute INIT_14 of inst : label is "1902249385253644C6009842309840A3540042309840A354C764D148A7342B09";
    attribute INIT_15 of inst : label is "1C984639611D07A0D6B5955A54B512AD2428854AAD255848850155D555801580";
    attribute INIT_16 of inst : label is "912193504890C988244864C4122432620912193104890C98D628570457580387";
    attribute INIT_17 of inst : label is "922358CACC832B159057400155609A4493D99255492AA4C122664D41224326A0";
    attribute INIT_18 of inst : label is "00000000000000000000000000000315C4624E490B03FB8B890E024AE480C961";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0D4CAE0200080018A20555550000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "20288014A40800801011004155208A90454A22A5115068C180C44C60200000A0";
    attribute INIT_1D of inst : label is "000000566200C1063041820C00608215988024001082000000029C0000000002";
    attribute INIT_1E of inst : label is "00000004007D0A560831804C006003041051D614DA52100C0342D4F090004A08";
    attribute INIT_1F of inst : label is "812448894813C4502D4D83018002194A0A2E1226705F4C9A8000000000000000";
    attribute INIT_20 of inst : label is "12CAD826C0B0224B2B6036B4959959959959912225204912225204F114448894";
    attribute INIT_21 of inst : label is "C0892CAD80F70C16C09004604C0B6048118862023026036B65B0240112594618";
    attribute INIT_22 of inst : label is "DC30CB02401181302D812046218808C0980DADB6C09004496518604B29609B02";
    attribute INIT_23 of inst : label is "8C6318C2308BD6B58C6316240D8A4D1A202445923203648C82748B3694B2A7B5";
    attribute INIT_24 of inst : label is "0CB0DE82C36120889032C36D068341A1D1B0D26C299A050A1521B0A2EA98C631";
    attribute INIT_25 of inst : label is "09960A504CB0584822240CB0DE82C36120889032C34A09960A504CB058482224";
    attribute INIT_26 of inst : label is "000236000C000000000000040404046D8C026012000B0018204A4A4A4A22244A";
    attribute INIT_27 of inst : label is "EA8829248C15011889274C92649D3248CC7489267773193319274B492C94CC00";
    attribute INIT_28 of inst : label is "000606C4A32400000180B128C9000000622C0A32500000189B02AF451C004540";
    attribute INIT_29 of inst : label is "8C9000002602C0A32500000189B028C9400000686C0AB25000001A1B028C9000";
    attribute INIT_2A of inst : label is "0000007C9400000686C0A325000001A1B02AC9000000606C4A32400000980B12";
    attribute INIT_2B of inst : label is "40C1208B72FD60C0154141414140154015414140154141541401414015401540";
    attribute INIT_2C of inst : label is "00808000080000000000000015D0000001A00001C631AD604B815B7814498090";
    attribute INIT_2D of inst : label is "0180008080000180008080000180008080000180008080000180008080000180";
    attribute INIT_2E of inst : label is "04CC1402011041080408088210081040402011099104201828044201820A4000";
    attribute INIT_2F of inst : label is "10420182C105104221008104044104201820A644104201008101104201008104";
    attribute INIT_30 of inst : label is "00400004049240492448840305322082100C14022100C10414C8821008104044";
    attribute INIT_31 of inst : label is "804C006011190040422000090910902009000900200404809140008001088400";
    attribute INIT_32 of inst : label is "C1B1FF7A03061FEFC4E9FFD00000000000000000000000000163041804A53041";
    attribute INIT_33 of inst : label is "00000000000000000000307FDD83060307F7638E19FEF000307FDD830783FBB0";
    attribute INIT_34 of inst : label is "4D36DB6CC0084980109803180002C0C60233FE000000082002800A04728D4170";
    attribute INIT_35 of inst : label is "00240015400504000000020000084000000DA69A6DB6DB49249A69B6DB6DB4DB";
    attribute INIT_36 of inst : label is "2080820208082100154020004004001000400100040010004001000410104100";
    attribute INIT_37 of inst : label is "0080080020808002000800200080020808202080820208082020808202080820";
    attribute INIT_38 of inst : label is "0808208208208208202082080820820208208080080020820008002004200401";
    attribute INIT_39 of inst : label is "0410600008008400020000000000000000000000082020008208208208208202";
    attribute INIT_3A of inst : label is "A800AA8000140002002A800AA2000100101000020000A0000000150000000000";
    attribute INIT_3B of inst : label is "51180D180B001A3200D26810C1608010A040B060C20190020100004428115000";
    attribute INIT_3C of inst : label is "2C7402945A327680A28D1468800006040200860A1A600C0080160C0000803000";
    attribute INIT_3D of inst : label is "9815300D1D2B05015555111415050000000000000000344288510290A428A347";
    attribute INIT_3E of inst : label is "03A500C070A8A8A2A50A0A9554A151530B0C050A01A74D34A946054A180D074A";
    attribute INIT_3F of inst : label is "554715531C3A3A7460D53438E9868A3450D050A3AD38382A70705282AA387066";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
