library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity eprom_5 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of eprom_5 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"06",X"0C",X"08",X"04",X"02",X"01",X"80",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",
		X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"04",X"C0",X"E0",X"F0",X"F8",X"EC",X"E6",X"E3",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",
		X"FF",X"0F",X"38",X"E0",X"80",X"00",X"00",X"00",X"FF",X"F0",X"FC",X"E7",X"E1",X"E0",X"E0",X"E0",
		X"FF",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"40",
		X"00",X"03",X"0F",X"1A",X"3B",X"60",X"5B",X"EA",X"E0",X"E0",X"F0",X"B8",X"BC",X"06",X"BA",X"AB",
		X"10",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"01",X"01",X"01",X"01",X"01",X"01",
		X"BB",X"80",X"BB",X"2A",X"3B",X"00",X"3B",X"2A",X"BB",X"01",X"BB",X"AA",X"BB",X"00",X"BB",X"AA",
		X"02",X"03",X"81",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"40",X"00",X"00",X"00",X"20",X"00",X"10",
		X"BB",X"80",X"9B",X"CA",X"4B",X"60",X"33",X"18",X"BB",X"01",X"BB",X"AB",X"BA",X"06",X"BC",X"B8",
		X"81",X"03",X"02",X"02",X"02",X"06",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"04",X"02",X"01",X"00",X"00",
		X"0E",X"03",X"00",X"00",X"00",X"00",X"80",X"20",X"70",X"E0",X"E0",X"E0",X"E0",X"E0",X"E1",X"E7",
		X"08",X"18",X"10",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"08",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"F0",X"FF",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"F0",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"01",X"03",X"06",X"0C",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E1",
		X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",
		X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"E3",X"E6",X"EC",X"F8",X"F0",X"FF",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"18",X"30",X"60",X"C0",X"80",X"FF",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"E0",X"E0",
		X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"F0",X"F8",
		X"01",X"01",X"01",X"01",X"01",X"FD",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"00",X"EC",X"E6",X"E3",X"E1",X"E0",X"E0",X"E0",X"60",
		X"60",X"C0",X"80",X"00",X"00",X"01",X"03",X"06",X"30",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",
		X"00",X"00",X"20",X"70",X"D8",X"8C",X"06",X"03",X"20",X"10",X"08",X"04",X"02",X"01",X"03",X"06",
		X"0C",X"18",X"30",X"70",X"D8",X"8C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"80",X"40",X"20",X"10",X"08",X"8C",X"D8",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"E1",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"80",X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"03",X"06",X"0C",X"18",X"30",
		X"00",X"DF",X"8C",X"06",X"03",X"01",X"00",X"00",X"E0",X"FF",X"01",X"03",X"06",X"8C",X"D8",X"F0",
		X"01",X"FF",X"8C",X"06",X"03",X"01",X"03",X"06",X"80",X"C0",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"40",X"20",X"11",X"7B",X"00",
		X"00",X"00",X"20",X"50",X"C8",X"84",X"FE",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E1",X"E0",X"E0",
		X"0C",X"18",X"30",X"60",X"C0",X"80",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"E0",
		X"30",X"18",X"0C",X"06",X"03",X"01",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"FF",X"F0",
		X"01",X"01",X"01",X"01",X"01",X"01",X"FD",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"00",X"F8",X"EC",X"E6",X"E3",X"E1",X"E0",X"E0",X"E0",
		X"30",X"60",X"C0",X"80",X"00",X"00",X"01",X"03",X"60",X"30",X"18",X"30",X"60",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"10",X"08",X"04",X"02",X"01",X"00",
		X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"00",X"7F",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"FE",X"AA",X"FF",X"AA",X"AA",X"FF",X"FF",X"55",X"AA",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"3F",X"40",X"3F",X"5E",X"5F",X"5F",X"5F",X"5F",X"60",X"3F",X"00",
		X"BF",X"BF",X"5E",X"00",X"5E",X"5E",X"5E",X"5E",X"72",X"BF",X"72",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"BF",X"BF",X"BF",X"BF",X"72",X"BF",X"72",X"BF",X"5E",X"5E",X"5E",X"00",X"7E",X"BF",X"BF",X"BF",
		X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"00",X"3F",X"6F",X"5F",X"5F",X"5F",X"5F",X"5E",
		X"00",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"FE",
		X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"AA",X"3F",X"FF",X"FF",X"FF",X"FF",X"BF",X"C0",X"3F",
		X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"80",X"DF",X"DF",X"DF",X"DF",X"C0",X"5F",X"80",
		X"BF",X"FF",X"BF",X"BF",X"FF",X"FF",X"40",X"BF",X"80",X"C1",X"80",X"80",X"C1",X"C1",X"41",X"80",
		X"FE",X"FF",X"FE",X"FE",X"FF",X"FF",X"01",X"FE",X"00",X"FD",X"FD",X"FD",X"FD",X"00",X"FD",X"00",
		X"E0",X"F7",X"F7",X"F7",X"F7",X"F0",X"17",X"E0",X"2F",X"7F",X"2F",X"2F",X"7F",X"7F",X"50",X"2F",
		X"FA",X"FF",X"FA",X"FA",X"FF",X"FF",X"05",X"FA",X"03",X"F7",X"F7",X"F7",X"F7",X"03",X"F4",X"03",
		X"F8",X"FD",X"FD",X"FD",X"FD",X"FC",X"05",X"F8",X"0B",X"1F",X"0B",X"0B",X"1F",X"1F",X"14",X"0B",
		X"E8",X"FC",X"E8",X"E8",X"FC",X"FC",X"14",X"E8",X"0F",X"DF",X"DF",X"DF",X"DF",X"0F",X"D0",X"0F",
		X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"02",X"FC",X"1F",X"BF",X"BF",X"BF",X"BF",X"1F",X"A0",X"1F",
		X"05",X"0F",X"C5",X"05",X"1F",X"0F",X"0A",X"05",X"00",X"00",X"C0",X"01",X"12",X"0C",X"00",X"00",
		X"D0",X"F8",X"D0",X"D1",X"FA",X"FC",X"28",X"D0",X"05",X"0F",X"15",X"45",X"8F",X"0F",X"0A",X"05",
		X"00",X"00",X"10",X"48",X"84",X"01",X"00",X"00",X"D0",X"F8",X"D0",X"D0",X"FC",X"F9",X"28",X"D0",
		X"05",X"0F",X"05",X"15",X"2F",X"CF",X"0A",X"05",X"00",X"00",X"0C",X"10",X"21",X"C0",X"00",X"00",
		X"D0",X"F8",X"D4",X"D0",X"F9",X"F8",X"28",X"D0",X"05",X"0F",X"05",X"85",X"4F",X"1F",X"0A",X"05",
		X"00",X"00",X"01",X"84",X"48",X"10",X"00",X"00",X"D0",X"F8",X"D1",X"D4",X"F8",X"F8",X"28",X"D0",
		X"A7",X"A7",X"46",X"00",X"5E",X"5E",X"5E",X"5E",X"62",X"A7",X"62",X"A7",X"A7",X"A7",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A7",X"62",X"A7",X"62",X"A7",X"5E",X"5E",X"5E",X"00",X"66",X"A7",X"A7",X"A7",
		X"83",X"83",X"46",X"00",X"5E",X"5E",X"5E",X"5E",X"42",X"83",X"42",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"42",X"83",X"42",X"83",X"5E",X"5E",X"5E",X"00",X"66",X"83",X"83",X"83",
		X"81",X"81",X"42",X"00",X"5E",X"5E",X"5E",X"5E",X"00",X"81",X"00",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"00",X"81",X"00",X"81",X"5E",X"5E",X"5E",X"00",X"42",X"81",X"81",X"81",
		X"81",X"81",X"42",X"00",X"5E",X"5E",X"5E",X"5E",X"00",X"81",X"00",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"00",X"81",X"00",X"81",X"5E",X"5E",X"5E",X"00",X"42",X"81",X"81",X"81",
		X"00",X"00",X"00",X"00",X"5E",X"5E",X"5E",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"5E",X"5E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"C0",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"7E",
		X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",X"0E",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"18",X"2C",X"7E",X"83",X"83",X"83",X"83",X"00",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"00",X"83",X"83",X"83",X"83",X"00",X"2C",X"18",
		X"F1",X"80",X"00",X"00",X"01",X"80",X"B0",X"B0",X"B0",X"B0",X"B1",X"80",X"00",X"00",X"01",X"8F",
		X"F1",X"80",X"00",X"00",X"01",X"80",X"B0",X"B0",X"B0",X"B0",X"B1",X"80",X"00",X"00",X"01",X"8F",
		X"F1",X"80",X"00",X"00",X"01",X"80",X"B0",X"B0",X"B0",X"B0",X"B1",X"80",X"00",X"00",X"01",X"8F",
		X"03",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",
		X"03",X"03",X"07",X"07",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",
		X"80",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"7E",X"78",X"E1",X"81",X"03",X"03",X"07",X"07",
		X"80",X"E0",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"7E",X"78",X"E1",X"81",X"03",X"03",X"07",X"07",
		X"1F",X"1F",X"3F",X"3F",X"7E",X"78",X"E1",X"81",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",
		X"1F",X"1F",X"3F",X"3F",X"7E",X"78",X"E1",X"81",X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",
		X"87",X"92",X"10",X"0C",X"C8",X"21",X"21",X"E1",X"19",X"21",X"41",X"8F",X"90",X"20",X"27",X"09",
		X"22",X"E6",X"39",X"11",X"93",X"F2",X"92",X"12",X"39",X"67",X"44",X"CC",X"43",X"40",X"44",X"4B",
		X"C9",X"09",X"1C",X"A4",X"26",X"49",X"48",X"7C",X"09",X"08",X"84",X"47",X"39",X"00",X"C6",X"F9",
		X"11",X"F9",X"C8",X"44",X"4C",X"32",X"31",X"C8",X"31",X"10",X"88",X"47",X"22",X"12",X"9E",X"F9",
		X"E3",X"C1",X"C8",X"5C",X"1C",X"18",X"C3",X"E6",X"91",X"92",X"DC",X"C0",X"01",X"1F",X"12",X"32",
		X"89",X"0F",X"11",X"70",X"92",X"0E",X"3F",X"4C",X"08",X"0C",X"D3",X"21",X"10",X"7C",X"83",X"81",
		X"3E",X"26",X"C2",X"03",X"34",X"CC",X"89",X"81",X"60",X"49",X"29",X"3F",X"E0",X"80",X"0E",X"1F",
		X"48",X"20",X"36",X"49",X"C8",X"0C",X"13",X"22",X"60",X"10",X"0F",X"88",X"40",X"F1",X"09",X"09",
		X"D0",X"D0",X"D0",X"D0",X"D7",X"D4",X"D4",X"D4",X"01",X"FF",X"81",X"81",X"FF",X"9F",X"90",X"90",
		X"25",X"E7",X"21",X"21",X"3F",X"FF",X"00",X"0E",X"6A",X"EF",X"42",X"42",X"7E",X"EE",X"2A",X"2A",
		X"D4",X"D4",X"94",X"94",X"94",X"9F",X"C4",X"FF",X"FF",X"90",X"90",X"90",X"91",X"91",X"91",X"D0",
		X"FF",X"21",X"71",X"A9",X"15",X"0F",X"05",X"89",X"7A",X"FB",X"FA",X"FA",X"7E",X"70",X"7F",X"F8",
		X"FC",X"7F",X"FE",X"42",X"FE",X"62",X"7B",X"4A",X"D0",X"D0",X"D0",X"D0",X"D7",X"D4",X"D4",X"FF",
		X"71",X"01",X"0D",X"01",X"BF",X"A1",X"A7",X"FF",X"28",X"FE",X"6B",X"6A",X"EB",X"4A",X"EA",X"6A",
		X"4A",X"DF",X"42",X"42",X"7F",X"50",X"50",X"FF",X"F5",X"FF",X"BD",X"81",X"FF",X"00",X"00",X"FF",
		X"24",X"FF",X"25",X"25",X"E5",X"25",X"25",X"25",X"6A",X"6B",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"24",X"12",X"01",X"01",X"19",X"A1",X"00",X"73",X"21",X"01",X"82",X"80",X"00",X"02",X"00",
		X"00",X"63",X"21",X"25",X"C4",X"00",X"01",X"03",X"00",X"80",X"80",X"A0",X"A4",X"78",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"05",X"1F",X"A1",X"00",X"7F",X"25",X"25",X"A2",X"80",X"00",X"23",X"21",
		X"25",X"67",X"25",X"25",X"FC",X"24",X"21",X"03",X"00",X"A0",X"A7",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"A5",X"7F",X"A5",X"00",X"FF",X"A5",X"25",X"FF",X"81",X"81",X"FB",X"A1",
		X"25",X"F7",X"25",X"A5",X"FD",X"A4",X"21",X"67",X"00",X"A5",X"EF",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"A5",X"FF",X"A5",X"00",X"FF",X"A5",X"A5",X"FF",X"A5",X"A5",X"FF",X"A5",
		X"A5",X"FF",X"A5",X"A5",X"FF",X"A5",X"A5",X"FF",X"00",X"A5",X"FF",X"A5",X"A5",X"7E",X"24",X"18",
		X"00",X"08",X"00",X"02",X"02",X"00",X"02",X"00",X"00",X"5A",X"5A",X"00",X"5A",X"5A",X"00",X"5A",
		X"5A",X"00",X"5A",X"5A",X"00",X"5A",X"5A",X"00",X"00",X"02",X"00",X"02",X"02",X"00",X"08",X"00",
		X"18",X"2C",X"7E",X"83",X"83",X"83",X"83",X"00",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"00",X"83",X"83",X"83",X"83",X"00",X"2C",X"18",
		X"00",X"00",X"00",X"18",X"2C",X"7E",X"83",X"83",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"83",X"83",X"00",X"2C",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"2C",X"7E",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"00",X"2C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"3E",X"00",X"D6",X"D6",X"D6",X"D6",X"D0",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"D0",X"D6",X"D6",X"D6",X"D6",X"3E",X"3E",X"1E",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"3E",X"3E",X"3E",X"3E",X"00",X"DE",X"DE",X"DE",X"DE",X"DF",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"DF",X"DE",X"DE",X"DE",X"DE",X"3E",X"3E",X"3E",X"3E",X"1E",X"0C",X"00",X"00",
		X"00",X"1C",X"3E",X"3E",X"3E",X"3E",X"3E",X"00",X"D6",X"D6",X"D6",X"D6",X"D0",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"D0",X"D6",X"D6",X"D6",X"D6",X"3E",X"3E",X"3E",X"3E",X"3E",X"1E",X"0C",X"00",
		X"0C",X"1E",X"38",X"77",X"2F",X"2F",X"2F",X"7E",X"D6",X"D6",X"D6",X"D6",X"D0",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"D0",X"D6",X"D6",X"D6",X"D6",X"7E",X"2F",X"2F",X"2F",X"77",X"38",X"0E",X"04",
		X"0C",X"1E",X"3E",X"7F",X"FF",X"BF",X"BF",X"00",X"D6",X"D6",X"D6",X"D6",X"D1",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"D1",X"D6",X"D6",X"D6",X"D6",X"00",X"BF",X"BF",X"FF",X"7F",X"2E",X"16",X"0C",
		X"0C",X"1E",X"3C",X"79",X"F3",X"B7",X"B7",X"00",X"D6",X"D6",X"D6",X"D6",X"D1",X"DE",X"DE",X"DE",
		X"DE",X"DE",X"DE",X"D1",X"D6",X"D6",X"D6",X"D6",X"00",X"B7",X"B7",X"F3",X"79",X"2C",X"16",X"0C",
		X"18",X"2C",X"5E",X"83",X"81",X"82",X"83",X"00",X"DE",X"9E",X"9E",X"D6",X"DA",X"D8",X"D6",X"DE",
		X"DE",X"DE",X"DE",X"1E",X"DE",X"CE",X"DC",X"DA",X"00",X"83",X"83",X"81",X"83",X"00",X"2C",X"18",
		X"18",X"2C",X"7E",X"A7",X"CB",X"D3",X"D3",X"7E",X"FE",X"DE",X"DE",X"FE",X"DE",X"DE",X"DF",X"DE",
		X"DE",X"DF",X"FE",X"DF",X"FE",X"DF",X"DE",X"DE",X"7E",X"97",X"A7",X"AB",X"D3",X"10",X"2C",X"18",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"00",X"01",X"31",X"38",X"98",X"40",X"80",X"03",X"01",X"00",X"40",X"21",X"11",X"00",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"80",X"80",
		X"00",X"40",X"88",X"18",X"30",X"02",X"01",X"00",X"80",X"88",X"04",X"04",X"08",X"03",X"07",X"07",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"02",X"04",X"00",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"1C",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"10",X"00",
		X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"10",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"06",X"0C",X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"38",X"10",X"00",X"00",X"00",X"00",X"10",X"38",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"7F",X"7F",X"5F",X"4F",X"3F",X"1E",X"02",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",X"2F",X"27",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",X"FC",X"FC",X"7C",X"3C",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"3F",X"3F",X"2F",X"27",X"1F",X"0F",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",X"FC",X"FC",X"7C",X"3C",X"F8",X"70",X"00",X"00",
		X"00",X"07",X"0F",X"1F",X"1F",X"17",X"13",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"F8",X"FC",X"FE",X"FE",X"BE",X"9E",X"7C",X"38",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"1F",X"1F",X"17",X"13",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"F8",X"FC",X"FE",X"FE",X"3E",X"1E",X"3C",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"07",X"0F",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"F0",X"F8",X"FC",X"FC",X"7C",X"3C",X"78",X"70",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"7C",X"3C",X"78",X"70",X"70",X"F0",X"E0",X"C0",X"00",
		X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"01",X"00",X"00",
		X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"C0",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"06",X"02",X"00",X"00",X"00",X"00",X"06",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"60",X"20",X"00",X"00",X"00",X"00",X"60",X"20",X"80",X"80",X"00",X"00",
		X"00",X"01",X"00",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"01",X"00",X"00",
		X"00",X"80",X"80",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"80",X"80",X"00",
		X"01",X"00",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"01",X"00",
		X"80",X"80",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"08",X"80",X"80",
		X"00",X"00",X"11",X"04",X"00",X"40",X"00",X"00",X"20",X"00",X"40",X"00",X"04",X"10",X"00",X"00",
		X"00",X"00",X"08",X"20",X"00",X"02",X"00",X"04",X"00",X"00",X"02",X"00",X"20",X"88",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"02",
		X"40",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"02",X"07",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",X"07",X"03",X"03",X"03",X"03",X"03",X"03",X"02",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"06",X"07",X"0F",X"1F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"F0",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",
		X"02",X"07",X"0F",X"1F",X"3F",X"7F",X"7D",X"78",X"70",X"60",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",
		X"00",X"80",X"C0",X"E0",X"F0",X"78",X"3C",X"3C",X"78",X"78",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",
		X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",
		X"00",X"80",X"C0",X"E0",X"F0",X"F0",X"78",X"78",X"78",X"70",X"F0",X"F0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"0F",X"1F",X"23",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"23",X"1F",X"0F",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"07",X"1F",X"3F",X"27",X"43",X"01",X"00",X"00",X"0C",X"0C",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"70",X"60",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"07",X"1F",X"3F",X"3F",X"67",X"43",X"41",X"40",X"40",X"20",X"20",X"19",X"07",X"00",
		X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",
		X"00",X"01",X"03",X"07",X"0C",X"18",X"20",X"43",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"A0",X"60",X"60",X"30",X"30",X"10",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"07",X"1C",X"30",X"43",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"1F",X"19",X"38",X"00",X"0C",X"04",X"04",X"06",X"02",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"1F",X"05",X"00",X"04",X"07",X"05",X"04",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"02",X"02",X"04",X"07",X"01",X"08",X"08",X"00",X"10",X"00",X"00",X"00",
		X"C0",X"C0",X"60",X"20",X"20",X"30",X"10",X"10",X"10",X"18",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"1D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"C0",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"18",X"0C",X"07",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"30",X"30",X"60",X"60",X"A0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"03",X"41",X"30",X"1C",X"07",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"06",X"04",X"07",X"0D",X"00",X"38",X"19",X"1F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"07",X"05",X"04",X"00",X"05",X"1F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"08",X"08",X"00",X"04",X"04",X"02",X"02",X"00",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"10",X"10",X"10",X"30",X"20",X"20",X"60",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"7F",X"80",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"7C",X"FC",X"FE",X"FE",X"FE",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"38",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"78",X"F8",X"FC",X"FC",X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"70",X"20",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"1C",X"3C",X"30",X"60",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"60",X"F0",X"F0",X"F0",X"78",X"78",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"1F",X"3F",X"63",X"83",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"78",X"F8",X"FC",X"FC",X"FC",X"FE",X"DE",X"1E",X"1E",X"0E",X"0E",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"1F",X"7F",X"86",X"06",X"06",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"7C",X"FC",X"FE",X"FE",X"FE",X"7E",X"7E",X"7E",X"7E",X"3C",X"3C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"1E",X"02",X"06",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"3E",X"3C",X"3C",X"3C",X"38",X"38",X"10",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"7C",X"1F",X"0F",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"1E",X"3C",X"3C",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"1F",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"7E",X"FE",X"FE",X"FE",X"FE",X"EE",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"7C",X"FE",X"BE",X"BE",X"9A",X"90",X"80",X"80",X"80",X"88",X"9A",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"B6",X"A4",X"A0",X"A0",X"A0",X"A2",X"B6",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"B8",X"B8",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BC",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"1E",X"1E",X"1E",X"1E",X"9E",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"2E",X"06",X"06",X"06",X"06",X"26",X"2E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"AA",X"80",X"90",X"98",X"80",X"82",X"86",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BA",X"B0",X"A4",X"A6",X"A0",X"A0",X"B0",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"B8",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"1E",X"1E",X"9E",X"1E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"AE",X"06",X"06",X"26",X"06",X"0E",X"1E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"80",X"80",X"82",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"B0",X"A0",X"A0",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BC",X"B8",X"B8",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"B6",X"A6",X"A6",X"A6",X"06",X"06",X"0E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"9C",X"90",X"80",X"80",X"80",X"80",X"82",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"B6",X"A4",X"A0",X"A0",X"A0",X"A0",X"A0",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BC",X"BC",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"9E",X"9E",X"9E",X"9E",X"1E",X"1E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"36",X"06",X"06",X"06",X"06",X"06",X"0E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"A2",X"80",X"80",X"98",X"80",X"80",X"82",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"B8",X"B0",X"A0",X"A6",X"A0",X"A0",X"A0",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"B8",X"B8",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BC",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"1E",X"1E",X"9E",X"1E",X"1E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"0E",X"06",X"06",X"26",X"06",X"06",X"0E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"AA",X"80",X"80",X"80",X"80",X"80",X"82",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BA",X"B0",X"A0",X"A0",X"A0",X"A0",X"A0",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BC",X"B8",X"B8",X"B8",X"B8",X"B8",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BC",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"1E",X"1E",X"1E",X"1E",X"1E",X"3E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"AE",X"06",X"06",X"06",X"06",X"06",X"0E",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"A6",X"B2",X"FA",X"FA",X"F8",X"FC",X"FE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"B8",X"BC",X"BE",X"B6",X"B2",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BC",X"BC",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"3E",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"3E",X"3E",X"BE",X"BE",X"9E",X"DE",X"FE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"7C",X"FE",X"BE",X"BE",X"1E",X"CE",X"EE",X"2E",X"26",X"F6",X"FE",X"BE",X"BE",X"BE",X"BE",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"60",X"60",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"CF",X"4F",X"7F",X"3F",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2A",X"55",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2A",X"55",X"2A",
		X"00",X"07",X"1F",X"13",X"17",X"38",X"28",X"38",X"34",X"20",X"20",X"1F",X"12",X"0F",X"07",X"00",
		X"00",X"C0",X"E0",X"30",X"B0",X"78",X"68",X"48",X"48",X"D8",X"B8",X"30",X"70",X"E0",X"80",X"00",
		X"00",X"21",X"1B",X"1F",X"0C",X"0A",X"18",X"10",X"14",X"1E",X"08",X"0D",X"0E",X"11",X"00",X"00",
		X"00",X"00",X"88",X"70",X"B0",X"50",X"18",X"08",X"48",X"58",X"10",X"30",X"F8",X"D8",X"84",X"00",
		X"81",X"63",X"3E",X"24",X"33",X"12",X"30",X"E0",X"34",X"14",X"12",X"10",X"36",X"2F",X"71",X"40",
		X"02",X"8E",X"F4",X"6C",X"08",X"48",X"08",X"2C",X"27",X"0C",X"48",X"0C",X"24",X"7C",X"C6",X"81",
		X"07",X"1F",X"1F",X"18",X"33",X"3E",X"68",X"6C",X"7C",X"78",X"76",X"33",X"38",X"0F",X"07",X"03",
		X"E0",X"F8",X"DC",X"E4",X"36",X"AE",X"16",X"16",X"1E",X"76",X"B6",X"EC",X"EC",X"F8",X"90",X"00",
		X"00",X"01",X"12",X"20",X"26",X"0C",X"08",X"00",X"20",X"20",X"34",X"12",X"08",X"03",X"00",X"00",
		X"00",X"90",X"18",X"08",X"28",X"10",X"02",X"06",X"14",X"14",X"28",X"00",X"18",X"30",X"00",X"00",
		X"03",X"00",X"06",X"28",X"40",X"40",X"00",X"00",X"00",X"40",X"40",X"10",X"00",X"00",X"04",X"03",
		X"40",X"00",X"00",X"08",X"04",X"00",X"08",X"08",X"00",X"00",X"04",X"04",X"28",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"0B",X"00",X"00",X"00",X"7E",X"42",X"02",X"12",X"A2",X"01",X"00",X"00",X"60",X"00",X"70",X"94",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"46",X"80",X"1E",X"B2",X"02",X"7E",X"00",
		X"10",X"90",X"90",X"14",X"80",X"00",X"4B",X"68",X"10",X"94",X"90",X"B4",X"00",X"00",X"A1",X"21",
		X"43",X"43",X"43",X"00",X"00",X"00",X"74",X"05",X"76",X"14",X"77",X"00",X"75",X"55",X"51",X"51",
		X"00",X"7D",X"45",X"45",X"7D",X"01",X"7D",X"45",X"00",X"E0",X"20",X"20",X"00",X"3C",X"00",X"28",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"00",X"0A",
		X"45",X"7D",X"01",X"5D",X"15",X"15",X"5D",X"01",X"28",X"28",X"28",X"28",X"00",X"3C",X"00",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"DD",X"55",X"DD",X"00",X"7E",X"42",X"02",X"12",X"22",X"61",X"E0",X"00",X"60",X"00",X"70",X"94",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"46",X"80",X"1E",X"B2",X"02",X"7E",X"00",
		X"10",X"90",X"90",X"14",X"80",X"00",X"4B",X"68",X"10",X"94",X"90",X"B4",X"00",X"00",X"A1",X"21",
		X"43",X"43",X"43",X"00",X"00",X"00",X"74",X"05",X"76",X"14",X"77",X"00",X"75",X"55",X"51",X"51",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A3",X"A3",X"20",X"A7",X"A7",X"27",X"07",X"07",
		X"62",X"62",X"06",X"F0",X"F7",X"F1",X"F1",X"F0",X"20",X"00",X"00",X"20",X"20",X"00",X"EA",X"20",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"07",X"27",X"A7",X"A7",X"27",X"A7",X"A7",X"27",
		X"F0",X"F0",X"F7",X"F0",X"F7",X"F1",X"F1",X"F7",X"2E",X"2A",X"EE",X"00",X"7E",X"42",X"4E",X"48",
		X"0B",X"00",X"00",X"00",X"7E",X"42",X"02",X"12",X"A3",X"03",X"03",X"03",X"63",X"01",X"71",X"95",
		X"60",X"60",X"60",X"60",X"B7",X"B7",X"B7",X"B3",X"48",X"78",X"00",X"78",X"08",X"C8",X"E0",X"F0",
		X"10",X"90",X"90",X"14",X"80",X"00",X"4B",X"68",X"11",X"94",X"90",X"B4",X"00",X"00",X"A1",X"21",
		X"DB",X"D9",X"D8",X"D8",X"D8",X"00",X"74",X"05",X"F8",X"F8",X"FC",X"7C",X"7E",X"3E",X"3E",X"00",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A0",X"A0",X"20",X"A0",X"A0",X"20",X"0F",X"0F",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E7",X"9E",X"7E",X"FC",X"F8",X"F2",X"E2",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"0F",X"2F",X"AF",X"AF",X"20",X"A7",X"AF",X"2F",
		X"FF",X"FE",X"F0",X"17",X"F1",X"F1",X"E1",X"EB",X"8A",X"0E",X"00",X"70",X"50",X"70",X"00",X"A8",
		X"0B",X"00",X"00",X"00",X"7E",X"42",X"02",X"12",X"AF",X"0F",X"1F",X"0E",X"68",X"00",X"70",X"94",
		X"C8",X"9B",X"1A",X"5A",X"DA",X"DB",X"D8",X"DB",X"00",X"F8",X"08",X"08",X"18",X"F8",X"00",X"78",
		X"10",X"90",X"90",X"14",X"80",X"00",X"4B",X"68",X"10",X"94",X"91",X"B5",X"01",X"01",X"A3",X"23",
		X"D9",X"DB",X"D8",X"B3",X"B1",X"B7",X"B0",X"66",X"48",X"78",X"00",X"70",X"50",X"70",X"00",X"60",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"0B",X"00",X"00",X"00",X"7E",X"42",X"02",X"12",X"A2",X"01",X"00",X"00",X"60",X"00",X"70",X"94",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"40",X"80",X"00",X"81",X"01",X"01",X"03",
		X"10",X"90",X"90",X"14",X"80",X"00",X"4B",X"68",X"10",X"94",X"90",X"B4",X"00",X"00",X"A0",X"20",
		X"43",X"43",X"43",X"00",X"01",X"07",X"0F",X"1F",X"03",X"03",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"0B",X"60",X"FE",X"FC",X"F8",X"F8",X"F1",X"F7",X"A2",X"01",X"08",X"1C",X"3E",X"7F",X"FF",X"FE",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"40",X"B0",X"3C",X"BF",X"3F",X"7F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E0",X"80",X"FC",X"F8",X"F0",X"C0",X"00",X"00",X"00",X"00",
		X"43",X"43",X"43",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"0B",X"00",X"00",X"00",X"00",X"E3",X"FF",X"FF",X"A2",X"01",X"08",X"1C",X"7E",X"FF",X"FE",X"FC",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"40",X"B0",X"3C",X"BF",X"3F",X"7F",X"3F",
		X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"F9",X"E1",X"05",X"77",X"00",X"00",X"00",X"00",
		X"43",X"43",X"43",X"00",X"06",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"12",
		X"0B",X"00",X"00",X"00",X"00",X"E3",X"FF",X"FF",X"A2",X"01",X"08",X"1C",X"7E",X"FF",X"FE",X"FC",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"22",X"4E",X"80",X"35",X"95",X"10",X"17",X"15",
		X"FF",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"F9",X"E1",X"05",X"77",X"00",X"00",X"00",X"00",
		X"43",X"43",X"43",X"00",X"06",X"00",X"00",X"00",X"77",X"00",X"07",X"05",X"BD",X"21",X"BF",X"00",
		X"4B",X"6B",X"C8",X"8B",X"6B",X"88",X"00",X"00",X"A1",X"A1",X"21",X"A1",X"80",X"3C",X"00",X"28",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"00",X"88",X"6B",X"8B",X"C8",X"6B",X"4B",X"28",X"28",X"28",X"A8",X"A8",X"00",X"BC",X"80",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"0B",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"A2",X"09",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"46",X"80",X"1E",X"B2",X"02",X"7E",X"00",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"FC",X"FC",X"FC",X"FE",X"FE",X"FC",X"FD",X"FD",
		X"43",X"43",X"43",X"00",X"00",X"00",X"74",X"05",X"76",X"14",X"77",X"00",X"75",X"55",X"51",X"51",
		X"0F",X"6F",X"4F",X"4F",X"47",X"77",X"07",X"77",X"FD",X"FD",X"FD",X"FD",X"80",X"BC",X"80",X"A8",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"47",X"47",X"43",X"7B",X"03",X"4B",X"03",X"01",X"A8",X"A8",X"A8",X"A8",X"80",X"BC",X"80",X"F4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"6D",X"29",X"6D",X"00",X"0E",X"08",X"08",X"0E",X"F2",X"F9",X"F8",X"FE",X"FF",X"FF",X"7F",X"7F",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"46",X"80",X"1E",X"B2",X"02",X"7E",X"00",
		X"03",X"0B",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"7F",X"7F",X"3F",X"BF",X"BF",X"BC",X"BD",X"9D",
		X"43",X"43",X"43",X"00",X"80",X"00",X"74",X"05",X"76",X"14",X"77",X"00",X"75",X"55",X"51",X"51",
		X"0F",X"0F",X"0F",X"07",X"02",X"01",X"03",X"01",X"DD",X"DD",X"DD",X"DD",X"00",X"BC",X"80",X"A8",
		X"74",X"75",X"04",X"74",X"00",X"00",X"00",X"00",X"95",X"B5",X"C0",X"5A",X"00",X"1E",X"00",X"0A",
		X"01",X"07",X"05",X"07",X"01",X"00",X"01",X"01",X"A8",X"A8",X"A8",X"A8",X"80",X"3C",X"80",X"C4",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"00",X"1E",X"00",X"10",
		X"01",X"00",X"07",X"07",X"0F",X"0F",X"0B",X"09",X"C2",X"09",X"EC",X"EE",X"EF",X"CF",X"1F",X"1F",
		X"00",X"00",X"80",X"00",X"43",X"00",X"43",X"43",X"20",X"46",X"80",X"1E",X"B2",X"02",X"7E",X"00",
		X"0F",X"00",X"6F",X"28",X"28",X"20",X"0B",X"28",X"1F",X"1F",X"9F",X"BF",X"BF",X"00",X"A1",X"21",
		X"43",X"43",X"43",X"00",X"00",X"00",X"74",X"05",X"76",X"14",X"77",X"00",X"75",X"55",X"51",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"DF",X"3F",X"FF",X"7F",X"FF",X"FF",
		X"5D",X"79",X"51",X"76",X"6A",X"F2",X"A4",X"A5",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",
		X"EE",X"B4",X"A4",X"E4",X"A7",X"BC",X"E4",X"A4",X"47",X"43",X"43",X"43",X"F3",X"4F",X"43",X"43",
		X"A4",X"E4",X"BC",X"A7",X"E4",X"A4",X"B4",X"EE",X"43",X"43",X"4F",X"F3",X"43",X"43",X"43",X"47",
		X"A5",X"A4",X"F2",X"6A",X"76",X"51",X"79",X"5D",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"FF",X"FF",X"7F",X"FF",X"3F",X"DF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",
		X"07",X"3F",X"D1",X"3F",X"C4",X"44",X"FE",X"89",X"FF",X"CB",X"2F",X"1F",X"BF",X"7F",X"7F",X"FF",
		X"5D",X"79",X"51",X"76",X"6A",X"F2",X"A4",X"A5",X"10",X"10",X"FD",X"23",X"21",X"21",X"21",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"B4",X"A4",X"E4",X"A7",X"BC",X"E4",X"A4",
		X"47",X"43",X"43",X"43",X"F3",X"4F",X"43",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",
		X"A4",X"E4",X"BC",X"A7",X"E4",X"A4",X"B4",X"EE",X"43",X"43",X"4F",X"F3",X"43",X"43",X"43",X"47",
		X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A5",X"A4",X"F2",X"6A",X"76",X"51",X"79",X"5D",
		X"FB",X"21",X"21",X"21",X"23",X"FD",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"89",X"FE",X"44",X"C4",X"3F",X"D1",X"3F",X"07",
		X"FF",X"7F",X"7F",X"BF",X"1F",X"2F",X"CB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"0B",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"DF",
		X"07",X"3F",X"D1",X"3F",X"C4",X"44",X"FE",X"89",X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",
		X"FC",X"37",X"2D",X"59",X"6F",X"5A",X"72",X"54",X"FF",X"BF",X"3F",X"3F",X"C8",X"88",X"88",X"9F",
		X"10",X"10",X"FD",X"23",X"21",X"21",X"21",X"FB",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A7",X"BD",X"E9",X"A9",X"A9",X"FF",X"A9",X"E9",X"F0",X"10",X"10",X"11",X"FF",X"1F",X"1F",X"1F",
		X"46",X"42",X"42",X"42",X"F2",X"4E",X"42",X"42",X"00",X"00",X"00",X"07",X"0F",X"12",X"1F",X"14",
		X"A9",X"9F",X"F7",X"78",X"88",X"9F",X"F1",X"91",X"FF",X"7F",X"FF",X"F7",X"E7",X"47",X"27",X"17",
		X"42",X"42",X"4E",X"F2",X"42",X"42",X"42",X"46",X"14",X"1F",X"12",X"0F",X"07",X"00",X"00",X"00",
		X"91",X"F1",X"9F",X"88",X"78",X"F7",X"9F",X"A9",X"17",X"27",X"47",X"E7",X"F7",X"FF",X"7F",X"FF",
		X"FB",X"21",X"21",X"21",X"23",X"FD",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"E9",X"A9",X"FF",X"A9",X"A9",X"E9",X"BD",X"A7",X"1F",X"1F",X"1F",X"FF",X"11",X"10",X"10",X"F0",
		X"89",X"FE",X"44",X"C4",X"3F",X"D1",X"3F",X"07",X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",
		X"54",X"72",X"5A",X"6F",X"59",X"2D",X"37",X"FC",X"9F",X"88",X"88",X"C8",X"3F",X"3F",X"BF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"DF",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"D5",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",
		X"FF",X"A4",X"24",X"3F",X"C8",X"88",X"88",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"10",X"10",X"11",X"FE",X"1A",X"11",X"11",X"FF",X"8F",X"8F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"EB",X"47",X"8F",X"97",X"A7",X"47",X"27",X"17",X"FF",X"FF",X"FE",X"FC",X"FC",X"FD",X"FE",X"FC",
		X"17",X"27",X"47",X"A7",X"97",X"8F",X"47",X"EB",X"FC",X"FE",X"FD",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"11",X"11",X"1A",X"FE",X"11",X"10",X"10",X"F0",X"FF",X"FF",X"FF",X"7F",X"FF",X"8F",X"8F",X"FF",
		X"9F",X"88",X"88",X"C8",X"3F",X"24",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D5",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"D5",X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"56",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",X"A4",X"24",X"3F",X"C8",X"88",X"88",X"9F",
		X"A9",X"FC",X"96",X"95",X"F2",X"9E",X"8B",X"89",X"7F",X"FF",X"7F",X"FF",X"7F",X"3F",X"BF",X"7F",
		X"F0",X"10",X"10",X"11",X"FE",X"1A",X"11",X"11",X"F9",X"8F",X"89",X"F9",X"65",X"82",X"02",X"03",
		X"3F",X"3F",X"DF",X"7F",X"7F",X"FF",X"FF",X"FF",X"EA",X"46",X"8C",X"94",X"A4",X"44",X"24",X"14",
		X"03",X"03",X"02",X"04",X"04",X"05",X"06",X"04",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"77",X"73",
		X"14",X"24",X"44",X"A4",X"94",X"8C",X"46",X"EA",X"04",X"06",X"05",X"04",X"04",X"02",X"03",X"03",
		X"73",X"77",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"11",X"11",X"1A",X"FE",X"11",X"10",X"10",X"F0",
		X"03",X"02",X"82",X"65",X"F9",X"89",X"8F",X"F9",X"FF",X"FF",X"FF",X"7F",X"7F",X"DF",X"3F",X"3F",
		X"9F",X"88",X"88",X"C8",X"3F",X"24",X"A4",X"FF",X"89",X"8B",X"9E",X"F2",X"95",X"96",X"FC",X"A9",
		X"7F",X"BF",X"3F",X"7F",X"FF",X"7F",X"FF",X"7F",X"D5",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"56",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",X"A9",X"FC",X"96",X"95",X"F2",X"9E",X"8B",X"89",
		X"5F",X"E7",X"5F",X"C7",X"7F",X"23",X"A3",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"F9",X"8F",X"89",X"F9",X"65",X"82",X"02",X"03",X"21",X"20",X"D0",X"6B",X"55",X"AD",X"AB",X"29",
		X"F8",X"F8",X"FF",X"FE",X"22",X"11",X"91",X"9F",X"03",X"03",X"02",X"04",X"04",X"05",X"06",X"04",
		X"49",X"56",X"D3",X"52",X"D2",X"5A",X"57",X"52",X"68",X"48",X"44",X"A4",X"7F",X"A4",X"24",X"24",
		X"04",X"06",X"05",X"04",X"04",X"02",X"03",X"03",X"52",X"57",X"5A",X"D2",X"52",X"D3",X"56",X"49",
		X"24",X"24",X"A4",X"7F",X"A4",X"44",X"48",X"68",X"03",X"02",X"82",X"65",X"F9",X"89",X"8F",X"F9",
		X"29",X"AB",X"AD",X"55",X"6B",X"D0",X"20",X"21",X"9F",X"91",X"11",X"22",X"FE",X"FF",X"F8",X"F8",
		X"89",X"8B",X"9E",X"F2",X"95",X"96",X"FC",X"A9",X"7F",X"A3",X"23",X"7F",X"C7",X"5F",X"E7",X"5F",
		X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"56",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"5F",X"E4",X"5F",X"C4",X"7F",X"22",X"A2",X"7F",
		X"CF",X"7F",X"C7",X"7F",X"C7",X"23",X"2F",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"03",
		X"21",X"20",X"D0",X"6B",X"55",X"AD",X"AB",X"29",X"08",X"88",X"87",X"FE",X"22",X"11",X"91",X"9F",
		X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",X"49",X"56",X"D3",X"52",X"D2",X"5A",X"57",X"52",
		X"68",X"48",X"44",X"A4",X"7F",X"A4",X"24",X"24",X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",
		X"52",X"57",X"5A",X"D2",X"52",X"D3",X"56",X"49",X"24",X"24",X"A4",X"7F",X"A4",X"44",X"48",X"68",
		X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",X"29",X"AB",X"AD",X"55",X"6B",X"D0",X"20",X"21",
		X"9F",X"91",X"11",X"22",X"FE",X"87",X"88",X"08",X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",
		X"7F",X"A2",X"22",X"7F",X"C4",X"5F",X"E4",X"5F",X"F1",X"2F",X"23",X"C7",X"7F",X"C7",X"7F",X"CF",
		X"03",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",X"00",X"00",X"00",X"00",X"00",X"0F",X"F7",X"17",
		X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",X"C8",X"7F",X"C4",X"7F",X"C4",X"22",X"2F",X"F1",
		X"79",X"8B",X"3D",X"C4",X"03",X"0E",X"F2",X"02",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"08",X"88",X"87",X"FE",X"22",X"11",X"91",X"9F",X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",
		X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",X"68",X"48",X"44",X"A4",X"7F",X"A4",X"24",X"24",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"24",X"24",X"A4",X"7F",X"A4",X"44",X"48",X"68",X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",
		X"BF",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"9F",X"91",X"11",X"22",X"FE",X"87",X"88",X"08",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"F1",X"2F",X"22",X"C4",X"7F",X"C4",X"7F",X"C8",X"02",X"F2",X"0E",X"03",X"C4",X"3D",X"8B",X"79",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"17",X"F7",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"79",X"8B",X"3D",X"C4",X"03",X"0E",X"F2",X"02",X"6F",X"FF",X"7F",X"BF",X"FF",X"BF",X"AF",X"9F",
		X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",X"F7",X"5F",X"57",X"4F",X"4F",X"EB",X"3B",X"2F",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"AB",X"AB",X"AB",X"FB",X"AF",X"AB",X"AB",X"AB",
		X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",X"AB",X"AB",X"AB",X"AF",X"FB",X"AB",X"AB",X"AB",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"2F",X"3B",X"EB",X"4F",X"4F",X"57",X"5F",X"F7",
		X"02",X"F2",X"0E",X"03",X"C4",X"3D",X"8B",X"79",X"9F",X"AF",X"BF",X"FF",X"BF",X"7F",X"FF",X"6F",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"6B",X"F4",X"7C",X"B3",X"F6",X"B9",X"A9",X"9B",X"FF",X"FF",X"FF",X"3F",X"3D",X"70",X"90",X"10",
		X"F4",X"5C",X"54",X"4D",X"4E",X"EA",X"3A",X"2E",X"8F",X"B8",X"C8",X"84",X"44",X"47",X"7C",X"C4",
		X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",X"44",X"44",X"44",X"45",X"7E",X"C4",X"44",X"44",
		X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",X"44",X"44",X"C4",X"7E",X"45",X"44",X"44",X"44",
		X"2E",X"3A",X"EA",X"4E",X"4D",X"54",X"5C",X"F4",X"C4",X"7C",X"47",X"44",X"84",X"C8",X"B8",X"8F",
		X"9B",X"A9",X"B9",X"F6",X"B3",X"7C",X"F4",X"6B",X"10",X"90",X"70",X"3D",X"3F",X"FF",X"FF",X"FF",
		X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",X"00",X"00",X"07",X"18",X"73",X"9C",X"28",X"C7",
		X"00",X"C0",X"40",X"60",X"A0",X"10",X"70",X"88",X"6B",X"F4",X"7C",X"B3",X"F6",X"B9",X"A9",X"9B",
		X"0E",X"B2",X"C1",X"23",X"3D",X"70",X"90",X"10",X"08",X"08",X"78",X"84",X"04",X"84",X"8E",X"F2",
		X"F4",X"5C",X"54",X"4D",X"4E",X"EA",X"3A",X"2E",X"8F",X"B8",X"C8",X"84",X"44",X"47",X"7C",X"C4",
		X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",
		X"44",X"44",X"44",X"45",X"7E",X"C4",X"44",X"44",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",X"44",X"44",X"C4",X"7E",X"45",X"44",X"44",X"44",
		X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"2E",X"3A",X"EA",X"4E",X"4D",X"54",X"5C",X"F4",
		X"C4",X"7C",X"47",X"44",X"84",X"C8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"9B",X"A9",X"B9",X"F6",X"B3",X"7C",X"F4",X"6B",X"10",X"90",X"70",X"3D",X"23",X"C1",X"B2",X"0E",
		X"F2",X"8E",X"84",X"04",X"84",X"78",X"08",X"08",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"28",X"9C",X"73",X"18",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"60",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1E",X"7F",X"3C",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"10",X"18",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"1C",X"0C",X"0E",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"1C",X"1E",X"1E",X"0E",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"14",X"22",X"41",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"C8",X"88",X"88",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"03",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"84",X"04",X"84",X"8E",X"F2",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"FE",X"FC",X"FD",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"E9",X"A9",X"A9",X"FF",X"A9",X"E9",
		X"F0",X"10",X"10",X"11",X"FF",X"1F",X"1F",X"1F",X"FF",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FF",X"FE",X"E2",X"F1",X"F1",X"FF",
		X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",
		X"FF",X"F8",X"C8",X"84",X"C4",X"C7",X"FC",X"C4",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"FE",X"F4",X"E4",X"E4",X"E7",X"FC",X"E4",X"E4",X"47",X"43",X"43",X"43",X"F3",X"4F",X"43",X"43",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"A9",X"9F",X"F7",X"FF",X"FF",X"FF",X"F1",X"91",
		X"FF",X"FF",X"FF",X"F7",X"E7",X"47",X"27",X"17",X"FF",X"FF",X"FE",X"FC",X"FC",X"FD",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"77",X"73",X"F8",X"F8",X"FC",X"FC",X"FF",X"FC",X"FC",X"FC",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"C5",X"FE",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"E4",X"E4",X"FC",X"E7",X"E4",X"E4",X"F4",X"FE",X"43",X"43",X"4F",X"F3",X"43",X"43",X"43",X"47",
		X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"91",X"F1",X"FF",X"FF",X"FF",X"F7",X"9F",X"A9",
		X"17",X"27",X"47",X"E7",X"F7",X"FF",X"FF",X"FF",X"FC",X"FE",X"FD",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"73",X"77",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FF",X"FC",X"FC",X"F8",X"F8",
		X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",X"BF",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"FE",X"C5",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"FD",X"FC",X"FE",X"7E",X"7E",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"A9",X"FF",X"A9",X"A9",X"E9",X"FD",X"FF",
		X"1F",X"1F",X"1F",X"FF",X"11",X"10",X"10",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F1",X"E2",X"FE",X"FF",X"F8",X"F8",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"C4",X"FC",X"C7",X"C4",X"84",X"C8",X"F8",X"FF",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9F",X"88",X"88",X"C8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"F0",X"F0",X"F0",X"FD",X"FF",X"FF",X"FF",X"FF",X"F2",X"8E",X"84",X"04",X"84",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"C8",X"90",X"90",X"7F",X"FF",X"FF",X"FF",X"FF",X"9F",X"8F",X"4F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"03",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"84",X"04",X"84",X"8E",X"F2",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"FE",X"FC",X"FD",X"FF",X"FF",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"E9",X"A9",X"AB",X"FD",X"A9",X"E9",
		X"90",X"10",X"10",X"11",X"FF",X"1F",X"1F",X"1F",X"4F",X"47",X"47",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FF",X"FE",X"F2",X"F9",X"F9",X"FF",
		X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",
		X"FF",X"F8",X"C8",X"84",X"C4",X"C7",X"FC",X"C4",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"FE",X"F4",X"E4",X"E4",X"E7",X"FC",X"E4",X"E4",X"47",X"43",X"43",X"43",X"F3",X"4F",X"43",X"43",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F4",X"A9",X"9F",X"F7",X"FF",X"FF",X"FF",X"F1",X"91",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"4F",X"2F",X"2F",X"FF",X"FF",X"FE",X"FC",X"FC",X"FD",X"FE",X"FC",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"7D",X"7D",X"7C",X"FC",X"FC",X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"C5",X"FE",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"E4",X"E4",X"FC",X"E7",X"E4",X"E4",X"F4",X"FE",X"43",X"43",X"4F",X"F3",X"43",X"43",X"43",X"47",
		X"F4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"91",X"F1",X"FF",X"FF",X"FF",X"F7",X"9F",X"A9",
		X"2F",X"2F",X"4F",X"EF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FD",X"FC",X"FC",X"FE",X"FF",X"FF",
		X"7C",X"7D",X"7D",X"FF",X"7F",X"7F",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",X"BF",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"FE",X"C5",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"FD",X"FC",X"FE",X"7E",X"7E",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",X"3F",X"3F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"A9",X"FD",X"AB",X"A9",X"E9",X"FD",X"FF",
		X"1F",X"1F",X"1F",X"FF",X"11",X"10",X"10",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"47",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"F2",X"FE",X"FF",X"F8",X"F8",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"C4",X"FC",X"C7",X"C4",X"84",X"C8",X"F8",X"FF",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"90",X"90",X"C8",X"FF",X"FF",X"FF",X"FF",X"FF",X"4F",X"8F",X"9F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"F0",X"F0",X"F0",X"FD",X"FF",X"FF",X"FF",X"FF",X"F2",X"8E",X"84",X"04",X"84",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"48",X"88",X"88",X"FF",X"10",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"FF",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"83",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"84",X"04",X"84",X"8E",X"F2",
		X"7F",X"7F",X"7F",X"7C",X"7C",X"FC",X"F8",X"F9",X"FF",X"FF",X"FF",X"3F",X"7F",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"E9",X"CA",X"D2",X"D3",X"FE",X"D2",X"D2",
		X"10",X"10",X"10",X"17",X"FF",X"3F",X"7F",X"7F",X"27",X"27",X"23",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FF",X"FE",X"E1",X"F1",X"F8",X"FF",
		X"43",X"2E",X"F1",X"11",X"09",X"09",X"BF",X"C9",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",
		X"FF",X"F8",X"C8",X"84",X"C4",X"C7",X"FC",X"C4",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"FE",X"F8",X"E8",X"E8",X"EF",X"F8",X"E8",X"E8",X"87",X"87",X"87",X"87",X"F7",X"8F",X"87",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"D2",X"DF",X"F7",X"FF",X"FE",X"FE",X"A2",X"22",
		X"FF",X"FF",X"FF",X"EF",X"CF",X"8F",X"4F",X"2F",X"FF",X"FE",X"FE",X"FC",X"FD",X"FE",X"FC",X"FC",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"44",X"44",X"24",X"3F",X"E2",X"22",X"22",X"22",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"C5",X"FE",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"E8",X"E8",X"F8",X"EF",X"E8",X"E8",X"F8",X"FE",X"87",X"87",X"8F",X"F7",X"87",X"87",X"87",X"87",
		X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"22",X"A2",X"FE",X"FE",X"FF",X"F7",X"DF",X"D2",
		X"2F",X"4F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FD",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",
		X"22",X"22",X"22",X"E2",X"3F",X"24",X"44",X"44",X"BF",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"FE",X"C5",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"F9",X"F8",X"FC",X"7C",X"7C",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"3F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D2",X"D2",X"FE",X"D3",X"D2",X"CA",X"E9",X"F9",
		X"7F",X"7F",X"3F",X"FF",X"17",X"10",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FB",X"23",X"27",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F1",X"E1",X"FE",X"FF",X"FC",X"F8",
		X"C9",X"BF",X"09",X"09",X"11",X"F1",X"2E",X"43",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"C4",X"FC",X"C7",X"C4",X"84",X"C8",X"F8",X"FF",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"10",X"FF",X"88",X"88",X"48",X"FF",X"FF",X"FF",X"27",X"FF",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"F0",X"F0",X"F0",X"FD",X"FF",X"FF",X"FF",X"FF",X"F2",X"8E",X"84",X"04",X"84",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"48",X"88",X"88",X"FF",X"10",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"FF",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"83",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"84",X"04",X"84",X"8E",X"F2",
		X"7F",X"7F",X"7F",X"7C",X"7C",X"FC",X"F8",X"F9",X"FF",X"FF",X"FF",X"3F",X"7F",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"E9",X"CA",X"D2",X"D3",X"FE",X"D2",X"D2",
		X"10",X"10",X"10",X"17",X"FF",X"3F",X"7F",X"7F",X"27",X"27",X"23",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FF",X"FD",X"F1",X"F8",X"F8",X"FF",
		X"43",X"2E",X"F1",X"11",X"09",X"89",X"BF",X"C9",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"3F",X"3F",
		X"FF",X"F8",X"C8",X"84",X"C4",X"C7",X"FC",X"C4",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"FE",X"F8",X"E8",X"E8",X"EF",X"F8",X"E8",X"E8",X"87",X"87",X"87",X"87",X"F7",X"8F",X"87",X"87",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"D2",X"DF",X"F7",X"FF",X"FE",X"FE",X"A2",X"22",
		X"FF",X"FF",X"FF",X"EF",X"CF",X"8F",X"4F",X"2F",X"FF",X"FE",X"FE",X"FC",X"FD",X"FE",X"FC",X"FC",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"24",X"24",X"3F",X"E2",X"92",X"92",X"92",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"C5",X"FE",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"E8",X"E8",X"F8",X"EF",X"E8",X"E8",X"F8",X"FE",X"87",X"87",X"8F",X"F7",X"87",X"87",X"87",X"87",
		X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"22",X"A2",X"FE",X"FE",X"FF",X"F7",X"DF",X"D2",
		X"2F",X"4F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FD",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"92",X"92",X"92",X"E2",X"3F",X"24",X"24",X"44",X"BF",X"BF",X"BF",X"BF",X"FF",X"BF",X"BF",X"BF",
		X"C4",X"C4",X"C4",X"FE",X"C5",X"C4",X"C4",X"C4",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"F9",X"F8",X"FC",X"7C",X"7C",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"3F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D2",X"D2",X"FE",X"D3",X"D2",X"CA",X"E9",X"F9",
		X"7F",X"7F",X"3F",X"FF",X"17",X"10",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FB",X"23",X"27",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F1",X"FD",X"FF",X"FC",X"F8",
		X"C9",X"BF",X"89",X"09",X"11",X"F1",X"2E",X"43",X"3F",X"3F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",
		X"C4",X"FC",X"C7",X"C4",X"84",X"C8",X"F8",X"FF",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"10",X"FF",X"88",X"88",X"48",X"FF",X"FF",X"FF",X"27",X"FF",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"F0",X"F0",X"F0",X"FD",X"FF",X"FF",X"FF",X"FF",X"F2",X"8E",X"84",X"04",X"84",X"F8",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",
		X"F1",X"80",X"F8",X"B8",X"B9",X"80",X"B0",X"B0",X"B0",X"B0",X"B1",X"80",X"B8",X"B8",X"B9",X"8F",
		X"00",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FE",X"36",X"00",X"C1",X"81",X"01",X"01",X"05",X"05",
		X"8F",X"01",X"01",X"FF",X"01",X"01",X"37",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"C6",
		X"7E",X"78",X"E1",X"81",X"01",X"01",X"05",X"05",X"7D",X"01",X"83",X"FF",X"1F",X"1F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"80",X"00",X"78",X"7C",X"6C",X"00",X"01",X"81",X"03",X"03",X"03",X"01",
		X"77",X"01",X"01",X"FF",X"1D",X"0D",X"2D",X"2D",X"00",X"00",X"00",X"00",X"80",X"00",X"60",X"72",
		X"31",X"00",X"80",X"47",X"22",X"12",X"9E",X"F9",X"31",X"01",X"40",X"CC",X"41",X"40",X"44",X"49",
		X"00",X"00",X"01",X"88",X"40",X"81",X"01",X"01",X"08",X"00",X"01",X"21",X"00",X"00",X"83",X"81",
		X"31",X"10",X"88",X"47",X"20",X"00",X"0C",X"69",X"39",X"01",X"00",X"CC",X"43",X"40",X"44",X"4B",
		X"60",X"00",X"0F",X"88",X"00",X"01",X"09",X"09",X"08",X"00",X"01",X"21",X"00",X"04",X"83",X"81",
		X"31",X"00",X"00",X"47",X"20",X"00",X"0C",X"69",X"39",X"67",X"44",X"CC",X"01",X"00",X"40",X"43",
		X"38",X"83",X"C2",X"FA",X"7E",X"70",X"7F",X"F8",X"22",X"81",X"40",X"42",X"60",X"60",X"28",X"28",
		X"0A",X"01",X"00",X"6A",X"40",X"00",X"22",X"62",X"28",X"00",X"01",X"6A",X"01",X"00",X"8A",X"42",
		X"7A",X"FB",X"FA",X"FA",X"7C",X"60",X"6D",X"68",X"68",X"01",X"02",X"42",X"7E",X"EE",X"2A",X"2A",
		X"62",X"03",X"0A",X"6A",X"02",X"00",X"68",X"68",X"28",X"00",X"01",X"6A",X"0B",X"02",X"E2",X"60",
		X"72",X"01",X"00",X"FA",X"7C",X"60",X"6D",X"68",X"6A",X"EF",X"42",X"42",X"0C",X"08",X"20",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"9F",
		X"FF",X"FF",X"FF",X"C5",X"91",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"3F",X"FF",X"FE",X"FD",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FE",
		X"FF",X"FF",X"F0",X"E7",X"FF",X"FF",X"F8",X"3F",X"F7",X"EF",X"3F",X"FF",X"FF",X"FF",X"5F",X"CF",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"FF",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"07",X"01",X"00",X"00",X"07",X"07",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"F1",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"DC",X"EC",X"FE",X"F7",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"57",X"07",X"04",X"FB",X"F7",X"06",X"17",X"17",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"FE",X"F8",
		X"7F",X"3F",X"BF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"F0",X"FF",X"FF",X"FF",
		X"07",X"00",X"07",X"1F",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FA",X"F8",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"DF",X"E7",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"BF",X"CF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"CF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"FF",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"DF",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"18",X"1F",X"7F",X"01",X"F0",X"FF",X"F9",X"E0",X"00",X"BF",
		X"FF",X"FF",X"7F",X"1F",X"8F",X"63",X"10",X"98",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"1F",X"03",
		X"FF",X"FF",X"FB",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"7F",X"10",X"04",X"05",X"00",X"03",X"00",X"FF",X"D7",X"FF",X"7C",X"7E",X"FF",X"FF",X"BE",
		X"FC",X"FD",X"7C",X"7B",X"F3",X"E7",X"0F",X"1E",X"00",X"00",X"80",X"80",X"C0",X"DC",X"9F",X"3F",
		X"FF",X"1F",X"01",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"80",X"C0",X"F0",X"F8",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"3F",X"FF",X"00",X"00",X"37",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"60",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"80",X"7F",X"FF",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"38",X"DB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E3",X"81",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"7F",
		X"BE",X"CF",X"FC",X"FF",X"F7",X"FF",X"FF",X"FF",X"00",X"C0",X"3C",X"83",X"F0",X"70",X"F0",X"FF",
		X"FF",X"FE",X"FE",X"FC",X"F8",X"F0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",
		X"1F",X"0F",X"00",X"00",X"1C",X"0F",X"4F",X"5F",X"FF",X"FF",X"3F",X"1F",X"03",X"F0",X"F8",X"98",
		X"FE",X"FF",X"FD",X"F8",X"F3",X"00",X"01",X"3F",X"FF",X"FF",X"DF",X"67",X"F7",X"FB",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"3E",X"3F",X"3F",X"1F",X"0F",X"00",X"00",X"02",
		X"7E",X"E0",X"FF",X"FE",X"78",X"5F",X"5F",X"1F",X"08",X"45",X"FF",X"FF",X"4F",X"CF",X"FE",X"F0",
		X"1F",X"0F",X"BF",X"3F",X"3F",X"0F",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F8",X"FC",X"FC",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C1",X"FF",X"FF",
		X"1F",X"3C",X"00",X"03",X"1F",X"FF",X"FF",X"FF",X"E0",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"C7",X"FE",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"3F",X"9C",X"DE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"40",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"3F",X"FF",X"80",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",
		X"78",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"03",X"03",X"83",X"C3",X"E3",X"E1",
		X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",
		X"F1",X"F1",X"F9",X"F9",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"1B",X"1B",X"17",X"17",X"0F",X"0E",X"00",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",
		X"3F",X"FB",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"1F",X"1C",X"3C",X"38",X"18",X"20",X"20",X"10",
		X"1F",X"8F",X"CF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"E3",X"E3",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"F7",X"F7",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"1F",X"1C",X"14",X"24",X"04",X"08",X"08",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"10",X"10",X"42",X"42",X"21",X"21",X"21",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"5E",
		X"C1",X"C1",X"C0",X"A0",X"20",X"10",X"50",X"48",X"FB",X"FB",X"FF",X"DD",X"5E",X"6E",X"2F",X"37",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"10",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"12",X"11",X"09",X"29",X"08",X"04",X"04",X"02",X"02",X"01",X"01",
		X"4C",X"24",X"20",X"28",X"28",X"04",X"04",X"04",X"28",X"24",X"14",X"12",X"22",X"25",X"45",X"42",
		X"17",X"1B",X"4B",X"8F",X"27",X"4F",X"1F",X"97",X"BF",X"BF",X"DF",X"DF",X"FF",X"FF",X"DF",X"CF",
		X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"10",X"10",X"00",X"41",X"41",X"29",
		X"81",X"81",X"81",X"81",X"82",X"02",X"12",X"12",X"05",X"09",X"48",X"48",X"20",X"20",X"10",X"90",
		X"02",X"04",X"84",X"80",X"40",X"40",X"20",X"20",X"A3",X"43",X"01",X"01",X"40",X"00",X"00",X"00",
		X"EF",X"E7",X"F7",X"F3",X"FB",X"F9",X"7D",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"BF",
		X"00",X"00",X"80",X"80",X"C0",X"C1",X"E7",X"EF",X"00",X"00",X"06",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"29",X"24",X"24",X"22",X"42",X"42",X"42",X"42",X"08",X"08",X"04",X"04",X"04",X"04",X"04",X"04",
		X"90",X"50",X"50",X"20",X"20",X"20",X"30",X"70",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"06",X"05",X"03",X"02",X"3E",X"3E",X"1F",X"1F",X"8F",X"8F",X"40",X"CF",
		X"BF",X"5F",X"5F",X"3F",X"BF",X"FF",X"00",X"FF",X"F7",X"F7",X"FB",X"FB",X"FD",X"FD",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"C0",X"E0",X"E0",X"F0",X"F0",X"E0",X"C0",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",
		X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"01",X"01",X"01",
		X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"BE",X"BC",X"D8",X"D0",X"E0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"0E",X"1E",X"1E",X"1E",X"1C",X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"81",X"C0",X"E0",X"F1",X"F9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"FF",X"FF",X"FF",X"FF",X"EF",X"CF",X"DF",X"DF",X"DF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"FD",X"FD",X"FD",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"FC",X"F8",X"F8",X"FC",X"FC",X"FF",X"3F",X"1F",X"11",X"18",X"18",X"30",X"70",X"E0",
		X"E2",X"C1",X"C1",X"81",X"81",X"43",X"47",X"3E",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",
		X"00",X"00",X"00",X"16",X"17",X"23",X"23",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",
		X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",X"FF",X"FF",X"FF",X"7F",X"3F",X"3F",X"3F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"FF",X"FF",X"F6",X"F6",X"F3",X"F3",X"E1",X"E1",X"FF",X"FF",X"FF",X"FF",X"7F",X"5F",X"BF",X"BF",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"3F",X"03",X"01",X"01",X"00",X"00",
		X"80",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"C0",
		X"BF",X"DF",X"7F",X"7F",X"7F",X"7F",X"77",X"77",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0E",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"77",X"77",X"F7",X"EF",X"EF",X"EF",X"EF",X"FF",
		X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"7F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"81",X"81",X"C1",X"C1",X"E1",X"E1",X"F3",X"F3",
		X"FF",X"FF",X"FF",X"DF",X"DF",X"DF",X"8F",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"87",X"87",X"87",X"CF",X"FF",X"77",X"07",X"07",
		X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8B",X"8B",X"D7",X"D7",X"DF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"4E",X"CF",X"A7",X"67",X"D0",X"B3",X"67",X"4F",
		X"1F",X"E1",X"FE",X"FF",X"00",X"FF",X"FF",X"FF",X"FD",X"FD",X"1D",X"E1",X"00",X"FF",X"FF",X"FF",
		X"00",X"80",X"80",X"C0",X"00",X"E0",X"E0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"1F",X"03",X"01",X"01",X"00",X"00",X"FB",X"F3",X"F7",X"F7",X"F7",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"07",X"BF",X"3F",X"7F",X"7F",X"7F",X"FF",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"04",X"06",X"06",X"0C",X"1C",X"F8",X"70",X"00",
		X"70",X"20",X"20",X"10",X"11",X"0F",X"07",X"00",X"40",X"60",X"60",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"13",X"0D",X"9E",X"A6",X"01",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"10",X"16",X"23",X"23",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"13",X"0D",X"9E",X"86",X"01",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"10",X"16",X"23",X"23",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"23",X"21",X"09",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"01",X"0D",X"86",X"87",X"06",X"0C",X"1C",X"3C",
		X"E0",X"E0",X"F0",X"60",X"E0",X"60",X"60",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"3E",X"3F",X"27",X"02",X"21",X"31",X"31",X"31",
		X"18",X"18",X"0C",X"8C",X"C6",X"F6",X"E6",X"F6",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"10",X"17",X"9F",X"BE",X"B2",X"B3",X"81",X"01",
		X"F6",X"94",X"1C",X"0C",X"0C",X"0C",X"8C",X"58",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"01",X"01",X"02",X"10",X"14",X"22",X"23",X"21",
		X"68",X"68",X"30",X"18",X"18",X"0C",X"10",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"09",X"0A",X"00",X"20",X"43",X"4D",X"CE",X"9F",X"1F",X"1D",X"9C",X"BE",
		X"E0",X"E0",X"F0",X"60",X"60",X"A4",X"A6",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2E",X"3F",X"3F",X"7F",X"7E",X"7E",X"3F",X"3F",X"3E",
		X"39",X"98",X"C0",X"F0",X"FA",X"FA",X"FA",X"F6",X"80",X"80",X"00",X"00",X"00",X"01",X"01",X"01",
		X"13",X"13",X"92",X"92",X"C0",X"C0",X"E0",X"E1",X"1E",X"9F",X"BF",X"BE",X"BE",X"FF",X"BF",X"3F",
		X"F6",X"F4",X"EC",X"E6",X"E3",X"C3",X"C2",X"64",X"01",X"03",X"03",X"43",X"67",X"67",X"67",X"27",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"23",X"27",X"27",X"11",X"16",X"23",X"23",X"20",
		X"68",X"F8",X"F0",X"A0",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"81",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"18",X"04",X"00",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"8F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"21",X"30",X"1C",X"08",X"08",X"00",X"20",X"83",X"0D",X"8E",X"9F",X"1F",X"1F",X"1F",X"3F",
		X"E0",X"30",X"32",X"33",X"19",X"99",X"8C",X"0C",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"3F",X"3F",X"3F",X"3E",X"7E",X"7F",X"3F",X"1E",
		X"48",X"F8",X"E0",X"F0",X"FA",X"FA",X"FA",X"F6",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"94",X"94",X"84",X"C0",X"E0",X"E1",X"0E",X"0F",X"BF",X"BE",X"BE",X"BF",X"9F",X"1F",
		X"F6",X"F4",X"EC",X"E8",X"E8",X"EC",X"EA",X"76",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"27",
		X"F1",X"F1",X"E3",X"C2",X"21",X"11",X"12",X"02",X"03",X"07",X"07",X"11",X"76",X"E3",X"E3",X"21",
		X"6E",X"EE",X"EE",X"AC",X"08",X"00",X"80",X"E0",X"27",X"27",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"04",X"04",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"02",X"8F",X"87",X"C3",X"C6",X"60",X"20",
		X"70",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"11",X"10",X"10",X"11",X"09",X"08",X"09",X"4B",X"C7",X"E7",X"AF",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"03",X"0D",X"8E",X"9F",X"1F",X"1F",X"1F",X"3F",
		X"E2",X"E3",X"F1",X"61",X"60",X"A0",X"A0",X"30",X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"C0",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"3F",X"3F",X"3F",X"3E",X"7E",X"7F",X"3F",X"1E",
		X"58",X"E8",X"E0",X"F0",X"FA",X"FA",X"FA",X"F6",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"13",X"96",X"96",X"C2",X"C0",X"E0",X"E1",X"0E",X"0F",X"BF",X"BE",X"BE",X"BF",X"9F",X"1F",
		X"F6",X"F4",X"EC",X"E8",X"E8",X"E8",X"E8",X"68",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C1",X"20",X"10",X"10",X"08",X"03",X"07",X"07",X"51",X"F6",X"63",X"23",X"21",
		X"68",X"E8",X"F0",X"A0",X"00",X"00",X"80",X"E0",X"07",X"07",X"4F",X"4E",X"6C",X"6C",X"6C",X"6E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C3",X"61",X"21",
		X"70",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"05",X"05",X"05",X"10",X"10",X"10",X"10",X"09",X"08",X"89",X"CB",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"03",X"0D",X"8E",X"9F",X"1F",X"1F",X"1F",X"3F",
		X"E0",X"E0",X"F0",X"60",X"60",X"A0",X"A0",X"30",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"3F",X"3F",X"3F",X"3E",X"7E",X"7F",X"3F",X"1E",
		X"58",X"E8",X"E0",X"F0",X"FA",X"FA",X"FA",X"F6",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"88",X"88",X"C0",X"C0",X"E0",X"E1",X"0E",X"0F",X"BF",X"BE",X"BE",X"BF",X"9F",X"1F",
		X"F6",X"F4",X"EC",X"E8",X"E8",X"E8",X"E8",X"68",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"03",X"07",X"07",X"11",X"16",X"23",X"23",X"61",
		X"68",X"E8",X"F0",X"A0",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"3C",X"3C",X"3C",X"3E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"30",X"00",X"80",X"80",X"C0",X"C0",X"63",X"21",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"03",X"0D",X"8E",X"9F",X"1F",X"1F",X"1F",X"3F",
		X"E0",X"E0",X"F0",X"60",X"60",X"A0",X"A0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"3F",X"3F",X"3F",X"3E",X"7E",X"7F",X"3F",X"1E",
		X"58",X"E8",X"E0",X"F0",X"FA",X"FA",X"FA",X"F6",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"0E",X"0F",X"BF",X"BE",X"BE",X"BF",X"9F",X"1F",
		X"F6",X"F4",X"EC",X"E8",X"E8",X"E8",X"E8",X"68",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"03",X"07",X"07",X"11",X"16",X"23",X"23",X"21",
		X"68",X"E8",X"F0",X"A0",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"16",X"17",X"23",X"23",X"21",
		X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"16",X"17",X"23",X"23",X"21",
		X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"02",X"00",X"00",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"00",X"00",X"08",X"18",X"1C",X"1C",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"1C",X"1C",X"8C",X"88",X"80",X"80",X"80",X"00",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"16",X"17",X"23",X"23",X"21",
		X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"02",X"00",X"08",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"18",X"18",X"18",X"18",X"18",X"1A",X"18",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"18",X"08",X"8C",X"8C",X"8C",X"86",X"84",X"00",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"16",X"17",X"23",X"23",X"21",
		X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"09",X"08",X"09",X"4B",X"47",X"27",X"2F",X"0F",
		X"F0",X"70",X"A0",X"C0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"30",X"1C",X"08",X"08",X"00",X"20",X"1F",X"1F",X"9F",X"A7",X"03",X"1A",X"10",X"30",
		X"E0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"10",X"08",X"48",X"48",X"2A",X"2A",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"24",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"11",X"11",X"90",X"90",X"C0",X"C0",X"E0",X"E1",X"30",X"30",X"98",X"98",X"98",X"98",X"8C",X"0C",
		X"24",X"3C",X"00",X"00",X"00",X"00",X"40",X"20",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"07",
		X"F1",X"F1",X"E1",X"C0",X"20",X"10",X"10",X"08",X"0C",X"06",X"00",X"16",X"17",X"23",X"23",X"21",
		X"10",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"07",X"07",X"0F",X"0E",X"0C",X"0C",X"0C",X"0E",
		X"00",X"00",X"00",X"01",X"23",X"27",X"3F",X"3F",X"20",X"00",X"80",X"80",X"C0",X"C0",X"60",X"20",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F1",X"F8",X"F8",X"F0",X"F0",X"E0",X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"07",X"07",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F3",X"F7",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"FC",X"FC",X"F8",X"70",X"00",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"00",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"01",X"06",X"18",X"01",X"02",X"04",X"08",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"74",X"BA",X"59",X"54",X"94",X"92",X"12",X"11",X"11",X"10",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"E0",X"18",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"18",X"07",X"00",X"1F",
		X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"48",X"49",X"29",X"2A",X"9A",X"5D",X"2E",X"FD",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"10",X"20",X"40",X"80",X"18",X"60",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"06",X"18",X"01",X"02",X"04",X"08",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"74",X"BA",X"59",X"54",X"94",X"92",X"12",X"11",X"11",X"10",X"00",X"00",X"00",X"00",
		X"FC",X"00",X"E0",X"18",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"18",X"07",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"48",X"49",X"29",X"2A",X"9A",X"5D",X"2E",X"FD",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"10",X"20",X"40",X"80",X"18",X"60",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"24",X"24",X"22",X"42",X"42",X"41",X"41",X"41",X"41",X"41",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"20",X"20",X"20",X"20",X"10",X"11",X"11",X"09",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"40",X"C0",X"C0",X"40",X"80",X"00",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"60",X"60",X"E0",X"E0",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"70",X"70",X"F0",X"F0",X"30",X"D0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"01",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"78",X"F0",X"F0",X"F0",X"70",X"10",X"C0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"04",
		X"18",X"3C",X"7E",X"FD",X"7C",X"38",X"98",X"C0",X"50",X"68",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"01",X"00",X"20",X"20",X"10",X"10",X"00",X"10",
		X"0C",X"3C",X"FE",X"FE",X"7D",X"7C",X"38",X"B8",X"C0",X"40",X"70",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"1C",X"FC",X"FC",X"FE",X"FE",X"7A",X"70",X"60",X"80",X"80",X"80",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"23",X"21",X"11",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"F8",X"7C",X"70",X"60",X"40",X"80",X"40",X"40",X"00",X"00",
		X"00",X"20",X"10",X"08",X"04",X"04",X"04",X"06",X"02",X"12",X"11",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E8",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"02",X"10",X"00",X"00",X"02",X"06",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"20",X"20",X"40",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"04",X"04",X"04",X"00",X"00",X"05",X"04",X"08",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"20",X"20",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"03",X"02",X"00",X"01",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"90",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"00",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"80",X"80",X"80",X"80",
		X"05",X"05",X"05",X"05",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"09",X"08",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"80",X"80",X"80",
		X"02",X"02",X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"A0",X"30",X"10",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"03",X"17",X"1B",X"0B",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"30",X"90",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"04",X"0E",X"0F",X"07",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"10",X"00",X"80",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"10",X"13",X"07",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"58",X"88",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"09",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"70",X"90",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"08",X"01",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"40",X"60",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"04",X"01",X"05",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",
		X"02",X"02",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"80",X"80",X"80",
		X"02",X"02",X"02",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"00",X"00",
		X"02",X"02",X"00",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"20",X"60",X"80",X"00",
		X"04",X"0A",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"A0",X"60",X"80",
		X"0D",X"0A",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"80",
		X"01",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"00",X"02",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"80",X"00",X"00",
		X"01",X"00",X"04",X"02",X"00",X"04",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"04",X"02",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"00",X"80",X"40",X"80",
		X"01",X"02",X"04",X"03",X"00",X"04",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"40",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"05",X"02",X"05",X"02",X"01",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"80",X"40",X"80",X"40",X"80",
		X"05",X"06",X"05",X"03",X"02",X"04",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"40",X"80",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"00",
		X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"04",X"00",X"05",X"05",X"05",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"80",X"80",X"80",X"80",
		X"05",X"05",X"05",X"05",X"00",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FB",
		X"FF",X"FF",X"FF",X"E0",X"C0",X"01",X"00",X"FF",X"FF",X"FF",X"80",X"00",X"07",X"00",X"00",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FD",X"F9",X"EF",X"DC",X"BF",X"1F",X"3C",X"A7",X"FF",X"FF",
		X"00",X"00",X"FF",X"FB",X"7D",X"04",X"87",X"C0",X"00",X"00",X"FF",X"FF",X"83",X"F4",X"08",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"FF",X"FF",X"FC",X"E0",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"0C",X"0E",X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",
		X"F0",X"FF",X"EF",X"CF",X"DF",X"07",X"40",X"03",X"03",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"F0",X"0F",X"E5",X"FC",X"EF",X"FD",X"FF",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"02",X"00",X"7F",X"1F",X"3F",X"7F",X"FF",X"7F",X"00",X"0F",X"E7",X"F3",X"F9",X"FD",X"FC",X"FE",
		X"2D",X"FE",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"3F",X"3F",X"7F",X"3F",X"9F",X"CF",
		X"FF",X"FF",X"FC",X"FF",X"FF",X"F8",X"FE",X"FF",X"F3",X"FD",X"7F",X"FF",X"C0",X"FF",X"00",X"FC",
		X"C0",X"C0",X"E0",X"E0",X"E0",X"F0",X"F8",X"FC",X"01",X"05",X"0F",X"1F",X"7E",X"3D",X"0D",X"00",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"FE",X"FF",X"FF",X"FE",X"BF",X"FF",X"FF",X"FF",
		X"FE",X"7F",X"78",X"00",X"67",X"BF",X"BF",X"FF",X"7F",X"FC",X"E1",X"7F",X"BF",X"BF",X"FC",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"04",X"FF",X"FF",X"FF",X"FE",X"80",X"DD",X"F0",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"FB",X"DF",X"F9",X"FF",X"F7",X"FF",X"FB",X"3F",X"FF",X"E8",X"FF",X"FF",X"C7",X"FF",X"FF",
		X"FF",X"FC",X"00",X"FF",X"80",X"FF",X"EF",X"FD",X"C4",X"4C",X"FF",X"FF",X"7F",X"C7",X"80",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"00",X"FF",X"FF",X"FF",X"FF",X"C0",X"1C",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"F0",X"E0",
		X"FF",X"FF",X"F8",X"80",X"00",X"00",X"00",X"00",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"C0",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"F8",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"00",X"00",X"00",X"36",X"0F",X"5F",X"5F",X"FF",X"FF",X"3F",X"1F",X"03",X"F0",X"FC",X"FE",
		X"FE",X"FC",X"F8",X"E0",X"C0",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"07",X"03",X"03",X"03",X"01",X"00",X"00",X"00",
		X"5F",X"F0",X"C7",X"FF",X"E0",X"FF",X"9F",X"9F",X"EF",X"67",X"EF",X"E7",X"67",X"EF",X"FF",X"FE",
		X"1F",X"1F",X"9F",X"9F",X"BF",X"3F",X"3F",X"7E",X"C0",X"E0",X"E0",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"E0",X"F8",X"FF",X"FF",
		X"5F",X"3F",X"30",X"00",X"01",X"1F",X"FF",X"FF",X"F8",X"C7",X"07",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"08",X"E0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"3B",X"37",X"6F",X"6D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"E0",X"FE",X"FF",X"FF",X"FF",X"1B",X"1B",X"1A",X"06",X"00",X"80",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"78",
		X"F0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",X"C0",X"00",X"00",X"01",X"00",X"02",X"19",X"0C",X"07",
		X"03",X"00",X"FE",X"FF",X"F9",X"86",X"17",X"64",X"FF",X"7E",X"1E",X"80",X"C0",X"DA",X"6E",X"CC",
		X"00",X"00",X"00",X"00",X"20",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"80",X"C0",X"C0",X"E0",X"F0",X"FC",X"FF",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"81",
		X"09",X"FF",X"7C",X"61",X"03",X"3F",X"3F",X"FF",X"9C",X"38",X"00",X"C0",X"F0",X"F0",X"F8",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"14",X"00",X"00",X"00",X"00",X"67",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"F0",X"E0",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"0C",
		X"FF",X"FF",X"FF",X"03",X"01",X"00",X"12",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"C0",X"81",X"81",X"81",X"81",X"81",X"80",X"38",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"7F",X"E5",X"FF",X"FF",X"F7",X"FF",X"F3",X"FB",X"7D",X"FD",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"F9",X"F0",X"E0",X"F0",X"FB",X"FF",X"FF",X"FC",X"80",X"00",X"00",X"E0",X"FF",
		X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"01",X"01",X"00",X"00",X"00",X"FF",
		X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"FE",X"FF",X"7D",X"3D",X"1C",X"0E",X"02",X"00",X"00",X"C1",
		X"7F",X"7F",X"BF",X"FE",X"02",X"03",X"0F",X"FF",X"F7",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"A1",X"FF",X"FC",X"00",X"00",X"00",X"F8",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F9",X"FA",X"F0",X"E0",X"C1",
		X"18",X"00",X"B6",X"E0",X"00",X"07",X"7F",X"E0",X"40",X"00",X"00",X"00",X"01",X"F0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"27",X"2F",X"01",X"00",X"04",X"00",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"07",X"00",X"00",X"07",X"9F",X"CF",X"C0",X"80",X"B0",X"09",X"00",X"E1",X"FC",X"FE",
		X"1F",X"67",X"1F",X"00",X"78",X"BF",X"FE",X"38",X"00",X"18",X"F8",X"FC",X"37",X"1F",X"06",X"E0",
		X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",X"07",X"07",X"13",X"0D",X"0F",X"1F",X"0E",X"0E",
		X"3F",X"B8",X"F7",X"FF",X"FA",X"7F",X"4F",X"4F",X"F7",X"77",X"FF",X"EF",X"FF",X"F7",X"FF",X"FF",
		X"C7",X"E7",X"F7",X"F7",X"F7",X"F7",X"EF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FC",
		X"1D",X"C9",X"E7",X"F7",X"9E",X"3C",X"1F",X"3F",X"18",X"81",X"FF",X"F9",X"0F",X"0F",X"C3",X"F0",
		X"F8",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"06",X"01",X"00",X"00",X"00",X"80",X"F8",X"FF",
		X"6F",X"0F",X"07",X"00",X"00",X"00",X"00",X"C1",X"FF",X"FE",X"F8",X"00",X"00",X"03",X"0F",X"FF",
		X"1F",X"3F",X"00",X"04",X"3F",X"FF",X"FF",X"FF",X"F4",X"E0",X"11",X"00",X"00",X"80",X"81",X"C0",
		X"FF",X"F2",X"01",X"00",X"7F",X"07",X"83",X"68",X"DC",X"02",X"FE",X"04",X"F0",X"9E",X"FF",X"7E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"EF",X"E6",X"F0",X"FB",X"F9",X"FD",X"FC",
		X"00",X"80",X"FF",X"78",X"C0",X"03",X"0F",X"FF",X"00",X"00",X"E0",X"70",X"00",X"80",X"E0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1C",X"01",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",X"80",X"E0",X"01",X"FC",X"78",X"87",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E4",X"9F",
		X"FF",X"FF",X"FE",X"F0",X"03",X"00",X"80",X"87",X"FF",X"F8",X"00",X"2C",X"98",X"00",X"00",X"D2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"03",X"7C",X"0C",X"25",X"71",X"8C",X"7E",X"00",
		X"B8",X"78",X"13",X"80",X"C6",X"70",X"01",X"00",X"07",X"80",X"18",X"42",X"00",X"C0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"E0",X"FF",X"FF",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"08",X"07",X"00",X"08",X"07",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"03",X"F8",
		X"F8",X"FA",X"F3",X"F0",X"F1",X"E4",X"E0",X"00",X"00",X"00",X"00",X"06",X"FF",X"08",X"03",X"5B",
		X"00",X"0E",X"7F",X"00",X"FF",X"3F",X"8C",X"8C",X"18",X"BF",X"C0",X"3F",X"BF",X"D8",X"47",X"37",
		X"E0",X"C0",X"80",X"80",X"80",X"C0",X"E0",X"F0",X"00",X"01",X"01",X"03",X"0F",X"0F",X"1F",X"3D",
		X"2F",X"2F",X"BF",X"F8",X"F7",X"FF",X"B0",X"3F",X"FC",X"EE",X"47",X"23",X"FF",X"FF",X"6F",X"E7",
		X"20",X"3C",X"9E",X"CF",X"DF",X"DF",X"DF",X"8F",X"0D",X"7E",X"00",X"80",X"80",X"FF",X"8F",X"7F",
		X"73",X"DF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"E6",X"E8",X"01",X"00",X"80",X"FD",X"FF",X"FF",
		X"F0",X"E0",X"E0",X"C0",X"C0",X"E0",X"FC",X"FF",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"4F",X"4F",X"0F",X"08",X"04",X"07",X"7F",X"FF",X"FF",X"F8",X"D0",X"0F",X"7F",X"FF",X"FF",X"FF",
		X"3E",X"78",X"00",X"C0",X"F0",X"F0",X"F0",X"F8",X"0E",X"0B",X"03",X"ED",X"6F",X"37",X"00",X"00",
		X"61",X"8E",X"8E",X"33",X"FF",X"DF",X"00",X"00",X"96",X"38",X"BA",X"D7",X"FD",X"F0",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"F8",X"FD",X"FC",X"FC",X"FE",X"FE",X"FF",X"3F",X"10",X"F7",X"7F",X"44",X"11",X"3D",X"4F",
		X"FC",X"1F",X"00",X"FF",X"F4",X"C7",X"D7",X"BF",X"FF",X"E0",X"3F",X"FF",X"C3",X"1C",X"D8",X"E3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"08",X"80",X"CE",X"F9",X"FC",X"FF",X"FF",
		X"6F",X"00",X"00",X"7F",X"80",X"60",X"80",X"FF",X"F4",X"02",X"E0",X"02",X"38",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FC",X"F8",X"F3",X"EC",X"DF",X"C7",X"FE",X"80",X"00",X"E0",X"00",X"80",X"F0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F8",X"FF",X"FF",X"F8",X"C0",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"03",X"FF",X"FF",X"FF",X"FE",X"3E",X"0D",X"00",X"80",
		X"BF",X"FF",X"79",X"FF",X"FF",X"FF",X"7F",X"1F",X"EF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"80",X"F8",X"FC",X"F9",X"7D",X"FC",X"EB",
		X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"09",X"05",X"01",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"61",X"0D",X"1F",X"05",X"E3",X"FF",X"C3",X"B9",X"8C",X"E1",X"E1",X"DD",X"FC",X"F3",
		X"CF",X"E7",X"EF",X"F7",X"73",X"FF",X"FF",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"FF",X"03",X"F8",X"FF",X"FF",X"F9",X"80",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"3B",X"07",X"04",X"00",X"01",X"07",X"1F",X"FF",X"C3",X"98",X"3E",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"E0",X"FC",X"FC",X"FD",X"FD",X"FD",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DF",X"EF",X"F7",X"FB",X"F8",X"FF",X"FF",X"FF",X"FC",X"FE",X"EC",X"F7",X"FF",X"6F",X"80",X"FC",
		X"0F",X"00",X"80",X"80",X"00",X"04",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"01",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E0",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"83",X"0F",X"FF",X"C0",X"81",X"07",X"0F",X"CF",X"C6",X"C3",X"AF",
		X"07",X"FF",X"FF",X"F8",X"8F",X"7F",X"FF",X"FF",X"C0",X"E1",X"83",X"5F",X"FF",X"FF",X"7C",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FF",X"FF",X"C7",X"BF",X"FF",X"AF",X"6F",X"57",X"50",X"01",
		X"FF",X"FE",X"F9",X"F7",X"EF",X"1F",X"FF",X"8F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FC",
		X"FF",X"F3",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"70",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FF",X"F8",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"F9",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"81",X"03",X"02",X"C0",X"C0",X"00",X"00",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"10",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",
		X"7F",X"FF",X"FF",X"FD",X"C6",X"C7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"43",X"D3",X"FB",
		X"F8",X"F8",X"F0",X"E0",X"E0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"06",X"06",X"05",X"04",X"02",X"00",X"FF",X"FF",X"FF",X"7F",X"F7",X"F7",X"7F",X"7F",
		X"E0",X"F2",X"F8",X"FC",X"FC",X"78",X"78",X"31",X"1F",X"9F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",
		X"F7",X"FF",X"FC",X"F2",X"F8",X"FF",X"FF",X"FF",X"FC",X"B0",X"3C",X"FF",X"BB",X"08",X"00",X"FF",
		X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"01",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"FD",X"DC",X"1C",X"03",X"38",X"10",X"0D",X"3B",
		X"23",X"07",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"E3",X"DF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
