library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity robotron_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of robotron_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7E",X"D1",X"06",X"7E",X"DE",X"0F",X"7E",X"D3",X"B6",X"7E",X"DC",X"11",X"7E",X"DB",X"9C",X"7E",
		X"DC",X"13",X"7E",X"DB",X"7C",X"7E",X"DB",X"03",X"7E",X"DA",X"F2",X"7E",X"DA",X"DF",X"7E",X"DA",
		X"BF",X"7E",X"DA",X"82",X"7E",X"D8",X"9E",X"7E",X"D7",X"C9",X"7E",X"D5",X"F5",X"7E",X"D5",X"E2",
		X"7E",X"D7",X"A5",X"7E",X"D7",X"95",X"7E",X"D6",X"EC",X"7E",X"D6",X"CD",X"7E",X"D6",X"C8",X"7E",
		X"D6",X"B6",X"7E",X"D6",X"AC",X"7E",X"D6",X"99",X"7E",X"D6",X"A8",X"7E",X"D3",X"C7",X"7E",X"D2",
		X"A7",X"7E",X"D2",X"8F",X"7E",X"D2",X"81",X"7E",X"D2",X"5A",X"7E",X"D2",X"43",X"7E",X"D2",X"18",
		X"7E",X"D1",X"FF",X"7E",X"D1",X"F3",X"7E",X"D1",X"E3",X"7E",X"D3",X"0E",X"7E",X"D3",X"2B",X"7E",
		X"D2",X"FD",X"7E",X"D3",X"06",X"7E",X"D3",X"1B",X"7E",X"D3",X"20",X"7E",X"D2",X"DA",X"7E",X"D2",
		X"C2",X"7E",X"D2",X"E7",X"7E",X"D2",X"CA",X"7E",X"D2",X"F2",X"7E",X"D2",X"D2",X"7E",X"DB",X"2F",
		X"7E",X"DA",X"9E",X"7E",X"DA",X"61",X"7E",X"D1",X"96",X"7E",X"D4",X"FC",X"7E",X"D5",X"03",X"7E",
		X"D5",X"C0",X"7E",X"D5",X"12",X"7E",X"D5",X"23",X"7E",X"D5",X"21",X"7E",X"D5",X"2B",X"7E",X"D5",
		X"39",X"7E",X"D5",X"37",X"7E",X"D5",X"E2",X"7E",X"DE",X"59",X"7E",X"D6",X"5B",X"7E",X"D6",X"55",
		X"7E",X"D1",X"8A",X"7E",X"DA",X"0D",X"7E",X"D5",X"D8",X"EF",X"01",X"20",X"1E",X"00",X"FF",X"01",
		X"20",X"0C",X"00",X"FF",X"01",X"20",X"20",X"00",X"FF",X"03",X"10",X"24",X"00",X"FF",X"01",X"20",
		X"27",X"00",X"FF",X"01",X"20",X"2D",X"00",X"FF",X"02",X"10",X"35",X"00",X"FF",X"01",X"20",X"3A",
		X"00",X"FF",X"01",X"20",X"3E",X"00",X"00",X"34",X"FF",X"35",X"00",X"34",X"00",X"3C",X"C8",X"0C",
		X"C8",X"0E",X"C8",X"04",X"C8",X"06",X"1A",X"FF",X"10",X"CE",X"BF",X"70",X"86",X"98",X"1F",X"8B",
		X"86",X"01",X"B7",X"C9",X"00",X"8E",X"D0",X"F6",X"4F",X"5F",X"ED",X"98",X"08",X"EC",X"81",X"ED",
		X"98",X"06",X"8C",X"D0",X"FE",X"26",X"F1",X"86",X"FF",X"B7",X"C8",X"0E",X"BD",X"D0",X"12",X"86",
		X"3F",X"B7",X"C8",X"0E",X"8E",X"98",X"00",X"6F",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",
		X"70",X"26",X"F4",X"CC",X"A5",X"5A",X"DD",X"85",X"86",X"60",X"97",X"41",X"BD",X"D0",X"99",X"BD",
		X"D0",X"36",X"8D",X"36",X"BD",X"6F",X"03",X"CC",X"FF",X"FF",X"DD",X"2F",X"DD",X"31",X"86",X"02",
		X"97",X"40",X"8E",X"CD",X"00",X"BD",X"D0",X"A2",X"1F",X"89",X"81",X"20",X"22",X"06",X"C4",X"0F",
		X"C1",X"09",X"25",X"04",X"4F",X"BD",X"D0",X"AB",X"97",X"51",X"BD",X"D0",X"54",X"77",X"A0",X"86",
		X"2C",X"B7",X"C8",X"0E",X"03",X"59",X"1C",X"00",X"20",X"0C",X"BD",X"D0",X"33",X"BD",X"5F",X"9C",
		X"BD",X"5B",X"40",X"7E",X"D0",X"30",X"8E",X"98",X"11",X"9F",X"15",X"96",X"10",X"81",X"02",X"25",
		X"FA",X"48",X"48",X"48",X"9B",X"42",X"44",X"97",X"42",X"0F",X"10",X"BD",X"D6",X"CD",X"96",X"59",
		X"85",X"04",X"26",X"03",X"BD",X"5B",X"49",X"9E",X"33",X"26",X"0C",X"9E",X"37",X"27",X"17",X"DC",
		X"39",X"0F",X"37",X"0F",X"38",X"20",X"06",X"DC",X"35",X"0F",X"33",X"0F",X"34",X"D4",X"59",X"26",
		X"E6",X"BD",X"D0",X"57",X"20",X"E1",X"DE",X"11",X"27",X"13",X"6A",X"44",X"26",X"0B",X"DF",X"15",
		X"6E",X"D8",X"02",X"DE",X"15",X"A7",X"44",X"AF",X"42",X"EE",X"C4",X"26",X"ED",X"10",X"CE",X"BF",
		X"70",X"20",X"A3",X"9E",X"15",X"10",X"CE",X"BF",X"70",X"8D",X"1D",X"33",X"84",X"20",X"EA",X"34",
		X"12",X"8E",X"98",X"11",X"AE",X"84",X"27",X"0E",X"9C",X"15",X"27",X"F8",X"A6",X"05",X"81",X"01",
		X"27",X"F2",X"8D",X"04",X"20",X"EE",X"35",X"92",X"34",X"46",X"CE",X"98",X"11",X"AC",X"C4",X"26",
		X"18",X"EC",X"84",X"ED",X"C4",X"A6",X"06",X"27",X"06",X"DC",X"1D",X"9F",X"1D",X"20",X"04",X"DC",
		X"13",X"9F",X"13",X"ED",X"84",X"30",X"C4",X"35",X"C6",X"EE",X"C4",X"26",X"E0",X"8D",X"00",X"1A",
		X"10",X"20",X"FE",X"34",X"62",X"DE",X"1D",X"26",X"01",X"BD",X"D2",X"3F",X"10",X"AE",X"C4",X"10",
		X"9F",X"1D",X"86",X"01",X"A7",X"46",X"A6",X"E4",X"20",X"11",X"34",X"62",X"DE",X"13",X"26",X"03",
		X"BD",X"D2",X"3F",X"10",X"AE",X"C4",X"10",X"9F",X"13",X"6F",X"46",X"AF",X"42",X"A7",X"45",X"86",
		X"01",X"A7",X"44",X"AE",X"9F",X"98",X"15",X"EF",X"9F",X"98",X"15",X"AF",X"C4",X"30",X"C4",X"35",
		X"E2",X"34",X"42",X"EE",X"63",X"37",X"10",X"EF",X"63",X"86",X"00",X"8D",X"CD",X"35",X"C2",X"34",
		X"06",X"9E",X"1B",X"26",X"03",X"BD",X"D2",X"3F",X"EC",X"84",X"DD",X"1B",X"C6",X"02",X"6F",X"85",
		X"5C",X"C1",X"18",X"26",X"F9",X"35",X"86",X"AC",X"C4",X"26",X"10",X"10",X"AE",X"D4",X"10",X"AF",
		X"C4",X"10",X"9E",X"1B",X"9F",X"1B",X"10",X"AF",X"84",X"35",X"F0",X"EE",X"C4",X"26",X"E8",X"BD",
		X"D2",X"3F",X"34",X"70",X"CE",X"98",X"21",X"7E",X"D0",X"4E",X"34",X"70",X"CE",X"98",X"23",X"7E",
		X"D0",X"4E",X"34",X"70",X"CE",X"98",X"1F",X"7E",X"D0",X"4E",X"34",X"06",X"BD",X"D0",X"51",X"DC",
		X"21",X"9F",X"21",X"ED",X"84",X"35",X"86",X"34",X"06",X"BD",X"D0",X"51",X"DC",X"23",X"9F",X"23",
		X"20",X"F1",X"34",X"06",X"BD",X"D0",X"51",X"DC",X"1F",X"9F",X"1F",X"20",X"E6",X"34",X"06",X"BD",
		X"D0",X"51",X"DC",X"17",X"20",X"DD",X"34",X"70",X"CE",X"98",X"17",X"7E",X"D0",X"4E",X"10",X"8E",
		X"AE",X"D9",X"BD",X"D0",X"54",X"D3",X"68",X"10",X"AF",X"09",X"39",X"8D",X"E9",X"7E",X"D0",X"15",
		X"34",X"10",X"8D",X"F7",X"AE",X"06",X"BD",X"D0",X"5D",X"35",X"90",X"34",X"26",X"9E",X"1B",X"27",
		X"2E",X"9E",X"13",X"27",X"2A",X"4F",X"EE",X"64",X"37",X"10",X"BD",X"D0",X"57",X"31",X"84",X"BD",
		X"D0",X"6F",X"EC",X"C1",X"ED",X"88",X"14",X"ED",X"02",X"37",X"06",X"ED",X"08",X"EF",X"64",X"33",
		X"A4",X"EF",X"06",X"AF",X"47",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"0E",X"43",X"35",X"A6",X"EE",
		X"64",X"33",X"48",X"EF",X"64",X"4F",X"35",X"A6",X"96",X"F2",X"26",X"47",X"0C",X"F2",X"86",X"03",
		X"AE",X"49",X"30",X"89",X"28",X"57",X"AF",X"49",X"A7",X"47",X"86",X"08",X"8E",X"D3",X"82",X"7E",
		X"D0",X"66",X"B6",X"C8",X"04",X"81",X"A1",X"27",X"0A",X"81",X"58",X"27",X"ED",X"6A",X"47",X"26",
		X"E9",X"20",X"1E",X"86",X"03",X"A7",X"47",X"86",X"08",X"8E",X"D3",X"9F",X"7E",X"D0",X"66",X"B6",
		X"C8",X"04",X"81",X"42",X"26",X"03",X"6E",X"D8",X"09",X"81",X"A1",X"27",X"EA",X"6A",X"47",X"26",
		X"E6",X"0F",X"F2",X"7E",X"D0",X"63",X"34",X"07",X"1A",X"FF",X"86",X"3F",X"B7",X"C8",X"0E",X"53",
		X"C4",X"3F",X"F7",X"C8",X"0E",X"35",X"87",X"34",X"17",X"1F",X"01",X"A6",X"84",X"91",X"56",X"25",
		X"0D",X"97",X"56",X"30",X"1E",X"1A",X"10",X"9F",X"54",X"CC",X"01",X"01",X"DD",X"57",X"35",X"97",
		X"96",X"57",X"27",X"1E",X"0A",X"57",X"26",X"1A",X"9E",X"54",X"0A",X"58",X"26",X"0E",X"30",X"03",
		X"9F",X"54",X"A6",X"84",X"26",X"04",X"97",X"56",X"20",X"08",X"97",X"58",X"EC",X"01",X"97",X"57",
		X"8D",X"B4",X"B6",X"C8",X"0C",X"85",X"40",X"27",X"04",X"86",X"3C",X"97",X"4B",X"96",X"4B",X"27",
		X"02",X"0A",X"4B",X"96",X"4C",X"27",X"02",X"0A",X"4C",X"96",X"4E",X"27",X"02",X"0A",X"4E",X"96",
		X"4D",X"27",X"02",X"0A",X"4D",X"96",X"59",X"2A",X"24",X"96",X"CE",X"26",X"6A",X"96",X"31",X"9A",
		X"32",X"43",X"D6",X"31",X"D7",X"32",X"F6",X"C8",X"04",X"D7",X"31",X"94",X"31",X"84",X"30",X"27",
		X"0C",X"8E",X"26",X"CC",X"85",X"10",X"26",X"03",X"8E",X"26",X"CF",X"8D",X"3B",X"96",X"CE",X"26",
		X"46",X"96",X"2F",X"9A",X"30",X"43",X"D6",X"2F",X"D7",X"30",X"F6",X"C8",X"0C",X"C4",X"3F",X"D7",
		X"2F",X"95",X"2F",X"27",X"32",X"8E",X"00",X"78",X"30",X"1F",X"26",X"FC",X"F6",X"C8",X"0C",X"D4",
		X"2F",X"D7",X"2F",X"94",X"2F",X"27",X"20",X"8E",X"D4",X"96",X"30",X"02",X"44",X"24",X"FB",X"AE",
		X"84",X"8D",X"05",X"86",X"01",X"A7",X"42",X"39",X"CE",X"98",X"33",X"EC",X"C4",X"27",X"02",X"33",
		X"44",X"AF",X"C4",X"6F",X"42",X"6F",X"43",X"39",X"00",X"00",X"F0",X"03",X"D6",X"15",X"E3",X"DF",
		X"D6",X"0C",X"D6",X"1E",X"00",X"00",X"00",X"00",X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",
		X"4E",X"3A",X"20",X"32",X"30",X"38",X"34",X"20",X"28",X"54",X"4D",X"29",X"20",X"20",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",
		X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"34",X"06",X"CC",X"01",
		X"3C",X"20",X"05",X"34",X"06",X"CC",X"03",X"34",X"97",X"45",X"B7",X"C9",X"00",X"F7",X"C8",X"07",
		X"35",X"86",X"A6",X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",
		X"39",X"8D",X"EF",X"34",X"02",X"8D",X"EB",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",
		X"44",X"44",X"44",X"A7",X"81",X"35",X"82",X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",
		X"82",X"34",X"12",X"9B",X"51",X"19",X"24",X"02",X"86",X"99",X"97",X"51",X"8E",X"CD",X"00",X"BD",
		X"D0",X"AB",X"35",X"92",X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",
		X"34",X"16",X"C6",X"01",X"BD",X"D0",X"BD",X"58",X"8E",X"CC",X"04",X"3A",X"BD",X"D0",X"A5",X"BD",
		X"D0",X"B4",X"96",X"4F",X"34",X"04",X"AB",X"E4",X"97",X"4F",X"96",X"50",X"AB",X"E0",X"97",X"50",
		X"8E",X"CC",X"10",X"BD",X"D0",X"A5",X"BD",X"D0",X"B4",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",
		X"96",X"8E",X"CC",X"0C",X"BD",X"D0",X"A5",X"BD",X"D0",X"B4",X"8D",X"24",X"34",X"02",X"D7",X"50",
		X"8E",X"CC",X"0E",X"BD",X"D0",X"A5",X"96",X"4F",X"8D",X"38",X"8D",X"14",X"4D",X"27",X"04",X"0F",
		X"50",X"0F",X"4F",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"D0",X"BA",X"BD",X"D5",X"41",X"35",X"96",
		X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",X"01",X"19",X"E0",
		X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"D8",X"3E",X"34",X"04",X"1F",X"89",X"8D",X"04",X"1F",X"98",
		X"35",X"84",X"34",X"02",X"4F",X"C1",X"10",X"25",X"06",X"8B",X"0A",X"C0",X"10",X"20",X"F6",X"34",
		X"02",X"EB",X"E0",X"35",X"82",X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",
		X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"8E",X"98",X"4C",X"10",
		X"8E",X"D5",X"60",X"20",X"10",X"8E",X"98",X"4D",X"10",X"8E",X"D5",X"54",X"20",X"07",X"8E",X"98",
		X"4E",X"10",X"8E",X"D5",X"5A",X"96",X"4B",X"26",X"27",X"A6",X"84",X"26",X"23",X"86",X"16",X"A7",
		X"84",X"10",X"AF",X"49",X"86",X"0A",X"8E",X"D6",X"3C",X"7E",X"D0",X"66",X"96",X"4B",X"26",X"10",
		X"86",X"05",X"D6",X"84",X"C4",X"07",X"3D",X"C3",X"D0",X"CE",X"BD",X"D0",X"4B",X"AD",X"D8",X"09",
		X"7E",X"D0",X"63",X"5E",X"31",X"34",X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"0F",X"58",
		X"34",X"04",X"58",X"EB",X"E0",X"8E",X"CC",X"FC",X"3A",X"BD",X"D0",X"A5",X"34",X"04",X"BD",X"D0",
		X"A5",X"34",X"04",X"BD",X"D0",X"A5",X"34",X"04",X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",X"89",
		X"00",X"19",X"A7",X"61",X"A6",X"62",X"89",X"00",X"19",X"30",X"1A",X"BD",X"D0",X"AB",X"35",X"04",
		X"35",X"02",X"BD",X"D0",X"B1",X"35",X"02",X"35",X"96",X"34",X"02",X"96",X"3F",X"8E",X"BD",X"E4",
		X"4A",X"27",X"03",X"8E",X"BE",X"20",X"35",X"82",X"34",X"02",X"20",X"F1",X"34",X"04",X"1F",X"89",
		X"8D",X"1B",X"3D",X"4C",X"35",X"84",X"34",X"02",X"8D",X"13",X"A1",X"E4",X"23",X"03",X"44",X"20",
		X"F9",X"4D",X"26",X"01",X"4C",X"32",X"61",X"39",X"8D",X"03",X"D6",X"86",X"39",X"34",X"04",X"D6",
		X"84",X"86",X"03",X"3D",X"CB",X"11",X"96",X"86",X"44",X"44",X"44",X"98",X"86",X"44",X"06",X"85",
		X"06",X"86",X"DB",X"86",X"D9",X"85",X"D7",X"84",X"96",X"84",X"35",X"84",X"34",X"56",X"4F",X"5F",
		X"8E",X"A9",X"E0",X"CE",X"97",X"6F",X"9F",X"13",X"30",X"0F",X"AF",X"11",X"8C",X"B0",X"D9",X"26",
		X"F7",X"ED",X"84",X"DD",X"11",X"8E",X"B0",X"E8",X"9F",X"1D",X"30",X"88",X"1F",X"AF",X"88",X"E1",
		X"8C",X"B3",X"35",X"26",X"F5",X"ED",X"84",X"8E",X"98",X"11",X"9F",X"15",X"C6",X"07",X"1F",X"01",
		X"AB",X"84",X"30",X"88",X"10",X"8C",X"89",X"35",X"25",X"F6",X"A7",X"C9",X"01",X"84",X"35",X"D6",
		X"BD",X"D0",X"60",X"86",X"FF",X"97",X"59",X"86",X"01",X"8E",X"D7",X"3F",X"7E",X"D0",X"66",X"BD",
		X"D0",X"12",X"BD",X"5F",X"9C",X"C6",X"7F",X"D7",X"01",X"10",X"BE",X"D5",X"D6",X"31",X"A5",X"A6",
		X"A0",X"27",X"2C",X"81",X"02",X"26",X"09",X"B6",X"C8",X"04",X"85",X"40",X"27",X"30",X"20",X"EF",
		X"81",X"01",X"26",X"06",X"AE",X"A1",X"0F",X"D0",X"20",X"E5",X"8B",X"2E",X"CE",X"D7",X"4F",X"34",
		X"40",X"FE",X"D6",X"53",X"F6",X"D7",X"ED",X"33",X"C5",X"33",X"C5",X"33",X"C5",X"6E",X"C4",X"86",
		X"01",X"8E",X"D7",X"87",X"7E",X"D0",X"66",X"B6",X"C8",X"04",X"85",X"40",X"26",X"F1",X"BD",X"D0",
		X"12",X"6E",X"9F",X"EF",X"FE",X"8E",X"DA",X"51",X"CE",X"98",X"00",X"C6",X"10",X"A6",X"80",X"A7",
		X"C0",X"5A",X"26",X"F9",X"39",X"34",X"17",X"1A",X"FF",X"8E",X"99",X"00",X"9F",X"1B",X"30",X"88",
		X"18",X"AF",X"88",X"E8",X"8C",X"A9",X"C8",X"26",X"F5",X"4F",X"5F",X"ED",X"84",X"DD",X"21",X"DD",
		X"17",X"DD",X"19",X"DD",X"23",X"DD",X"1F",X"35",X"97",X"DD",X"7C",X"E3",X"C4",X"DD",X"7E",X"20",
		X"17",X"EC",X"04",X"27",X"13",X"91",X"7E",X"24",X"0F",X"D1",X"7F",X"24",X"0B",X"E3",X"98",X"02",
		X"91",X"7C",X"23",X"04",X"D1",X"7D",X"22",X"06",X"AE",X"84",X"26",X"E5",X"39",X"76",X"DF",X"82",
		X"0D",X"48",X"26",X"06",X"10",X"AE",X"88",X"16",X"26",X"03",X"10",X"AE",X"02",X"A3",X"A4",X"10",
		X"9F",X"2D",X"DD",X"2B",X"4F",X"5F",X"DD",X"76",X"DD",X"78",X"DC",X"2B",X"D0",X"7D",X"22",X"05",
		X"50",X"D7",X"77",X"20",X"02",X"D7",X"79",X"90",X"7C",X"22",X"05",X"40",X"97",X"76",X"20",X"02",
		X"97",X"78",X"DC",X"2B",X"E3",X"A4",X"D0",X"7F",X"22",X"01",X"5F",X"90",X"7E",X"22",X"01",X"4F",
		X"DD",X"80",X"EC",X"A4",X"93",X"76",X"93",X"80",X"DD",X"74",X"A6",X"C4",X"97",X"7B",X"D6",X"79",
		X"3D",X"EE",X"42",X"33",X"CB",X"A6",X"A4",X"97",X"7A",X"D6",X"77",X"3D",X"10",X"AE",X"22",X"31",
		X"AB",X"96",X"76",X"31",X"A6",X"96",X"78",X"33",X"C6",X"D6",X"74",X"5A",X"A6",X"C5",X"27",X"2C",
		X"A6",X"A5",X"27",X"28",X"31",X"A5",X"1F",X"20",X"DE",X"2D",X"A3",X"42",X"10",X"AE",X"04",X"E0",
		X"C4",X"82",X"00",X"25",X"08",X"31",X"21",X"E0",X"C4",X"82",X"00",X"24",X"F8",X"EB",X"C4",X"1F",
		X"98",X"5F",X"33",X"AB",X"DF",X"A6",X"AD",X"98",X"08",X"86",X"01",X"39",X"5A",X"2A",X"CD",X"DC",
		X"7A",X"31",X"A6",X"33",X"C5",X"0A",X"75",X"26",X"C0",X"DE",X"82",X"7E",X"D7",X"E8",X"BD",X"D0",
		X"54",X"D9",X"DF",X"BD",X"D0",X"54",X"D9",X"D2",X"BD",X"D0",X"54",X"DA",X"0D",X"BD",X"D0",X"54",
		X"D9",X"81",X"BD",X"D0",X"54",X"D9",X"AE",X"BD",X"D0",X"54",X"D9",X"8E",X"39",X"01",X"0C",X"28",
		X"26",X"1A",X"1B",X"25",X"0C",X"1B",X"25",X"0C",X"24",X"21",X"14",X"21",X"26",X"24",X"21",X"20",
		X"11",X"0C",X"04",X"21",X"0A",X"06",X"02",X"01",X"0C",X"58",X"16",X"17",X"25",X"1B",X"19",X"20",
		X"17",X"16",X"0C",X"17",X"2A",X"15",X"1E",X"27",X"25",X"1B",X"28",X"17",X"1E",X"2B",X"0C",X"18",
		X"21",X"24",X"01",X"0C",X"68",X"29",X"1B",X"1E",X"1E",X"1B",X"13",X"1F",X"25",X"0C",X"17",X"1E",
		X"17",X"15",X"26",X"24",X"21",X"20",X"1B",X"15",X"25",X"0C",X"1B",X"20",X"15",X"0F",X"02",X"01",
		X"0C",X"78",X"14",X"2B",X"0C",X"17",X"27",X"19",X"17",X"20",X"17",X"0C",X"22",X"0F",X"0C",X"1C",
		X"13",X"24",X"28",X"1B",X"25",X"0C",X"13",X"20",X"16",X"0C",X"1E",X"13",X"29",X"24",X"17",X"20",
		X"15",X"17",X"0C",X"17",X"0F",X"0C",X"16",X"17",X"1F",X"13",X"24",X"02",X"01",X"0C",X"A8",X"15",
		X"21",X"22",X"2B",X"24",X"1B",X"19",X"1A",X"26",X"0C",X"03",X"0B",X"0A",X"04",X"0C",X"29",X"1B",
		X"1E",X"1E",X"1B",X"13",X"1F",X"25",X"0C",X"17",X"1E",X"17",X"15",X"26",X"24",X"21",X"20",X"1B",
		X"15",X"25",X"0C",X"1B",X"20",X"15",X"0F",X"01",X"0C",X"B8",X"13",X"1E",X"1E",X"0C",X"24",X"1B",
		X"19",X"1A",X"26",X"25",X"0C",X"24",X"17",X"25",X"17",X"24",X"28",X"17",X"16",X"00",X"17",X"22",
		X"30",X"BD",X"D9",X"E8",X"D9",X"8A",X"98",X"0B",X"00",X"08",X"38",X"07",X"C0",X"00",X"BD",X"D9",
		X"E8",X"D9",X"97",X"98",X"0C",X"00",X"02",X"C0",X"C0",X"D0",X"E0",X"F0",X"F8",X"FA",X"BA",X"7A",
		X"3A",X"34",X"2D",X"1F",X"17",X"0F",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"BD",X"D9",
		X"E8",X"D9",X"B7",X"98",X"0E",X"00",X"01",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"87",
		X"87",X"47",X"47",X"07",X"07",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",
		X"C1",X"00",X"BD",X"D9",X"E8",X"D9",X"DB",X"98",X"0F",X"00",X"06",X"07",X"07",X"2F",X"00",X"BD",
		X"D9",X"E8",X"DA",X"2C",X"98",X"0D",X"00",X"02",X"AE",X"E1",X"EC",X"81",X"ED",X"47",X"EC",X"81",
		X"ED",X"4B",X"EC",X"81",X"ED",X"49",X"6F",X"49",X"AE",X"47",X"E6",X"49",X"6C",X"49",X"A6",X"85",
		X"27",X"F4",X"A7",X"D8",X"0B",X"A6",X"4A",X"8E",X"D9",X"F8",X"7E",X"D0",X"66",X"86",X"FF",X"97",
		X"0A",X"86",X"02",X"8E",X"DA",X"19",X"7E",X"D0",X"66",X"96",X"84",X"84",X"1F",X"8E",X"DA",X"2C",
		X"A6",X"86",X"97",X"0A",X"86",X"06",X"8E",X"DA",X"0D",X"7E",X"D0",X"66",X"38",X"39",X"3A",X"3B",
		X"3C",X"3D",X"3E",X"3F",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",
		X"C5",X"CC",X"CB",X"CA",X"DA",X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"3C",
		X"00",X"00",X"07",X"17",X"C7",X"1F",X"3F",X"38",X"C0",X"A4",X"FF",X"38",X"17",X"CC",X"81",X"81",
		X"07",X"34",X"07",X"1A",X"10",X"FD",X"CA",X"04",X"EC",X"A4",X"88",X"04",X"C8",X"04",X"FD",X"CA",
		X"06",X"EC",X"22",X"FD",X"CA",X"02",X"D6",X"2D",X"F7",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",
		X"35",X"87",X"34",X"07",X"1A",X"10",X"FD",X"CA",X"04",X"EC",X"A4",X"88",X"04",X"C8",X"04",X"FD",
		X"CA",X"06",X"EC",X"22",X"FD",X"CA",X"02",X"86",X"02",X"B7",X"CA",X"00",X"35",X"87",X"34",X"07",
		X"1A",X"10",X"FD",X"CA",X"04",X"EC",X"A4",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"22",
		X"FD",X"CA",X"02",X"D6",X"2D",X"F7",X"CA",X"01",X"86",X"1A",X"B7",X"CA",X"00",X"35",X"87",X"34",
		X"07",X"1A",X"10",X"FD",X"CA",X"04",X"EC",X"A4",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",
		X"22",X"FD",X"CA",X"02",X"CC",X"12",X"00",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"87",X"34",
		X"07",X"1A",X"10",X"BF",X"CA",X"04",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"CC",X"00",X"00",
		X"20",X"DF",X"34",X"47",X"EE",X"02",X"EC",X"C4",X"88",X"04",X"C8",X"04",X"1A",X"10",X"FD",X"CA",
		X"06",X"20",X"58",X"34",X"47",X"EE",X"88",X"14",X"EC",X"C4",X"EE",X"42",X"88",X"04",X"C8",X"04",
		X"1A",X"10",X"FD",X"CA",X"06",X"EC",X"04",X"FD",X"CA",X"04",X"FF",X"CA",X"02",X"CC",X"1A",X"00",
		X"F7",X"CA",X"01",X"E6",X"88",X"12",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"35",X"C7",X"34",
		X"47",X"EE",X"88",X"14",X"EC",X"C4",X"EE",X"42",X"88",X"04",X"C8",X"04",X"1A",X"10",X"FD",X"CA",
		X"06",X"EC",X"04",X"FD",X"CA",X"04",X"FF",X"CA",X"02",X"CC",X"1A",X"00",X"F7",X"CA",X"01",X"E6",
		X"88",X"12",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"EE",X"02",X"EF",X"88",X"14",X"EE",X"42",
		X"FF",X"CA",X"02",X"A6",X"0A",X"E6",X"0C",X"ED",X"04",X"FD",X"CA",X"04",X"86",X"0A",X"E6",X"0B",
		X"E7",X"88",X"12",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"35",X"C7",X"34",X"76",X"CE",X"98",
		X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",
		X"36",X"36",X"36",X"10",X"11",X"83",X"00",X"00",X"26",X"EE",X"35",X"F6",X"34",X"76",X"0C",X"F0",
		X"44",X"34",X"02",X"86",X"00",X"24",X"08",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"BD",
		X"D0",X"45",X"DD",X"2B",X"C6",X"03",X"E0",X"E0",X"A6",X"85",X"9B",X"2C",X"19",X"A7",X"85",X"5A",
		X"2B",X"0E",X"A6",X"85",X"99",X"2B",X"19",X"A7",X"85",X"86",X"00",X"97",X"2B",X"5A",X"2A",X"F2",
		X"DC",X"46",X"27",X"38",X"31",X"04",X"EC",X"84",X"10",X"A3",X"A4",X"26",X"05",X"EC",X"02",X"10",
		X"A3",X"22",X"25",X"28",X"A6",X"22",X"9B",X"47",X"19",X"A7",X"22",X"A6",X"21",X"99",X"46",X"19",
		X"A7",X"21",X"A6",X"A4",X"89",X"00",X"19",X"A7",X"A4",X"CC",X"D0",X"C9",X"BD",X"D0",X"4B",X"BD",
		X"D0",X"45",X"6C",X"08",X"BD",X"26",X"C9",X"C6",X"05",X"BD",X"D0",X"BD",X"8D",X"03",X"35",X"76",
		X"39",X"96",X"3F",X"C6",X"11",X"91",X"3F",X"26",X"02",X"C6",X"AA",X"34",X"02",X"D7",X"CF",X"4A",
		X"26",X"08",X"8E",X"18",X"0E",X"CE",X"BD",X"E4",X"20",X"06",X"8E",X"58",X"0E",X"CE",X"BE",X"20",
		X"CC",X"15",X"06",X"BD",X"D0",X"1B",X"30",X"89",X"FD",X"00",X"0F",X"D6",X"A6",X"C4",X"84",X"0F",
		X"BD",X"5F",X"9F",X"A6",X"41",X"BD",X"5F",X"9F",X"A6",X"42",X"BD",X"5F",X"9F",X"0C",X"D6",X"A6",
		X"43",X"BD",X"5F",X"9F",X"35",X"82",X"B6",X"C8",X"0E",X"86",X"01",X"9A",X"45",X"B7",X"C9",X"00",
		X"B6",X"CB",X"00",X"81",X"80",X"25",X"32",X"96",X"43",X"26",X"20",X"0C",X"43",X"0C",X"10",X"BD",
		X"D3",X"E0",X"BD",X"26",X"C0",X"B6",X"CB",X"00",X"7F",X"CA",X"01",X"D6",X"45",X"C5",X"02",X"27",
		X"0C",X"8B",X"10",X"97",X"41",X"BD",X"DC",X"FF",X"BD",X"DD",X"4E",X"20",X"54",X"80",X"10",X"97",
		X"41",X"BD",X"DD",X"90",X"BD",X"DD",X"3E",X"20",X"48",X"D6",X"43",X"27",X"44",X"0F",X"43",X"0C",
		X"10",X"C6",X"39",X"F7",X"CB",X"FF",X"81",X"04",X"22",X"1B",X"CE",X"C0",X"10",X"DC",X"0A",X"9E",
		X"0C",X"10",X"9E",X"0E",X"36",X"36",X"DC",X"04",X"9E",X"06",X"10",X"9E",X"08",X"36",X"36",X"DC",
		X"00",X"9E",X"02",X"36",X"16",X"0C",X"44",X"BD",X"D4",X"4D",X"7F",X"CA",X"01",X"D6",X"45",X"C5",
		X"02",X"27",X"08",X"BD",X"DC",X"E7",X"BD",X"DD",X"3E",X"20",X"06",X"BD",X"DD",X"60",X"BD",X"DD",
		X"4E",X"96",X"45",X"B7",X"C9",X"00",X"3B",X"96",X"59",X"85",X"08",X"26",X"11",X"9E",X"17",X"27",
		X"0D",X"EC",X"04",X"D1",X"41",X"22",X"03",X"BD",X"DD",X"CE",X"AE",X"84",X"26",X"F3",X"39",X"96",
		X"59",X"85",X"08",X"26",X"72",X"9E",X"17",X"27",X"34",X"EC",X"0A",X"EE",X"02",X"E3",X"0E",X"81",
		X"07",X"25",X"0A",X"AB",X"C4",X"81",X"90",X"22",X"04",X"A0",X"C4",X"ED",X"0A",X"EC",X"0C",X"E3",
		X"88",X"10",X"81",X"18",X"25",X"0A",X"AB",X"41",X"81",X"EB",X"22",X"04",X"A0",X"41",X"ED",X"0C",
		X"EC",X"04",X"D1",X"41",X"23",X"03",X"BD",X"DD",X"CE",X"AE",X"84",X"26",X"CC",X"39",X"96",X"59",
		X"85",X"10",X"26",X"09",X"8E",X"98",X"5A",X"DC",X"5E",X"D1",X"41",X"23",X"11",X"39",X"96",X"59",
		X"85",X"10",X"26",X"F9",X"8E",X"98",X"5A",X"DC",X"5E",X"D1",X"41",X"22",X"71",X"39",X"20",X"6E",
		X"96",X"59",X"85",X"08",X"26",X"10",X"9E",X"17",X"27",X"0C",X"EC",X"04",X"D1",X"41",X"23",X"02",
		X"8D",X"5C",X"AE",X"84",X"26",X"F4",X"39",X"96",X"59",X"85",X"02",X"26",X"12",X"96",X"44",X"84",
		X"07",X"26",X"0C",X"9E",X"17",X"27",X"08",X"EC",X"04",X"8D",X"43",X"AE",X"84",X"26",X"F8",X"39",
		X"96",X"59",X"85",X"08",X"26",X"E1",X"9E",X"17",X"27",X"33",X"EC",X"0A",X"EE",X"02",X"E3",X"0E",
		X"81",X"07",X"25",X"0A",X"AB",X"C4",X"81",X"90",X"22",X"04",X"A0",X"C4",X"ED",X"0A",X"EC",X"0C",
		X"E3",X"88",X"10",X"81",X"18",X"25",X"0A",X"AB",X"41",X"81",X"EB",X"22",X"04",X"A0",X"41",X"ED",
		X"0C",X"EC",X"04",X"D1",X"41",X"22",X"02",X"8D",X"05",X"AE",X"84",X"26",X"CD",X"39",X"FD",X"CA",
		X"04",X"EE",X"88",X"14",X"37",X"26",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"10",X"BF",X"CA",
		X"02",X"86",X"1A",X"E6",X"88",X"12",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"A6",X"0A",X"E6",
		X"0C",X"ED",X"04",X"FD",X"CA",X"04",X"EE",X"02",X"EF",X"88",X"14",X"EC",X"42",X"FD",X"CA",X"02",
		X"86",X"0A",X"E6",X"0B",X"E7",X"88",X"12",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"39",X"34",
		X"56",X"8E",X"DA",X"05",X"34",X"06",X"C6",X"FE",X"D4",X"45",X"D7",X"45",X"F7",X"C9",X"00",X"5F",
		X"6A",X"61",X"A6",X"61",X"EA",X"C6",X"4A",X"2A",X"FB",X"86",X"37",X"33",X"C9",X"01",X"00",X"6A",
		X"E4",X"26",X"EF",X"A1",X"89",X"BE",X"EE",X"27",X"12",X"96",X"86",X"81",X"01",X"22",X"0C",X"34",
		X"04",X"D6",X"85",X"86",X"98",X"1F",X"01",X"6A",X"84",X"35",X"04",X"86",X"01",X"9A",X"45",X"97",
		X"45",X"B7",X"C9",X"00",X"5D",X"32",X"62",X"35",X"D6",X"34",X"36",X"34",X"16",X"D6",X"45",X"C4",
		X"FE",X"D7",X"45",X"F7",X"C9",X"00",X"E6",X"84",X"E7",X"A0",X"30",X"89",X"01",X"00",X"4A",X"26",
		X"F5",X"AE",X"62",X"30",X"01",X"AF",X"62",X"A6",X"E4",X"6A",X"61",X"26",X"E9",X"32",X"64",X"96",
		X"45",X"8A",X"01",X"97",X"45",X"B7",X"C9",X"00",X"35",X"B6",X"20",X"52",X"4F",X"42",X"4F",X"54",
		X"52",X"4F",X"4E",X"3A",X"20",X"32",X"30",X"38",X"34",X"20",X"28",X"54",X"4D",X"29",X"20",X"20",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",
		X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",
		X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"35",X"06",X"DE",X"15",X"ED",X"C8",X"19",X"BD",X"D0",X"54",X"E2",X"6F",X"BD",X"E1",X"E3",X"86",
		X"99",X"97",X"D8",X"86",X"CC",X"97",X"D9",X"10",X"8E",X"CF",X"6E",X"DE",X"15",X"86",X"07",X"A7",
		X"47",X"CC",X"05",X"02",X"ED",X"48",X"CC",X"09",X"34",X"ED",X"4A",X"86",X"01",X"A7",X"4D",X"8E",
		X"1A",X"35",X"BD",X"E0",X"5C",X"86",X"AA",X"97",X"D8",X"86",X"DD",X"97",X"D9",X"10",X"8E",X"CD",
		X"5A",X"BD",X"E0",X"E9",X"8E",X"CD",X"5E",X"BD",X"D0",X"A2",X"30",X"1C",X"81",X"3A",X"26",X"05",
		X"8C",X"CD",X"38",X"24",X"F2",X"30",X"02",X"34",X"10",X"8E",X"15",X"7A",X"86",X"31",X"BD",X"5F",
		X"93",X"86",X"5C",X"BD",X"5F",X"93",X"30",X"89",X"03",X"00",X"10",X"8E",X"CD",X"38",X"1E",X"12",
		X"BD",X"D0",X"A2",X"1E",X"12",X"BD",X"5F",X"93",X"10",X"AC",X"E4",X"23",X"F1",X"30",X"89",X"02",
		X"00",X"10",X"8E",X"CD",X"60",X"BD",X"E1",X"37",X"9F",X"2B",X"8E",X"CC",X"16",X"BD",X"D0",X"A2",
		X"81",X"03",X"27",X"23",X"9E",X"2B",X"30",X"89",X"05",X"00",X"86",X"5B",X"BD",X"5F",X"93",X"10",
		X"8E",X"CD",X"32",X"C6",X"03",X"1E",X"12",X"BD",X"D0",X"A2",X"1E",X"12",X"BD",X"5F",X"93",X"5A",
		X"26",X"F3",X"86",X"5C",X"BD",X"5F",X"93",X"DE",X"15",X"86",X"05",X"A7",X"47",X"CC",X"0C",X"03",
		X"ED",X"48",X"CC",X"07",X"28",X"ED",X"4A",X"86",X"02",X"A7",X"4D",X"8E",X"14",X"88",X"10",X"8E",
		X"CD",X"68",X"8D",X"48",X"86",X"6E",X"BD",X"5F",X"99",X"BD",X"D0",X"54",X"E2",X"E0",X"BD",X"D0",
		X"54",X"E2",X"9A",X"BD",X"D0",X"54",X"E2",X"E9",X"BD",X"D0",X"54",X"E2",X"F5",X"DE",X"15",X"86",
		X"C8",X"A7",X"47",X"86",X"03",X"8E",X"E0",X"3B",X"7E",X"D0",X"66",X"6A",X"47",X"26",X"F4",X"86",
		X"FF",X"A7",X"47",X"86",X"04",X"8E",X"E0",X"4B",X"7E",X"D0",X"66",X"B6",X"C8",X"06",X"84",X"03",
		X"BA",X"C8",X"04",X"27",X"04",X"6A",X"47",X"26",X"EA",X"6E",X"D8",X"19",X"35",X"06",X"DE",X"15",
		X"ED",X"C8",X"12",X"AF",X"C8",X"16",X"AF",X"4E",X"10",X"AF",X"C8",X"10",X"A6",X"48",X"A7",X"4C",
		X"86",X"04",X"A7",X"C8",X"18",X"AE",X"4E",X"10",X"AE",X"C8",X"10",X"8D",X"6C",X"E6",X"4D",X"86",
		X"6F",X"BD",X"E1",X"6E",X"34",X"10",X"C6",X"03",X"1E",X"12",X"BD",X"D0",X"A2",X"1E",X"12",X"BD",
		X"E1",X"84",X"5A",X"26",X"F3",X"35",X"10",X"A6",X"47",X"C6",X"03",X"3D",X"54",X"5C",X"1F",X"98",
		X"E6",X"47",X"C1",X"05",X"26",X"01",X"4C",X"5F",X"30",X"8B",X"BD",X"E1",X"37",X"A6",X"4D",X"8B",
		X"01",X"19",X"A7",X"4D",X"1F",X"10",X"A6",X"C8",X"16",X"EB",X"4A",X"1F",X"01",X"6A",X"4C",X"27",
		X"13",X"6A",X"C8",X"18",X"26",X"B5",X"AF",X"4E",X"10",X"AF",X"C8",X"10",X"86",X"01",X"8E",X"E0",
		X"70",X"7E",X"D0",X"66",X"EC",X"C8",X"16",X"AB",X"4B",X"A7",X"C8",X"16",X"1F",X"01",X"A6",X"48",
		X"A7",X"4C",X"6A",X"49",X"26",X"DB",X"6E",X"D8",X"12",X"34",X"36",X"31",X"26",X"8E",X"BD",X"E4",
		X"8D",X"1C",X"27",X"0C",X"D6",X"40",X"5A",X"27",X"0F",X"8E",X"BE",X"20",X"8D",X"10",X"26",X"08",
		X"8D",X"23",X"27",X"04",X"96",X"D9",X"20",X"02",X"96",X"D8",X"97",X"CF",X"35",X"B6",X"34",X"20",
		X"1E",X"12",X"BD",X"D0",X"A2",X"84",X"0F",X"C6",X"04",X"A1",X"A0",X"26",X"06",X"BD",X"D0",X"A2",
		X"5A",X"26",X"F6",X"35",X"A0",X"31",X"21",X"30",X"2E",X"C6",X"07",X"A6",X"80",X"A8",X"A0",X"84",
		X"0F",X"26",X"03",X"5A",X"26",X"F5",X"39",X"1E",X"12",X"BD",X"D0",X"A2",X"BD",X"D0",X"A5",X"1E",
		X"12",X"84",X"0F",X"26",X"07",X"5D",X"26",X"04",X"86",X"63",X"20",X"0D",X"34",X"20",X"1F",X"02",
		X"86",X"62",X"BD",X"E1",X"6E",X"35",X"20",X"86",X"2A",X"34",X"02",X"1E",X"12",X"BD",X"D0",X"A8",
		X"1E",X"12",X"34",X"20",X"1F",X"02",X"A6",X"62",X"8D",X"04",X"35",X"20",X"35",X"82",X"34",X"52",
		X"8E",X"5F",X"99",X"A6",X"47",X"81",X"07",X"27",X"03",X"8E",X"5F",X"96",X"1F",X"13",X"35",X"12",
		X"AD",X"C4",X"35",X"C0",X"34",X"52",X"8E",X"5F",X"93",X"A6",X"47",X"81",X"07",X"27",X"ED",X"8E",
		X"5F",X"90",X"20",X"E8",X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",X"3A",X"20",X"32",
		X"30",X"38",X"34",X"20",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",
		X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",
		X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",
		X"45",X"44",X"20",X"35",X"06",X"DE",X"15",X"ED",X"4F",X"8E",X"98",X"00",X"CC",X"00",X"00",X"ED",
		X"81",X"8C",X"98",X"10",X"25",X"F9",X"8E",X"06",X"0D",X"AF",X"C8",X"17",X"86",X"11",X"A7",X"C8",
		X"15",X"8E",X"3E",X"7D",X"AF",X"C8",X"11",X"10",X"8E",X"59",X"7F",X"10",X"AF",X"C8",X"13",X"86",
		X"02",X"A7",X"C8",X"16",X"AE",X"C8",X"11",X"10",X"AE",X"C8",X"13",X"A6",X"C8",X"15",X"BD",X"E3",
		X"13",X"AC",X"C8",X"17",X"27",X"32",X"30",X"89",X"FE",X"FE",X"31",X"A9",X"01",X"02",X"8D",X"17",
		X"6A",X"C8",X"16",X"26",X"E9",X"A7",X"C8",X"15",X"AF",X"C8",X"11",X"10",X"AF",X"C8",X"13",X"86",
		X"01",X"8E",X"E2",X"0F",X"7E",X"D0",X"66",X"34",X"04",X"E6",X"C8",X"17",X"C1",X"06",X"26",X"06",
		X"80",X"11",X"26",X"02",X"86",X"88",X"35",X"84",X"AE",X"C8",X"17",X"8C",X"06",X"0D",X"27",X"03",
		X"6E",X"D8",X"0F",X"8E",X"0E",X"1D",X"AF",X"C8",X"17",X"6F",X"C8",X"15",X"7E",X"E2",X"01",X"8E",
		X"E2",X"FE",X"A6",X"80",X"8D",X"13",X"AF",X"47",X"86",X"03",X"8E",X"E2",X"80",X"7E",X"D0",X"66",
		X"AE",X"47",X"8C",X"E3",X"13",X"25",X"EB",X"20",X"E6",X"10",X"8E",X"98",X"01",X"E6",X"21",X"E7",
		X"A0",X"10",X"8C",X"98",X"08",X"25",X"F6",X"A7",X"A4",X"39",X"10",X"8E",X"98",X"0A",X"8E",X"E2",
		X"C2",X"CC",X"E2",X"C2",X"ED",X"4B",X"10",X"AF",X"49",X"20",X"02",X"AE",X"4B",X"AF",X"47",X"AE",
		X"47",X"A6",X"80",X"27",X"F6",X"A7",X"D8",X"09",X"AF",X"47",X"86",X"04",X"8E",X"E2",X"AF",X"7E",
		X"D0",X"66",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"57",X"A7",X"FF",X"FF",X"A7",X"57",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"D2",X"C0",X"C0",X"C0",X"D2",X"E4",X"00",
		X"8E",X"E2",X"C9",X"10",X"8E",X"98",X"09",X"20",X"B8",X"8E",X"E2",X"D8",X"10",X"8E",X"98",X"0C",
		X"CC",X"E2",X"D1",X"20",X"AF",X"8E",X"E2",X"D1",X"10",X"8E",X"98",X"0D",X"20",X"F2",X"37",X"2F",
		X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",X"CA",X"C0",X"D0",
		X"98",X"38",X"33",X"34",X"36",X"DE",X"15",X"84",X"F0",X"A7",X"4B",X"A6",X"E4",X"84",X"0F",X"A7",
		X"4C",X"1F",X"10",X"A7",X"49",X"E7",X"47",X"1F",X"20",X"A7",X"4A",X"E7",X"48",X"E0",X"47",X"56",
		X"24",X"02",X"6A",X"48",X"A6",X"47",X"8D",X"3B",X"4C",X"8D",X"4A",X"A6",X"48",X"8D",X"34",X"4A",
		X"8D",X"43",X"A6",X"49",X"8D",X"0B",X"8D",X"17",X"A6",X"4A",X"8D",X"05",X"4A",X"8D",X"10",X"35",
		X"B6",X"34",X"16",X"8D",X"14",X"5C",X"A6",X"4B",X"A7",X"81",X"5A",X"26",X"FB",X"35",X"96",X"34",
		X"16",X"8D",X"06",X"30",X"01",X"A6",X"4C",X"20",X"EF",X"E6",X"47",X"1F",X"01",X"E6",X"48",X"E0",
		X"47",X"54",X"39",X"34",X"16",X"8D",X"16",X"5C",X"A6",X"4B",X"A7",X"84",X"30",X"89",X"01",X"00",
		X"5A",X"26",X"F7",X"35",X"96",X"34",X"16",X"8D",X"04",X"A6",X"4C",X"20",X"ED",X"1F",X"89",X"A6",
		X"49",X"1F",X"01",X"E6",X"4A",X"E0",X"49",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"E5",X"F5",X"7E",X"E6",X"F7",X"7E",X"E8",X"A5",X"7E",X"E4",X"33",X"7E",X"E4",X"13",X"7E",
		X"E3",X"E2",X"86",X"18",X"A7",X"47",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"08",X"8E",X"E3",X"F3",
		X"7E",X"D0",X"66",X"B6",X"C8",X"0C",X"85",X"08",X"27",X"16",X"6A",X"47",X"26",X"ED",X"10",X"8E",
		X"CD",X"32",X"8E",X"E4",X"6C",X"C6",X"17",X"BD",X"6F",X"0C",X"BD",X"E5",X"BC",X"7F",X"C8",X"0E",
		X"7E",X"D0",X"63",X"10",X"8E",X"CD",X"68",X"C6",X"08",X"BD",X"E5",X"E3",X"A8",X"26",X"84",X"0F",
		X"27",X"03",X"5A",X"27",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"6E",
		X"25",X"E7",X"39",X"86",X"39",X"B7",X"CB",X"FF",X"8E",X"E4",X"6C",X"10",X"8E",X"CD",X"32",X"C6",
		X"92",X"BD",X"6F",X"0C",X"8E",X"E4",X"FE",X"10",X"8E",X"CE",X"56",X"C6",X"8C",X"BD",X"6F",X"0C",
		X"BD",X"E5",X"BC",X"10",X"8E",X"CD",X"68",X"BD",X"E5",X"DB",X"86",X"39",X"B7",X"CB",X"FF",X"31",
		X"2E",X"10",X"8C",X"CF",X"6E",X"25",X"F0",X"86",X"5D",X"7E",X"5F",X"99",X"42",X"49",X"4C",X"57",
		X"49",X"4C",X"4C",X"59",X"3A",X"45",X"4C",X"4B",X"54",X"52",X"49",X"58",X"3A",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"00",X"15",X"17",X"82",X"56",X"49",X"44",X"00",X"12",X"21",X"45",X"4B",X"49",
		X"44",X"00",X"12",X"21",X"35",X"44",X"52",X"4A",X"00",X"05",X"21",X"27",X"4C",X"45",X"44",X"00",
		X"05",X"02",X"18",X"45",X"50",X"4A",X"00",X"04",X"12",X"55",X"4A",X"45",X"52",X"00",X"04",X"12",
		X"50",X"4B",X"49",X"44",X"00",X"03",X"19",X"20",X"4D",X"4C",X"47",X"00",X"03",X"19",X"19",X"53",
		X"53",X"52",X"00",X"02",X"66",X"45",X"55",X"4E",X"41",X"00",X"02",X"66",X"35",X"4A",X"52",X"53",
		X"00",X"02",X"52",X"50",X"43",X"4A",X"4D",X"00",X"02",X"41",X"10",X"4B",X"4A",X"46",X"00",X"02",
		X"30",X"20",X"4D",X"52",X"53",X"00",X"02",X"20",X"35",X"50",X"47",X"44",X"00",X"02",X"10",X"90",
		X"4E",X"4A",X"4D",X"00",X"02",X"09",X"65",X"4E",X"48",X"44",X"00",X"02",X"09",X"60",X"44",X"4F",
		X"4E",X"00",X"01",X"82",X"80",X"56",X"49",X"56",X"00",X"01",X"82",X"80",X"47",X"57",X"57",X"00",
		X"01",X"81",X"05",X"43",X"52",X"42",X"00",X"01",X"80",X"55",X"4D",X"44",X"52",X"00",X"01",X"75",
		X"65",X"42",X"41",X"43",X"00",X"01",X"72",X"56",X"57",X"3A",X"52",X"00",X"01",X"70",X"70",X"4D",
		X"50",X"54",X"00",X"01",X"60",X"60",X"53",X"55",X"45",X"00",X"01",X"55",X"20",X"4D",X"4F",X"4D",
		X"00",X"01",X"44",X"80",X"44",X"41",X"44",X"00",X"01",X"44",X"79",X"53",X"46",X"44",X"00",X"01",
		X"44",X"78",X"41",X"4B",X"44",X"00",X"01",X"44",X"77",X"43",X"57",X"4B",X"00",X"01",X"33",X"30",
		X"54",X"4D",X"48",X"00",X"01",X"32",X"70",X"45",X"4A",X"53",X"00",X"01",X"31",X"20",X"52",X"41",
		X"59",X"00",X"01",X"30",X"65",X"47",X"41",X"59",X"00",X"01",X"29",X"65",X"52",X"4B",X"4D",X"00",
		X"01",X"28",X"55",X"43",X"4E",X"53",X"00",X"01",X"27",X"55",X"3A",X"3A",X"3A",X"00",X"01",X"00",
		X"00",X"C0",X"01",X"01",X"1B",X"01",X"01",X"02",X"00",X"C0",X"01",X"FF",X"3C",X"01",X"FF",X"00",
		X"01",X"20",X"00",X"01",X"C0",X"36",X"01",X"60",X"3D",X"02",X"0A",X"11",X"02",X"40",X"3E",X"00",
		X"34",X"34",X"8E",X"E5",X"8A",X"C6",X"07",X"BD",X"6F",X"0C",X"35",X"B4",X"34",X"02",X"8D",X"05",
		X"B7",X"CD",X"60",X"35",X"82",X"34",X"10",X"8E",X"CD",X"32",X"4F",X"AB",X"84",X"30",X"01",X"8C",
		X"CD",X"60",X"27",X"F9",X"8C",X"CD",X"68",X"26",X"F2",X"35",X"90",X"34",X"02",X"8D",X"04",X"A7",
		X"26",X"35",X"82",X"34",X"24",X"C6",X"0E",X"4F",X"C1",X"08",X"27",X"02",X"AB",X"A4",X"31",X"21",
		X"5A",X"26",X"F5",X"35",X"A4",X"86",X"32",X"34",X"02",X"10",X"8E",X"CD",X"68",X"8D",X"E4",X"A8",
		X"26",X"84",X"0F",X"27",X"0F",X"BD",X"E6",X"CC",X"7F",X"CD",X"00",X"7F",X"CD",X"01",X"6A",X"E4",
		X"27",X"12",X"20",X"E9",X"86",X"03",X"C6",X"04",X"8D",X"68",X"25",X"E9",X"31",X"2E",X"10",X"8C",
		X"CF",X"6E",X"25",X"D9",X"35",X"02",X"8E",X"E4",X"95",X"10",X"8E",X"CF",X"6E",X"C6",X"46",X"BD",
		X"6F",X"0C",X"8D",X"91",X"B8",X"CD",X"60",X"84",X"0F",X"27",X"02",X"8D",X"0F",X"10",X"8E",X"CD",
		X"32",X"86",X"17",X"C6",X"04",X"8D",X"3B",X"24",X"02",X"8D",X"01",X"39",X"8E",X"CD",X"38",X"86",
		X"3A",X"BD",X"D0",X"AB",X"8C",X"CD",X"60",X"25",X"F8",X"8E",X"CD",X"68",X"10",X"8E",X"CD",X"38",
		X"86",X"06",X"BD",X"E6",X"EC",X"10",X"8E",X"CD",X"32",X"BD",X"E6",X"EC",X"8E",X"CD",X"6E",X"10",
		X"8E",X"CD",X"60",X"86",X"08",X"BD",X"E6",X"EC",X"BD",X"E5",X"BC",X"10",X"8E",X"CD",X"68",X"7E",
		X"E6",X"CC",X"34",X"16",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"21",X"BD",X"D0",X"A5",X"C1",X"41",
		X"24",X"04",X"C1",X"3A",X"26",X"32",X"C1",X"5A",X"22",X"2E",X"4A",X"26",X"EE",X"A6",X"61",X"BD",
		X"D0",X"A5",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",X"D0",X"A5",X"34",X"04",X"C4",X"0F",
		X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",X"22",X"0C",X"4A",X"26",X"EA",X"1C",
		X"FE",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"96",X"1A",X"01",X"20",X"F5",X"34",X"36",X"30",X"2E",
		X"8C",X"CF",X"6E",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",X"2E",X"30",X"0E",X"86",X"39",X"B7",
		X"CB",X"FF",X"20",X"EC",X"BD",X"E5",X"B0",X"BD",X"E5",X"DB",X"35",X"B6",X"34",X"36",X"E6",X"80",
		X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"BD",X"D0",X"60",X"BD",X"D0",X"12",X"BD",X"D0",X"33",
		X"BD",X"D0",X"99",X"8E",X"BD",X"E4",X"C6",X"01",X"8D",X"20",X"D6",X"40",X"5A",X"27",X"18",X"BD",
		X"D0",X"12",X"B6",X"C8",X"06",X"2A",X"03",X"BD",X"D0",X"9C",X"8E",X"BE",X"20",X"C6",X"02",X"8D",
		X"09",X"BD",X"D0",X"12",X"BD",X"D0",X"99",X"7E",X"77",X"A0",X"35",X"20",X"10",X"BF",X"B3",X"E4",
		X"BF",X"B3",X"E8",X"D7",X"3F",X"BD",X"E9",X"0E",X"24",X"5B",X"BD",X"E8",X"B5",X"10",X"8E",X"CD",
		X"68",X"8E",X"CF",X"60",X"BD",X"E8",X"8F",X"8E",X"CD",X"60",X"10",X"8E",X"CD",X"6E",X"86",X"08",
		X"BD",X"E6",X"EC",X"8E",X"CD",X"32",X"10",X"8E",X"CD",X"68",X"86",X"06",X"BD",X"E6",X"EC",X"10",
		X"8E",X"CD",X"68",X"BD",X"E5",X"DB",X"BE",X"B3",X"E8",X"10",X"8E",X"CD",X"60",X"C6",X"04",X"BD",
		X"6F",X"0C",X"BD",X"E5",X"BC",X"8E",X"E5",X"8A",X"10",X"8E",X"CD",X"32",X"C6",X"03",X"BD",X"6F",
		X"0C",X"BD",X"D0",X"12",X"86",X"60",X"B7",X"B3",X"E6",X"8E",X"CC",X"16",X"BD",X"D0",X"A5",X"C1",
		X"03",X"27",X"42",X"20",X"22",X"BD",X"E9",X"1B",X"25",X"09",X"BD",X"E9",X"38",X"25",X"04",X"6E",
		X"9F",X"B3",X"E4",X"7F",X"B3",X"E6",X"CC",X"E5",X"91",X"10",X"8C",X"CF",X"6E",X"26",X"03",X"CC",
		X"E5",X"99",X"BD",X"E9",X"71",X"86",X"5F",X"D6",X"3F",X"BD",X"D0",X"12",X"BD",X"5F",X"99",X"CC",
		X"3A",X"3A",X"FD",X"B3",X"EA",X"B7",X"B3",X"EC",X"CC",X"03",X"00",X"8E",X"46",X"80",X"10",X"8E",
		X"B3",X"EA",X"BD",X"6F",X"09",X"BD",X"E9",X"1B",X"24",X"06",X"8E",X"CF",X"EC",X"BD",X"E8",X"75",
		X"BD",X"E9",X"38",X"24",X"43",X"7D",X"B3",X"E6",X"27",X"1C",X"8E",X"B3",X"EA",X"10",X"8E",X"CD",
		X"32",X"C6",X"03",X"BD",X"6F",X"0C",X"BD",X"E5",X"BC",X"86",X"05",X"8D",X"2F",X"24",X"29",X"1F",
		X"12",X"BD",X"E6",X"CC",X"20",X"12",X"BD",X"E8",X"30",X"34",X"01",X"34",X"10",X"10",X"AC",X"E1",
		X"22",X"02",X"8D",X"61",X"35",X"01",X"24",X"10",X"BD",X"D0",X"12",X"86",X"64",X"BD",X"5F",X"99",
		X"86",X"60",X"8E",X"E8",X"28",X"7E",X"D0",X"66",X"6E",X"9F",X"B3",X"E4",X"34",X"26",X"20",X"0C",
		X"34",X"26",X"8E",X"CD",X"32",X"8D",X"24",X"86",X"04",X"25",X"01",X"4C",X"97",X"2B",X"8E",X"CD",
		X"68",X"8D",X"18",X"24",X"04",X"0A",X"2B",X"27",X"0E",X"30",X"0E",X"8C",X"CF",X"6E",X"25",X"F1",
		X"8E",X"CF",X"60",X"1C",X"FE",X"35",X"A6",X"1A",X"01",X"35",X"A6",X"34",X"10",X"10",X"8E",X"B3",
		X"EA",X"C6",X"03",X"BD",X"D0",X"A2",X"A1",X"A0",X"26",X"07",X"5A",X"26",X"F6",X"1A",X"01",X"35",
		X"90",X"1C",X"FE",X"35",X"90",X"34",X"20",X"BD",X"E8",X"8F",X"8E",X"B3",X"EA",X"C6",X"03",X"BD",
		X"6F",X"0C",X"BE",X"B3",X"E8",X"C6",X"04",X"BD",X"6F",X"0C",X"35",X"20",X"7E",X"E5",X"DB",X"34",
		X"30",X"1F",X"12",X"10",X"AC",X"62",X"27",X"0B",X"30",X"32",X"86",X"0E",X"BD",X"E6",X"EC",X"31",
		X"32",X"20",X"F0",X"35",X"B0",X"35",X"06",X"FD",X"B3",X"E4",X"C6",X"01",X"8D",X"07",X"BD",X"E5",
		X"BC",X"6E",X"9F",X"B3",X"E4",X"35",X"20",X"10",X"BF",X"B3",X"E6",X"4F",X"1F",X"02",X"CC",X"E5",
		X"99",X"BD",X"E9",X"71",X"8E",X"CC",X"16",X"BD",X"D0",X"A5",X"BD",X"D0",X"12",X"C1",X"03",X"26",
		X"0E",X"D6",X"3F",X"86",X"5F",X"BD",X"5F",X"99",X"86",X"03",X"8E",X"46",X"80",X"20",X"0D",X"86",
		X"5E",X"BD",X"5F",X"99",X"1F",X"98",X"BD",X"D0",X"C6",X"8E",X"2D",X"80",X"10",X"8E",X"B3",X"FE",
		X"C6",X"3A",X"E7",X"A2",X"10",X"8C",X"B3",X"EA",X"22",X"F8",X"5F",X"BD",X"6F",X"09",X"8E",X"B3",
		X"EA",X"10",X"8E",X"CD",X"38",X"C6",X"14",X"BD",X"6F",X"0C",X"6E",X"9F",X"B3",X"E6",X"34",X"30",
		X"10",X"8E",X"CD",X"60",X"BE",X"B3",X"E8",X"8D",X"38",X"35",X"B0",X"34",X"10",X"10",X"8E",X"CF",
		X"74",X"BE",X"B3",X"E8",X"8D",X"2B",X"25",X"0C",X"31",X"2E",X"10",X"8C",X"CF",X"FA",X"25",X"F4",
		X"1C",X"FE",X"35",X"90",X"31",X"3A",X"35",X"90",X"34",X"10",X"10",X"8E",X"CD",X"60",X"BE",X"B3",
		X"E8",X"8D",X"0E",X"25",X"EF",X"31",X"2E",X"10",X"8C",X"CF",X"60",X"25",X"F4",X"1C",X"FE",X"35",
		X"90",X"34",X"36",X"1E",X"12",X"C6",X"04",X"BD",X"D0",X"A2",X"C1",X"04",X"26",X"02",X"84",X"0F",
		X"A1",X"A0",X"22",X"05",X"25",X"07",X"5A",X"26",X"EE",X"1C",X"FE",X"35",X"B6",X"1A",X"01",X"35",
		X"B6",X"0F",X"56",X"7E",X"D0",X"4B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"CC",X"EC",X"34",X"EA",X"2A",X"EA",X"35",
		X"EA",X"40",X"EA",X"4B",X"EA",X"56",X"EA",X"61",X"EA",X"6C",X"EA",X"77",X"EA",X"82",X"EA",X"8D",
		X"EA",X"98",X"EA",X"9E",X"EA",X"A4",X"EA",X"AF",X"EA",X"B5",X"EA",X"C5",X"EA",X"CB",X"EA",X"D6",
		X"EA",X"E1",X"EA",X"EC",X"EA",X"F7",X"EB",X"02",X"EB",X"0D",X"EB",X"18",X"EB",X"23",X"EB",X"2E",
		X"EB",X"39",X"EB",X"44",X"EB",X"4F",X"EB",X"5A",X"EB",X"6A",X"EB",X"75",X"EB",X"80",X"EB",X"8B",
		X"EB",X"96",X"EB",X"A1",X"EB",X"AC",X"EB",X"B7",X"EB",X"C2",X"EB",X"CD",X"EB",X"DD",X"EB",X"E8",
		X"EB",X"F3",X"EB",X"FE",X"EC",X"09",X"EC",X"14",X"EC",X"29",X"03",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"F0",X"03",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"03",X"FF",X"F0",X"00",X"F0",X"FF",X"F0",X"F0",X"00",X"FF",X"F0",X"03",X"FF",X"F0",X"00",X"F0",
		X"0F",X"F0",X"00",X"F0",X"FF",X"F0",X"03",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"00",X"F0",X"00",
		X"F0",X"03",X"FF",X"F0",X"F0",X"00",X"FF",X"F0",X"00",X"F0",X"FF",X"F0",X"03",X"FF",X"F0",X"F0",
		X"00",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"03",X"FF",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",
		X"00",X"F0",X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"03",X"FF",X"F0",
		X"F0",X"F0",X"FF",X"F0",X"00",X"F0",X"00",X"F0",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"F0",
		X"F0",X"F0",X"00",X"F0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"00",X"01",
		X"00",X"00",X"00",X"00",X"F0",X"05",X"00",X"F0",X"00",X"0F",X"FF",X"00",X"FF",X"FF",X"F0",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"01",X"00",X"F0",X"00",X"F0",X"00",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"F0",X"00",X"00",X"00",X"00",X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"FF",X"F0",X"03",X"FF",X"F0",X"F0",
		X"00",X"F0",X"00",X"F0",X"00",X"FF",X"F0",X"03",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"00",X"03",X"FF",X"F0",X"F0",X"00",X"FF",X"00",X"F0",X"00",X"FF",X"F0",X"03",X"FF",X"F0",
		X"F0",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"00",X"03",X"FF",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",
		X"F0",X"FF",X"F0",X"03",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"FF",
		X"F0",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"FF",X"F0",X"03",X"00",X"F0",X"00",X"F0",X"00",X"F0",
		X"F0",X"F0",X"FF",X"F0",X"03",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"03",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"F0",X"05",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"00",X"F0",X"03",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"03",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",
		X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"00",X"F0",X"00",X"03",X"FF",X"F0",X"F0",X"F0",
		X"FF",X"F0",X"00",X"F0",X"00",X"F0",X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",
		X"F0",X"03",X"FF",X"F0",X"F0",X"00",X"FF",X"F0",X"00",X"F0",X"FF",X"F0",X"03",X"FF",X"F0",X"0F",
		X"00",X"0F",X"00",X"0F",X"00",X"0F",X"00",X"03",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"F0",X"03",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"00",X"0F",X"00",X"05",X"F0",X"00",
		X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"03",X"F0",X"F0",
		X"F0",X"F0",X"0F",X"00",X"F0",X"F0",X"F0",X"F0",X"03",X"F0",X"F0",X"F0",X"F0",X"FF",X"F0",X"0F",
		X"00",X"0F",X"00",X"03",X"FF",X"F0",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"FF",X"F0",X"03",X"0F",
		X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"03",X"0F",X"00",X"00",X"F0",X"00",X"F0",
		X"00",X"F0",X"0F",X"00",X"07",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"03",X"00",X"F0",X"00",X"F0",X"0F",X"00",
		X"F0",X"00",X"F0",X"00",X"EC",X"92",X"EC",X"A5",X"EC",X"B8",X"EC",X"CB",X"EC",X"DE",X"EC",X"F1",
		X"ED",X"04",X"ED",X"17",X"ED",X"2A",X"ED",X"3D",X"ED",X"50",X"ED",X"5D",X"ED",X"6C",X"ED",X"79",
		X"ED",X"86",X"ED",X"A5",X"ED",X"B2",X"ED",X"BF",X"ED",X"D2",X"ED",X"E5",X"ED",X"F8",X"EE",X"0B",
		X"EE",X"1E",X"EE",X"31",X"EE",X"44",X"EE",X"57",X"EE",X"6A",X"EE",X"7D",X"EE",X"90",X"EE",X"A3",
		X"EE",X"B6",X"EE",X"C9",X"EE",X"DC",X"EE",X"EF",X"EF",X"02",X"EF",X"15",X"EF",X"28",X"EF",X"3B",
		X"EF",X"4E",X"EF",X"61",X"EF",X"74",X"EF",X"87",X"EF",X"9A",X"EF",X"AD",X"EF",X"BA",X"EF",X"C7",
		X"EF",X"DA",X"05",X"99",X"99",X"90",X"90",X"00",X"90",X"90",X"00",X"90",X"90",X"00",X"90",X"90",
		X"00",X"90",X"99",X"99",X"90",X"05",X"00",X"99",X"00",X"00",X"09",X"00",X"00",X"09",X"00",X"00",
		X"09",X"00",X"00",X"09",X"00",X"09",X"99",X"90",X"05",X"09",X"99",X"90",X"00",X"00",X"90",X"99",
		X"99",X"90",X"90",X"00",X"00",X"90",X"00",X"00",X"99",X"99",X"00",X"05",X"09",X"99",X"90",X"00",
		X"00",X"90",X"09",X"99",X"90",X"00",X"00",X"90",X"00",X"00",X"90",X"99",X"99",X"90",X"05",X"90",
		X"00",X"00",X"90",X"09",X"00",X"90",X"09",X"00",X"99",X"99",X"90",X"00",X"09",X"00",X"00",X"09",
		X"00",X"05",X"99",X"99",X"00",X"90",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"90",X"00",X"00",
		X"90",X"99",X"99",X"90",X"05",X"99",X"99",X"00",X"90",X"00",X"00",X"99",X"99",X"90",X"90",X"00",
		X"90",X"90",X"00",X"90",X"99",X"99",X"90",X"05",X"99",X"99",X"90",X"00",X"00",X"90",X"00",X"09",
		X"00",X"00",X"90",X"00",X"09",X"00",X"00",X"90",X"00",X"00",X"05",X"99",X"99",X"90",X"90",X"00",
		X"90",X"99",X"99",X"90",X"90",X"00",X"90",X"90",X"00",X"90",X"99",X"99",X"90",X"05",X"99",X"99",
		X"90",X"90",X"00",X"90",X"99",X"99",X"90",X"00",X"00",X"90",X"00",X"00",X"90",X"09",X"99",X"90",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"FF",X"00",X"09",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"02",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"00",X"05",
		X"66",X"66",X"60",X"60",X"06",X"60",X"66",X"66",X"60",X"60",X"06",X"60",X"60",X"06",X"60",X"60",
		X"06",X"60",X"05",X"66",X"66",X"00",X"60",X"06",X"00",X"66",X"66",X"60",X"66",X"00",X"60",X"66",
		X"00",X"60",X"66",X"66",X"60",X"05",X"66",X"66",X"60",X"66",X"00",X"00",X"66",X"00",X"00",X"66",
		X"00",X"00",X"66",X"00",X"00",X"66",X"66",X"60",X"05",X"66",X"66",X"00",X"66",X"00",X"60",X"66",
		X"00",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"66",X"00",X"05",X"66",X"66",X"60",X"60",
		X"00",X"00",X"66",X"66",X"60",X"66",X"00",X"00",X"66",X"00",X"00",X"66",X"66",X"60",X"05",X"66",
		X"66",X"60",X"60",X"00",X"00",X"66",X"66",X"60",X"66",X"00",X"00",X"66",X"00",X"00",X"66",X"00",
		X"00",X"05",X"66",X"66",X"60",X"66",X"06",X"60",X"66",X"00",X"00",X"66",X"06",X"60",X"66",X"00",
		X"60",X"66",X"66",X"60",X"05",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"66",X"60",X"66",X"00",
		X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"04",X"06",X"60",X"00",X"06",X"60",X"00",X"06",X"60",
		X"00",X"06",X"60",X"00",X"06",X"60",X"00",X"06",X"60",X"00",X"05",X"00",X"00",X"60",X"00",X"00",
		X"60",X"00",X"00",X"60",X"00",X"00",X"60",X"66",X"00",X"60",X"66",X"66",X"60",X"05",X"66",X"00",
		X"60",X"66",X"06",X"00",X"66",X"60",X"00",X"66",X"60",X"00",X"66",X"06",X"00",X"66",X"00",X"60",
		X"05",X"60",X"00",X"00",X"60",X"00",X"00",X"60",X"00",X"00",X"60",X"00",X"00",X"66",X"66",X"60",
		X"66",X"66",X"60",X"05",X"66",X"66",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"60",X"00",X"60",
		X"60",X"00",X"60",X"60",X"00",X"60",X"05",X"66",X"66",X"60",X"60",X"00",X"60",X"66",X"00",X"60",
		X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"05",X"66",X"66",X"60",X"60",X"06",X"60",
		X"60",X"00",X"60",X"60",X"00",X"60",X"60",X"00",X"60",X"66",X"66",X"60",X"05",X"66",X"66",X"60",
		X"60",X"00",X"60",X"66",X"66",X"60",X"66",X"00",X"00",X"66",X"00",X"00",X"66",X"00",X"00",X"05",
		X"66",X"66",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"06",X"00",X"66",
		X"60",X"60",X"05",X"66",X"66",X"00",X"60",X"06",X"00",X"66",X"66",X"60",X"66",X"00",X"60",X"66",
		X"00",X"60",X"66",X"00",X"60",X"05",X"66",X"66",X"60",X"60",X"00",X"00",X"66",X"66",X"60",X"00",
		X"00",X"60",X"66",X"00",X"60",X"66",X"66",X"60",X"05",X"66",X"66",X"60",X"00",X"60",X"00",X"00",
		X"66",X"00",X"00",X"66",X"00",X"00",X"66",X"00",X"00",X"66",X"00",X"05",X"60",X"06",X"60",X"60",
		X"06",X"60",X"60",X"06",X"60",X"60",X"06",X"60",X"60",X"06",X"60",X"66",X"66",X"60",X"05",X"66",
		X"00",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"00",X"60",X"06",X"06",X"00",X"00",X"60",
		X"00",X"05",X"60",X"00",X"60",X"60",X"00",X"60",X"60",X"00",X"60",X"60",X"60",X"60",X"60",X"60",
		X"60",X"66",X"66",X"60",X"05",X"60",X"00",X"60",X"06",X"06",X"00",X"00",X"60",X"00",X"00",X"60",
		X"00",X"06",X"06",X"00",X"60",X"00",X"60",X"05",X"66",X"00",X"60",X"66",X"00",X"60",X"66",X"66",
		X"60",X"00",X"60",X"00",X"00",X"60",X"00",X"00",X"60",X"00",X"05",X"66",X"66",X"60",X"00",X"06",
		X"00",X"00",X"60",X"00",X"06",X"00",X"00",X"66",X"66",X"60",X"66",X"66",X"60",X"03",X"00",X"F0",
		X"0F",X"00",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"00",X"F0",X"03",X"F0",X"00",X"0F",X"00",X"00",
		X"F0",X"00",X"F0",X"0F",X"00",X"F0",X"00",X"04",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"F0",
		X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"05",X"00",X"F0",X"00",X"0F",X"F0",
		X"00",X"FF",X"FF",X"F0",X"0F",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"D1",X"06",X"D1",X"06",X"D1",X"06",X"D1",X"06",X"DC",X"56",X"D1",X"06",X"D1",X"06",X"D1",X"06",
		X"7E",X"F4",X"31",X"7E",X"F4",X"A0",X"7E",X"F6",X"1B",X"7E",X"F0",X"1D",X"7E",X"F0",X"D7",X"7E",
		X"F0",X"66",X"7E",X"F3",X"4A",X"F1",X"24",X"F1",X"D5",X"F3",X"68",X"F3",X"EB",X"34",X"16",X"8E",
		X"B3",X"E4",X"9F",X"AD",X"30",X"89",X"00",X"F2",X"AF",X"89",X"FF",X"0E",X"8C",X"BA",X"82",X"CC",
		X"00",X"00",X"ED",X"84",X"DD",X"A9",X"DD",X"AB",X"35",X"96",X"34",X"10",X"DE",X"AD",X"27",X"0E",
		X"AE",X"C4",X"9F",X"AD",X"9E",X"A9",X"AF",X"C4",X"DF",X"A9",X"1C",X"FE",X"35",X"90",X"1A",X"01",
		X"35",X"90",X"34",X"10",X"DE",X"AD",X"27",X"F6",X"AE",X"C4",X"9F",X"AD",X"9E",X"AB",X"AF",X"C4",
		X"DF",X"AB",X"1C",X"FE",X"35",X"90",X"34",X"76",X"BD",X"F0",X"52",X"25",X"66",X"EC",X"04",X"AE",
		X"02",X"ED",X"49",X"D6",X"A6",X"E7",X"44",X"E0",X"49",X"25",X"04",X"E1",X"84",X"25",X"0A",X"E6",
		X"84",X"E7",X"45",X"EB",X"49",X"E7",X"44",X"20",X"03",X"58",X"E7",X"45",X"CC",X"46",X"46",X"ED",
		X"4F",X"EC",X"84",X"ED",X"4B",X"86",X"01",X"A7",X"C8",X"11",X"88",X"04",X"C8",X"04",X"ED",X"4D",
		X"AE",X"02",X"AF",X"42",X"CC",X"10",X"00",X"ED",X"46",X"30",X"C8",X"11",X"9F",X"B0",X"10",X"AE",
		X"42",X"E6",X"4C",X"D7",X"B3",X"9E",X"B0",X"30",X"01",X"9F",X"B0",X"A6",X"4B",X"97",X"B2",X"A6",
		X"A0",X"A7",X"84",X"3A",X"48",X"48",X"48",X"48",X"A7",X"84",X"3A",X"0A",X"B2",X"26",X"F0",X"0A",
		X"B3",X"26",X"E2",X"1C",X"FE",X"35",X"F6",X"34",X"76",X"BD",X"D0",X"15",X"BD",X"F0",X"3A",X"25",
		X"F2",X"EC",X"04",X"AE",X"02",X"ED",X"49",X"D6",X"A6",X"E7",X"44",X"E0",X"49",X"25",X"04",X"E1",
		X"84",X"25",X"0A",X"E6",X"84",X"E7",X"45",X"EB",X"49",X"E7",X"44",X"20",X"03",X"58",X"E7",X"45",
		X"CC",X"46",X"46",X"ED",X"4F",X"EC",X"84",X"ED",X"4B",X"48",X"A7",X"C8",X"11",X"86",X"01",X"88",
		X"04",X"C8",X"04",X"ED",X"4D",X"AE",X"02",X"AF",X"42",X"CC",X"00",X"00",X"ED",X"46",X"86",X"10",
		X"A7",X"48",X"20",X"85",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",
		X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",
		X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",
		X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",
		X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",
		X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",
		X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",
		X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",
		X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",
		X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",
		X"BF",X"CA",X"02",X"FF",X"CA",X"00",X"3A",X"9B",X"A8",X"A7",X"A4",X"BF",X"CA",X"02",X"FF",X"CA",
		X"00",X"1C",X"EF",X"35",X"A0",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",
		X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",
		X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",
		X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",
		X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",
		X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",X"C4",X"E7",X"84",X"9B",X"A8",X"A7",
		X"C4",X"E7",X"84",X"1C",X"EF",X"39",X"E6",X"A8",X"11",X"C0",X"10",X"50",X"86",X"06",X"3D",X"8E",
		X"F1",X"D5",X"3A",X"34",X"10",X"A6",X"26",X"97",X"A8",X"EC",X"29",X"1A",X"10",X"F7",X"CA",X"05",
		X"E6",X"2F",X"CA",X"10",X"C4",X"F7",X"CE",X"00",X"00",X"FF",X"CA",X"01",X"F7",X"CA",X"03",X"EE",
		X"2D",X"FF",X"CA",X"06",X"CE",X"CA",X"04",X"8E",X"CA",X"00",X"39",X"CE",X"98",X"A9",X"10",X"AC",
		X"C4",X"27",X"08",X"EE",X"C4",X"26",X"F7",X"1A",X"10",X"20",X"FE",X"EC",X"A4",X"ED",X"C4",X"DC",
		X"AD",X"ED",X"A4",X"10",X"9F",X"AD",X"31",X"C4",X"39",X"EC",X"26",X"83",X"00",X"80",X"A1",X"26",
		X"26",X"03",X"E7",X"27",X"39",X"BD",X"F2",X"36",X"96",X"59",X"26",X"0B",X"D6",X"5F",X"E7",X"2A",
		X"E6",X"25",X"54",X"DB",X"5E",X"E7",X"24",X"A6",X"2B",X"48",X"4A",X"97",X"AF",X"EC",X"26",X"83",
		X"00",X"80",X"4D",X"22",X"15",X"CE",X"98",X"AB",X"7E",X"F2",X"6E",X"6A",X"28",X"27",X"AC",X"A6",
		X"2B",X"48",X"4A",X"97",X"AF",X"EC",X"26",X"C3",X"01",X"00",X"ED",X"26",X"97",X"A8",X"44",X"E6",
		X"25",X"26",X"01",X"4F",X"97",X"B2",X"30",X"A8",X"12",X"96",X"A8",X"E6",X"25",X"3D",X"DD",X"B0",
		X"E6",X"24",X"4F",X"93",X"B0",X"DB",X"B2",X"89",X"00",X"26",X"04",X"C1",X"07",X"22",X"16",X"0A",
		X"AF",X"DB",X"A8",X"89",X"00",X"26",X"F8",X"C1",X"07",X"23",X"F4",X"E7",X"29",X"EC",X"2B",X"90",
		X"AF",X"3D",X"3A",X"20",X"02",X"E7",X"29",X"96",X"AF",X"4A",X"D6",X"A8",X"3D",X"EB",X"29",X"89",
		X"00",X"27",X"08",X"0A",X"AF",X"D0",X"A8",X"82",X"00",X"26",X"F8",X"C1",X"8F",X"24",X"F4",X"96",
		X"AF",X"10",X"27",X"FF",X"46",X"A7",X"A8",X"11",X"80",X"10",X"40",X"C6",X"0B",X"3D",X"C3",X"F1",
		X"24",X"34",X"26",X"EE",X"2F",X"EC",X"2D",X"1A",X"10",X"FD",X"CA",X"06",X"A6",X"2A",X"B7",X"CA",
		X"05",X"E6",X"2C",X"A6",X"29",X"10",X"8E",X"CA",X"04",X"39",X"10",X"9E",X"A9",X"27",X"0B",X"BD",
		X"F2",X"36",X"BD",X"F2",X"BB",X"10",X"AE",X"A4",X"26",X"F5",X"10",X"9E",X"AB",X"27",X"08",X"BD",
		X"F2",X"89",X"10",X"AE",X"A4",X"26",X"F8",X"39",X"17",X"21",X"90",X"0D",X"21",X"08",X"22",X"90",
		X"0C",X"22",X"07",X"21",X"41",X"21",X"90",X"0B",X"21",X"41",X"21",X"06",X"21",X"42",X"21",X"90",
		X"0A",X"21",X"42",X"21",X"05",X"21",X"43",X"21",X"90",X"09",X"21",X"43",X"21",X"04",X"21",X"44",
		X"21",X"90",X"08",X"21",X"44",X"21",X"03",X"21",X"45",X"21",X"90",X"08",X"21",X"44",X"21",X"02",
		X"21",X"46",X"21",X"90",X"08",X"21",X"44",X"21",X"01",X"21",X"43",X"21",X"43",X"21",X"90",X"08",
		X"21",X"43",X"21",X"01",X"21",X"43",X"22",X"43",X"21",X"90",X"08",X"21",X"43",X"21",X"01",X"21",
		X"42",X"21",X"01",X"21",X"43",X"21",X"90",X"C4",X"08",X"21",X"43",X"23",X"42",X"21",X"01",X"21",
		X"43",X"21",X"90",X"08",X"21",X"48",X"21",X"01",X"21",X"43",X"21",X"90",X"C2",X"08",X"2A",X"01",
		X"21",X"43",X"21",X"90",X"12",X"21",X"44",X"21",X"90",X"C3",X"A0",X"0B",X"28",X"44",X"21",X"90",
		X"0A",X"21",X"4A",X"23",X"90",X"09",X"21",X"4B",X"21",X"90",X"08",X"21",X"4D",X"21",X"90",X"07",
		X"21",X"44",X"27",X"44",X"21",X"90",X"06",X"21",X"44",X"21",X"07",X"21",X"44",X"21",X"90",X"05",
		X"21",X"44",X"21",X"09",X"21",X"44",X"21",X"90",X"04",X"21",X"44",X"2D",X"44",X"21",X"90",X"03",
		X"21",X"57",X"21",X"90",X"02",X"21",X"59",X"21",X"90",X"01",X"21",X"5B",X"21",X"90",X"3F",X"90",
		X"A0",X"1A",X"FF",X"10",X"CE",X"BF",X"70",X"7F",X"C8",X"0D",X"7F",X"C8",X"0C",X"86",X"3C",X"B7",
		X"C8",X"0D",X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",X"B7",X"C8",X"0F",X"86",
		X"C0",X"B7",X"C8",X"0E",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"F6",X"0B",X"10",X"8E",X"C0",X"00",
		X"EC",X"81",X"ED",X"A1",X"8C",X"F6",X"1B",X"25",X"F7",X"86",X"02",X"10",X"8E",X"F4",X"75",X"8E",
		X"00",X"00",X"7E",X"FD",X"65",X"10",X"8E",X"F4",X"7C",X"7E",X"FF",X"3F",X"86",X"34",X"B7",X"C8",
		X"0D",X"B7",X"C8",X"0F",X"7F",X"C8",X"0E",X"86",X"98",X"1F",X"8B",X"10",X"CE",X"BF",X"70",X"BD",
		X"D0",X"12",X"86",X"01",X"BD",X"5F",X"99",X"10",X"8E",X"D0",X"00",X"86",X"07",X"7E",X"FE",X"7F",
		X"86",X"00",X"A7",X"45",X"96",X"CE",X"26",X"0F",X"86",X"02",X"8E",X"F4",X"B0",X"7E",X"D0",X"66",
		X"B6",X"C8",X"0C",X"85",X"02",X"26",X"03",X"7E",X"D0",X"63",X"BD",X"D0",X"60",X"BD",X"D0",X"99",
		X"86",X"FF",X"97",X"CE",X"97",X"59",X"BD",X"F5",X"F5",X"BD",X"D0",X"12",X"B6",X"C8",X"0C",X"46",
		X"10",X"25",X"06",X"1A",X"1A",X"BF",X"10",X"8E",X"F4",X"DD",X"7E",X"FF",X"0D",X"86",X"39",X"B7",
		X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"10",X"8E",X"F4",X"F0",X"7E",X"FF",X"3F",
		X"86",X"98",X"1F",X"8B",X"BD",X"D0",X"12",X"86",X"04",X"BD",X"5F",X"99",X"C6",X"03",X"8E",X"70",
		X"00",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"16",X"30",X"1F",X"8C",
		X"00",X"00",X"26",X"ED",X"5A",X"26",X"E7",X"10",X"8E",X"F5",X"23",X"8E",X"00",X"00",X"86",X"FF",
		X"7E",X"FD",X"65",X"86",X"01",X"B7",X"C9",X"00",X"86",X"98",X"1F",X"8B",X"BD",X"D0",X"12",X"86",
		X"05",X"BD",X"5F",X"99",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",
		X"8E",X"98",X"00",X"4F",X"A7",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",X"71",X"25",X"F4",
		X"BD",X"F5",X"F5",X"CC",X"A5",X"5A",X"DD",X"85",X"97",X"CE",X"BD",X"D0",X"36",X"BD",X"D0",X"C0",
		X"BD",X"D0",X"99",X"86",X"FF",X"97",X"59",X"BD",X"D0",X"54",X"F5",X"73",X"8D",X"7A",X"1C",X"00",
		X"7E",X"D0",X"96",X"BD",X"FA",X"AF",X"BD",X"FD",X"00",X"1C",X"01",X"86",X"06",X"24",X"28",X"C6",
		X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",X"1A",X"10",X"10",X"CE",X"F5",X"93",X"86",X"03",
		X"7E",X"FE",X"93",X"10",X"CE",X"BF",X"70",X"8D",X"4F",X"86",X"98",X"1F",X"8B",X"1C",X"EF",X"86",
		X"07",X"C1",X"1F",X"22",X"02",X"86",X"08",X"BD",X"D0",X"12",X"BD",X"5F",X"99",X"BD",X"FA",X"AF",
		X"DE",X"15",X"6F",X"49",X"BD",X"FC",X"90",X"BD",X"FC",X"99",X"BD",X"FA",X"DD",X"24",X"F8",X"86",
		X"3F",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"F5",X"CC",X"7E",X"D0",X"66",X"86",X"2C",X"B7",X"C8",
		X"0E",X"BD",X"FA",X"AF",X"BD",X"F9",X"28",X"BD",X"FA",X"AF",X"BD",X"F8",X"88",X"BD",X"FA",X"DD",
		X"24",X"03",X"BD",X"FA",X"AF",X"7E",X"F6",X"77",X"7F",X"C8",X"0E",X"86",X"34",X"B7",X"C8",X"0D",
		X"4C",X"B7",X"C8",X"0F",X"39",X"8E",X"F6",X"0B",X"10",X"8E",X"98",X"00",X"CE",X"C0",X"00",X"EC",
		X"81",X"ED",X"A1",X"ED",X"C1",X"8C",X"F6",X"1B",X"25",X"F5",X"39",X"00",X"07",X"17",X"C7",X"1F",
		X"3F",X"38",X"C0",X"A4",X"FF",X"38",X"17",X"CC",X"81",X"81",X"07",X"86",X"3F",X"1F",X"8A",X"8D",
		X"D4",X"86",X"85",X"BE",X"B9",X"EA",X"30",X"89",X"12",X"34",X"10",X"8E",X"F6",X"31",X"7E",X"FD",
		X"65",X"10",X"8E",X"F6",X"38",X"7E",X"FF",X"3F",X"86",X"98",X"1F",X"8B",X"10",X"CE",X"BF",X"70",
		X"BD",X"FD",X"00",X"24",X"1F",X"86",X"03",X"8D",X"26",X"86",X"08",X"8C",X"CD",X"00",X"23",X"02",
		X"86",X"07",X"C6",X"39",X"F7",X"CB",X"FF",X"BD",X"D0",X"12",X"BD",X"5F",X"99",X"86",X"39",X"B7",
		X"CB",X"FF",X"20",X"F9",X"8D",X"47",X"10",X"8E",X"F6",X"1B",X"86",X"04",X"7E",X"FE",X"7F",X"10",
		X"8E",X"F6",X"76",X"BD",X"FF",X"1D",X"39",X"BD",X"F6",X"FE",X"BD",X"FA",X"AF",X"BD",X"D0",X"12",
		X"86",X"07",X"97",X"00",X"BD",X"FA",X"AF",X"86",X"38",X"97",X"00",X"BD",X"FA",X"AF",X"86",X"C0",
		X"97",X"00",X"BD",X"FA",X"AF",X"8D",X"16",X"BD",X"FA",X"AF",X"7E",X"FA",X"EE",X"9F",X"2B",X"30",
		X"89",X"10",X"00",X"30",X"89",X"FF",X"00",X"8C",X"98",X"00",X"22",X"F7",X"39",X"8E",X"98",X"00",
		X"10",X"8E",X"F6",X"EE",X"CE",X"C0",X"00",X"EC",X"A1",X"ED",X"81",X"ED",X"C1",X"86",X"39",X"B7",
		X"CB",X"FF",X"8C",X"98",X"10",X"25",X"F0",X"CC",X"00",X"00",X"8E",X"00",X"00",X"8D",X"CE",X"ED",
		X"83",X"34",X"02",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"02",X"9C",X"2B",X"26",X"F1",X"30",X"89",
		X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",X"E0",X"39",X"05",X"05",
		X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",X"BD",X"D0",
		X"12",X"4F",X"BD",X"F9",X"1D",X"86",X"FF",X"97",X"01",X"86",X"C0",X"97",X"02",X"86",X"38",X"97",
		X"03",X"86",X"07",X"97",X"04",X"10",X"8E",X"F8",X"10",X"CC",X"01",X"01",X"AE",X"A4",X"ED",X"81",
		X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"F8",X"38",X"26",X"F0",X"86",X"11",X"10",X"8E",
		X"F7",X"F0",X"AE",X"A4",X"9F",X"2B",X"A7",X"84",X"0C",X"2B",X"9E",X"2B",X"AC",X"22",X"26",X"F6",
		X"31",X"24",X"10",X"8C",X"F8",X"10",X"26",X"EA",X"10",X"8E",X"F8",X"38",X"AE",X"A4",X"9F",X"2B",
		X"A6",X"24",X"A7",X"84",X"0C",X"2B",X"9E",X"2B",X"AC",X"22",X"26",X"F6",X"31",X"25",X"10",X"8C",
		X"F8",X"74",X"26",X"E8",X"10",X"8E",X"F8",X"74",X"AE",X"A4",X"A6",X"24",X"A7",X"80",X"AC",X"22",
		X"26",X"FA",X"31",X"25",X"10",X"8C",X"F8",X"88",X"26",X"EE",X"86",X"21",X"B7",X"43",X"7E",X"86",
		X"20",X"B7",X"93",X"7E",X"8E",X"4B",X"0A",X"1A",X"10",X"7F",X"C9",X"00",X"A6",X"84",X"C6",X"01",
		X"F7",X"C9",X"00",X"1C",X"EF",X"84",X"F0",X"8A",X"02",X"A7",X"80",X"8C",X"4B",X"6D",X"26",X"E7",
		X"8E",X"4B",X"90",X"1A",X"10",X"7F",X"C9",X"00",X"A6",X"84",X"C6",X"01",X"F7",X"C9",X"00",X"1C",
		X"EF",X"84",X"F0",X"8A",X"02",X"A7",X"80",X"8C",X"4B",X"F3",X"26",X"E7",X"8E",X"0B",X"18",X"9F",
		X"2B",X"9E",X"2B",X"1A",X"10",X"7F",X"C9",X"00",X"A6",X"84",X"C6",X"01",X"F7",X"C9",X"00",X"1C",
		X"EF",X"84",X"F0",X"8A",X"01",X"A7",X"84",X"D6",X"2C",X"CB",X"22",X"25",X"04",X"D7",X"2C",X"20",
		X"E0",X"C6",X"18",X"D7",X"2C",X"D6",X"2B",X"CB",X"10",X"D7",X"2B",X"C1",X"9B",X"26",X"D2",X"39",
		X"04",X"07",X"94",X"07",X"04",X"29",X"94",X"29",X"04",X"4B",X"94",X"4B",X"04",X"6D",X"94",X"6D",
		X"04",X"8F",X"94",X"8F",X"04",X"B1",X"94",X"B1",X"04",X"D3",X"94",X"D3",X"04",X"F5",X"94",X"F5",
		X"03",X"07",X"03",X"F5",X"13",X"07",X"13",X"F5",X"23",X"07",X"23",X"F5",X"33",X"07",X"33",X"F5",
		X"43",X"07",X"43",X"F5",X"53",X"07",X"53",X"F5",X"63",X"07",X"63",X"F5",X"73",X"07",X"73",X"F5",
		X"83",X"07",X"83",X"F5",X"93",X"07",X"93",X"F5",X"45",X"05",X"52",X"05",X"44",X"45",X"06",X"52",
		X"06",X"44",X"45",X"07",X"52",X"07",X"00",X"45",X"08",X"52",X"08",X"33",X"45",X"09",X"52",X"09",
		X"33",X"45",X"F3",X"52",X"F3",X"33",X"45",X"F4",X"52",X"F4",X"33",X"45",X"F5",X"52",X"F5",X"00",
		X"45",X"F6",X"52",X"F6",X"44",X"45",X"F7",X"52",X"F7",X"44",X"04",X"7E",X"43",X"7E",X"22",X"54",
		X"7E",X"93",X"7E",X"22",X"02",X"6F",X"02",X"8E",X"04",X"03",X"6F",X"03",X"8E",X"30",X"93",X"6F",
		X"93",X"8E",X"00",X"94",X"6F",X"94",X"8E",X"34",X"35",X"06",X"DE",X"15",X"ED",X"4D",X"BD",X"D0",
		X"12",X"86",X"1E",X"BD",X"5F",X"99",X"86",X"80",X"A7",X"47",X"86",X"01",X"8E",X"F8",X"A2",X"7E",
		X"D0",X"66",X"BD",X"FA",X"DD",X"25",X"34",X"6A",X"47",X"26",X"EF",X"B6",X"F9",X"05",X"8D",X"6D",
		X"8D",X"2E",X"8E",X"F9",X"05",X"A6",X"80",X"DE",X"15",X"AF",X"49",X"8D",X"60",X"86",X"80",X"A7",
		X"47",X"86",X"01",X"8E",X"F8",X"C9",X"7E",X"D0",X"66",X"BD",X"FA",X"DD",X"25",X"0D",X"6A",X"47",
		X"26",X"EF",X"AE",X"49",X"8C",X"F9",X"0D",X"25",X"DC",X"20",X"D7",X"DE",X"15",X"6E",X"D8",X"0D",
		X"8E",X"00",X"00",X"10",X"8E",X"F9",X"0D",X"BD",X"F6",X"9D",X"A6",X"A0",X"1F",X"89",X"ED",X"83",
		X"9C",X"2B",X"26",X"FA",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"10",X"8C",
		X"F9",X"1D",X"26",X"E3",X"39",X"02",X"03",X"04",X"10",X"18",X"20",X"40",X"80",X"00",X"FF",X"11",
		X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",X"8E",X"98",X"00",
		X"A7",X"80",X"8C",X"98",X"10",X"25",X"F9",X"39",X"35",X"06",X"DE",X"15",X"ED",X"4D",X"86",X"0A",
		X"A7",X"4B",X"BD",X"D0",X"12",X"86",X"0C",X"BD",X"5F",X"99",X"CE",X"B3",X"EA",X"6F",X"C0",X"11",
		X"83",X"B3",X"F4",X"23",X"F8",X"CE",X"F9",X"E1",X"8D",X"26",X"86",X"34",X"B7",X"C8",X"07",X"8D",
		X"1F",X"86",X"3C",X"B7",X"C8",X"07",X"8D",X"28",X"BD",X"FA",X"DD",X"24",X"06",X"DE",X"15",X"6A",
		X"4B",X"27",X"08",X"86",X"01",X"8E",X"F9",X"45",X"7E",X"D0",X"66",X"DE",X"15",X"6E",X"D8",X"0D",
		X"AE",X"C1",X"27",X"0B",X"10",X"AE",X"C1",X"A6",X"84",X"A8",X"A4",X"A7",X"21",X"20",X"F1",X"39",
		X"CE",X"F9",X"F9",X"10",X"8E",X"B3",X"EA",X"C6",X"01",X"E5",X"21",X"27",X"02",X"8D",X"19",X"33",
		X"43",X"58",X"24",X"F5",X"31",X"22",X"10",X"8C",X"B3",X"F3",X"22",X"0B",X"B6",X"C8",X"06",X"2B",
		X"E6",X"10",X"8C",X"B3",X"EF",X"23",X"E0",X"39",X"34",X"14",X"86",X"3F",X"B7",X"C8",X"0E",X"E8",
		X"A4",X"E7",X"A4",X"E6",X"E4",X"E5",X"A4",X"26",X"10",X"E6",X"42",X"27",X"22",X"86",X"40",X"1F",
		X"01",X"CC",X"30",X"06",X"BD",X"D0",X"1B",X"35",X"94",X"E6",X"42",X"27",X"12",X"86",X"40",X"1F",
		X"01",X"C6",X"BB",X"D7",X"CF",X"EC",X"C4",X"BD",X"5F",X"96",X"86",X"37",X"B7",X"C8",X"0E",X"35",
		X"94",X"C8",X"0C",X"B3",X"EA",X"C8",X"04",X"B3",X"EC",X"C8",X"06",X"B3",X"EE",X"00",X"00",X"C8",
		X"04",X"B3",X"F0",X"C8",X"06",X"B3",X"F2",X"00",X"00",X"0D",X"00",X"2C",X"0E",X"00",X"33",X"0F",
		X"00",X"3A",X"10",X"00",X"41",X"11",X"00",X"48",X"12",X"00",X"4F",X"13",X"00",X"56",X"00",X"00",
		X"00",X"14",X"01",X"5D",X"15",X"01",X"64",X"16",X"01",X"6B",X"17",X"01",X"72",X"18",X"00",X"79",
		X"19",X"00",X"80",X"1A",X"01",X"87",X"1B",X"01",X"8E",X"1C",X"01",X"95",X"1D",X"01",X"9C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"14",X"02",X"A3",X"15",X"02",X"AA",X"16",X"02",X"B1",X"17",X"02",X"B8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1A",X"02",X"BF",X"1B",X"02",X"C6",X"1C",X"02",X"CD",X"1D",X"02",X"D4",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CE",X"F5",X"40",X"20",X"03",X"CE",X"F5",X"17",X"10",X"CE",X"BF",X"70",X"10",X"8E",X"FA",
		X"86",X"86",X"01",X"7E",X"FE",X"7F",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"10",X"8E",X"FA",
		X"96",X"86",X"01",X"7E",X"FE",X"7F",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F0",X"10",X"8E",X"FA",
		X"A6",X"86",X"01",X"7E",X"FE",X"7F",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"6E",X"C4",X"35",
		X"06",X"DE",X"15",X"ED",X"4D",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"08",X"86",X"01",X"8E",X"FA",
		X"B5",X"7E",X"D0",X"66",X"0F",X"00",X"BD",X"D0",X"12",X"20",X"07",X"B6",X"C8",X"0C",X"85",X"02",
		X"27",X"08",X"86",X"02",X"8E",X"FA",X"CB",X"7E",X"D0",X"66",X"6E",X"D8",X"0D",X"34",X"02",X"B6",
		X"C8",X"0C",X"85",X"02",X"27",X"04",X"1A",X"01",X"35",X"82",X"1C",X"FE",X"35",X"82",X"86",X"FF",
		X"97",X"59",X"BD",X"F5",X"F5",X"8D",X"E6",X"24",X"02",X"8D",X"B4",X"86",X"1F",X"BD",X"5F",X"99",
		X"CE",X"CD",X"02",X"86",X"20",X"34",X"02",X"BD",X"5F",X"99",X"1E",X"31",X"BD",X"D0",X"A5",X"34",
		X"04",X"BD",X"D0",X"A8",X"1F",X"02",X"35",X"04",X"1E",X"31",X"8D",X"71",X"35",X"02",X"4C",X"11",
		X"83",X"CD",X"32",X"25",X"E0",X"86",X"6A",X"BD",X"5F",X"99",X"34",X"10",X"8E",X"CD",X"20",X"10",
		X"8E",X"CD",X"2C",X"BD",X"FB",X"BF",X"35",X"10",X"F6",X"B4",X"18",X"10",X"BE",X"B4",X"19",X"8D",
		X"4C",X"B6",X"B4",X"1B",X"84",X"0F",X"B7",X"B4",X"1C",X"B6",X"B4",X"1B",X"85",X"10",X"27",X"08",
		X"84",X"EF",X"44",X"8B",X"05",X"19",X"20",X"01",X"44",X"BB",X"B4",X"1C",X"19",X"1F",X"89",X"86",
		X"6B",X"BD",X"5F",X"99",X"86",X"6C",X"BD",X"5F",X"99",X"34",X"10",X"8E",X"CD",X"26",X"10",X"8E",
		X"CD",X"2C",X"8D",X"4B",X"35",X"10",X"F6",X"B4",X"18",X"10",X"BE",X"B4",X"19",X"8D",X"0E",X"F6",
		X"B4",X"1B",X"86",X"6D",X"BD",X"5F",X"99",X"BD",X"FA",X"AF",X"7E",X"6F",X"00",X"5D",X"27",X"0C",
		X"86",X"29",X"BD",X"5F",X"99",X"86",X"2A",X"BD",X"5F",X"99",X"20",X"05",X"86",X"2B",X"BD",X"5F",
		X"99",X"39",X"34",X"04",X"BD",X"D0",X"A2",X"1F",X"89",X"84",X"0F",X"81",X"09",X"23",X"02",X"86",
		X"09",X"C4",X"F0",X"C1",X"90",X"23",X"02",X"C6",X"90",X"34",X"04",X"AA",X"E0",X"35",X"84",X"34",
		X"76",X"CC",X"00",X"00",X"FD",X"B4",X"18",X"FD",X"B4",X"1A",X"8D",X"D6",X"B7",X"B4",X"06",X"8D",
		X"D1",X"B7",X"B4",X"07",X"8D",X"CC",X"B7",X"B4",X"08",X"CC",X"00",X"00",X"B7",X"B4",X"09",X"FD",
		X"B4",X"0A",X"B7",X"B4",X"15",X"FD",X"B4",X"16",X"1F",X"21",X"BD",X"FB",X"A2",X"B7",X"B4",X"12",
		X"BD",X"FB",X"A2",X"B7",X"B4",X"13",X"BD",X"FB",X"A2",X"B7",X"B4",X"14",X"26",X"05",X"FC",X"B4",
		X"12",X"27",X"3A",X"CE",X"B4",X"1A",X"7D",X"B4",X"12",X"26",X"12",X"33",X"5F",X"C6",X"05",X"8E",
		X"B4",X"12",X"A6",X"01",X"A7",X"80",X"5A",X"26",X"F9",X"6F",X"84",X"20",X"E9",X"8E",X"B4",X"06",
		X"8D",X"1D",X"24",X"FC",X"10",X"8E",X"B4",X"17",X"C6",X"05",X"A6",X"3F",X"A7",X"A4",X"31",X"3F",
		X"5A",X"26",X"F7",X"6F",X"A4",X"33",X"41",X"11",X"83",X"B4",X"1B",X"23",X"E3",X"35",X"F6",X"10",
		X"8E",X"B4",X"12",X"86",X"00",X"E6",X"86",X"E0",X"A0",X"22",X"07",X"25",X"40",X"4C",X"81",X"06",
		X"25",X"F3",X"C6",X"06",X"10",X"8E",X"B4",X"0C",X"86",X"99",X"A0",X"26",X"A7",X"A0",X"5A",X"26",
		X"F7",X"C6",X"06",X"1C",X"FE",X"86",X"01",X"A9",X"A2",X"19",X"A7",X"A4",X"86",X"00",X"5A",X"26",
		X"F6",X"C6",X"05",X"10",X"8E",X"B4",X"12",X"1C",X"FE",X"A6",X"A2",X"A9",X"85",X"19",X"A7",X"85",
		X"5A",X"2A",X"F6",X"A6",X"C4",X"8B",X"01",X"19",X"A7",X"C4",X"1C",X"FE",X"39",X"1A",X"01",X"39",
		X"BD",X"D0",X"12",X"CC",X"FE",X"01",X"ED",X"47",X"39",X"35",X"06",X"ED",X"4D",X"86",X"3F",X"B7",
		X"C8",X"0E",X"86",X"01",X"8E",X"FC",X"AA",X"7E",X"D0",X"66",X"86",X"2C",X"B7",X"C8",X"0E",X"86",
		X"01",X"8E",X"FC",X"B7",X"7E",X"D0",X"66",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"FC",
		X"C4",X"7E",X"D0",X"66",X"EC",X"47",X"84",X"3F",X"B7",X"C8",X"0E",X"86",X"09",X"BD",X"5F",X"99",
		X"86",X"40",X"A7",X"4B",X"86",X"01",X"8E",X"FC",X"DC",X"7E",X"D0",X"66",X"BD",X"FA",X"DD",X"25",
		X"04",X"6A",X"4B",X"26",X"EF",X"A6",X"49",X"26",X"06",X"B6",X"C8",X"0C",X"46",X"24",X"0E",X"EC",
		X"47",X"1A",X"01",X"49",X"5C",X"C1",X"07",X"25",X"02",X"8D",X"98",X"ED",X"47",X"6E",X"D8",X"0D",
		X"8E",X"CC",X"00",X"10",X"8E",X"B3",X"EA",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",
		X"C6",X"06",X"1A",X"3F",X"DE",X"85",X"10",X"9E",X"84",X"8E",X"CC",X"00",X"BD",X"D0",X"39",X"A7",
		X"80",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"F1",X"10",X"9F",X"84",X"DF",X"85",
		X"8E",X"CC",X"00",X"BD",X"D0",X"39",X"A8",X"80",X"84",X"0F",X"26",X"24",X"86",X"39",X"B7",X"CB",
		X"FF",X"8C",X"D0",X"00",X"26",X"ED",X"5A",X"26",X"CB",X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"B3",
		X"EA",X"10",X"8E",X"CC",X"00",X"A6",X"C0",X"A7",X"A0",X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",
		X"8D",X"EC",X"1A",X"01",X"39",X"1A",X"3F",X"7F",X"C9",X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",
		X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",
		X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"ED",X"81",X"1E",X"10",X"5D",X"26",X"15",X"C6",
		X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",
		X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",X"C8",X"1F",X"30",X"8E",X"00",X"00",
		X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",
		X"56",X"20",X"02",X"44",X"56",X"10",X"A3",X"81",X"26",X"43",X"1E",X"10",X"5D",X"26",X"15",X"C6",
		X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",
		X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",X"C5",X"1F",X"03",X"1F",X"B8",X"81",
		X"FF",X"26",X"05",X"1F",X"30",X"7E",X"FD",X"70",X"4A",X"1F",X"8B",X"81",X"80",X"27",X"07",X"4D",
		X"1F",X"30",X"10",X"26",X"FF",X"6A",X"C6",X"01",X"F7",X"C9",X"00",X"6E",X"A4",X"30",X"1E",X"A8",
		X"84",X"E8",X"01",X"4D",X"26",X"07",X"5D",X"26",X"04",X"30",X"02",X"20",X"AD",X"CE",X"00",X"30",
		X"1E",X"10",X"5F",X"1E",X"10",X"8C",X"00",X"00",X"27",X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",
		X"10",X"11",X"83",X"00",X"30",X"23",X"EE",X"CE",X"00",X"10",X"20",X"E9",X"33",X"41",X"47",X"25",
		X"05",X"57",X"25",X"02",X"20",X"F6",X"1F",X"30",X"86",X"01",X"B7",X"C9",X"00",X"10",X"CE",X"FE",
		X"53",X"20",X"40",X"86",X"98",X"1F",X"8B",X"1F",X"A8",X"43",X"85",X"C0",X"27",X"04",X"86",X"0B",
		X"20",X"02",X"86",X"02",X"10",X"CE",X"BF",X"70",X"BD",X"D0",X"12",X"BD",X"5F",X"99",X"1F",X"A8",
		X"85",X"40",X"26",X"03",X"7E",X"FA",X"71",X"10",X"8E",X"D0",X"00",X"20",X"00",X"86",X"20",X"8E",
		X"58",X"00",X"30",X"1F",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",
		X"EE",X"6E",X"A4",X"1F",X"03",X"86",X"02",X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"FE",X"A1",X"20",
		X"7C",X"86",X"02",X"10",X"8E",X"FE",X"A9",X"20",X"D6",X"10",X"8E",X"FE",X"AF",X"20",X"5E",X"86",
		X"01",X"10",X"8E",X"FE",X"B7",X"20",X"C8",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",
		X"8E",X"FE",X"C5",X"20",X"58",X"86",X"02",X"10",X"8E",X"FE",X"CD",X"20",X"B2",X"10",X"8E",X"FE",
		X"D3",X"20",X"3A",X"86",X"01",X"10",X"8E",X"FE",X"DB",X"20",X"A4",X"1F",X"30",X"1F",X"98",X"10",
		X"8E",X"FE",X"E5",X"20",X"38",X"86",X"02",X"10",X"8E",X"FE",X"ED",X"20",X"92",X"10",X"8E",X"FE",
		X"F3",X"20",X"1A",X"86",X"05",X"10",X"8E",X"FE",X"FC",X"7E",X"FE",X"7F",X"1F",X"B8",X"4A",X"1F",
		X"8B",X"26",X"96",X"10",X"8E",X"FF",X"09",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",X"B7",
		X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",X"46",
		X"46",X"46",X"84",X"C0",X"B7",X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",X"B7",
		X"C8",X"0F",X"86",X"34",X"C5",X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",X"1A",
		X"3F",X"8E",X"FF",X"B5",X"8C",X"FF",X"D5",X"27",X"6A",X"A6",X"01",X"27",X"18",X"A6",X"84",X"5F",
		X"1F",X"03",X"86",X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",X"1E",X"03",X"26",
		X"F3",X"E1",X"01",X"26",X"04",X"30",X"02",X"20",X"DB",X"A6",X"84",X"44",X"44",X"44",X"44",X"81",
		X"0D",X"25",X"02",X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",X"CE",X"FF",X"83",
		X"7E",X"FE",X"93",X"86",X"98",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"BF",X"70",
		X"BD",X"D0",X"12",X"1F",X"A8",X"43",X"85",X"C0",X"27",X"04",X"86",X"0A",X"20",X"02",X"86",X"03",
		X"BD",X"5F",X"99",X"1F",X"A9",X"C5",X"40",X"26",X"03",X"7E",X"FA",X"76",X"10",X"8E",X"D0",X"00",
		X"7E",X"FE",X"7D",X"6E",X"A4",X"00",X"73",X"10",X"EA",X"20",X"1A",X"30",X"6C",X"40",X"B3",X"50",
		X"23",X"60",X"A3",X"70",X"3B",X"80",X"63",X"90",X"00",X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",
		X"5C",X"E0",X"82",X"F0",X"01",X"00",X"3D",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"2E",X"49",X"4E",X"43",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"DC",X"56",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"7E",X"01",X"6D",X"7E",X"02",X"B2",X"7E",X"00",X"9E",X"7E",X"03",X"51",X"04",X"85",X"05",X"2F",
		X"07",X"FF",X"0B",X"3B",X"0C",X"F9",X"01",X"CC",X"03",X"CF",X"04",X"37",X"D0",X"01",X"10",X"06",
		X"00",X"D0",X"03",X"04",X"17",X"00",X"E0",X"01",X"20",X"0D",X"00",X"E0",X"01",X"18",X"1A",X"00",
		X"96",X"59",X"85",X"7F",X"27",X"08",X"86",X"08",X"8E",X"00",X"30",X"7E",X"D0",X"66",X"AE",X"47",
		X"10",X"AE",X"4D",X"A6",X"4B",X"31",X"A6",X"E6",X"A4",X"2A",X"04",X"6F",X"4B",X"20",X"F1",X"8B",
		X"03",X"A7",X"4B",X"4F",X"C3",X"0C",X"F9",X"ED",X"02",X"A6",X"21",X"5F",X"47",X"56",X"E3",X"0A",
		X"34",X"06",X"E6",X"22",X"EB",X"0C",X"8D",X"36",X"27",X"04",X"32",X"62",X"20",X"22",X"E7",X"0C",
		X"35",X"06",X"ED",X"0A",X"E6",X"0C",X"EE",X"02",X"8E",X"98",X"23",X"34",X"46",X"BD",X"D0",X"27",
		X"35",X"46",X"8E",X"98",X"1F",X"BD",X"D0",X"27",X"DE",X"15",X"AE",X"47",X"6A",X"4C",X"26",X"02",
		X"8D",X"74",X"BD",X"D0",X"8D",X"8E",X"00",X"3E",X"B6",X"BE",X"61",X"7E",X"D0",X"66",X"34",X"06",
		X"81",X"07",X"25",X"10",X"C1",X"18",X"25",X"0C",X"E3",X"98",X"02",X"81",X"8F",X"22",X"05",X"C1",
		X"EA",X"22",X"01",X"4F",X"35",X"86",X"96",X"48",X"26",X"49",X"96",X"88",X"5F",X"0D",X"84",X"2B",
		X"01",X"48",X"E3",X"0A",X"34",X"06",X"D6",X"89",X"96",X"86",X"81",X"C0",X"24",X"01",X"58",X"EB",
		X"0C",X"A6",X"E4",X"8D",X"C9",X"27",X"04",X"32",X"62",X"20",X"21",X"E7",X"0C",X"35",X"06",X"ED",
		X"0A",X"E6",X"0C",X"EE",X"02",X"34",X"10",X"8E",X"98",X"23",X"34",X"46",X"BD",X"D0",X"27",X"35",
		X"46",X"8E",X"98",X"1F",X"BD",X"D0",X"27",X"35",X"10",X"BD",X"D0",X"8D",X"CC",X"00",X"1C",X"BD",
		X"D0",X"4B",X"39",X"7E",X"D0",X"18",X"96",X"86",X"84",X"1F",X"4C",X"A7",X"4C",X"10",X"AE",X"D8",
		X"09",X"26",X"04",X"10",X"8E",X"98",X"5A",X"EC",X"4D",X"10",X"83",X"01",X"CC",X"27",X"26",X"10",
		X"83",X"01",X"D9",X"27",X"20",X"96",X"84",X"84",X"1F",X"8B",X"F0",X"AB",X"24",X"81",X"8F",X"23",
		X"06",X"81",X"CF",X"23",X"02",X"86",X"07",X"A1",X"04",X"23",X"05",X"CC",X"01",X"D9",X"20",X"1F",
		X"CC",X"01",X"CC",X"20",X"1A",X"96",X"85",X"84",X"1F",X"8B",X"F0",X"AB",X"25",X"81",X"06",X"24",
		X"02",X"86",X"EA",X"A1",X"05",X"23",X"05",X"CC",X"01",X"E6",X"20",X"03",X"CC",X"01",X"F3",X"ED",
		X"4D",X"4F",X"A7",X"4B",X"E6",X"D8",X"0D",X"C3",X"0C",X"F9",X"ED",X"02",X"39",X"B6",X"BE",X"6D",
		X"34",X"02",X"27",X"06",X"8D",X"06",X"6A",X"E4",X"26",X"FA",X"35",X"82",X"BD",X"D0",X"54",X"00",
		X"30",X"33",X"84",X"BD",X"D0",X"7B",X"CC",X"0C",X"F9",X"ED",X"02",X"ED",X"88",X"14",X"EF",X"06",
		X"AF",X"47",X"CC",X"00",X"B6",X"ED",X"08",X"BD",X"38",X"8E",X"BD",X"26",X"C3",X"D1",X"2B",X"23",
		X"0C",X"D1",X"2C",X"24",X"08",X"91",X"2D",X"23",X"04",X"91",X"2E",X"23",X"ED",X"ED",X"04",X"A7",
		X"0A",X"E7",X"0C",X"96",X"84",X"81",X"C0",X"23",X"05",X"CC",X"B3",X"A2",X"20",X"02",X"8D",X"77",
		X"ED",X"49",X"BD",X"01",X"06",X"BD",X"38",X"8B",X"6F",X"88",X"13",X"39",X"00",X"FD",X"00",X"04",
		X"FC",X"00",X"00",X"FD",X"00",X"08",X"FC",X"00",X"FF",X"0C",X"03",X"00",X"10",X"04",X"00",X"0C",
		X"03",X"00",X"14",X"04",X"00",X"FF",X"18",X"00",X"02",X"1C",X"00",X"02",X"18",X"00",X"02",X"20",
		X"00",X"02",X"FF",X"18",X"00",X"FE",X"1C",X"00",X"FE",X"18",X"00",X"FE",X"20",X"00",X"FE",X"FF",
		X"8E",X"B3",X"54",X"9F",X"49",X"6F",X"80",X"8C",X"B3",X"A4",X"26",X"F9",X"39",X"34",X"16",X"8E",
		X"B3",X"54",X"EC",X"81",X"26",X"FC",X"EC",X"62",X"ED",X"1E",X"35",X"96",X"34",X"16",X"8E",X"B3",
		X"54",X"EC",X"62",X"10",X"A3",X"81",X"27",X"09",X"8C",X"B3",X"A4",X"26",X"F6",X"1A",X"10",X"20",
		X"FE",X"4F",X"5F",X"ED",X"1E",X"35",X"96",X"34",X"10",X"9E",X"49",X"8C",X"B3",X"A4",X"25",X"09",
		X"8E",X"B3",X"54",X"20",X"04",X"9C",X"49",X"27",X"14",X"EC",X"81",X"26",X"0A",X"8C",X"B3",X"A4",
		X"25",X"F3",X"8E",X"B3",X"54",X"20",X"EE",X"9F",X"49",X"30",X"1E",X"1F",X"10",X"35",X"90",X"AE",
		X"47",X"10",X"AE",X"4D",X"A6",X"4B",X"31",X"A6",X"E6",X"A4",X"2A",X"04",X"6F",X"4B",X"20",X"F1",
		X"8B",X"03",X"A7",X"4B",X"4F",X"E3",X"49",X"ED",X"02",X"A6",X"21",X"5F",X"47",X"56",X"E3",X"0A",
		X"34",X"06",X"E6",X"22",X"EB",X"0C",X"34",X"40",X"CE",X"98",X"23",X"BD",X"26",X"C6",X"35",X"40",
		X"26",X"05",X"BD",X"00",X"06",X"27",X"04",X"32",X"62",X"20",X"0A",X"E7",X"0C",X"35",X"06",X"ED",
		X"0A",X"6A",X"4C",X"26",X"02",X"8D",X"6B",X"BD",X"D0",X"8D",X"86",X"08",X"8E",X"02",X"5F",X"7E",
		X"D0",X"66",X"BD",X"02",X"00",X"8E",X"0B",X"3B",X"CE",X"03",X"30",X"B6",X"BE",X"6C",X"8D",X"14",
		X"8E",X"05",X"2F",X"CE",X"03",X"35",X"B6",X"BE",X"6A",X"8D",X"09",X"8E",X"07",X"FF",X"CE",X"03",
		X"3A",X"B6",X"BE",X"6B",X"34",X"52",X"4D",X"27",X"37",X"BD",X"D0",X"54",X"02",X"5F",X"33",X"84",
		X"BD",X"D0",X"87",X"EC",X"61",X"ED",X"02",X"ED",X"88",X"14",X"ED",X"49",X"EF",X"06",X"AF",X"47",
		X"EC",X"63",X"ED",X"08",X"BD",X"26",X"C3",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"96",X"84",X"84",
		X"07",X"4C",X"A7",X"44",X"8D",X"0C",X"BD",X"D0",X"18",X"BD",X"02",X"0D",X"6A",X"E4",X"26",X"C9",
		X"35",X"D2",X"96",X"86",X"84",X"7F",X"4C",X"A7",X"4C",X"96",X"84",X"84",X"07",X"C6",X"0D",X"3D",
		X"C3",X"03",X"CF",X"ED",X"4D",X"4F",X"A7",X"4B",X"E6",X"D8",X"0D",X"E3",X"49",X"ED",X"02",X"39",
		X"7A",X"BE",X"6C",X"20",X"08",X"7A",X"BE",X"6A",X"20",X"03",X"7A",X"BE",X"6B",X"BD",X"02",X"1C",
		X"BD",X"D0",X"8A",X"BD",X"D0",X"15",X"EC",X"04",X"AE",X"06",X"BD",X"D0",X"5D",X"0D",X"95",X"26",
		X"51",X"BD",X"D0",X"6C",X"03",X"A3",X"04",X"7D",X"03",X"90",X"81",X"89",X"25",X"02",X"86",X"89",
		X"ED",X"04",X"0D",X"95",X"26",X"2D",X"0D",X"48",X"27",X"29",X"86",X"3C",X"A7",X"49",X"0C",X"8D",
		X"96",X"8D",X"81",X"05",X"23",X"02",X"86",X"05",X"48",X"48",X"CE",X"04",X"81",X"33",X"C6",X"EF",
		X"02",X"CE",X"03",X"C3",X"44",X"EC",X"C6",X"BD",X"D0",X"0C",X"CC",X"00",X"26",X"BD",X"D0",X"4B",
		X"4F",X"35",X"86",X"86",X"5A",X"A7",X"49",X"CC",X"04",X"37",X"ED",X"02",X"CC",X"00",X"2B",X"BD",
		X"D0",X"4B",X"39",X"AE",X"47",X"EC",X"04",X"10",X"AE",X"02",X"BD",X"D0",X"21",X"6A",X"49",X"27",
		X"08",X"86",X"01",X"8E",X"03",X"A3",X"7E",X"D0",X"66",X"BD",X"D0",X"1E",X"DC",X"1B",X"ED",X"84",
		X"9F",X"1B",X"7E",X"D0",X"63",X"02",X"10",X"02",X"20",X"02",X"30",X"02",X"40",X"02",X"50",X"00",
		X"FE",X"00",X"04",X"FF",X"00",X"00",X"FE",X"00",X"08",X"FF",X"00",X"FF",X"0C",X"02",X"00",X"10",
		X"01",X"00",X"0C",X"02",X"00",X"14",X"01",X"00",X"FF",X"18",X"00",X"01",X"1C",X"00",X"01",X"18",
		X"00",X"01",X"20",X"00",X"01",X"FF",X"24",X"00",X"FF",X"28",X"00",X"FF",X"24",X"00",X"FF",X"2C",
		X"00",X"FF",X"FF",X"00",X"FE",X"FF",X"08",X"FF",X"FF",X"00",X"FE",X"FF",X"08",X"FF",X"FF",X"FF",
		X"0C",X"02",X"FF",X"10",X"01",X"FF",X"0C",X"02",X"FF",X"14",X"01",X"FF",X"FF",X"0C",X"02",X"01",
		X"10",X"01",X"01",X"0C",X"02",X"01",X"14",X"01",X"01",X"FF",X"00",X"FE",X"01",X"04",X"FF",X"01",
		X"00",X"FE",X"01",X"08",X"FF",X"01",X"FF",X"06",X"0B",X"04",X"3B",X"00",X"00",X"AA",X"A0",X"00",
		X"00",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"0A",X"0F",X"FA",X"FF",X"0A",X"00",X"AA",X"0A",X"A0",
		X"AA",X"0A",X"A0",X"00",X"A0",X"AA",X"A0",X"A0",X"00",X"00",X"0A",X"0A",X"0A",X"00",X"00",X"00",
		X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"0A",X"A0",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"02",X"02",X"04",
		X"81",X"00",X"00",X"00",X"00",X"06",X"05",X"04",X"99",X"06",X"05",X"04",X"B7",X"06",X"05",X"04",
		X"D5",X"06",X"05",X"04",X"F3",X"06",X"05",X"05",X"11",X"0F",X"F0",X"FF",X"FF",X"FF",X"F0",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"0F",X"FF",X"FF",X"FF",X"FF",X"F0",X"0F",X"FF",X"BB",X"BB",X"BB",X"B0",X"00",X"0F",X"B0",
		X"B0",X"B0",X"B0",X"0F",X"FF",X"B0",X"B0",X"B0",X"B0",X"0F",X"00",X"B0",X"B0",X"B0",X"B0",X"0F",
		X"FF",X"BB",X"BB",X"BB",X"B0",X"0F",X"FF",X"EE",X"EE",X"EE",X"E0",X"00",X"0F",X"E0",X"E0",X"E0",
		X"E0",X"0F",X"FF",X"E0",X"E0",X"E0",X"E0",X"00",X"0F",X"E0",X"E0",X"E0",X"E0",X"0F",X"FF",X"EE",
		X"EE",X"EE",X"E0",X"0F",X"0F",X"BB",X"BB",X"BB",X"B0",X"0F",X"0F",X"B0",X"B0",X"B0",X"B0",X"0F",
		X"FF",X"B0",X"B0",X"B0",X"B0",X"00",X"0F",X"B0",X"B0",X"B0",X"B0",X"00",X"0F",X"BB",X"BB",X"BB",
		X"B0",X"0A",X"AA",X"EE",X"EE",X"EE",X"E0",X"0A",X"00",X"E0",X"E0",X"E0",X"E0",X"0A",X"AA",X"E0",
		X"E0",X"E0",X"E0",X"00",X"0A",X"E0",X"E0",X"E0",X"E0",X"0A",X"AA",X"EE",X"EE",X"EE",X"E0",X"04",
		X"0E",X"05",X"5F",X"04",X"0E",X"05",X"97",X"04",X"0E",X"05",X"CF",X"04",X"0E",X"06",X"07",X"04",
		X"0E",X"06",X"3F",X"04",X"0E",X"06",X"77",X"04",X"0E",X"06",X"AF",X"04",X"0E",X"06",X"E7",X"04",
		X"0E",X"07",X"1F",X"04",X"0E",X"07",X"57",X"04",X"0E",X"07",X"8F",X"04",X"0E",X"07",X"C7",X"00",
		X"55",X"00",X"00",X"00",X"25",X"50",X"00",X"00",X"62",X"50",X"00",X"00",X"22",X"55",X"00",X"00",
		X"03",X"30",X"00",X"00",X"34",X"30",X"00",X"00",X"04",X"30",X"00",X"00",X"39",X"30",X"00",X"03",
		X"33",X"33",X"00",X"00",X"69",X"60",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"25",X"50",X"00",X"00",
		X"62",X"50",X"00",X"00",X"22",X"55",X"00",X"00",X"03",X"30",X"00",X"00",X"33",X"34",X"00",X"00",
		X"03",X"34",X"00",X"09",X"33",X"39",X"00",X"63",X"33",X"33",X"00",X"66",X"90",X"90",X"00",X"09",
		X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"33",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"25",X"50",X"00",X"00",X"62",X"50",X"00",X"00",X"22",X"55",X"00",X"00",
		X"03",X"30",X"00",X"00",X"43",X"34",X"00",X"04",X"43",X"34",X"00",X"09",X"33",X"39",X"00",X"03",
		X"33",X"33",X"60",X"00",X"90",X"96",X"60",X"09",X"00",X"90",X"00",X"09",X"00",X"90",X"00",X"33",
		X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"55",X"20",X"00",X"00",
		X"52",X"60",X"00",X"05",X"52",X"20",X"00",X"00",X"33",X"00",X"00",X"00",X"34",X"30",X"00",X"00",
		X"34",X"00",X"00",X"00",X"39",X"30",X"00",X"03",X"66",X"63",X"00",X"00",X"66",X"60",X"00",X"00",
		X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"50",X"00",X"00",X"55",X"20",X"00",X"00",X"52",X"60",X"00",X"05",X"52",X"20",X"00",X"00",
		X"33",X"00",X"00",X"04",X"33",X"30",X"00",X"04",X"33",X"00",X"00",X"09",X"33",X"39",X"00",X"66",
		X"63",X"33",X"00",X"66",X"60",X"90",X"00",X"00",X"90",X"09",X"00",X"00",X"90",X"09",X"00",X"00",
		X"33",X"03",X"30",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"55",X"20",X"00",X"00",
		X"52",X"60",X"00",X"05",X"52",X"20",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"40",X"00",X"00",
		X"33",X"44",X"00",X"09",X"33",X"39",X"00",X"03",X"33",X"66",X"60",X"00",X"90",X"66",X"60",X"00",
		X"90",X"09",X"00",X"00",X"90",X"09",X"00",X"00",X"33",X"03",X"30",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"00",X"05",X"22",X"25",X"00",X"05",X"62",X"65",X"00",X"55",X"22",X"25",X"50",X"33",
		X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"40",X"03",X"00",X"40",X"90",X"33",X"30",X"90",X"63",
		X"33",X"33",X"00",X"60",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"03",
		X"30",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"05",X"22",X"25",X"00",X"05",
		X"62",X"65",X"00",X"55",X"22",X"25",X"50",X"33",X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"90",
		X"03",X"00",X"40",X"60",X"33",X"30",X"90",X"63",X"33",X"33",X"00",X"00",X"90",X"90",X"00",X"00",
		X"90",X"90",X"00",X"00",X"90",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"55",X"50",X"00",X"05",X"22",X"25",X"00",X"05",X"62",X"65",X"00",X"55",X"22",X"25",X"50",X"33",
		X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"40",X"03",X"00",X"90",X"90",X"33",X"30",X"00",X"63",
		X"33",X"33",X"00",X"60",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"03",X"30",X"90",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"55",X"50",X"00",X"05",X"55",X"55",X"00",X"05",
		X"55",X"55",X"00",X"55",X"55",X"55",X"50",X"33",X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"40",
		X"03",X"00",X"40",X"90",X"33",X"30",X"90",X"03",X"33",X"33",X"60",X"00",X"90",X"90",X"60",X"00",
		X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"03",X"30",X"33",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"50",X"00",X"05",X"55",X"55",X"00",X"05",X"55",X"55",X"00",X"55",X"55",X"55",X"50",X"33",
		X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"90",X"03",X"00",X"40",X"00",X"33",X"30",X"90",X"03",
		X"33",X"33",X"60",X"00",X"90",X"90",X"60",X"00",X"90",X"90",X"00",X"00",X"90",X"33",X"00",X"00",
		X"90",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"55",X"50",X"00",X"05",X"55",X"55",X"00",X"05",
		X"55",X"55",X"00",X"55",X"55",X"55",X"50",X"33",X"33",X"33",X"30",X"40",X"33",X"30",X"40",X"40",
		X"03",X"00",X"90",X"90",X"33",X"30",X"60",X"03",X"33",X"33",X"60",X"00",X"90",X"90",X"00",X"00",
		X"90",X"90",X"00",X"03",X"30",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"30",X"00",X"05",
		X"0D",X"08",X"2F",X"05",X"0D",X"08",X"70",X"05",X"0D",X"08",X"B1",X"05",X"0D",X"08",X"F2",X"05",
		X"0D",X"09",X"33",X"05",X"0D",X"09",X"74",X"05",X"0D",X"09",X"B5",X"05",X"0D",X"09",X"F6",X"05",
		X"0D",X"0A",X"37",X"05",X"0D",X"0A",X"78",X"05",X"0D",X"0A",X"B9",X"05",X"0D",X"0A",X"FA",X"00",
		X"02",X"55",X"00",X"00",X"00",X"09",X"25",X"00",X"00",X"00",X"02",X"25",X"00",X"00",X"00",X"07",
		X"77",X"00",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"07",X"77",
		X"00",X"00",X"00",X"07",X"27",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"88",X"88",X"00",
		X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"55",X"00",X"00",X"00",X"09",X"25",X"00",X"00",X"00",X"02",X"25",X"00",X"00",X"00",
		X"07",X"77",X"00",X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"07",
		X"77",X"70",X"00",X"00",X"27",X"77",X"20",X"00",X"00",X"07",X"88",X"88",X"00",X"00",X"70",X"88",
		X"88",X"00",X"00",X"70",X"88",X"88",X"00",X"02",X"20",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"55",X"00",X"00",X"00",X"09",X"25",X"00",X"00",X"00",X"02",X"25",X"00",X"00",
		X"00",X"07",X"77",X"00",X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"07",X"77",X"70",X"00",X"00",
		X"77",X"77",X"70",X"00",X"00",X"27",X"77",X"20",X"00",X"88",X"88",X"07",X"00",X"00",X"88",X"88",
		X"07",X"00",X"00",X"88",X"88",X"07",X"00",X"00",X"02",X"20",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"20",X"00",X"00",X"00",X"52",X"90",X"00",X"00",X"00",X"52",X"20",X"00",
		X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"77",X"70",X"00",X"00",X"00",X"77",X"70",X"00",X"00",
		X"00",X"77",X"70",X"00",X"00",X"00",X"72",X"70",X"00",X"00",X"00",X"87",X"88",X"00",X"00",X"00",
		X"87",X"88",X"00",X"00",X"00",X"87",X"88",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"20",X"00",X"00",X"00",X"52",X"90",X"00",X"00",X"00",X"52",X"20",
		X"00",X"00",X"00",X"77",X"70",X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"07",X"77",X"70",X"00",
		X"00",X"07",X"77",X"70",X"00",X"00",X"02",X"77",X"72",X"00",X"00",X"00",X"77",X"78",X"88",X"00",
		X"00",X"70",X"87",X"88",X"00",X"00",X"70",X"87",X"88",X"00",X"00",X"22",X"02",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"20",X"00",X"00",X"00",X"52",X"90",X"00",X"00",X"00",X"52",
		X"20",X"00",X"00",X"00",X"77",X"70",X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"07",X"77",X"70",
		X"00",X"00",X"07",X"77",X"77",X"00",X"00",X"02",X"77",X"72",X"00",X"00",X"88",X"77",X"70",X"00",
		X"00",X"88",X"78",X"07",X"00",X"00",X"88",X"78",X"07",X"00",X"00",X"00",X"22",X"02",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"92",X"90",X"00",X"00",X"00",
		X"22",X"20",X"00",X"00",X"77",X"81",X"87",X"70",X"00",X"77",X"71",X"77",X"70",X"00",X"70",X"71",
		X"70",X"70",X"00",X"70",X"71",X"70",X"70",X"00",X"20",X"77",X"70",X"20",X"00",X"00",X"70",X"70",
		X"88",X"00",X"00",X"70",X"70",X"88",X"00",X"00",X"70",X"70",X"88",X"00",X"02",X"20",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"92",X"90",X"00",X"00",
		X"00",X"22",X"20",X"00",X"00",X"77",X"81",X"87",X"70",X"00",X"77",X"71",X"77",X"70",X"00",X"70",
		X"71",X"70",X"70",X"00",X"20",X"71",X"70",X"70",X"00",X"00",X"77",X"70",X"20",X"00",X"00",X"70",
		X"70",X"88",X"00",X"00",X"70",X"70",X"88",X"00",X"00",X"70",X"22",X"88",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"92",X"90",X"00",
		X"00",X"00",X"22",X"20",X"00",X"00",X"77",X"81",X"87",X"70",X"00",X"77",X"71",X"77",X"70",X"00",
		X"70",X"71",X"70",X"70",X"00",X"70",X"71",X"70",X"20",X"00",X"20",X"77",X"70",X"88",X"00",X"00",
		X"70",X"70",X"88",X"00",X"00",X"70",X"70",X"88",X"00",X"02",X"20",X"70",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",X"55",
		X"50",X"00",X"00",X"00",X"45",X"40",X"00",X"00",X"77",X"77",X"77",X"70",X"00",X"77",X"77",X"77",
		X"70",X"00",X"70",X"77",X"70",X"70",X"00",X"70",X"77",X"70",X"70",X"00",X"20",X"77",X"70",X"20",
		X"08",X"80",X"70",X"70",X"00",X"08",X"80",X"70",X"70",X"00",X"08",X"80",X"70",X"70",X"00",X"00",
		X"02",X"20",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"00",
		X"55",X"50",X"00",X"00",X"00",X"45",X"40",X"00",X"00",X"77",X"77",X"77",X"70",X"00",X"77",X"77",
		X"77",X"70",X"00",X"70",X"77",X"70",X"70",X"00",X"20",X"77",X"70",X"70",X"08",X"80",X"77",X"70",
		X"20",X"08",X"80",X"70",X"70",X"00",X"08",X"80",X"70",X"70",X"00",X"00",X"00",X"70",X"22",X"00",
		X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"55",X"50",X"00",X"00",
		X"00",X"55",X"50",X"00",X"00",X"00",X"45",X"40",X"00",X"00",X"77",X"77",X"77",X"70",X"00",X"77",
		X"77",X"77",X"70",X"00",X"70",X"77",X"70",X"70",X"00",X"70",X"77",X"70",X"20",X"00",X"20",X"77",
		X"70",X"00",X"08",X"80",X"70",X"70",X"00",X"08",X"80",X"70",X"70",X"00",X"08",X"82",X"20",X"70",
		X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"20",X"00",X"03",X"0B",X"0B",X"6B",X"03",
		X"0B",X"0B",X"8C",X"03",X"0B",X"0B",X"AD",X"03",X"0B",X"0B",X"CE",X"03",X"0B",X"0B",X"EF",X"03",
		X"0B",X"0C",X"10",X"03",X"0B",X"0C",X"31",X"03",X"0B",X"0C",X"52",X"03",X"0B",X"0C",X"73",X"03",
		X"0B",X"0C",X"94",X"03",X"0B",X"0C",X"B5",X"03",X"0B",X"0C",X"D6",X"02",X"22",X"00",X"09",X"22",
		X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"01",X"91",X"00",X"01",X"91",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"09",X"90",X"00",X"00",X"00",X"00",X"02",X"22",X"00",X"09",
		X"22",X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"09",X"11",X"00",X"90",X"10",
		X"90",X"01",X"01",X"00",X"01",X"00",X"10",X"99",X"09",X"90",X"00",X"00",X"00",X"02",X"22",X"00",
		X"09",X"22",X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"01",X"11",X"90",X"90",
		X"10",X"90",X"01",X"01",X"00",X"01",X"00",X"10",X"99",X"09",X"90",X"00",X"00",X"00",X"02",X"22",
		X"00",X"02",X"29",X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"01",X"91",X"00",
		X"01",X"91",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"02",
		X"22",X"00",X"02",X"29",X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"91",X"11",
		X"00",X"90",X"10",X"90",X"01",X"01",X"00",X"10",X"01",X"00",X"99",X"09",X"90",X"00",X"00",X"00",
		X"02",X"22",X"00",X"02",X"29",X"00",X"02",X"22",X"00",X"00",X"20",X"00",X"01",X"11",X"00",X"01",
		X"19",X"00",X"90",X"10",X"90",X"01",X"01",X"00",X"10",X"01",X"00",X"99",X"09",X"90",X"00",X"00",
		X"00",X"02",X"22",X"00",X"09",X"29",X"00",X"02",X"92",X"00",X"00",X"20",X"00",X"11",X"11",X"10",
		X"91",X"11",X"90",X"91",X"11",X"90",X"01",X"01",X"00",X"01",X"01",X"00",X"99",X"09",X"90",X"00",
		X"00",X"00",X"02",X"22",X"00",X"09",X"29",X"00",X"02",X"92",X"00",X"00",X"20",X"00",X"91",X"11",
		X"10",X"91",X"11",X"90",X"01",X"11",X"90",X"01",X"01",X"00",X"01",X"09",X"90",X"01",X"00",X"00",
		X"99",X"00",X"00",X"02",X"22",X"00",X"09",X"29",X"00",X"02",X"92",X"00",X"00",X"20",X"00",X"11",
		X"11",X"90",X"91",X"11",X"90",X"91",X"11",X"00",X"01",X"01",X"00",X"99",X"01",X"00",X"00",X"01",
		X"00",X"00",X"09",X"90",X"02",X"22",X"00",X"02",X"22",X"00",X"02",X"22",X"00",X"00",X"20",X"00",
		X"11",X"11",X"10",X"91",X"11",X"90",X"91",X"11",X"90",X"01",X"01",X"00",X"01",X"01",X"00",X"99",
		X"09",X"90",X"00",X"00",X"00",X"02",X"22",X"00",X"02",X"22",X"00",X"02",X"22",X"00",X"00",X"20",
		X"00",X"91",X"11",X"10",X"91",X"11",X"90",X"01",X"11",X"90",X"01",X"01",X"00",X"01",X"09",X"90",
		X"01",X"00",X"00",X"99",X"00",X"00",X"02",X"22",X"00",X"02",X"22",X"00",X"02",X"22",X"00",X"00",
		X"20",X"00",X"11",X"11",X"90",X"91",X"11",X"90",X"91",X"11",X"00",X"01",X"01",X"00",X"99",X"01",
		X"00",X"00",X"01",X"00",X"00",X"09",X"90",X"07",X"10",X"07",X"10",X"0D",X"1D",X"07",X"10",X"0D",
		X"8D",X"07",X"10",X"0D",X"FD",X"07",X"10",X"0F",X"BD",X"07",X"10",X"10",X"2D",X"07",X"10",X"10",
		X"9D",X"07",X"10",X"0E",X"6D",X"07",X"10",X"0E",X"DD",X"07",X"10",X"0F",X"4D",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",
		X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",
		X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"6A",X"AA",
		X"66",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"66",X"AA",X"A6",X"00",X"00",
		X"00",X"06",X"66",X"6A",X"AA",X"00",X"00",X"00",X"06",X"66",X"66",X"AA",X"A0",X"00",X"00",X"A6",
		X"66",X"66",X"6A",X"A0",X"00",X"0A",X"A6",X"66",X"66",X"A6",X"00",X"00",X"00",X"06",X"66",X"66",
		X"66",X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"10",X"01",X"10",X"00",X"11",X"10",
		X"00",X"01",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"11",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"06",X"66",X"AA",X"66",X"00",X"00",X"00",X"06",X"6A",X"AA",X"66",X"00",X"00",
		X"00",X"06",X"AA",X"A6",X"66",X"00",X"00",X"00",X"0A",X"AA",X"66",X"66",X"00",X"00",X"A0",X"AA",
		X"A6",X"66",X"66",X"A0",X"00",X"0A",X"A6",X"66",X"66",X"66",X"AA",X"00",X"00",X"06",X"66",X"66",
		X"66",X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"10",X"01",X"10",X"00",X"11",X"10",
		X"00",X"01",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"11",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",
		X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",
		X"66",X"66",X"66",X"0A",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"A0",X"A6",X"66",X"66",
		X"66",X"A0",X"A0",X"A0",X"A0",X"11",X"01",X"10",X"A0",X"A0",X"00",X"00",X"11",X"01",X"10",X"00",
		X"00",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"00",X"11",X"11",X"01",X"11",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",
		X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",
		X"66",X"66",X"66",X"0A",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"A0",X"A6",X"66",X"66",
		X"66",X"A0",X"A0",X"A0",X"A0",X"11",X"01",X"10",X"A0",X"A0",X"00",X"11",X"11",X"01",X"10",X"00",
		X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"10",X"00",X"00",X"00",X"0B",
		X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",
		X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",X"66",X"66",X"66",X"0A",X"A0",X"AA",X"06",
		X"66",X"66",X"66",X"0A",X"A0",X"AA",X"A6",X"66",X"66",X"66",X"AA",X"A0",X"A0",X"A6",X"66",X"66",
		X"66",X"A0",X"A0",X"A0",X"A0",X"11",X"01",X"10",X"A0",X"A0",X"00",X"00",X"11",X"01",X"11",X"10",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",
		X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"66",
		X"AA",X"66",X"60",X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"66",X"AA",X"A6",
		X"60",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"6A",X"AA",X"66",X"60",X"00",X"00",
		X"00",X"AA",X"A6",X"66",X"60",X"00",X"00",X"0A",X"AA",X"66",X"66",X"60",X"00",X"00",X"0A",X"A6",
		X"66",X"66",X"6A",X"00",X"00",X"00",X"6A",X"66",X"66",X"6A",X"A0",X"00",X"00",X"66",X"66",X"66",
		X"60",X"00",X"00",X"00",X"01",X"10",X"11",X"00",X"00",X"00",X"01",X"11",X"00",X"01",X"10",X"01",
		X"00",X"11",X"00",X"00",X"00",X"11",X"10",X"00",X"01",X"11",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"66",X"AA",X"66",X"60",X"00",X"00",X"00",X"66",X"AA",X"A6",X"60",X"00",X"00",
		X"00",X"66",X"6A",X"AA",X"60",X"00",X"00",X"00",X"66",X"66",X"AA",X"A0",X"A0",X"00",X"0A",X"66",
		X"66",X"6A",X"AA",X"00",X"00",X"AA",X"66",X"66",X"66",X"60",X"00",X"00",X"00",X"66",X"66",X"66",
		X"60",X"00",X"00",X"00",X"01",X"10",X"11",X"00",X"00",X"00",X"01",X"11",X"00",X"01",X"10",X"01",
		X"00",X"11",X"00",X"00",X"00",X"11",X"10",X"00",X"01",X"11",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"11",X"68",X"7E",X"12",X"FA",X"14",X"F2",X"18",X"D2",X"18",X"E6",X"D8",X"01",X"08",X"18",
		X"00",X"D1",X"01",X"08",X"08",X"00",X"D0",X"01",X"08",X"1D",X"00",X"D0",X"03",X"04",X"17",X"00",
		X"D0",X"01",X"04",X"15",X"01",X"08",X"14",X"00",X"B6",X"BE",X"6F",X"34",X"02",X"27",X"3E",X"BD",
		X"D0",X"6C",X"11",X"AF",X"15",X"02",X"12",X"C8",X"27",X"33",X"BD",X"26",X"C3",X"86",X"09",X"0D",
		X"84",X"2B",X"02",X"86",X"87",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"B6",X"BE",X"60",X"BD",X"D0",
		X"3F",X"A7",X"49",X"B6",X"BE",X"5E",X"BD",X"D0",X"3F",X"44",X"89",X"00",X"A7",X"4A",X"BD",X"12",
		X"5F",X"CC",X"15",X"02",X"ED",X"88",X"16",X"9F",X"17",X"6A",X"E4",X"26",X"C2",X"35",X"82",X"AE",
		X"47",X"EC",X"02",X"C3",X"00",X"04",X"10",X"83",X"15",X"02",X"23",X"0B",X"CC",X"14",X"F2",X"0D",
		X"59",X"26",X"04",X"6A",X"49",X"27",X"14",X"ED",X"02",X"6A",X"4E",X"26",X"03",X"BD",X"12",X"5F",
		X"BD",X"12",X"79",X"86",X"02",X"8E",X"11",X"AF",X"7E",X"D0",X"66",X"B6",X"BE",X"60",X"44",X"44",
		X"BD",X"D0",X"3F",X"A7",X"49",X"AE",X"47",X"EC",X"02",X"C3",X"00",X"04",X"10",X"83",X"15",X"0E",
		X"23",X"1C",X"6A",X"49",X"26",X"15",X"96",X"ED",X"81",X"08",X"24",X"DF",X"96",X"42",X"81",X"11",
		X"24",X"D9",X"BD",X"13",X"54",X"6A",X"4A",X"27",X"19",X"20",X"D0",X"CC",X"14",X"F2",X"ED",X"02",
		X"6A",X"4E",X"26",X"03",X"BD",X"12",X"5F",X"BD",X"12",X"79",X"86",X"02",X"8E",X"11",X"E5",X"7E",
		X"D0",X"66",X"CC",X"00",X"00",X"ED",X"88",X"10",X"CC",X"01",X"00",X"0D",X"84",X"2A",X"01",X"40",
		X"ED",X"0E",X"AE",X"47",X"EC",X"02",X"C3",X"00",X"04",X"10",X"83",X"15",X"02",X"23",X"0D",X"A6",
		X"0A",X"81",X"0A",X"23",X"11",X"81",X"85",X"24",X"0D",X"CC",X"14",X"F2",X"ED",X"02",X"86",X"02",
		X"8E",X"12",X"32",X"7E",X"D0",X"66",X"BD",X"D0",X"75",X"7A",X"BE",X"6F",X"7E",X"D0",X"63",X"96",
		X"85",X"84",X"1F",X"8B",X"F0",X"A7",X"4C",X"96",X"86",X"98",X"84",X"84",X"3F",X"8B",X"E0",X"A7",
		X"4D",X"86",X"0F",X"BD",X"D0",X"42",X"A7",X"4E",X"39",X"E6",X"4C",X"1D",X"E3",X"0E",X"10",X"83",
		X"01",X"00",X"2D",X"03",X"CC",X"01",X"00",X"10",X"83",X"FF",X"00",X"2E",X"03",X"CC",X"FF",X"00",
		X"ED",X"0E",X"43",X"53",X"58",X"49",X"58",X"49",X"1F",X"89",X"1D",X"E3",X"0E",X"ED",X"0E",X"E6",
		X"4D",X"1D",X"E3",X"88",X"10",X"10",X"83",X"02",X"00",X"2D",X"03",X"CC",X"02",X"00",X"10",X"83",
		X"FE",X"00",X"2E",X"03",X"CC",X"FE",X"00",X"ED",X"88",X"10",X"43",X"53",X"58",X"49",X"1F",X"89",
		X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"39",X"96",X"48",X"26",X"24",X"BD",X"D0",X"78",X"DE",
		X"1B",X"EC",X"C4",X"DD",X"1B",X"BD",X"D0",X"54",X"12",X"F1",X"EF",X"07",X"CC",X"14",X"F6",X"ED",
		X"42",X"7A",X"BE",X"6F",X"CC",X"02",X"10",X"BD",X"D0",X"0C",X"CC",X"11",X"51",X"7E",X"D0",X"4B",
		X"39",X"CC",X"FF",X"AA",X"ED",X"4B",X"86",X"07",X"A7",X"4D",X"AE",X"47",X"10",X"AE",X"02",X"EC",
		X"04",X"BD",X"D0",X"1E",X"31",X"24",X"10",X"AF",X"02",X"6A",X"4D",X"27",X"11",X"A6",X"4C",X"97",
		X"2D",X"EC",X"04",X"BD",X"D0",X"90",X"86",X"02",X"8E",X"12",X"FA",X"7E",X"D0",X"66",X"EC",X"04",
		X"C3",X"01",X"05",X"ED",X"04",X"86",X"1E",X"A7",X"49",X"FC",X"00",X"0C",X"ED",X"02",X"AE",X"47",
		X"A6",X"4B",X"97",X"2D",X"10",X"AE",X"02",X"EC",X"04",X"BD",X"D0",X"90",X"6A",X"49",X"27",X"08",
		X"86",X"02",X"8E",X"13",X"2E",X"7E",X"D0",X"66",X"BD",X"D0",X"1E",X"DC",X"1B",X"ED",X"84",X"9F",
		X"1B",X"7E",X"D0",X"63",X"34",X"76",X"1F",X"12",X"BD",X"D0",X"6C",X"13",X"90",X"18",X"D2",X"14",
		X"83",X"27",X"1C",X"A6",X"2A",X"E6",X"2C",X"A7",X"0A",X"E7",X"0C",X"ED",X"04",X"B6",X"BE",X"5F",
		X"BD",X"D0",X"3F",X"A7",X"4D",X"9F",X"17",X"CC",X"11",X"4C",X"BD",X"D0",X"4B",X"0C",X"ED",X"35",
		X"F6",X"AE",X"47",X"EC",X"02",X"C3",X"00",X"04",X"10",X"83",X"18",X"E6",X"24",X"0A",X"ED",X"02",
		X"86",X"08",X"8E",X"13",X"81",X"7E",X"D0",X"66",X"ED",X"02",X"BD",X"13",X"B5",X"AE",X"47",X"6A",
		X"4E",X"26",X"03",X"BD",X"13",X"B5",X"6A",X"4D",X"26",X"03",X"BD",X"14",X"04",X"86",X"03",X"8E",
		X"13",X"9D",X"7E",X"D0",X"66",X"BD",X"D0",X"3C",X"84",X"1F",X"A7",X"4E",X"4F",X"57",X"57",X"57",
		X"DB",X"5E",X"C1",X"07",X"24",X"02",X"C6",X"07",X"81",X"8F",X"23",X"0A",X"C1",X"CF",X"24",X"04",
		X"C6",X"8F",X"20",X"02",X"C6",X"07",X"E0",X"0A",X"82",X"00",X"58",X"49",X"ED",X"0E",X"4F",X"D6",
		X"85",X"57",X"57",X"57",X"DB",X"5F",X"C1",X"EA",X"23",X"02",X"C6",X"EA",X"C1",X"18",X"24",X"0A",
		X"C1",X"0C",X"24",X"04",X"C6",X"EA",X"20",X"02",X"C6",X"18",X"E0",X"0C",X"82",X"00",X"58",X"49",
		X"ED",X"88",X"10",X"39",X"34",X"50",X"1F",X"12",X"B6",X"BE",X"5F",X"BD",X"D0",X"3F",X"A7",X"4D",
		X"96",X"8A",X"81",X"14",X"24",X"6B",X"96",X"42",X"81",X"11",X"24",X"65",X"BD",X"D0",X"6C",X"14",
		X"A8",X"1A",X"34",X"14",X"DC",X"27",X"5A",X"0C",X"8A",X"EC",X"24",X"A7",X"0A",X"E7",X"0C",X"ED",
		X"04",X"D6",X"84",X"C4",X"1F",X"CB",X"F0",X"96",X"5E",X"81",X"17",X"24",X"01",X"5F",X"DB",X"5E",
		X"4F",X"E0",X"04",X"82",X"00",X"58",X"49",X"58",X"49",X"ED",X"0E",X"D6",X"86",X"C4",X"1F",X"CB",
		X"F0",X"DB",X"5F",X"4F",X"E0",X"05",X"82",X"00",X"58",X"49",X"58",X"49",X"ED",X"88",X"10",X"D6",
		X"86",X"C4",X"1F",X"CB",X"F0",X"1D",X"ED",X"49",X"D6",X"85",X"C4",X"1F",X"CB",X"F0",X"1D",X"ED",
		X"4B",X"9F",X"17",X"96",X"85",X"84",X"0F",X"8B",X"14",X"A7",X"4E",X"CC",X"11",X"56",X"BD",X"D0",
		X"4B",X"35",X"D0",X"96",X"48",X"26",X"20",X"BD",X"D0",X"78",X"9E",X"1B",X"EC",X"84",X"DD",X"1B",
		X"BD",X"5B",X"43",X"DC",X"1B",X"ED",X"84",X"9F",X"1B",X"0A",X"ED",X"CC",X"01",X"15",X"BD",X"D0",
		X"0C",X"CC",X"11",X"5B",X"7E",X"D0",X"4B",X"39",X"AE",X"47",X"EC",X"02",X"C3",X"00",X"04",X"10",
		X"83",X"1A",X"40",X"23",X"03",X"CC",X"1A",X"34",X"ED",X"02",X"EC",X"0E",X"E3",X"49",X"ED",X"0E",
		X"EC",X"88",X"10",X"E3",X"4B",X"ED",X"88",X"10",X"6A",X"4E",X"27",X"08",X"86",X"04",X"8E",X"14",
		X"A8",X"7E",X"D0",X"66",X"BD",X"D0",X"75",X"0A",X"8A",X"7E",X"D0",X"63",X"96",X"48",X"26",X"11",
		X"BD",X"D0",X"78",X"0A",X"8A",X"CC",X"00",X"25",X"BD",X"D0",X"0C",X"CC",X"11",X"60",X"7E",X"D0",
		X"4B",X"39",X"08",X"0F",X"15",X"12",X"08",X"0F",X"15",X"8A",X"08",X"0F",X"16",X"02",X"08",X"0F",
		X"16",X"7A",X"08",X"0F",X"16",X"F2",X"08",X"0F",X"17",X"6A",X"08",X"0F",X"17",X"E2",X"08",X"0F",
		X"18",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"F0",
		X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"FF",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"FF",X"00",X"0F",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",
		X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",
		X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"FF",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"05",X"0B",X"19",X"21",X"05",X"0B",X"19",X"58",X"05",X"0B",X"19",X"8F",X"05",X"0B",
		X"19",X"C6",X"05",X"0B",X"19",X"FD",X"05",X"0B",X"18",X"EA",X"00",X"00",X"80",X"00",X"00",X"00",
		X"08",X"88",X"00",X"00",X"00",X"8A",X"AA",X"80",X"00",X"08",X"FF",X"FF",X"F8",X"00",X"00",X"08",
		X"88",X"00",X"00",X"90",X"88",X"78",X"80",X"90",X"09",X"97",X"77",X"99",X"00",X"90",X"77",X"77",
		X"70",X"90",X"00",X"00",X"80",X"00",X"00",X"00",X"DD",X"DD",X"D0",X"00",X"0D",X"DD",X"DD",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"08",X"F8",X"00",X"00",X"00",
		X"00",X"70",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"08",X"F8",X"00",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"09",X"79",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"00",X"00",X"00",X"08",X"FF",X"80",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"09",X"77",
		X"90",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"08",X"A8",X"00",X"00",X"00",X"8F",X"FF",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"08",X"78",X"00",X"00",X"09",X"97",X"77",X"99",X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"0D",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"08",X"AA",X"80",X"00",X"00",X"8F",X"FF",X"F8",
		X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"98",X"88",X"89",X"00",X"00",X"09",X"77",X"90",X"00",
		X"00",X"97",X"77",X"79",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"0D",X"DD",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"07",X"1A",X"44",X"04",X"07",X"1A",X"60",X"04",X"07",X"1A",X"7C",
		X"04",X"07",X"1A",X"98",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"FF",X"FB",X"FF",X"F0",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"0B",X"00",X"00",X"F0",X"B0",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"B0",X"F0",X"00",X"0B",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"BB",X"BB",X"BB",X"B0",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0F",X"00",
		X"00",X"B0",X"F0",X"00",X"00",X"0B",X"00",X"00",X"00",X"F0",X"B0",X"00",X"0F",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"1A",X"F4",X"21",X"41",X"7E",X"1D",X"AF",X"7E",X"1D",X"C2",X"1F",X"68",X"D0",X"01",X"04",
		X"14",X"01",X"08",X"11",X"00",X"D0",X"02",X"04",X"17",X"00",X"D0",X"01",X"04",X"14",X"02",X"04",
		X"17",X"00",X"C8",X"01",X"08",X"15",X"01",X"08",X"14",X"00",X"D0",X"02",X"03",X"12",X"00",X"D8",
		X"01",X"08",X"11",X"00",X"0F",X"95",X"B6",X"BE",X"6E",X"34",X"02",X"27",X"58",X"D6",X"95",X"10",
		X"8E",X"D0",X"15",X"EB",X"A4",X"31",X"28",X"10",X"8C",X"EA",X"B1",X"25",X"F6",X"C1",X"4A",X"27",
		X"0E",X"96",X"85",X"81",X"20",X"24",X"08",X"86",X"98",X"D6",X"86",X"1F",X"02",X"63",X"A4",X"BD",
		X"D0",X"54",X"1B",X"D8",X"33",X"84",X"BD",X"D0",X"7B",X"CC",X"21",X"59",X"ED",X"02",X"ED",X"88",
		X"14",X"EF",X"06",X"AF",X"47",X"CC",X"1C",X"B2",X"ED",X"4D",X"6F",X"4B",X"CC",X"1D",X"D6",X"ED",
		X"08",X"8D",X"14",X"BD",X"1B",X"95",X"B6",X"BE",X"62",X"BD",X"D0",X"3F",X"A7",X"4C",X"BD",X"D0",
		X"18",X"6A",X"E4",X"26",X"CA",X"35",X"82",X"BD",X"26",X"C3",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",
		X"10",X"AE",X"02",X"0D",X"84",X"2B",X"17",X"86",X"10",X"BD",X"D0",X"42",X"0D",X"85",X"2B",X"04",
		X"8B",X"07",X"20",X"05",X"AB",X"A4",X"40",X"8B",X"8F",X"A7",X"04",X"A7",X"0A",X"39",X"86",X"20",
		X"BD",X"D0",X"42",X"0D",X"86",X"2B",X"04",X"8B",X"18",X"20",X"05",X"AB",X"21",X"40",X"8B",X"EA",
		X"A7",X"05",X"A7",X"0C",X"39",X"CC",X"FF",X"FF",X"10",X"8E",X"B3",X"54",X"34",X"66",X"EE",X"A4",
		X"27",X"28",X"4F",X"E6",X"44",X"E0",X"04",X"82",X"00",X"2A",X"04",X"43",X"50",X"82",X"FF",X"DD",
		X"2B",X"4F",X"E6",X"45",X"E0",X"05",X"82",X"00",X"2A",X"04",X"43",X"50",X"82",X"FF",X"D3",X"2B",
		X"10",X"A3",X"E4",X"22",X"05",X"ED",X"E4",X"10",X"AF",X"62",X"31",X"22",X"10",X"8C",X"B3",X"A4",
		X"26",X"CC",X"35",X"66",X"10",X"AF",X"49",X"39",X"96",X"59",X"85",X"7F",X"27",X"08",X"86",X"04",
		X"8E",X"1B",X"D8",X"7E",X"D0",X"66",X"86",X"0C",X"8E",X"1B",X"EE",X"7E",X"D0",X"66",X"AE",X"47",
		X"CC",X"00",X"00",X"DD",X"2B",X"10",X"AE",X"D8",X"09",X"26",X"14",X"10",X"8E",X"98",X"5A",X"B6",
		X"BE",X"6A",X"BB",X"BE",X"6B",X"BB",X"BE",X"6C",X"27",X"05",X"BD",X"1B",X"95",X"20",X"E6",X"A6",
		X"24",X"A0",X"04",X"8B",X"02",X"81",X"04",X"23",X"0B",X"C6",X"01",X"A6",X"24",X"A1",X"04",X"24",
		X"01",X"50",X"D7",X"2B",X"A6",X"25",X"C6",X"01",X"A1",X"05",X"24",X"01",X"50",X"D7",X"2C",X"EC",
		X"04",X"9B",X"2B",X"DB",X"2C",X"BD",X"00",X"06",X"27",X"04",X"90",X"2B",X"D0",X"2C",X"A7",X"0A",
		X"E7",X"0C",X"10",X"8C",X"98",X"5A",X"27",X"10",X"E0",X"25",X"CB",X"03",X"C1",X"06",X"22",X"08",
		X"A0",X"24",X"8B",X"03",X"81",X"06",X"23",X"6A",X"96",X"2B",X"27",X"0C",X"2B",X"05",X"CC",X"1C",
		X"AA",X"20",X"11",X"CC",X"1C",X"A2",X"20",X"0C",X"96",X"2C",X"2B",X"05",X"CC",X"1C",X"B2",X"20",
		X"03",X"CC",X"1C",X"BA",X"10",X"A3",X"4D",X"27",X"04",X"ED",X"4D",X"20",X"08",X"E6",X"4B",X"CB",
		X"02",X"C1",X"08",X"25",X"01",X"5F",X"E7",X"4B",X"10",X"AE",X"4D",X"EC",X"A5",X"ED",X"02",X"BD",
		X"D0",X"8D",X"6A",X"4C",X"26",X"03",X"BD",X"20",X"06",X"8E",X"1B",X"EE",X"B6",X"BE",X"63",X"7E",
		X"D0",X"66",X"21",X"41",X"21",X"45",X"21",X"41",X"21",X"49",X"21",X"4D",X"21",X"51",X"21",X"4D",
		X"21",X"55",X"21",X"59",X"21",X"5D",X"21",X"59",X"21",X"61",X"21",X"65",X"21",X"69",X"21",X"65",
		X"21",X"6D",X"A6",X"0A",X"A1",X"24",X"25",X"12",X"A6",X"0A",X"A0",X"B8",X"02",X"80",X"01",X"81",
		X"07",X"25",X"07",X"A7",X"2A",X"CC",X"21",X"41",X"20",X"0D",X"A6",X"0A",X"8B",X"08",X"81",X"8B",
		X"24",X"E6",X"A7",X"2A",X"CC",X"21",X"4D",X"ED",X"02",X"A6",X"0C",X"8B",X"02",X"A7",X"2C",X"BD",
		X"D0",X"15",X"6F",X"0B",X"6F",X"88",X"12",X"BD",X"1D",X"AF",X"AE",X"D8",X"09",X"34",X"50",X"86",
		X"01",X"97",X"95",X"AD",X"98",X"08",X"35",X"50",X"0F",X"95",X"EC",X"84",X"DD",X"1B",X"AF",X"49",
		X"6F",X"0B",X"6F",X"88",X"12",X"10",X"AE",X"06",X"EC",X"29",X"ED",X"02",X"86",X"14",X"A7",X"4B",
		X"AE",X"47",X"CC",X"1A",X"EA",X"BD",X"D0",X"4B",X"BD",X"1D",X"AF",X"AE",X"49",X"EC",X"04",X"10",
		X"AE",X"02",X"BD",X"D0",X"1E",X"A6",X"0A",X"D6",X"84",X"C4",X"07",X"EB",X"0C",X"C1",X"DC",X"23",
		X"02",X"C6",X"DC",X"ED",X"04",X"CC",X"AA",X"BB",X"8D",X"78",X"86",X"02",X"8E",X"1D",X"52",X"7E",
		X"D0",X"66",X"AE",X"49",X"EC",X"04",X"10",X"AE",X"02",X"BD",X"D0",X"1E",X"A6",X"0A",X"D6",X"84",
		X"C4",X"07",X"50",X"EB",X"0C",X"C1",X"18",X"24",X"02",X"C6",X"18",X"ED",X"04",X"CC",X"AA",X"BB",
		X"8D",X"50",X"86",X"02",X"8E",X"1D",X"7A",X"7E",X"D0",X"66",X"6A",X"4B",X"26",X"A2",X"CC",X"1A",
		X"EF",X"BD",X"D0",X"4B",X"AE",X"49",X"DC",X"1B",X"ED",X"84",X"9F",X"1B",X"EC",X"04",X"10",X"AE",
		X"02",X"BD",X"D0",X"1E",X"EC",X"04",X"10",X"AE",X"02",X"BD",X"1E",X"19",X"AE",X"47",X"EC",X"04",
		X"10",X"AE",X"02",X"BD",X"D0",X"1E",X"BD",X"D0",X"18",X"BD",X"1B",X"95",X"7E",X"1B",X"EE",X"C6",
		X"BB",X"D7",X"2D",X"A6",X"0A",X"E6",X"0C",X"ED",X"04",X"10",X"AE",X"02",X"BD",X"D0",X"93",X"7E",
		X"D0",X"18",X"34",X"06",X"97",X"2D",X"EC",X"04",X"BD",X"D0",X"93",X"A6",X"61",X"97",X"2D",X"A6",
		X"04",X"BD",X"D0",X"90",X"35",X"86",X"96",X"48",X"26",X"3C",X"7A",X"BE",X"6E",X"BD",X"5B",X"4F",
		X"BD",X"D0",X"7E",X"AE",X"06",X"33",X"84",X"BD",X"D0",X"5D",X"EC",X"42",X"10",X"83",X"1D",X"52",
		X"25",X"17",X"AE",X"49",X"DC",X"1B",X"ED",X"84",X"9F",X"1B",X"10",X"AE",X"02",X"EC",X"04",X"BD",
		X"D0",X"1E",X"0C",X"95",X"BD",X"00",X"09",X"0F",X"95",X"CC",X"1A",X"CD",X"BD",X"D0",X"4B",X"CC",
		X"01",X"50",X"BD",X"D0",X"0C",X"39",X"7E",X"D0",X"18",X"34",X"56",X"DC",X"1D",X"27",X"34",X"4F",
		X"8E",X"1E",X"AB",X"BD",X"D0",X"5A",X"33",X"84",X"BD",X"1F",X"FC",X"86",X"11",X"A7",X"4F",X"BD",
		X"D0",X"7B",X"AF",X"47",X"EF",X"06",X"10",X"AF",X"49",X"10",X"AF",X"02",X"10",X"AF",X"88",X"14",
		X"EC",X"E4",X"A7",X"0A",X"E7",X"0C",X"CC",X"1F",X"1F",X"ED",X"08",X"8D",X"08",X"8D",X"22",X"4F",
		X"5F",X"ED",X"04",X"35",X"D6",X"86",X"0F",X"BD",X"D0",X"3F",X"8B",X"F0",X"40",X"48",X"48",X"8B",
		X"E0",X"A7",X"4B",X"86",X"12",X"BD",X"D0",X"3F",X"8B",X"ED",X"40",X"48",X"8B",X"EE",X"A7",X"4C",
		X"39",X"96",X"85",X"2B",X"18",X"96",X"64",X"AB",X"4B",X"81",X"BF",X"23",X"02",X"86",X"07",X"A1",
		X"0A",X"23",X"05",X"CC",X"1F",X"D8",X"20",X"1B",X"CC",X"1F",X"CC",X"20",X"16",X"96",X"66",X"AB",
		X"4C",X"81",X"FC",X"23",X"02",X"86",X"18",X"A1",X"0C",X"23",X"05",X"CC",X"1F",X"E4",X"20",X"03",
		X"CC",X"1F",X"F0",X"ED",X"4D",X"86",X"FD",X"A7",X"88",X"13",X"39",X"AE",X"47",X"10",X"AE",X"4D",
		X"A6",X"88",X"13",X"8B",X"03",X"81",X"09",X"23",X"01",X"4F",X"A7",X"88",X"13",X"31",X"A6",X"E6",
		X"A4",X"4F",X"E3",X"49",X"ED",X"02",X"EC",X"21",X"AB",X"0A",X"EB",X"0C",X"BD",X"00",X"06",X"26",
		X"13",X"A7",X"0A",X"E7",X"0C",X"96",X"84",X"81",X"F8",X"23",X"03",X"BD",X"1E",X"55",X"96",X"86",
		X"81",X"E4",X"23",X"03",X"BD",X"1E",X"71",X"10",X"AE",X"02",X"A6",X"4F",X"EC",X"C6",X"BD",X"D0",
		X"1E",X"CC",X"EE",X"00",X"BD",X"1D",X"C2",X"A6",X"0A",X"E6",X"0C",X"ED",X"04",X"1F",X"02",X"A6",
		X"4F",X"10",X"AF",X"C6",X"8B",X"02",X"81",X"1F",X"25",X"02",X"86",X"11",X"A7",X"4F",X"10",X"AE",
		X"02",X"CC",X"00",X"AA",X"BD",X"1D",X"C2",X"86",X"03",X"8E",X"1E",X"AB",X"7E",X"D0",X"66",X"96",
		X"48",X"26",X"44",X"34",X"10",X"10",X"AE",X"02",X"AE",X"06",X"86",X"11",X"34",X"02",X"EC",X"86",
		X"BD",X"D0",X"1E",X"35",X"02",X"8B",X"02",X"81",X"1F",X"25",X"F1",X"BD",X"D0",X"5D",X"35",X"10",
		X"CC",X"1F",X"68",X"ED",X"02",X"86",X"8A",X"A1",X"04",X"24",X"02",X"A7",X"04",X"86",X"DB",X"A1",
		X"05",X"24",X"02",X"A7",X"05",X"BD",X"5B",X"43",X"BD",X"D0",X"7E",X"CC",X"1A",X"DA",X"BD",X"D0",
		X"4B",X"CC",X"01",X"10",X"BD",X"D0",X"0C",X"39",X"06",X"10",X"1F",X"6C",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"A0",X"AA",X"00",X"00",X"00",X"0A",X"A0",X"AA",X"0B",X"B0",X"BB",X"0A",X"A0",X"AA",X"0B",
		X"B0",X"BB",X"0A",X"A0",X"AA",X"0B",X"B0",X"BB",X"0A",X"A0",X"AA",X"00",X"00",X"00",X"0A",X"A0",
		X"AA",X"AA",X"A0",X"AA",X"AA",X"A0",X"AA",X"A0",X"00",X"00",X"AA",X"A0",X"AA",X"00",X"00",X"00",
		X"0A",X"A0",X"AA",X"0A",X"00",X"0A",X"0A",X"A0",X"AA",X"0A",X"00",X"0A",X"0A",X"A0",X"AA",X"AA",
		X"0A",X"0A",X"AA",X"A0",X"AA",X"AA",X"0A",X"0A",X"AA",X"A0",X"AA",X"AA",X"0A",X"0A",X"AA",X"A0",
		X"AA",X"00",X"0A",X"00",X"0A",X"A0",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"FE",X"00",X"04",
		X"FE",X"00",X"00",X"FE",X"00",X"08",X"FE",X"00",X"0C",X"02",X"00",X"10",X"02",X"00",X"0C",X"02",
		X"00",X"14",X"02",X"00",X"18",X"00",X"04",X"1C",X"00",X"04",X"18",X"00",X"04",X"20",X"00",X"04",
		X"24",X"00",X"FC",X"28",X"00",X"FC",X"24",X"00",X"FC",X"2C",X"00",X"FC",X"86",X"07",X"6F",X"C6",
		X"4C",X"81",X"1F",X"25",X"F9",X"39",X"34",X"50",X"B6",X"BE",X"62",X"BD",X"D0",X"3F",X"A7",X"4C",
		X"96",X"8E",X"81",X"08",X"24",X"43",X"DC",X"1D",X"27",X"3F",X"31",X"84",X"4F",X"8E",X"20",X"B0",
		X"BD",X"D0",X"5A",X"33",X"84",X"8D",X"D5",X"BD",X"D0",X"7B",X"CC",X"20",X"5B",X"ED",X"88",X"16",
		X"CC",X"20",X"6B",X"ED",X"02",X"ED",X"88",X"14",X"CC",X"21",X"19",X"ED",X"08",X"EF",X"06",X"AF",
		X"47",X"EC",X"24",X"C3",X"03",X"04",X"ED",X"04",X"ED",X"0A",X"BD",X"20",X"7B",X"0C",X"8E",X"86",
		X"0D",X"A7",X"4C",X"CC",X"1A",X"E2",X"BD",X"D0",X"4B",X"35",X"D0",X"03",X"04",X"20",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"04",X"20",X"6F",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"CC",X"00",X"00",X"ED",X"49",
		X"96",X"84",X"2A",X"13",X"84",X"0F",X"8B",X"FA",X"9B",X"64",X"C6",X"01",X"A1",X"0A",X"24",X"01",
		X"50",X"E7",X"49",X"96",X"86",X"2B",X"11",X"96",X"85",X"84",X"0F",X"8B",X"FA",X"C6",X"01",X"9B",
		X"66",X"A1",X"0B",X"24",X"01",X"50",X"E7",X"4A",X"86",X"07",X"BD",X"D0",X"3F",X"A7",X"4B",X"39",
		X"AE",X"47",X"6A",X"4B",X"26",X"03",X"BD",X"20",X"7B",X"BD",X"20",X"C7",X"BD",X"20",X"C7",X"86",
		X"02",X"8E",X"20",X"B0",X"7E",X"D0",X"66",X"EC",X"0A",X"AB",X"49",X"81",X"07",X"24",X"06",X"A0",
		X"49",X"60",X"49",X"20",X"F4",X"81",X"8E",X"22",X"F6",X"EB",X"4A",X"C1",X"18",X"24",X"06",X"E0",
		X"4A",X"60",X"4A",X"20",X"F4",X"C1",X"EA",X"22",X"F6",X"10",X"8E",X"DD",X"DD",X"10",X"AF",X"98",
		X"0A",X"ED",X"0A",X"83",X"01",X"01",X"ED",X"04",X"10",X"8E",X"00",X"00",X"A6",X"4C",X"10",X"AF",
		X"D6",X"CC",X"AA",X"AA",X"10",X"AE",X"0A",X"ED",X"A4",X"A6",X"4C",X"10",X"AF",X"C6",X"8B",X"02",
		X"81",X"1F",X"25",X"02",X"86",X"0D",X"A7",X"4C",X"39",X"0A",X"8E",X"96",X"48",X"26",X"21",X"BD",
		X"D0",X"7E",X"AE",X"06",X"CE",X"00",X"00",X"86",X"0D",X"EF",X"96",X"8B",X"02",X"81",X"1F",X"26",
		X"F8",X"BD",X"D0",X"5D",X"CC",X"00",X"25",X"BD",X"D0",X"0C",X"CC",X"1A",X"D5",X"BD",X"D0",X"4B",
		X"39",X"07",X"10",X"21",X"71",X"07",X"10",X"21",X"E1",X"07",X"10",X"22",X"51",X"07",X"10",X"22",
		X"C1",X"07",X"10",X"23",X"31",X"07",X"10",X"23",X"A1",X"07",X"10",X"24",X"11",X"07",X"10",X"24",
		X"81",X"07",X"10",X"24",X"F1",X"07",X"10",X"25",X"61",X"07",X"10",X"25",X"D1",X"07",X"10",X"26",
		X"41",X"00",X"00",X"7C",X"7C",X"70",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"7C",X"00",X"00",X"00",
		X"7C",X"7C",X"C0",X"CC",X"70",X"00",X"07",X"0C",X"C0",X"C7",X"C0",X"C7",X"00",X"0C",X"CC",X"7C",
		X"CC",X"C7",X"C7",X"00",X"07",X"77",X"7C",X"C7",X"C0",X"CC",X"00",X"00",X"07",X"77",X"CC",X"0C",
		X"C7",X"00",X"00",X"7A",X"A7",X"77",X"0C",X"70",X"00",X"00",X"77",X"77",X"7C",X"C0",X"00",X"00",
		X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"00",X"66",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"04",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"7C",X"7C",X"70",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"7C",X"00",X"00",X"00",
		X"7C",X"7C",X"C0",X"CC",X"70",X"00",X"07",X"0C",X"C0",X"C7",X"C0",X"C7",X"00",X"0C",X"CC",X"7C",
		X"CC",X"C7",X"C7",X"00",X"07",X"77",X"7C",X"C7",X"C0",X"CC",X"00",X"00",X"07",X"77",X"CC",X"0C",
		X"C7",X"00",X"00",X"7A",X"A7",X"77",X"0C",X"70",X"00",X"00",X"77",X"77",X"7C",X"C0",X"00",X"00",
		X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"00",X"66",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"40",X"40",X"06",
		X"00",X"00",X"00",X"00",X"04",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"7C",X"7C",X"70",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"7C",X"00",X"00",X"00",
		X"7C",X"7C",X"C0",X"CC",X"70",X"00",X"07",X"0C",X"C0",X"C7",X"C0",X"C7",X"00",X"0C",X"CC",X"7C",
		X"CC",X"C7",X"C7",X"00",X"07",X"77",X"7C",X"C7",X"C0",X"CC",X"00",X"00",X"07",X"77",X"CC",X"0C",
		X"C7",X"00",X"00",X"7A",X"A7",X"77",X"0C",X"70",X"00",X"00",X"77",X"77",X"7C",X"C0",X"00",X"00",
		X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"00",X"06",X"70",X"00",X"00",X"00",X"00",X"66",
		X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"40",X"00",X"00",X"00",X"00",X"60",X"60",X"04",
		X"00",X"00",X"00",X"00",X"06",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"CC",X"7C",X"00",X"00",X"00",X"00",X"CC",X"7C",X"CC",X"70",X"00",X"00",X"07",
		X"C7",X"0C",X"70",X"7C",X"00",X"00",X"77",X"CC",X"7C",X"7C",X"CC",X"70",X"00",X"CC",X"0C",X"CC",
		X"0C",X"70",X"70",X"00",X"7C",X"C0",X"7C",X"CC",X"CC",X"70",X"00",X"77",X"CC",X"CC",X"77",X"70",
		X"00",X"00",X"0C",X"C7",X"C7",X"7A",X"A7",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"00",
		X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"CC",X"7C",X"00",X"00",X"00",X"00",X"CC",X"7C",X"CC",X"70",X"00",X"00",X"07",
		X"C7",X"0C",X"70",X"7C",X"00",X"00",X"77",X"CC",X"7C",X"7C",X"CC",X"70",X"00",X"CC",X"0C",X"CC",
		X"0C",X"70",X"70",X"00",X"7C",X"C0",X"7C",X"CC",X"CC",X"70",X"00",X"77",X"CC",X"CC",X"77",X"70",
		X"00",X"00",X"0C",X"C7",X"C7",X"7A",X"A7",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"00",
		X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"60",X"04",
		X"04",X"00",X"00",X"00",X"00",X"06",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"CC",X"7C",X"00",X"00",X"00",X"00",X"CC",X"7C",X"CC",X"70",X"00",X"00",X"07",
		X"C7",X"0C",X"70",X"7C",X"00",X"00",X"77",X"CC",X"7C",X"7C",X"CC",X"70",X"00",X"CC",X"0C",X"CC",
		X"0C",X"70",X"70",X"00",X"7C",X"C0",X"7C",X"CC",X"CC",X"70",X"00",X"77",X"CC",X"CC",X"77",X"70",
		X"00",X"00",X"0C",X"C7",X"C7",X"7A",X"A7",X"00",X"00",X"00",X"07",X"77",X"77",X"77",X"00",X"00",
		X"00",X"00",X"07",X"77",X"70",X"00",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"04",X"60",X"00",X"00",X"00",X"00",X"00",X"40",X"06",
		X"06",X"00",X"00",X"00",X"00",X"04",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"70",X"00",X"00",X"00",X"00",X"7C",X"C7",X"7C",X"7C",X"70",X"00",X"07",
		X"CC",X"0C",X"CC",X"0C",X"77",X"00",X"77",X"C7",X"C7",X"C0",X"C0",X"CC",X"70",X"CC",X"C0",X"CC",
		X"C7",X"CC",X"0C",X"70",X"C7",X"C7",X"7C",X"0C",X"77",X"C7",X"C0",X"70",X"C7",X"77",X"C7",X"70",
		X"7C",X"70",X"0C",X"CA",X"AA",X"7A",X"AA",X"77",X"00",X"07",X"77",X"77",X"77",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"00",X"60",X"06",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"70",X"00",X"00",X"00",X"00",X"7C",X"C7",X"7C",X"7C",X"70",X"00",X"07",
		X"CC",X"0C",X"CC",X"0C",X"77",X"00",X"77",X"C7",X"C7",X"C0",X"C0",X"CC",X"70",X"CC",X"C0",X"CC",
		X"C7",X"CC",X"0C",X"70",X"C7",X"C7",X"7C",X"0C",X"77",X"C7",X"C0",X"70",X"C7",X"77",X"C7",X"70",
		X"7C",X"70",X"0C",X"CA",X"AA",X"7A",X"AA",X"77",X"00",X"07",X"77",X"77",X"77",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"06",X"06",
		X"60",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"70",X"00",X"00",X"00",X"00",X"7C",X"C7",X"7C",X"7C",X"70",X"00",X"07",
		X"CC",X"0C",X"CC",X"0C",X"77",X"00",X"77",X"C7",X"C7",X"C0",X"C0",X"CC",X"70",X"CC",X"C0",X"CC",
		X"C7",X"CC",X"0C",X"70",X"C7",X"C7",X"7C",X"0C",X"77",X"C7",X"C0",X"70",X"C7",X"77",X"C7",X"70",
		X"7C",X"70",X"0C",X"CA",X"AA",X"7A",X"AA",X"77",X"00",X"07",X"77",X"77",X"77",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"06",X"60",X"06",X"00",X"00",X"00",X"00",X"66",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",
		X"00",X"00",X"00",X"07",X"C0",X"00",X"00",X"00",X"00",X"7C",X"70",X"C7",X"C7",X"70",X"00",X"0C",
		X"70",X"C7",X"CC",X"C7",X"C7",X"00",X"7C",X"00",X"C7",X"0C",X"0C",X"07",X"70",X"7C",X"C7",X"7C",
		X"CC",X"7C",X"7C",X"C0",X"77",X"7C",X"C0",X"C0",X"C7",X"C7",X"70",X"77",X"00",X"CC",X"0C",X"07",
		X"C7",X"70",X"07",X"7C",X"77",X"CC",X"CC",X"77",X"00",X"00",X"C7",X"70",X"C7",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"00",X"60",X"06",X"00",X"00",X"00",X"00",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"66",X"06",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"C0",X"00",X"00",X"00",X"00",X"7C",X"70",X"C7",X"C7",X"70",X"00",X"0C",
		X"70",X"C7",X"CC",X"C7",X"C7",X"00",X"7C",X"00",X"C7",X"0C",X"0C",X"07",X"70",X"7C",X"C7",X"7C",
		X"CC",X"7C",X"7C",X"C0",X"77",X"7C",X"C0",X"C0",X"C7",X"C7",X"70",X"77",X"00",X"CC",X"0C",X"07",
		X"C7",X"70",X"07",X"7C",X"77",X"CC",X"CC",X"77",X"00",X"00",X"C7",X"70",X"C7",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"00",X"66",X"06",X"00",X"00",X"00",X"00",X"06",X"06",
		X"60",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"C0",X"00",X"00",X"00",X"00",X"7C",X"70",X"C7",X"C7",X"70",X"00",X"0C",
		X"70",X"C7",X"CC",X"C7",X"C7",X"00",X"7C",X"00",X"C7",X"0C",X"0C",X"07",X"70",X"7C",X"C7",X"7C",
		X"CC",X"7C",X"7C",X"C0",X"77",X"7C",X"C0",X"C0",X"C7",X"C7",X"70",X"77",X"00",X"CC",X"0C",X"07",
		X"C7",X"70",X"07",X"7C",X"77",X"CC",X"CC",X"77",X"00",X"00",X"C7",X"70",X"C7",X"77",X"70",X"00",
		X"00",X"00",X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"67",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"60",X"00",X"00",X"00",X"06",X"06",X"60",X"06",X"00",X"00",X"00",X"00",X"66",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"60",X"00",
		X"00",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"2F",X"C2",X"7E",X"31",X"99",X"7E",X"30",X"85",X"7E",X"34",X"E0",X"7E",X"26",X"FC",X"7E",
		X"26",X"F5",X"7E",X"34",X"AF",X"35",X"EB",X"35",X"AE",X"EE",X"02",X"08",X"11",X"01",X"20",X"17",
		X"00",X"F0",X"01",X"10",X"28",X"00",X"F0",X"01",X"10",X"25",X"00",X"E0",X"1D",X"04",X"0E",X"00",
		X"D0",X"01",X"08",X"01",X"00",X"86",X"02",X"20",X"05",X"7E",X"D0",X"63",X"86",X"01",X"10",X"8E",
		X"C3",X"B3",X"0D",X"59",X"2A",X"F3",X"F6",X"CC",X"05",X"C4",X"0F",X"C1",X"09",X"26",X"02",X"97",
		X"51",X"91",X"51",X"22",X"E4",X"97",X"40",X"0F",X"4F",X"0F",X"50",X"C6",X"08",X"BD",X"D0",X"BA",
		X"CE",X"D0",X"15",X"40",X"8B",X"9A",X"9B",X"51",X"19",X"97",X"51",X"8E",X"CD",X"00",X"BD",X"D0",
		X"AB",X"96",X"40",X"80",X"02",X"CC",X"26",X"E1",X"25",X"03",X"CC",X"26",X"E6",X"BD",X"D0",X"4B",
		X"4F",X"AB",X"C4",X"33",X"48",X"11",X"83",X"EA",X"B1",X"25",X"F6",X"A7",X"A9",X"FA",X"BF",X"86",
		X"7F",X"97",X"59",X"BD",X"D0",X"12",X"8E",X"BD",X"E4",X"6F",X"80",X"8C",X"BE",X"5C",X"26",X"F9",
		X"8E",X"CC",X"02",X"BD",X"D0",X"A2",X"BD",X"D0",X"C6",X"B7",X"BD",X"EC",X"86",X"01",X"97",X"3F",
		X"86",X"01",X"B7",X"BD",X"ED",X"97",X"48",X"8E",X"CC",X"00",X"BD",X"D0",X"A2",X"5F",X"44",X"56",
		X"44",X"56",X"44",X"56",X"44",X"56",X"DD",X"46",X"FD",X"BD",X"E9",X"BD",X"2B",X"7C",X"8E",X"BD",
		X"E4",X"A6",X"80",X"A7",X"88",X"3B",X"8C",X"BE",X"20",X"26",X"F6",X"96",X"40",X"4A",X"26",X"03",
		X"7F",X"BE",X"28",X"86",X"7F",X"97",X"59",X"BD",X"D0",X"45",X"6A",X"08",X"BD",X"D0",X"12",X"BD",
		X"D0",X"60",X"AE",X"9F",X"98",X"11",X"26",X"0B",X"BD",X"D0",X"36",X"BD",X"D0",X"54",X"27",X"C3",
		X"7E",X"D0",X"96",X"BD",X"D0",X"33",X"BD",X"5B",X"40",X"BD",X"D0",X"30",X"BD",X"2A",X"21",X"BD",
		X"D0",X"99",X"B6",X"C8",X"06",X"2A",X"08",X"96",X"3F",X"4A",X"27",X"03",X"BD",X"D0",X"9C",X"BD",
		X"34",X"AF",X"BD",X"D0",X"24",X"0F",X"F2",X"96",X"48",X"26",X"05",X"BD",X"34",X"C0",X"20",X"36",
		X"FC",X"BD",X"E5",X"26",X"0B",X"86",X"11",X"97",X"CF",X"86",X"71",X"BD",X"5F",X"96",X"20",X"03",
		X"BD",X"34",X"C0",X"0F",X"48",X"96",X"40",X"4A",X"27",X"1C",X"96",X"90",X"97",X"CF",X"D6",X"3F",
		X"86",X"67",X"BD",X"5F",X"99",X"86",X"73",X"8E",X"28",X"1D",X"7E",X"D0",X"66",X"0F",X"CF",X"D6",
		X"3F",X"86",X"67",X"BD",X"5F",X"99",X"BD",X"2B",X"0B",X"BD",X"2F",X"8C",X"0F",X"06",X"7F",X"C0",
		X"06",X"BD",X"00",X"00",X"BD",X"1A",X"C0",X"BD",X"4B",X"00",X"BD",X"00",X"03",X"BD",X"38",X"83",
		X"BD",X"38",X"80",X"BD",X"29",X"A4",X"86",X"08",X"97",X"92",X"BD",X"D0",X"54",X"35",X"4B",X"BD",
		X"29",X"8F",X"BD",X"D0",X"33",X"BD",X"11",X"40",X"BD",X"4B",X"03",X"86",X"19",X"97",X"59",X"B6",
		X"BE",X"6E",X"27",X"0D",X"BD",X"D0",X"54",X"41",X"40",X"86",X"96",X"8E",X"28",X"74",X"7E",X"D0",
		X"66",X"7E",X"28",X"FE",X"BD",X"29",X"F5",X"BD",X"29",X"8F",X"86",X"06",X"8E",X"28",X"82",X"7E",
		X"D0",X"66",X"BD",X"29",X"D2",X"86",X"04",X"8E",X"28",X"8D",X"7E",X"D0",X"66",X"BD",X"29",X"83",
		X"BD",X"D0",X"54",X"31",X"B5",X"BD",X"D0",X"54",X"30",X"B3",X"0F",X"59",X"86",X"0C",X"8E",X"28",
		X"A4",X"7E",X"D0",X"66",X"BD",X"29",X"83",X"BD",X"29",X"8F",X"86",X"0A",X"8E",X"28",X"B2",X"7E",
		X"D0",X"66",X"BD",X"29",X"83",X"BD",X"29",X"8F",X"86",X"04",X"97",X"92",X"0F",X"CF",X"86",X"71",
		X"BD",X"5F",X"96",X"BD",X"34",X"C0",X"8E",X"20",X"FB",X"CE",X"2C",X"03",X"A6",X"C0",X"88",X"5A",
		X"27",X"05",X"BD",X"5F",X"90",X"20",X"F5",X"7E",X"2A",X"85",X"20",X"28",X"43",X"29",X"20",X"31",
		X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"DE",X"15",
		X"6F",X"47",X"8E",X"98",X"21",X"AF",X"49",X"9E",X"21",X"AF",X"4B",X"AF",X"4D",X"86",X"01",X"34",
		X"02",X"AE",X"49",X"AE",X"84",X"27",X"15",X"BD",X"29",X"B5",X"A6",X"47",X"84",X"03",X"81",X"03",
		X"26",X"05",X"BD",X"5B",X"58",X"20",X"03",X"BD",X"5B",X"46",X"AF",X"49",X"6C",X"47",X"A6",X"47",
		X"81",X"20",X"23",X"0D",X"10",X"AE",X"4D",X"27",X"18",X"10",X"AE",X"A4",X"27",X"13",X"10",X"AF",
		X"4D",X"6A",X"E4",X"26",X"CC",X"35",X"02",X"8D",X"1C",X"86",X"01",X"8E",X"29",X"0D",X"7E",X"D0",
		X"66",X"35",X"02",X"86",X"02",X"8E",X"29",X"5B",X"7E",X"D0",X"66",X"8D",X"26",X"86",X"0A",X"8E",
		X"28",X"74",X"7E",X"D0",X"66",X"34",X"10",X"86",X"04",X"97",X"2B",X"AE",X"4B",X"AC",X"4D",X"26",
		X"05",X"8E",X"98",X"21",X"20",X"03",X"BD",X"D0",X"18",X"AE",X"84",X"0A",X"2B",X"26",X"EE",X"AF",
		X"4B",X"35",X"90",X"9E",X"21",X"27",X"07",X"BD",X"D0",X"18",X"AE",X"84",X"26",X"F9",X"39",X"9E",
		X"23",X"27",X"0C",X"96",X"90",X"BD",X"38",X"88",X"AF",X"98",X"06",X"AE",X"84",X"26",X"F4",X"39",
		X"9E",X"23",X"20",X"02",X"9E",X"21",X"27",X"0C",X"EC",X"04",X"10",X"AE",X"02",X"BD",X"D0",X"1E",
		X"AE",X"84",X"26",X"F4",X"39",X"34",X"46",X"EE",X"02",X"E6",X"C4",X"A6",X"04",X"48",X"24",X"02",
		X"86",X"FF",X"3D",X"AB",X"04",X"97",X"A6",X"E6",X"41",X"A6",X"05",X"3D",X"AB",X"05",X"97",X"A7",
		X"35",X"C6",X"8E",X"98",X"5A",X"10",X"AE",X"02",X"A6",X"21",X"34",X"02",X"A6",X"E4",X"9B",X"5F",
		X"4A",X"97",X"A7",X"4F",X"BD",X"46",X"86",X"43",X"BD",X"46",X"86",X"A6",X"E4",X"80",X"03",X"A7",
		X"E4",X"2A",X"E9",X"35",X"82",X"8E",X"98",X"5A",X"10",X"AE",X"02",X"A6",X"21",X"34",X"02",X"A6",
		X"E4",X"9B",X"5F",X"4A",X"97",X"A7",X"BD",X"5B",X"46",X"6A",X"E4",X"26",X"F2",X"A6",X"A4",X"A7",
		X"E4",X"A6",X"E4",X"9B",X"5E",X"4A",X"97",X"A6",X"BD",X"5B",X"58",X"6A",X"E4",X"26",X"F2",X"35",
		X"82",X"BD",X"D0",X"45",X"CE",X"2A",X"4B",X"A6",X"09",X"4A",X"81",X"09",X"23",X"04",X"80",X"0A",
		X"20",X"F8",X"33",X"C6",X"A6",X"C4",X"97",X"8F",X"A6",X"4A",X"97",X"90",X"E6",X"C8",X"14",X"BE",
		X"38",X"86",X"3A",X"9F",X"93",X"A6",X"C8",X"1E",X"97",X"91",X"39",X"22",X"55",X"11",X"EE",X"77",
		X"33",X"44",X"88",X"00",X"CC",X"FF",X"EE",X"BB",X"DD",X"EE",X"FF",X"11",X"BB",X"DD",X"AA",X"00",
		X"10",X"20",X"30",X"40",X"50",X"70",X"80",X"00",X"60",X"99",X"00",X"99",X"66",X"99",X"99",X"99",
		X"11",X"AA",X"99",X"B6",X"BE",X"68",X"BB",X"BE",X"6F",X"9B",X"ED",X"BB",X"BE",X"6E",X"BB",X"BE",
		X"71",X"BB",X"BE",X"70",X"39",X"DE",X"15",X"86",X"12",X"A7",X"47",X"0F",X"F0",X"8D",X"E4",X"26",
		X"24",X"BD",X"D0",X"45",X"6C",X"09",X"26",X"02",X"6C",X"09",X"6C",X"08",X"CC",X"26",X"EB",X"BD",
		X"D0",X"4B",X"BD",X"2B",X"7C",X"BD",X"D0",X"60",X"86",X"7F",X"97",X"59",X"BD",X"D0",X"12",X"BD",
		X"57",X"00",X"7E",X"27",X"A3",X"B6",X"C8",X"04",X"81",X"58",X"26",X"03",X"BD",X"D0",X"69",X"6A",
		X"47",X"26",X"31",X"86",X"0F",X"A7",X"47",X"B6",X"BE",X"68",X"81",X"1E",X"24",X"26",X"CC",X"FF",
		X"FE",X"0D",X"F0",X"26",X"03",X"CC",X"FE",X"FC",X"BB",X"BE",X"5D",X"0F",X"F0",X"81",X"01",X"2C",
		X"02",X"86",X"01",X"B7",X"BE",X"5D",X"FB",X"BE",X"5C",X"F1",X"BE",X"5D",X"2C",X"03",X"F6",X"BE",
		X"5D",X"F7",X"BE",X"5C",X"96",X"EE",X"4C",X"81",X"96",X"25",X"06",X"C6",X"06",X"BD",X"D0",X"BD",
		X"4F",X"97",X"EE",X"86",X"0F",X"8E",X"2A",X"8D",X"7E",X"D0",X"66",X"BD",X"D0",X"45",X"30",X"0A",
		X"CE",X"BE",X"5C",X"A6",X"80",X"A7",X"C0",X"11",X"83",X"BE",X"72",X"26",X"F6",X"BD",X"D0",X"45",
		X"A6",X"09",X"81",X"04",X"22",X"32",X"E6",X"08",X"DD",X"2B",X"5D",X"27",X"12",X"81",X"02",X"22",
		X"27",X"8E",X"CC",X"02",X"BD",X"D0",X"A2",X"BD",X"D0",X"C6",X"4A",X"91",X"2C",X"23",X"19",X"96",
		X"2B",X"8E",X"2B",X"55",X"48",X"48",X"30",X"86",X"EC",X"81",X"B7",X"BE",X"60",X"F7",X"BE",X"5F",
		X"EC",X"84",X"B7",X"BE",X"5C",X"F7",X"BE",X"5D",X"39",X"26",X"60",X"1E",X"0F",X"26",X"60",X"19",
		X"0C",X"24",X"30",X"14",X"0A",X"1E",X"1E",X"0F",X"07",X"BD",X"D0",X"45",X"30",X"0A",X"CE",X"BE",
		X"5C",X"A6",X"C0",X"A7",X"80",X"11",X"83",X"BE",X"72",X"26",X"F6",X"39",X"8E",X"CC",X"14",X"BD",
		X"D0",X"A5",X"BD",X"D0",X"B4",X"BD",X"D0",X"45",X"C1",X"05",X"24",X"14",X"A6",X"09",X"81",X"0E",
		X"25",X"02",X"C6",X"05",X"81",X"05",X"25",X"08",X"A6",X"08",X"81",X"03",X"25",X"02",X"C6",X"05",
		X"C0",X"05",X"D7",X"2C",X"2A",X"01",X"50",X"D7",X"2B",X"E6",X"09",X"CE",X"2C",X"22",X"30",X"0A",
		X"C1",X"28",X"23",X"04",X"C0",X"14",X"20",X"F8",X"11",X"83",X"2E",X"24",X"25",X"06",X"33",X"5D",
		X"A6",X"C5",X"20",X"31",X"A6",X"C5",X"34",X"06",X"E6",X"5E",X"C4",X"1F",X"96",X"2B",X"3D",X"35",
		X"02",X"3D",X"89",X"00",X"D6",X"2C",X"E8",X"5E",X"35",X"04",X"2A",X"09",X"40",X"27",X"06",X"AB",
		X"C5",X"25",X"06",X"20",X"08",X"AB",X"C5",X"25",X"0A",X"A1",X"5F",X"24",X"02",X"A6",X"5F",X"A1",
		X"C4",X"23",X"02",X"A6",X"C4",X"A7",X"80",X"33",X"C8",X"2B",X"11",X"83",X"2F",X"8B",X"25",X"B8",
		X"6F",X"80",X"39",X"01",X"19",X"06",X"7A",X"6B",X"63",X"62",X"68",X"7A",X"0D",X"13",X"16",X"16",
		X"13",X"1B",X"17",X"09",X"7A",X"1F",X"16",X"1F",X"19",X"67",X"7A",X"13",X"14",X"19",X"67",X"5A",
		X"8E",X"0A",X"14",X"14",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"0D",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",X"0C",X"8E",X"03",X"0A",X"09",X"07",
		X"06",X"05",X"05",X"05",X"05",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"03",X"04",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"04",X"03",X"0E",X"08",X"0C",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0B",X"8E",X"0D",X"28",X"1E",X"1C",X"1A",X"18",X"16",X"14",X"12",X"12",X"10",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"8E",X"0C",X"28",X"1E",
		X"1C",X"1A",X"18",X"1E",X"14",X"12",X"10",X"12",X"19",X"0C",X"0C",X"0C",X"19",X"19",X"0C",X"0C",
		X"0C",X"12",X"14",X"0E",X"0E",X"0E",X"0E",X"0E",X"19",X"0E",X"0E",X"12",X"19",X"0C",X"0C",X"0C",
		X"0C",X"19",X"0C",X"0C",X"0C",X"12",X"14",X"8E",X"05",X"09",X"08",X"08",X"07",X"07",X"07",X"07",
		X"07",X"06",X"06",X"06",X"06",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",
		X"05",X"05",X"8E",X"19",X"50",X"40",X"40",X"40",X"40",X"40",X"28",X"28",X"26",X"26",X"26",X"26",
		X"26",X"26",X"26",X"26",X"26",X"24",X"24",X"24",X"24",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"8E",X"06",X"0A",
		X"08",X"08",X"08",X"08",X"08",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"8E",X"14",X"28",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1E",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"1C",X"1C",X"1C",X"1C",X"1C",X"1A",X"1A",X"1A",X"1A",X"1A",X"18",
		X"18",X"18",X"18",X"0E",X"A0",X"FF",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",
		X"B8",X"B8",X"B8",X"B8",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"8E",X"0C",
		X"30",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"28",X"44",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"3C",X"3C",X"3C",X"3C",X"0F",X"11",X"16",X"22",X"14",X"20",X"00",X"23",X"3C",X"19",X"23",X"00",
		X"23",X"1B",X"19",X"23",X"00",X"23",X"46",X"19",X"23",X"00",X"23",X"00",X"19",X"23",X"00",X"23",
		X"4B",X"19",X"23",X"00",X"23",X"1E",X"1B",X"23",X"00",X"23",X"50",X"1E",X"05",X"0F",X"19",X"19",
		X"14",X"19",X"00",X"19",X"00",X"14",X"19",X"00",X"19",X"05",X"14",X"19",X"00",X"19",X"00",X"14",
		X"19",X"00",X"19",X"00",X"14",X"19",X"00",X"19",X"00",X"14",X"19",X"00",X"19",X"00",X"0F",X"19",
		X"00",X"19",X"00",X"0F",X"01",X"01",X"02",X"02",X"0F",X"03",X"04",X"03",X"03",X"00",X"03",X"03",
		X"03",X"05",X"00",X"03",X"03",X"03",X"03",X"08",X"03",X"03",X"03",X"03",X"19",X"03",X"03",X"03",
		X"03",X"00",X"03",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"03",X"0A",X"01",X"01",X"02",X"02",
		X"00",X"03",X"04",X"03",X"03",X"16",X"03",X"03",X"03",X"05",X"00",X"03",X"03",X"03",X"03",X"08",
		X"03",X"03",X"03",X"03",X"00",X"03",X"03",X"03",X"03",X"19",X"03",X"03",X"03",X"03",X"00",X"03",
		X"03",X"03",X"03",X"0A",X"00",X"01",X"02",X"02",X"01",X"03",X"04",X"03",X"03",X"00",X"03",X"03",
		X"03",X"05",X"16",X"03",X"03",X"03",X"03",X"08",X"03",X"03",X"03",X"03",X"01",X"03",X"03",X"03",
		X"03",X"00",X"03",X"03",X"03",X"03",X"19",X"03",X"03",X"03",X"03",X"0A",X"00",X"05",X"06",X"07",
		X"00",X"07",X"0C",X"08",X"04",X"00",X"08",X"0D",X"08",X"14",X"02",X"03",X"0E",X"08",X"03",X"02",
		X"08",X"0F",X"08",X"0D",X"01",X"08",X"10",X"08",X"04",X"01",X"08",X"10",X"08",X"19",X"02",X"08",
		X"10",X"08",X"06",X"02",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"14",X"00",X"00",
		X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"00",X"16",X"00",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"00",X"19",X"00",X"01",X"03",X"04",
		X"01",X"04",X"00",X"05",X"05",X"01",X"05",X"00",X"05",X"02",X"01",X"05",X"00",X"05",X"05",X"02",
		X"05",X"00",X"05",X"06",X"01",X"05",X"00",X"05",X"05",X"01",X"05",X"00",X"05",X"02",X"01",X"05",
		X"00",X"05",X"05",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"0C",X"00",X"07",X"00",X"00",X"0C",X"01",
		X"01",X"01",X"01",X"0D",X"01",X"02",X"02",X"02",X"0E",X"02",X"01",X"01",X"8E",X"98",X"5A",X"CC",
		X"36",X"03",X"ED",X"02",X"ED",X"88",X"14",X"0F",X"70",X"0F",X"71",X"CC",X"30",X"7B",X"DD",X"72",
		X"CC",X"4A",X"7C",X"ED",X"04",X"A7",X"0A",X"6F",X"0B",X"E7",X"0C",X"6F",X"0D",X"0F",X"87",X"0F",
		X"48",X"0F",X"8D",X"0F",X"8E",X"0F",X"8A",X"0F",X"95",X"0F",X"ED",X"86",X"02",X"97",X"EF",X"0F",
		X"F1",X"39",X"96",X"59",X"85",X"01",X"27",X"01",X"39",X"4D",X"2A",X"04",X"96",X"52",X"20",X"03",
		X"B6",X"C8",X"04",X"8E",X"98",X"5A",X"CE",X"30",X"31",X"84",X"0F",X"48",X"48",X"33",X"C6",X"EC",
		X"C4",X"DB",X"66",X"C1",X"18",X"25",X"06",X"C1",X"DF",X"22",X"02",X"D7",X"66",X"5F",X"47",X"56",
		X"D3",X"64",X"81",X"07",X"25",X"06",X"81",X"8C",X"22",X"02",X"DD",X"64",X"EC",X"42",X"27",X"30",
		X"10",X"93",X"72",X"27",X"06",X"DD",X"72",X"0F",X"71",X"0F",X"70",X"D6",X"70",X"26",X"17",X"DE",
		X"72",X"96",X"71",X"E6",X"C6",X"26",X"04",X"0F",X"71",X"E6",X"C4",X"0C",X"71",X"5A",X"58",X"58",
		X"4F",X"C3",X"35",X"EB",X"DD",X"5C",X"96",X"70",X"4C",X"81",X"02",X"25",X"01",X"4F",X"97",X"70",
		X"39",X"00",X"00",X"00",X"00",X"00",X"FF",X"30",X"80",X"00",X"01",X"30",X"7B",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"30",X"71",X"FF",X"FF",X"30",X"71",X"FF",X"01",X"30",X"71",X"00",X"00",X"00",
		X"00",X"01",X"00",X"30",X"76",X"01",X"FF",X"30",X"76",X"01",X"01",X"30",X"76",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"02",X"01",X"03",X"00",X"04",X"05",X"04",X"06",X"00",X"07",X"08",X"07",X"09",X"00",
		X"0A",X"0B",X"0A",X"0C",X"00",X"34",X"46",X"34",X"06",X"E3",X"98",X"02",X"34",X"06",X"20",X"1B",
		X"EC",X"44",X"A1",X"E4",X"24",X"15",X"E1",X"61",X"24",X"11",X"E3",X"D8",X"02",X"A1",X"62",X"23",
		X"0A",X"E1",X"63",X"23",X"06",X"34",X"40",X"AC",X"E1",X"26",X"04",X"EE",X"C4",X"26",X"E1",X"32",
		X"64",X"35",X"C6",X"86",X"01",X"97",X"48",X"DC",X"5E",X"DE",X"6E",X"8E",X"98",X"21",X"BD",X"D0",
		X"27",X"26",X"2C",X"DC",X"5E",X"DE",X"6E",X"8E",X"98",X"23",X"BD",X"D0",X"27",X"26",X"20",X"DC",
		X"5E",X"DE",X"6E",X"8E",X"98",X"17",X"BD",X"D0",X"27",X"26",X"14",X"DC",X"5E",X"DE",X"6E",X"8E",
		X"98",X"1F",X"BD",X"D0",X"27",X"0F",X"48",X"86",X"01",X"8E",X"30",X"B3",X"7E",X"D0",X"66",X"CC",
		X"26",X"D9",X"BD",X"D0",X"4B",X"86",X"1B",X"97",X"59",X"BD",X"D0",X"60",X"C6",X"07",X"BD",X"D0",
		X"BD",X"BD",X"D0",X"24",X"BD",X"5B",X"4C",X"BD",X"D0",X"45",X"B6",X"BD",X"EC",X"BA",X"BE",X"28",
		X"26",X"1E",X"86",X"FF",X"97",X"59",X"CC",X"1C",X"0A",X"8E",X"3C",X"7E",X"BD",X"D0",X"1B",X"86",
		X"28",X"C6",X"AA",X"D7",X"CF",X"BD",X"5F",X"99",X"86",X"78",X"8E",X"E3",X"D3",X"7E",X"D0",X"66",
		X"BD",X"D0",X"45",X"A6",X"0B",X"B7",X"BE",X"5D",X"B1",X"BE",X"5C",X"23",X"03",X"B7",X"BE",X"5C",
		X"4F",X"D6",X"ED",X"27",X"1E",X"C0",X"04",X"2B",X"03",X"4C",X"20",X"F9",X"4D",X"26",X"06",X"7D",
		X"BE",X"6F",X"26",X"01",X"4C",X"BB",X"BE",X"6F",X"A1",X"88",X"1D",X"23",X"03",X"A6",X"88",X"1D",
		X"B7",X"BE",X"6F",X"BD",X"2B",X"69",X"BD",X"D0",X"45",X"E6",X"08",X"26",X"1C",X"CC",X"1C",X"20",
		X"8E",X"3C",X"77",X"BD",X"D0",X"1B",X"86",X"4B",X"C6",X"AA",X"D7",X"CF",X"D6",X"3F",X"BD",X"5F",
		X"99",X"86",X"60",X"8E",X"31",X"89",X"7E",X"D0",X"66",X"96",X"3F",X"88",X"03",X"BD",X"D0",X"48",
		X"E6",X"08",X"27",X"F7",X"97",X"3F",X"7E",X"27",X"A3",X"EC",X"98",X"02",X"34",X"06",X"86",X"88",
		X"A0",X"E0",X"BD",X"D0",X"42",X"8B",X"06",X"1F",X"89",X"86",X"D2",X"A0",X"E0",X"BD",X"D0",X"42",
		X"8B",X"17",X"1E",X"89",X"39",X"6F",X"47",X"6F",X"48",X"96",X"59",X"2A",X"04",X"DC",X"52",X"20",
		X"06",X"B6",X"C8",X"04",X"F6",X"C8",X"06",X"54",X"46",X"54",X"46",X"84",X"F0",X"E6",X"47",X"A7",
		X"47",X"E1",X"47",X"26",X"54",X"6C",X"48",X"E6",X"48",X"C1",X"02",X"27",X"04",X"C4",X"07",X"26",
		X"4E",X"D6",X"87",X"C1",X"04",X"24",X"46",X"0D",X"13",X"27",X"44",X"44",X"44",X"34",X"02",X"44",
		X"AB",X"E0",X"10",X"8E",X"32",X"37",X"31",X"A6",X"81",X"42",X"24",X"33",X"AE",X"A4",X"27",X"2F",
		X"4F",X"BD",X"D0",X"57",X"1F",X"13",X"BD",X"D0",X"51",X"AF",X"47",X"EC",X"24",X"C3",X"35",X"AE",
		X"ED",X"02",X"ED",X"88",X"14",X"DC",X"5E",X"AB",X"22",X"A7",X"0A",X"EB",X"23",X"E7",X"0C",X"0C",
		X"87",X"CC",X"26",X"F0",X"BD",X"D0",X"4B",X"20",X"06",X"6F",X"48",X"20",X"02",X"6A",X"48",X"86",
		X"01",X"8E",X"31",X"B9",X"7E",X"D0",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"AD",X"02",
		X"FF",X"00",X"04",X"32",X"C7",X"02",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"32",
		X"93",X"00",X"04",X"00",X"00",X"33",X"FF",X"00",X"00",X"00",X"0C",X"33",X"DC",X"00",X"04",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"32",X"79",X"02",X"04",X"00",X"00",X"34",X"22",X"02",
		X"00",X"00",X"08",X"34",X"45",X"02",X"04",X"00",X"0C",X"AE",X"47",X"A6",X"0A",X"8B",X"03",X"81",
		X"8D",X"22",X"5E",X"A7",X"0A",X"CC",X"01",X"00",X"BD",X"34",X"6B",X"86",X"01",X"8E",X"32",X"79",
		X"7E",X"D0",X"66",X"AE",X"47",X"A6",X"0A",X"80",X"03",X"81",X"07",X"25",X"48",X"A7",X"0A",X"CC",
		X"FF",X"00",X"BD",X"34",X"6B",X"86",X"01",X"8E",X"32",X"93",X"7E",X"D0",X"66",X"AE",X"47",X"A6",
		X"0C",X"8B",X"FA",X"81",X"18",X"25",X"34",X"A7",X"0C",X"CC",X"00",X"FF",X"BD",X"34",X"6B",X"86",
		X"01",X"8E",X"32",X"AD",X"7E",X"D0",X"66",X"AE",X"47",X"A6",X"0C",X"8B",X"06",X"81",X"E5",X"22",
		X"1E",X"A7",X"0C",X"CC",X"00",X"01",X"BD",X"34",X"6B",X"86",X"01",X"8E",X"32",X"C7",X"7E",X"D0",
		X"66",X"86",X"90",X"20",X"02",X"86",X"06",X"E6",X"0C",X"20",X"0A",X"C6",X"17",X"20",X"02",X"C6",
		X"EB",X"A6",X"0A",X"20",X"2F",X"ED",X"49",X"BD",X"34",X"A3",X"AE",X"49",X"96",X"91",X"D6",X"91",
		X"ED",X"1F",X"A7",X"01",X"86",X"02",X"8E",X"33",X"0C",X"7E",X"D0",X"66",X"96",X"8F",X"AE",X"49",
		X"A7",X"1F",X"A7",X"01",X"86",X"01",X"8E",X"33",X"1C",X"7E",X"D0",X"66",X"96",X"8F",X"A7",X"D8",
		X"09",X"7E",X"D0",X"63",X"C1",X"EA",X"24",X"02",X"C6",X"16",X"81",X"06",X"22",X"01",X"4C",X"ED",
		X"49",X"BD",X"34",X"A3",X"96",X"91",X"D6",X"91",X"AE",X"49",X"ED",X"84",X"96",X"8F",X"84",X"F0",
		X"34",X"02",X"96",X"91",X"84",X"0F",X"AB",X"E0",X"1F",X"89",X"ED",X"89",X"FF",X"00",X"86",X"02",
		X"8E",X"33",X"56",X"7E",X"D0",X"66",X"AE",X"49",X"96",X"8F",X"D6",X"8F",X"ED",X"89",X"FF",X"00",
		X"84",X"0F",X"C4",X"0F",X"34",X"06",X"96",X"91",X"D6",X"91",X"84",X"F0",X"C4",X"F0",X"E3",X"E1",
		X"ED",X"84",X"86",X"01",X"8E",X"33",X"7A",X"7E",X"D0",X"66",X"96",X"8F",X"D6",X"8F",X"ED",X"D8",
		X"09",X"7E",X"D0",X"63",X"7E",X"32",X"F5",X"20",X"9B",X"D7",X"2C",X"5F",X"47",X"56",X"DD",X"2D",
		X"1F",X"20",X"AB",X"0A",X"EB",X"0C",X"A7",X"0A",X"E7",X"0C",X"DC",X"2D",X"E3",X"0A",X"ED",X"0A",
		X"E6",X"0C",X"DB",X"2C",X"E7",X"0C",X"C1",X"EA",X"22",X"DD",X"C1",X"18",X"25",X"D9",X"81",X"8F",
		X"22",X"D2",X"81",X"07",X"25",X"CE",X"20",X"E2",X"10",X"8E",X"00",X"05",X"CC",X"FF",X"01",X"20",
		X"C8",X"10",X"8E",X"00",X"00",X"CC",X"FF",X"FF",X"20",X"BF",X"10",X"8E",X"02",X"00",X"CC",X"01",
		X"FF",X"20",X"B6",X"10",X"8E",X"02",X"05",X"CC",X"01",X"01",X"20",X"AD",X"AE",X"47",X"A6",X"0A",
		X"80",X"03",X"E6",X"0C",X"CB",X"06",X"81",X"07",X"25",X"CE",X"C1",X"E5",X"22",X"CA",X"A7",X"0A",
		X"E7",X"0C",X"CC",X"FF",X"01",X"8D",X"74",X"86",X"01",X"8E",X"33",X"DC",X"7E",X"D0",X"66",X"AE",
		X"47",X"A6",X"0A",X"80",X"03",X"81",X"07",X"25",X"B8",X"E6",X"0C",X"C0",X"06",X"C1",X"18",X"25",
		X"B0",X"A7",X"0A",X"E7",X"0C",X"CC",X"FF",X"FF",X"8D",X"51",X"86",X"01",X"8E",X"33",X"FF",X"7E",
		X"D0",X"66",X"AE",X"47",X"A6",X"0A",X"8B",X"03",X"81",X"8D",X"22",X"9E",X"E6",X"0C",X"C0",X"06",
		X"C1",X"18",X"25",X"96",X"A7",X"0A",X"E7",X"0C",X"CC",X"01",X"FF",X"8D",X"2E",X"86",X"01",X"8E",
		X"34",X"22",X"7E",X"D0",X"66",X"AE",X"47",X"A6",X"0A",X"8B",X"03",X"81",X"8D",X"22",X"84",X"E6",
		X"0C",X"CB",X"06",X"C1",X"E5",X"23",X"03",X"7E",X"33",X"D3",X"A7",X"0A",X"E7",X"0C",X"CC",X"01",
		X"01",X"8D",X"08",X"86",X"01",X"8E",X"34",X"45",X"7E",X"D0",X"66",X"DD",X"88",X"BD",X"D0",X"8D",
		X"34",X"50",X"EE",X"02",X"EC",X"04",X"8E",X"98",X"23",X"BD",X"D0",X"27",X"26",X"1E",X"AE",X"E4",
		X"EE",X"02",X"EC",X"04",X"8E",X"98",X"21",X"BD",X"D0",X"27",X"26",X"10",X"AE",X"E4",X"EE",X"02",
		X"EC",X"04",X"8E",X"98",X"17",X"BD",X"D0",X"27",X"26",X"02",X"35",X"D0",X"35",X"50",X"8D",X"03",
		X"7E",X"D0",X"63",X"BD",X"D0",X"15",X"DC",X"1B",X"ED",X"84",X"9F",X"1B",X"0A",X"87",X"39",X"34",
		X"76",X"96",X"40",X"BD",X"D0",X"0F",X"4A",X"26",X"FA",X"8D",X"6B",X"BD",X"26",X"C9",X"35",X"F6",
		X"B6",X"BD",X"ED",X"BD",X"D0",X"2A",X"1F",X"89",X"86",X"68",X"BD",X"5F",X"96",X"96",X"40",X"4A",
		X"27",X"0D",X"B6",X"BE",X"29",X"BD",X"D0",X"2A",X"1F",X"89",X"86",X"72",X"BD",X"5F",X"96",X"39",
		X"8E",X"2E",X"0E",X"CC",X"15",X"08",X"BD",X"D0",X"1B",X"8E",X"6E",X"0E",X"BD",X"D0",X"1B",X"10",
		X"8E",X"35",X"92",X"B6",X"BD",X"EC",X"27",X"14",X"81",X"07",X"23",X"02",X"86",X"07",X"97",X"2B",
		X"CC",X"2E",X"0E",X"BD",X"D0",X"21",X"8B",X"04",X"0A",X"2B",X"26",X"F7",X"B6",X"BE",X"28",X"27",
		X"14",X"81",X"07",X"23",X"02",X"86",X"07",X"97",X"2B",X"CC",X"6E",X"0E",X"BD",X"D0",X"21",X"8B",
		X"04",X"0A",X"2B",X"26",X"F7",X"39",X"8E",X"06",X"16",X"96",X"8F",X"A7",X"89",X"8A",X"00",X"A7",
		X"80",X"8C",X"06",X"EC",X"23",X"F5",X"8E",X"07",X"16",X"D6",X"8F",X"ED",X"84",X"ED",X"89",X"00",
		X"D5",X"30",X"89",X"01",X"00",X"8C",X"8F",X"16",X"23",X"F1",X"39",X"DE",X"27",X"11",X"83",X"B3",
		X"E4",X"25",X"03",X"CE",X"B3",X"A4",X"96",X"92",X"34",X"02",X"10",X"9E",X"93",X"AE",X"C1",X"27",
		X"21",X"EC",X"A4",X"88",X"04",X"C8",X"04",X"1A",X"10",X"FD",X"CA",X"06",X"D6",X"90",X"F7",X"CA",
		X"01",X"EC",X"22",X"FD",X"CA",X"02",X"EC",X"04",X"FD",X"CA",X"04",X"C6",X"1A",X"F7",X"CA",X"00",
		X"1C",X"EF",X"6A",X"E4",X"26",X"D7",X"32",X"61",X"DF",X"27",X"86",X"02",X"8E",X"35",X"4B",X"7E",
		X"D0",X"66",X"03",X"08",X"35",X"96",X"02",X"22",X"00",X"BB",X"0B",X"B0",X"BB",X"0B",X"B0",X"00",
		X"20",X"00",X"88",X"08",X"80",X"30",X"80",X"30",X"08",X"08",X"00",X"88",X"08",X"80",X"03",X"01",
		X"35",X"BE",X"01",X"06",X"35",X"C1",X"03",X"06",X"35",X"C7",X"03",X"06",X"35",X"D9",X"AA",X"AA",
		X"AA",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"00",X"00",X"0A",X"00",X"00",X"A0",X"00",X"0A",X"00",
		X"00",X"A0",X"00",X"0A",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"04",X"0C",X"36",X"1B",X"04",
		X"0C",X"36",X"4B",X"04",X"0C",X"36",X"7B",X"04",X"0C",X"36",X"AB",X"04",X"0C",X"36",X"DB",X"04",
		X"0C",X"37",X"0B",X"04",X"0C",X"37",X"3B",X"04",X"0C",X"37",X"6B",X"04",X"0C",X"37",X"9B",X"04",
		X"0C",X"37",X"CB",X"04",X"0C",X"37",X"FB",X"04",X"0C",X"38",X"2B",X"0B",X"22",X"20",X"00",X"0B",
		X"BB",X"BB",X"00",X"0B",X"22",X"2B",X"00",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"93",X"90",X"00",X"00",X"93",X"90",X"00",X"00",X"03",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"22",X"20",X"00",X"0B",
		X"BB",X"BB",X"00",X"0B",X"22",X"2B",X"00",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"90",X"00",X"03",X"33",X"93",X"00",X"00",X"09",X"93",X"00",X"00",X"90",X"93",X"00",X"00",
		X"90",X"90",X"00",X"09",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"0B",X"22",X"20",X"00",X"0B",
		X"BB",X"BB",X"00",X"0B",X"22",X"2B",X"00",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"90",X"00",X"03",X"39",X"93",X"00",X"00",X"09",X"93",X"00",X"00",X"90",X"93",X"00",X"00",
		X"90",X"90",X"00",X"09",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"B0",X"00",X"BB",
		X"BB",X"B0",X"00",X"B2",X"22",X"B0",X"00",X"02",X"22",X"00",X"00",X"00",X"90",X"00",X"00",X"09",
		X"99",X"00",X"00",X"09",X"39",X"00",X"00",X"09",X"39",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"B0",X"00",X"BB",
		X"BB",X"B0",X"00",X"B2",X"22",X"B0",X"00",X"02",X"22",X"00",X"00",X"00",X"90",X"00",X"00",X"09",
		X"90",X"00",X"00",X"39",X"93",X"30",X"00",X"39",X"90",X"00",X"00",X"39",X"09",X"00",X"00",X"09",
		X"09",X"00",X"00",X"09",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"02",X"22",X"B0",X"00",X"BB",
		X"BB",X"B0",X"00",X"B2",X"22",X"B0",X"00",X"02",X"22",X"00",X"00",X"00",X"90",X"00",X"00",X"09",
		X"90",X"00",X"00",X"39",X"33",X"30",X"00",X"39",X"90",X"00",X"00",X"39",X"09",X"00",X"00",X"09",
		X"09",X"00",X"00",X"09",X"09",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"BB",
		X"B2",X"BB",X"B0",X"B0",X"B0",X"B0",X"B0",X"0B",X"22",X"2B",X"00",X"00",X"09",X"00",X"00",X"09",
		X"93",X"99",X"00",X"39",X"93",X"99",X"30",X"30",X"93",X"90",X"30",X"30",X"90",X"90",X"30",X"00",
		X"90",X"90",X"00",X"09",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"BB",
		X"B2",X"BB",X"B0",X"B0",X"B0",X"B0",X"B0",X"0B",X"22",X"2B",X"00",X"00",X"09",X"00",X"00",X"09",
		X"93",X"99",X"00",X"39",X"93",X"99",X"30",X"30",X"93",X"90",X"30",X"30",X"90",X"90",X"00",X"09",
		X"90",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"22",X"20",X"00",X"BB",
		X"B2",X"BB",X"B0",X"B0",X"B0",X"B0",X"B0",X"0B",X"22",X"2B",X"00",X"00",X"09",X"00",X"00",X"09",
		X"93",X"99",X"00",X"39",X"93",X"99",X"30",X"30",X"93",X"90",X"30",X"00",X"90",X"90",X"30",X"00",
		X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"BB",X"22",X"2B",X"B0",X"B2",
		X"22",X"22",X"B0",X"B2",X"22",X"22",X"B0",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"09",
		X"99",X"99",X"00",X"39",X"99",X"99",X"30",X"30",X"99",X"90",X"30",X"30",X"90",X"90",X"30",X"00",
		X"90",X"90",X"00",X"09",X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"BB",X"22",X"2B",X"B0",X"B2",
		X"22",X"22",X"B0",X"B2",X"22",X"22",X"B0",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"09",
		X"99",X"99",X"00",X"39",X"99",X"99",X"30",X"30",X"99",X"90",X"30",X"30",X"90",X"90",X"00",X"09",
		X"90",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"BB",X"22",X"2B",X"B0",X"B2",
		X"22",X"22",X"B0",X"B2",X"22",X"22",X"B0",X"00",X"22",X"20",X"00",X"00",X"09",X"00",X"00",X"09",
		X"99",X"99",X"00",X"39",X"99",X"99",X"30",X"30",X"99",X"90",X"30",X"00",X"90",X"90",X"30",X"00",
		X"90",X"99",X"00",X"00",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"38",X"AA",X"7E",X"39",X"50",X"3B",X"05",X"7E",X"39",X"42",X"7E",X"39",X"3C",X"7E",X"38",
		X"FE",X"40",X"63",X"3B",X"05",X"7E",X"3A",X"D9",X"D0",X"01",X"0C",X"14",X"01",X"08",X"17",X"00",
		X"C0",X"01",X"0A",X"06",X"00",X"D0",X"01",X"08",X"17",X"00",X"B6",X"BE",X"68",X"34",X"02",X"27",
		X"4B",X"BD",X"D0",X"7B",X"CC",X"40",X"63",X"ED",X"02",X"ED",X"88",X"14",X"8D",X"D0",X"BD",X"26",
		X"C3",X"D1",X"2B",X"23",X"0C",X"D1",X"2C",X"24",X"08",X"91",X"2D",X"23",X"04",X"91",X"2E",X"25",
		X"ED",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"1F",X"03",X"EC",X"98",X"02",X"BD",X"D0",X"03",X"26",
		X"DD",X"B6",X"BE",X"5C",X"BD",X"D0",X"42",X"A7",X"88",X"13",X"CC",X"3A",X"76",X"ED",X"08",X"8D",
		X"9A",X"6A",X"E4",X"26",X"BC",X"9F",X"8B",X"BD",X"D0",X"54",X"39",X"B7",X"35",X"82",X"34",X"56",
		X"BD",X"D0",X"45",X"A6",X"09",X"81",X"0A",X"25",X"04",X"86",X"06",X"20",X"06",X"81",X"05",X"23",
		X"02",X"86",X"05",X"8E",X"39",X"20",X"48",X"48",X"30",X"86",X"EC",X"84",X"DD",X"2B",X"EC",X"02",
		X"DD",X"2D",X"35",X"D6",X"40",X"B0",X"1A",X"7A",X"48",X"A8",X"1A",X"7A",X"50",X"A0",X"2A",X"6A",
		X"54",X"9D",X"30",X"60",X"5D",X"96",X"35",X"59",X"62",X"94",X"38",X"5C",X"34",X"26",X"86",X"66",
		X"20",X"02",X"34",X"26",X"97",X"2D",X"EC",X"04",X"10",X"AE",X"02",X"BD",X"D0",X"90",X"35",X"A6",
		X"34",X"70",X"8E",X"B3",X"A4",X"9F",X"27",X"31",X"84",X"6F",X"80",X"8C",X"B3",X"E4",X"25",X"F9",
		X"B6",X"BE",X"69",X"34",X"02",X"27",X"4E",X"BD",X"D0",X"81",X"DC",X"93",X"ED",X"02",X"ED",X"88",
		X"14",X"8D",X"8B",X"DC",X"2B",X"C3",X"03",X"FC",X"DD",X"2B",X"DC",X"2D",X"C3",X"02",X"FD",X"DD",
		X"2D",X"BD",X"26",X"C3",X"D1",X"2B",X"23",X"0C",X"D1",X"2C",X"24",X"08",X"91",X"2D",X"23",X"04",
		X"91",X"2E",X"25",X"ED",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"EE",X"04",X"EC",X"98",X"02",X"BD",
		X"D0",X"03",X"26",X"DD",X"CC",X"3A",X"A9",X"ED",X"08",X"10",X"AF",X"06",X"31",X"22",X"BD",X"38",
		X"8B",X"6A",X"E4",X"26",X"B2",X"35",X"F2",X"96",X"59",X"85",X"7F",X"27",X"08",X"86",X"02",X"8E",
		X"39",X"B7",X"7E",X"D0",X"66",X"86",X"0A",X"8E",X"39",X"CD",X"7E",X"D0",X"66",X"5F",X"B6",X"BE",
		X"68",X"34",X"06",X"27",X"0F",X"9E",X"8B",X"20",X"02",X"AE",X"84",X"6A",X"88",X"13",X"27",X"06",
		X"6A",X"E4",X"26",X"F5",X"20",X"7E",X"B6",X"BE",X"5C",X"BD",X"D0",X"42",X"A7",X"88",X"13",X"E6",
		X"0C",X"D0",X"66",X"22",X"08",X"C1",X"FE",X"22",X"16",X"C6",X"04",X"20",X"06",X"C1",X"02",X"25",
		X"0E",X"C6",X"FC",X"EB",X"0C",X"C1",X"DE",X"22",X"06",X"C1",X"18",X"25",X"02",X"E7",X"0C",X"E6",
		X"0A",X"D0",X"64",X"22",X"04",X"C6",X"02",X"20",X"06",X"C1",X"01",X"25",X"0E",X"C6",X"FE",X"EB",
		X"0A",X"C1",X"8A",X"22",X"06",X"C1",X"07",X"25",X"02",X"E7",X"0A",X"EC",X"02",X"C3",X"00",X"04",
		X"10",X"83",X"40",X"6F",X"23",X"03",X"CC",X"40",X"63",X"ED",X"02",X"BD",X"D0",X"8D",X"6C",X"61",
		X"EE",X"02",X"EC",X"04",X"34",X"10",X"8E",X"98",X"23",X"BD",X"D0",X"27",X"35",X"10",X"27",X"0E",
		X"10",X"AE",X"84",X"8D",X"21",X"6A",X"E4",X"27",X"0B",X"30",X"A4",X"7E",X"39",X"DB",X"6A",X"E4",
		X"10",X"26",X"FF",X"75",X"EC",X"E1",X"27",X"06",X"CC",X"38",X"A0",X"BD",X"D0",X"4B",X"86",X"04",
		X"8E",X"39",X"CD",X"7E",X"D0",X"66",X"96",X"48",X"26",X"2C",X"BD",X"5B",X"43",X"9C",X"8B",X"26",
		X"04",X"EC",X"84",X"DD",X"8B",X"BD",X"D0",X"7E",X"CC",X"01",X"10",X"BD",X"D0",X"0C",X"CC",X"38",
		X"98",X"BD",X"D0",X"4B",X"C6",X"E0",X"B6",X"BE",X"5C",X"3D",X"B1",X"BE",X"5D",X"25",X"03",X"B7",
		X"BE",X"5C",X"7A",X"BE",X"68",X"39",X"7E",X"D0",X"18",X"96",X"48",X"26",X"27",X"BD",X"D0",X"84",
		X"CC",X"00",X"00",X"ED",X"98",X"06",X"BD",X"D0",X"15",X"7A",X"BE",X"69",X"DC",X"13",X"27",X"13",
		X"33",X"84",X"AE",X"84",X"9F",X"1B",X"BD",X"D0",X"54",X"3A",X"D9",X"EF",X"07",X"CC",X"38",X"A5",
		X"7E",X"D0",X"4B",X"39",X"96",X"90",X"7E",X"38",X"88",X"AE",X"47",X"10",X"AE",X"02",X"20",X"17",
		X"AE",X"47",X"10",X"AE",X"02",X"31",X"25",X"A6",X"A4",X"26",X"0C",X"BD",X"D0",X"15",X"DC",X"1B",
		X"ED",X"84",X"9F",X"1B",X"7E",X"D0",X"63",X"10",X"AF",X"02",X"BD",X"D0",X"8D",X"A6",X"24",X"8E",
		X"3A",X"E0",X"7E",X"D0",X"66",X"05",X"09",X"3B",X"95",X"06",X"05",X"09",X"3B",X"C2",X"03",X"05",
		X"09",X"3B",X"EF",X"02",X"00",X"05",X"09",X"3C",X"1C",X"06",X"05",X"09",X"3C",X"49",X"03",X"05",
		X"09",X"3C",X"76",X"02",X"00",X"05",X"09",X"3C",X"A3",X"06",X"05",X"09",X"3C",X"D0",X"03",X"05",
		X"09",X"3C",X"FD",X"02",X"00",X"05",X"09",X"3D",X"2A",X"06",X"05",X"09",X"3D",X"57",X"03",X"05",
		X"09",X"3D",X"84",X"02",X"00",X"03",X"09",X"3D",X"B1",X"06",X"03",X"09",X"3D",X"CC",X"03",X"03",
		X"09",X"3D",X"E7",X"02",X"00",X"05",X"09",X"3E",X"02",X"06",X"05",X"09",X"3E",X"2F",X"03",X"05",
		X"09",X"3E",X"5C",X"02",X"00",X"09",X"07",X"3E",X"89",X"06",X"09",X"07",X"3E",X"C8",X"03",X"09",
		X"07",X"3F",X"07",X"02",X"00",X"05",X"09",X"3F",X"46",X"06",X"05",X"09",X"3F",X"73",X"03",X"05",
		X"09",X"3F",X"A0",X"02",X"00",X"05",X"0A",X"3F",X"CD",X"06",X"05",X"0A",X"3F",X"FF",X"03",X"05",
		X"0A",X"40",X"31",X"02",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"90",X"09",X"00",X"00",
		X"90",X"90",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"99",X"99",X"90",X"00",X"09",
		X"99",X"00",X"00",X"00",X"90",X"90",X"90",X"00",X"09",X"00",X"90",X"09",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"A0",X"A0",
		X"00",X"00",X"0A",X"AA",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"AA",X"00",X"00",
		X"00",X"A0",X"A0",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"09",X"09",X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"09",X"00",
		X"90",X"90",X"00",X"90",X"90",X"09",X"09",X"09",X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"09",
		X"09",X"09",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"0A",X"0A",X"0A",
		X"0A",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",
		X"99",X"90",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",
		X"90",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"99",X"90",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"0A",
		X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"0A",X"AA",
		X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"99",X"90",X"00",X"00",
		X"99",X"99",X"90",X"00",X"09",X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"90",X"09",X"99",X"99",
		X"99",X"90",X"99",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"AA",X"00",
		X"00",X"00",X"AA",X"AA",X"00",X"00",X"0A",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",
		X"A0",X"00",X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"90",X"99",X"99",X"90",X"99",X"99",X"90",X"99",X"99",X"90",X"99",X"99",X"90",
		X"99",X"99",X"90",X"99",X"99",X"90",X"99",X"99",X"90",X"99",X"99",X"90",X"00",X"00",X"00",X"0A",
		X"AA",X"00",X"0A",X"AA",X"00",X"0A",X"AA",X"00",X"0A",X"AA",X"00",X"0A",X"AA",X"00",X"0A",X"AA",
		X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",X"99",X"90",
		X"00",X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"90",X"09",X"99",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"AA",
		X"AA",X"A0",X"00",X"0A",X"AA",X"AA",X"AA",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"00",X"0A",X"AA",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"90",X"90",X"00",X"90",X"00",X"90",X"00",X"90",X"90",X"90",X"99",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"00",X"90",X"90",X"99",X"90",
		X"90",X"90",X"90",X"99",X"90",X"90",X"90",X"00",X"90",X"00",X"90",X"00",X"99",X"90",X"90",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"0A",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"AA",X"00",X"0A",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"0A",X"00",X"0A",X"AA",X"A0",X"A0",
		X"A0",X"A0",X"AA",X"AA",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"99",X"99",X"00",
		X"09",X"99",X"09",X"99",X"00",X"09",X"90",X"00",X"99",X"00",X"99",X"00",X"00",X"09",X"90",X"09",
		X"90",X"00",X"99",X"00",X"09",X"99",X"09",X"99",X"00",X"09",X"99",X"99",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"AA",
		X"A0",X"00",X"00",X"AA",X"0A",X"A0",X"00",X"0A",X"A0",X"00",X"AA",X"00",X"00",X"AA",X"0A",X"A0",
		X"00",X"00",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"0A",X"AA",X"00",X"00",X"00",X"AA",X"0A",X"A0",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",
		X"99",X"90",X"90",X"00",X"00",X"00",X"90",X"90",X"99",X"99",X"90",X"90",X"90",X"90",X"00",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"99",X"90",X"90",X"90",X"90",X"00",X"00",X"90",X"90",
		X"99",X"99",X"99",X"90",X"90",X"00",X"00",X"00",X"00",X"90",X"09",X"99",X"99",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"00",X"A0",
		X"00",X"A0",X"00",X"A0",X"A0",X"A0",X"A0",X"00",X"A0",X"AA",X"A0",X"A0",X"00",X"A0",X"00",X"00",
		X"A0",X"00",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A0",X"00",
		X"00",X"A0",X"00",X"A0",X"00",X"00",X"A0",X"A0",X"A0",X"00",X"00",X"AA",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"0D",X"40",X"73",X"05",X"0D",X"40",X"B4",X"05",X"0D",X"40",X"73",X"05",
		X"0D",X"40",X"F5",X"00",X"01",X"11",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"CC",X"CC",
		X"C0",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"91",X"11",X"91",X"10",X"51",X"19",X"99",X"11",
		X"50",X"50",X"11",X"91",X"10",X"50",X"50",X"01",X"11",X"00",X"50",X"00",X"01",X"11",X"00",X"00",
		X"00",X"11",X"01",X"10",X"00",X"00",X"11",X"01",X"10",X"00",X"05",X"55",X"05",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",X"CC",
		X"CC",X"C0",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"91",X"11",X"91",X"10",X"51",X"19",X"99",
		X"11",X"50",X"50",X"11",X"91",X"10",X"50",X"50",X"01",X"11",X"00",X"50",X"00",X"11",X"11",X"00",
		X"00",X"00",X"11",X"01",X"10",X"00",X"05",X"55",X"01",X"10",X"00",X"00",X"00",X"01",X"10",X"00",
		X"00",X"00",X"05",X"55",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"66",X"66",X"60",X"00",X"00",
		X"CC",X"CC",X"C0",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"91",X"11",X"91",X"10",X"51",X"19",
		X"99",X"11",X"50",X"50",X"11",X"91",X"10",X"50",X"50",X"01",X"11",X"00",X"50",X"00",X"01",X"11",
		X"10",X"00",X"00",X"11",X"01",X"10",X"00",X"00",X"11",X"05",X"55",X"00",X"00",X"11",X"00",X"00",
		X"00",X"05",X"55",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"45",X"9B",X"FF",X"01",X"01",X"13",X"00",X"99",X"22",X"55",X"11",X"99",X"22",X"55",X"11",
		X"99",X"22",X"55",X"11",X"99",X"22",X"55",X"11",X"99",X"22",X"55",X"11",X"AA",X"CC",X"AA",X"CC",
		X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",X"AA",X"CC",
		X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",X"99",X"77",
		X"99",X"77",X"99",X"77",X"11",X"55",X"11",X"55",X"11",X"55",X"11",X"55",X"11",X"55",X"11",X"55",
		X"11",X"55",X"11",X"55",X"11",X"55",X"11",X"55",X"FF",X"EE",X"DD",X"CC",X"BB",X"AA",X"FF",X"EE",
		X"DD",X"CC",X"BB",X"AA",X"FF",X"EE",X"DD",X"CC",X"BB",X"AA",X"FF",X"EE",X"11",X"66",X"77",X"BB",
		X"AA",X"11",X"66",X"77",X"BB",X"AA",X"11",X"66",X"77",X"BB",X"AA",X"11",X"66",X"77",X"BB",X"AA",
		X"33",X"55",X"33",X"55",X"AA",X"33",X"55",X"33",X"55",X"AA",X"33",X"55",X"33",X"55",X"AA",X"33",
		X"55",X"33",X"55",X"AA",X"41",X"48",X"41",X"5C",X"41",X"70",X"41",X"84",X"41",X"98",X"41",X"AC",
		X"41",X"C0",X"41",X"98",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",
		X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"34",X"30",
		X"8E",X"B3",X"ED",X"BF",X"B3",X"E4",X"31",X"89",X"00",X"81",X"10",X"AF",X"84",X"10",X"8C",X"B8",
		X"F7",X"24",X"04",X"30",X"A4",X"20",X"EF",X"10",X"8E",X"00",X"00",X"10",X"AF",X"84",X"10",X"BF",
		X"B3",X"E6",X"35",X"B0",X"34",X"66",X"8D",X"37",X"25",X"27",X"10",X"BF",X"B3",X"E6",X"AF",X"26",
		X"EC",X"84",X"ED",X"22",X"3D",X"E7",X"28",X"33",X"2D",X"EF",X"24",X"8D",X"16",X"CE",X"43",X"38",
		X"EF",X"29",X"BD",X"D0",X"39",X"84",X"07",X"48",X"CE",X"41",X"D4",X"EC",X"C6",X"ED",X"2B",X"30",
		X"22",X"35",X"E6",X"34",X"26",X"10",X"AE",X"24",X"6F",X"A0",X"5A",X"26",X"FB",X"35",X"A6",X"34",
		X"10",X"10",X"BE",X"B3",X"E4",X"27",X"0E",X"AE",X"A4",X"BF",X"B3",X"E4",X"BE",X"B3",X"E6",X"AF",
		X"A4",X"1C",X"FE",X"35",X"90",X"1A",X"01",X"35",X"90",X"AE",X"29",X"34",X"10",X"30",X"01",X"AF",
		X"29",X"96",X"84",X"84",X"07",X"AE",X"2B",X"30",X"86",X"BF",X"B3",X"E8",X"AE",X"26",X"E6",X"28",
		X"35",X"C0",X"34",X"76",X"AE",X"02",X"10",X"AE",X"24",X"A6",X"C4",X"2A",X"13",X"84",X"7F",X"BD",
		X"42",X"F5",X"EC",X"C1",X"B1",X"B3",X"EA",X"24",X"1C",X"53",X"E4",X"A6",X"E7",X"A6",X"20",X"F2",
		X"85",X"40",X"26",X"13",X"8D",X"2F",X"EC",X"C1",X"B1",X"B3",X"EA",X"24",X"08",X"E4",X"86",X"EA",
		X"A6",X"E7",X"A6",X"20",X"F1",X"35",X"F6",X"84",X"3F",X"8D",X"1A",X"EC",X"C1",X"B1",X"B3",X"EA",
		X"24",X"F3",X"E4",X"86",X"27",X"F5",X"E6",X"9F",X"B3",X"E8",X"7C",X"B3",X"E9",X"E4",X"5F",X"EA",
		X"A6",X"E7",X"A6",X"20",X"E6",X"CE",X"43",X"BB",X"4A",X"48",X"EE",X"C6",X"F7",X"B3",X"EA",X"39",
		X"34",X"10",X"AE",X"A4",X"AF",X"9F",X"B3",X"EB",X"BE",X"B3",X"E4",X"AF",X"A4",X"10",X"BF",X"B3",
		X"E4",X"10",X"BE",X"B3",X"EB",X"35",X"90",X"10",X"8E",X"B3",X"E6",X"20",X"0C",X"BD",X"42",X"89",
		X"11",X"83",X"43",X"BA",X"27",X"0D",X"BD",X"42",X"A2",X"10",X"BF",X"B3",X"EB",X"10",X"AE",X"A4",
		X"26",X"EB",X"39",X"BD",X"43",X"00",X"20",X"F1",X"43",X"83",X"46",X"86",X"44",X"84",X"42",X"82",
		X"41",X"81",X"47",X"87",X"44",X"46",X"84",X"42",X"86",X"43",X"82",X"41",X"83",X"45",X"81",X"48",
		X"85",X"47",X"88",X"44",X"87",X"45",X"42",X"84",X"46",X"85",X"47",X"82",X"48",X"86",X"43",X"87",
		X"41",X"88",X"42",X"83",X"44",X"81",X"45",X"47",X"82",X"46",X"84",X"85",X"48",X"87",X"43",X"86",
		X"44",X"42",X"88",X"45",X"83",X"41",X"84",X"43",X"82",X"47",X"46",X"85",X"48",X"81",X"42",X"83",
		X"44",X"87",X"41",X"86",X"45",X"88",X"43",X"46",X"84",X"48",X"81",X"47",X"85",X"44",X"82",X"41",
		X"45",X"83",X"42",X"86",X"88",X"43",X"87",X"46",X"84",X"48",X"85",X"07",X"81",X"04",X"05",X"82",
		X"01",X"83",X"02",X"86",X"03",X"88",X"06",X"87",X"08",X"84",X"07",X"85",X"04",X"81",X"05",X"01",
		X"82",X"83",X"02",X"03",X"88",X"08",X"84",X"87",X"07",X"04",X"00",X"43",X"CB",X"44",X"05",X"44",
		X"3F",X"44",X"79",X"44",X"B3",X"44",X"ED",X"45",X"27",X"45",X"61",X"00",X"F0",X"06",X"0F",X"09",
		X"0F",X"0C",X"F0",X"13",X"F0",X"17",X"0F",X"18",X"0F",X"1D",X"F0",X"22",X"F0",X"25",X"0F",X"2B",
		X"F0",X"2E",X"0F",X"30",X"F0",X"32",X"0F",X"3C",X"F0",X"3E",X"0F",X"43",X"0F",X"45",X"F0",X"48",
		X"F0",X"4C",X"0F",X"50",X"0F",X"51",X"F0",X"5A",X"F0",X"5D",X"0F",X"60",X"0F",X"65",X"F0",X"6A",
		X"0F",X"6E",X"0F",X"73",X"F0",X"01",X"0F",X"03",X"F0",X"08",X"F0",X"0F",X"0F",X"12",X"F0",X"14",
		X"0F",X"1B",X"0F",X"1E",X"F0",X"20",X"F0",X"22",X"0F",X"2D",X"F0",X"2F",X"0F",X"33",X"0F",X"35",
		X"F0",X"39",X"0F",X"3D",X"F0",X"43",X"F0",X"47",X"0F",X"4A",X"0F",X"4E",X"F0",X"53",X"F0",X"55",
		X"0F",X"5B",X"0F",X"5B",X"F0",X"63",X"0F",X"68",X"F0",X"6D",X"F0",X"71",X"0F",X"73",X"0F",X"04",
		X"0F",X"07",X"F0",X"09",X"F0",X"0A",X"0F",X"14",X"F0",X"15",X"0F",X"1C",X"0F",X"1F",X"F0",X"21",
		X"F0",X"23",X"0F",X"29",X"0F",X"2E",X"F0",X"34",X"0F",X"36",X"F0",X"3A",X"F0",X"3D",X"0F",X"42",
		X"F0",X"44",X"0F",X"49",X"0F",X"4D",X"F0",X"55",X"F0",X"57",X"0F",X"59",X"0F",X"5C",X"F0",X"61",
		X"F0",X"68",X"0F",X"6A",X"F0",X"6D",X"0F",X"72",X"0F",X"00",X"0F",X"02",X"F0",X"0A",X"F0",X"0C",
		X"0F",X"10",X"F0",X"16",X"0F",X"1A",X"F0",X"1E",X"0F",X"21",X"0F",X"23",X"F0",X"2C",X"0F",X"2F",
		X"F0",X"33",X"F0",X"36",X"0F",X"38",X"F0",X"3B",X"0F",X"42",X"0F",X"46",X"F0",X"49",X"F0",X"4D",
		X"0F",X"52",X"F0",X"54",X"0F",X"5A",X"0F",X"5D",X"F0",X"61",X"0F",X"64",X"F0",X"69",X"0F",X"6C",
		X"F0",X"70",X"F0",X"02",X"0F",X"06",X"F0",X"08",X"0F",X"0E",X"F0",X"13",X"0F",X"16",X"F0",X"19",
		X"F0",X"1D",X"0F",X"24",X"0F",X"27",X"F0",X"29",X"F0",X"2B",X"0F",X"30",X"0F",X"31",X"F0",X"3C",
		X"0F",X"3E",X"F0",X"40",X"0F",X"41",X"F0",X"4B",X"F0",X"4E",X"0F",X"52",X"0F",X"57",X"F0",X"59",
		X"F0",X"5E",X"0F",X"62",X"F0",X"65",X"0F",X"67",X"F0",X"6B",X"0F",X"6F",X"F0",X"01",X"F0",X"07",
		X"0F",X"0B",X"0F",X"0D",X"F0",X"11",X"0F",X"15",X"F0",X"1A",X"0F",X"1C",X"F0",X"20",X"0F",X"25",
		X"F0",X"2A",X"F0",X"2D",X"0F",X"31",X"0F",X"32",X"F0",X"38",X"0F",X"3F",X"F0",X"44",X"F0",X"46",
		X"0F",X"4B",X"0F",X"4F",X"F0",X"54",X"F0",X"56",X"0F",X"58",X"0F",X"5F",X"F0",X"60",X"F0",X"66",
		X"F0",X"6C",X"0F",X"6F",X"0F",X"71",X"F0",X"03",X"0F",X"04",X"F0",X"0D",X"0F",X"0F",X"F0",X"11",
		X"F0",X"12",X"0F",X"18",X"F0",X"1F",X"0F",X"26",X"F0",X"27",X"0F",X"28",X"0F",X"2C",X"F0",X"34",
		X"F0",X"37",X"0F",X"3B",X"F0",X"3F",X"0F",X"40",X"F0",X"45",X"0F",X"48",X"0F",X"4A",X"F0",X"53",
		X"0F",X"56",X"F0",X"58",X"F0",X"5C",X"0F",X"62",X"0F",X"64",X"0F",X"6B",X"F0",X"70",X"0F",X"72",
		X"F0",X"05",X"F0",X"05",X"0F",X"0B",X"F0",X"0E",X"0F",X"10",X"0F",X"17",X"F0",X"19",X"0F",X"1B",
		X"F0",X"24",X"F0",X"26",X"0F",X"28",X"F0",X"2A",X"0F",X"35",X"0F",X"37",X"F0",X"39",X"F0",X"3A",
		X"0F",X"41",X"0F",X"47",X"F0",X"4C",X"F0",X"4F",X"0F",X"50",X"F0",X"51",X"0F",X"5E",X"F0",X"5F",
		X"0F",X"63",X"F0",X"66",X"0F",X"67",X"0F",X"69",X"F0",X"6E",X"F0",X"BD",X"42",X"0E",X"9E",X"21",
		X"27",X"52",X"BD",X"D0",X"54",X"46",X"07",X"9E",X"21",X"CC",X"00",X"00",X"10",X"8E",X"00",X"00",
		X"34",X"06",X"34",X"06",X"EC",X"02",X"ED",X"88",X"14",X"31",X"21",X"10",X"8C",X"00",X"0F",X"22",
		X"05",X"10",X"A3",X"E4",X"27",X"11",X"10",X"8E",X"00",X"00",X"ED",X"E4",X"34",X"10",X"AE",X"02",
		X"BD",X"42",X"34",X"AF",X"64",X"35",X"10",X"EC",X"62",X"ED",X"02",X"AE",X"84",X"26",X"D5",X"32",
		X"64",X"BD",X"46",X"39",X"BD",X"43",X"17",X"BE",X"B3",X"E6",X"27",X"08",X"86",X"01",X"8E",X"45",
		X"E1",X"7E",X"D0",X"66",X"9E",X"21",X"27",X"09",X"EC",X"88",X"14",X"ED",X"02",X"AE",X"84",X"26",
		X"F7",X"BD",X"F0",X"09",X"7E",X"D0",X"63",X"CC",X"41",X"43",X"BD",X"D0",X"4B",X"86",X"48",X"A7",
		X"47",X"C6",X"12",X"BD",X"D0",X"06",X"6A",X"47",X"27",X"08",X"86",X"01",X"8E",X"46",X"11",X"7E",
		X"D0",X"66",X"86",X"24",X"A7",X"47",X"C6",X"12",X"BD",X"D0",X"06",X"6A",X"47",X"10",X"27",X"8A",
		X"32",X"86",X"02",X"8E",X"46",X"26",X"7E",X"D0",X"66",X"9E",X"21",X"27",X"23",X"10",X"AE",X"02",
		X"EC",X"A4",X"88",X"04",X"C8",X"04",X"1A",X"10",X"FD",X"CA",X"06",X"EE",X"22",X"FF",X"CA",X"02",
		X"EC",X"04",X"FD",X"CA",X"04",X"86",X"06",X"B7",X"CA",X"00",X"1C",X"EF",X"AE",X"84",X"26",X"DD",
		X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"46",X"8C",X"7E",X"47",X"3F",X"7E",X"46",X"E6",X"7E",X"4A",X"79",X"34",X"30",X"8E",X"BB",
		X"E4",X"9F",X"C0",X"31",X"88",X"33",X"10",X"AF",X"84",X"10",X"8C",X"BD",X"E2",X"24",X"04",X"30",
		X"A4",X"20",X"F0",X"10",X"8E",X"00",X"00",X"10",X"AF",X"84",X"10",X"9F",X"BC",X"10",X"9F",X"BE",
		X"35",X"B0",X"34",X"20",X"DE",X"C0",X"27",X"12",X"10",X"AE",X"C4",X"10",X"9F",X"C0",X"10",X"9E",
		X"BC",X"10",X"AF",X"C4",X"DF",X"BC",X"1C",X"FE",X"35",X"A0",X"1A",X"01",X"35",X"A0",X"34",X"20",
		X"DE",X"C0",X"27",X"F6",X"10",X"AE",X"C4",X"10",X"9F",X"C0",X"10",X"9E",X"BE",X"10",X"AF",X"C4",
		X"DF",X"BE",X"1C",X"FE",X"35",X"A0",X"34",X"76",X"BD",X"46",X"CE",X"25",X"40",X"A7",X"C8",X"12",
		X"EC",X"04",X"AE",X"02",X"ED",X"4B",X"A7",X"44",X"D6",X"A7",X"E7",X"45",X"E0",X"4C",X"25",X"04",
		X"E1",X"01",X"25",X"0B",X"E6",X"84",X"54",X"E7",X"46",X"EB",X"4C",X"E7",X"45",X"20",X"02",X"E7",
		X"46",X"EC",X"84",X"ED",X"4D",X"C6",X"01",X"E7",X"C8",X"11",X"88",X"04",X"C8",X"04",X"ED",X"4F",
		X"AE",X"02",X"AF",X"42",X"CC",X"10",X"00",X"ED",X"48",X"6F",X"47",X"8D",X"02",X"35",X"F6",X"AE",
		X"42",X"E6",X"4D",X"A6",X"4E",X"33",X"C8",X"13",X"AF",X"C1",X"3A",X"4A",X"26",X"FA",X"39",X"34",
		X"76",X"BD",X"46",X"B2",X"25",X"44",X"A7",X"C8",X"12",X"EC",X"04",X"AE",X"02",X"ED",X"4B",X"A7",
		X"44",X"D6",X"A7",X"E7",X"45",X"E0",X"4C",X"25",X"04",X"E1",X"01",X"25",X"0B",X"E6",X"84",X"54",
		X"E7",X"46",X"EB",X"4C",X"E7",X"45",X"20",X"02",X"E7",X"46",X"EC",X"84",X"ED",X"4D",X"E7",X"C8",
		X"11",X"C6",X"01",X"88",X"04",X"C8",X"04",X"ED",X"4F",X"AE",X"02",X"AF",X"42",X"CC",X"01",X"00",
		X"ED",X"48",X"6F",X"47",X"86",X"10",X"A7",X"4A",X"8D",X"A5",X"35",X"F6",X"AE",X"A1",X"BF",X"CA",
		X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",
		X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",
		X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",
		X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",
		X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",
		X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",
		X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",
		X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",
		X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",
		X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",
		X"FF",X"CA",X"00",X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",
		X"D3",X"BA",X"AE",X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"D3",X"BA",X"AE",
		X"A1",X"BF",X"CA",X"02",X"FD",X"CA",X"04",X"FF",X"CA",X"00",X"1C",X"EF",X"35",X"A0",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",
		X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"FD",X"CA",X"04",X"FF",X"C9",X"FF",X"D3",X"BA",X"1C",X"EF",
		X"39",X"E6",X"A8",X"11",X"C0",X"10",X"50",X"58",X"58",X"58",X"8E",X"48",X"5E",X"3A",X"EC",X"27",
		X"DD",X"BA",X"96",X"45",X"C6",X"12",X"1F",X"03",X"CC",X"00",X"00",X"1A",X"10",X"FD",X"CA",X"01",
		X"EC",X"2F",X"FD",X"CA",X"06",X"EC",X"2B",X"6E",X"84",X"CE",X"98",X"BC",X"10",X"AC",X"C4",X"27",
		X"08",X"EE",X"C4",X"26",X"F7",X"1A",X"10",X"20",X"FE",X"EC",X"A4",X"ED",X"C4",X"DC",X"C0",X"ED",
		X"A4",X"10",X"9F",X"C0",X"31",X"C4",X"39",X"EC",X"28",X"83",X"01",X"00",X"A1",X"28",X"26",X"03",
		X"E7",X"29",X"39",X"BD",X"48",X"E1",X"96",X"59",X"26",X"08",X"DC",X"5E",X"A7",X"24",X"EB",X"26",
		X"E7",X"25",X"A6",X"2E",X"97",X"C2",X"EC",X"28",X"83",X"01",X"00",X"81",X"01",X"22",X"12",X"CE",
		X"98",X"BE",X"20",X"B8",X"6A",X"2A",X"27",X"B1",X"A6",X"2E",X"97",X"C2",X"EC",X"28",X"C3",X"01",
		X"00",X"97",X"BB",X"ED",X"28",X"44",X"97",X"C5",X"E6",X"A8",X"12",X"2A",X"01",X"40",X"A7",X"27",
		X"97",X"BA",X"E6",X"26",X"26",X"02",X"D7",X"C5",X"96",X"BB",X"E6",X"26",X"D7",X"B9",X"3D",X"DD",
		X"C3",X"E6",X"25",X"4F",X"93",X"C3",X"DB",X"C5",X"89",X"00",X"26",X"04",X"C1",X"18",X"22",X"0E",
		X"0A",X"C2",X"0A",X"B9",X"DB",X"BB",X"89",X"00",X"26",X"F6",X"C1",X"18",X"23",X"F2",X"E7",X"2C",
		X"96",X"B9",X"D6",X"BA",X"2B",X"2C",X"3D",X"DD",X"C3",X"E6",X"24",X"4F",X"93",X"C3",X"4D",X"26",
		X"04",X"C1",X"07",X"22",X"41",X"0F",X"B8",X"0A",X"C2",X"0C",X"B8",X"DB",X"BA",X"89",X"00",X"26",
		X"F6",X"C1",X"07",X"23",X"F2",X"E7",X"2B",X"D6",X"B8",X"96",X"BB",X"3D",X"EB",X"2C",X"E7",X"2C",
		X"20",X"26",X"50",X"3D",X"EB",X"2D",X"EB",X"24",X"89",X"00",X"26",X"04",X"C1",X"8F",X"23",X"14",
		X"0F",X"B8",X"0A",X"C2",X"0C",X"B8",X"DB",X"BA",X"89",X"FF",X"26",X"F6",X"C1",X"8F",X"22",X"F2",
		X"E0",X"2D",X"20",X"D1",X"E0",X"2D",X"E7",X"2B",X"30",X"A8",X"13",X"E6",X"2E",X"D0",X"C2",X"58",
		X"3A",X"96",X"C2",X"4A",X"D6",X"BB",X"3D",X"EB",X"2C",X"89",X"00",X"27",X"0A",X"0A",X"C2",X"27",
		X"48",X"D0",X"BB",X"82",X"00",X"26",X"F6",X"C1",X"EA",X"24",X"F2",X"96",X"C2",X"4A",X"D6",X"BA",
		X"2B",X"19",X"3D",X"EB",X"2D",X"EB",X"2B",X"89",X"00",X"27",X"0A",X"0A",X"C2",X"27",X"2A",X"D0",
		X"BA",X"82",X"00",X"26",X"F6",X"C1",X"8F",X"22",X"F2",X"20",X"1A",X"50",X"3D",X"DD",X"C3",X"E6",
		X"2B",X"4F",X"93",X"C3",X"4D",X"27",X"0A",X"0A",X"C2",X"27",X"0E",X"D0",X"BA",X"82",X"FF",X"26",
		X"F6",X"C1",X"07",X"23",X"F2",X"96",X"C2",X"26",X"03",X"7E",X"49",X"09",X"A7",X"A8",X"11",X"80",
		X"10",X"40",X"C6",X"0D",X"3D",X"C3",X"47",X"8C",X"34",X"26",X"CE",X"0A",X"0A",X"EC",X"2F",X"1A",
		X"10",X"FD",X"CA",X"06",X"EC",X"2B",X"31",X"84",X"39",X"10",X"9E",X"BC",X"27",X"0B",X"BD",X"48",
		X"E1",X"BD",X"49",X"54",X"10",X"AE",X"A4",X"26",X"F5",X"10",X"9E",X"BE",X"27",X"08",X"BD",X"49",
		X"27",X"10",X"AE",X"A4",X"26",X"F8",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"4D",X"10",X"7E",X"4B",X"36",X"50",X"C2",X"50",X"0E",X"50",X"26",X"D0",X"01",X"08",X"11",
		X"00",X"C8",X"01",X"08",X"04",X"00",X"C8",X"01",X"04",X"14",X"01",X"01",X"13",X"00",X"D0",X"01",
		X"03",X"01",X"01",X"04",X"15",X"01",X"04",X"13",X"00",X"D0",X"01",X"04",X"15",X"01",X"08",X"11",
		X"00",X"D0",X"01",X"08",X"19",X"00",X"B6",X"BE",X"70",X"34",X"02",X"27",X"43",X"BD",X"D0",X"6C",
		X"4B",X"FB",X"50",X"C6",X"4B",X"C9",X"27",X"38",X"C6",X"1A",X"BD",X"D0",X"39",X"2A",X"02",X"C6",
		X"DC",X"86",X"7E",X"BD",X"D0",X"42",X"8B",X"06",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"B6",X"BE",
		X"66",X"BD",X"D0",X"3F",X"A7",X"49",X"B6",X"BE",X"5E",X"BD",X"D0",X"3F",X"44",X"89",X"00",X"A7",
		X"4A",X"CC",X"50",X"D2",X"ED",X"88",X"16",X"9F",X"17",X"BD",X"4B",X"82",X"6A",X"E4",X"26",X"BD",
		X"35",X"82",X"B6",X"BE",X"67",X"BD",X"D0",X"3F",X"E6",X"0A",X"C1",X"0C",X"23",X"09",X"C1",X"83",
		X"24",X"04",X"D6",X"86",X"2A",X"01",X"40",X"1F",X"89",X"1D",X"58",X"49",X"58",X"49",X"ED",X"0E",
		X"B6",X"BE",X"67",X"BD",X"D0",X"3F",X"E6",X"0C",X"C1",X"1D",X"23",X"09",X"C1",X"D6",X"24",X"04",
		X"D6",X"85",X"2B",X"01",X"40",X"1F",X"89",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"ED",X"88",
		X"10",X"96",X"84",X"84",X"1F",X"4C",X"A7",X"4E",X"39",X"96",X"48",X"26",X"2D",X"BD",X"D0",X"78",
		X"DE",X"1B",X"EC",X"C4",X"DD",X"1B",X"BD",X"D0",X"54",X"11",X"43",X"EF",X"07",X"CC",X"50",X"C6",
		X"ED",X"42",X"CC",X"DD",X"DD",X"ED",X"0B",X"86",X"08",X"A7",X"0D",X"CC",X"4B",X"29",X"BD",X"D0",
		X"4B",X"CC",X"02",X"10",X"BD",X"D0",X"0C",X"7A",X"BE",X"70",X"39",X"AE",X"47",X"EC",X"02",X"C3",
		X"00",X"04",X"10",X"83",X"50",X"D2",X"23",X"0B",X"CC",X"50",X"C2",X"0D",X"59",X"26",X"04",X"6A",
		X"49",X"27",X"11",X"ED",X"02",X"6A",X"4E",X"26",X"03",X"BD",X"4B",X"82",X"86",X"03",X"8E",X"4B",
		X"FB",X"7E",X"D0",X"66",X"B6",X"BE",X"66",X"44",X"4C",X"BD",X"D0",X"3F",X"A7",X"49",X"AE",X"47",
		X"6A",X"49",X"26",X"1C",X"96",X"42",X"81",X"11",X"24",X"EA",X"96",X"13",X"9A",X"1B",X"27",X"E4",
		X"B6",X"BE",X"71",X"81",X"14",X"24",X"DD",X"BD",X"4C",X"AC",X"6A",X"4A",X"27",X"21",X"20",X"D4",
		X"EC",X"02",X"C3",X"00",X"04",X"10",X"83",X"50",X"E2",X"23",X"03",X"CC",X"50",X"C2",X"ED",X"02",
		X"6A",X"4E",X"26",X"03",X"BD",X"4B",X"82",X"86",X"03",X"8E",X"4C",X"2E",X"7E",X"D0",X"66",X"CC",
		X"00",X"00",X"ED",X"0E",X"CC",X"02",X"00",X"0D",X"84",X"2A",X"01",X"40",X"ED",X"88",X"10",X"AE",
		X"47",X"EC",X"02",X"83",X"00",X"04",X"10",X"83",X"50",X"C2",X"24",X"0D",X"A6",X"0C",X"81",X"1A",
		X"23",X"11",X"81",X"DA",X"24",X"0D",X"CC",X"50",X"E2",X"ED",X"02",X"86",X"03",X"8E",X"4C",X"7F",
		X"7E",X"D0",X"66",X"BD",X"D0",X"75",X"7A",X"BE",X"70",X"7E",X"D0",X"63",X"34",X"76",X"31",X"84",
		X"BD",X"D0",X"54",X"4D",X"83",X"33",X"84",X"BD",X"D0",X"7B",X"7C",X"BE",X"71",X"CC",X"50",X"0E",
		X"ED",X"02",X"ED",X"88",X"14",X"EF",X"06",X"AF",X"47",X"CC",X"4D",X"F2",X"ED",X"08",X"CC",X"4B",
		X"31",X"BD",X"D0",X"4B",X"EC",X"24",X"C1",X"18",X"27",X"01",X"5A",X"C3",X"02",X"06",X"ED",X"04",
		X"A7",X"0A",X"E7",X"0C",X"BD",X"4E",X"11",X"B6",X"BE",X"64",X"A7",X"4D",X"BD",X"D0",X"18",X"35",
		X"F6",X"20",X"28",X"43",X"29",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",
		X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",
		X"B6",X"BE",X"71",X"34",X"02",X"27",X"4A",X"BD",X"D0",X"54",X"4D",X"8B",X"33",X"84",X"BD",X"D0",
		X"7B",X"CC",X"50",X"26",X"ED",X"02",X"ED",X"88",X"14",X"EF",X"06",X"AF",X"47",X"CC",X"4D",X"F2",
		X"ED",X"08",X"BD",X"38",X"8E",X"BD",X"26",X"C3",X"D1",X"2B",X"23",X"0C",X"D1",X"2C",X"24",X"08",
		X"91",X"2D",X"23",X"04",X"91",X"2E",X"23",X"ED",X"ED",X"04",X"A7",X"0A",X"E7",X"0C",X"BD",X"4E",
		X"11",X"96",X"84",X"84",X"1F",X"BB",X"BE",X"64",X"A7",X"4D",X"BD",X"38",X"8B",X"6A",X"E4",X"26",
		X"B6",X"35",X"82",X"AE",X"47",X"BD",X"D0",X"15",X"EC",X"04",X"10",X"AE",X"02",X"AB",X"24",X"EB",
		X"25",X"A7",X"0A",X"E7",X"0C",X"31",X"26",X"10",X"AF",X"02",X"BD",X"D0",X"18",X"10",X"8C",X"50",
		X"26",X"24",X"08",X"86",X"0C",X"8E",X"4D",X"63",X"7E",X"D0",X"66",X"96",X"59",X"85",X"7F",X"27",
		X"08",X"86",X"0F",X"8E",X"4D",X"8B",X"7E",X"D0",X"66",X"AE",X"47",X"6A",X"4D",X"26",X"03",X"BD",
		X"4E",X"46",X"A6",X"4B",X"5F",X"47",X"56",X"E3",X"0A",X"34",X"06",X"E6",X"4C",X"EB",X"0C",X"BD",
		X"00",X"06",X"27",X"04",X"32",X"62",X"20",X"2F",X"E7",X"0C",X"35",X"06",X"ED",X"0A",X"EC",X"02",
		X"6D",X"4B",X"2A",X"0E",X"83",X"00",X"04",X"10",X"83",X"50",X"26",X"24",X"11",X"CC",X"50",X"32",
		X"20",X"0C",X"C3",X"00",X"04",X"10",X"83",X"50",X"32",X"23",X"03",X"CC",X"50",X"26",X"ED",X"02",
		X"BD",X"D0",X"8D",X"6A",X"4E",X"26",X"03",X"BD",X"4E",X"11",X"96",X"EF",X"8E",X"4D",X"99",X"7E",
		X"D0",X"66",X"96",X"48",X"26",X"1A",X"7A",X"BE",X"71",X"BD",X"5B",X"4F",X"BD",X"D0",X"7E",X"AE",
		X"06",X"BD",X"D0",X"5D",X"CC",X"01",X"20",X"BD",X"D0",X"0C",X"CC",X"4B",X"0C",X"BD",X"D0",X"4B",
		X"39",X"96",X"84",X"81",X"60",X"23",X"05",X"BD",X"26",X"C3",X"20",X"02",X"DC",X"5E",X"DD",X"2B",
		X"E0",X"05",X"24",X"01",X"50",X"C1",X"10",X"24",X"03",X"5F",X"20",X"09",X"DC",X"2B",X"E1",X"05",
		X"C6",X"01",X"24",X"01",X"50",X"A1",X"04",X"86",X"01",X"24",X"01",X"40",X"ED",X"4B",X"96",X"84",
		X"84",X"1F",X"4C",X"A7",X"4E",X"39",X"34",X"50",X"31",X"84",X"B6",X"BE",X"64",X"A7",X"4D",X"96",
		X"42",X"81",X"11",X"10",X"24",X"01",X"3B",X"96",X"F1",X"81",X"14",X"10",X"22",X"01",X"33",X"0C",
		X"F1",X"BD",X"D0",X"6C",X"4F",X"94",X"4F",X"EE",X"4F",X"D5",X"10",X"27",X"01",X"24",X"EC",X"24",
		X"C3",X"01",X"00",X"A7",X"0A",X"E7",X"0C",X"ED",X"04",X"C6",X"80",X"D1",X"84",X"23",X"55",X"D6",
		X"86",X"C4",X"1F",X"CB",X"F0",X"96",X"5E",X"81",X"11",X"24",X"01",X"5F",X"DB",X"5E",X"4F",X"E0",
		X"04",X"82",X"00",X"34",X"02",X"2A",X"01",X"50",X"B6",X"BE",X"65",X"3D",X"1F",X"89",X"A6",X"E0",
		X"2A",X"01",X"53",X"58",X"49",X"58",X"49",X"58",X"49",X"ED",X"0E",X"D6",X"86",X"C4",X"1F",X"CB",
		X"F0",X"DB",X"5F",X"4F",X"E0",X"05",X"82",X"00",X"34",X"02",X"2A",X"01",X"50",X"B6",X"BE",X"65",
		X"3D",X"1F",X"89",X"A6",X"E0",X"2A",X"01",X"53",X"58",X"49",X"58",X"49",X"58",X"49",X"ED",X"88",
		X"10",X"7E",X"4F",X"82",X"BD",X"D0",X"39",X"44",X"25",X"29",X"4F",X"D6",X"84",X"C4",X"1F",X"CB",
		X"F0",X"EB",X"05",X"DB",X"5F",X"89",X"00",X"44",X"56",X"96",X"86",X"84",X"07",X"27",X"0A",X"96",
		X"5E",X"81",X"4B",X"25",X"0A",X"86",X"8F",X"20",X"33",X"96",X"5E",X"81",X"4B",X"23",X"F6",X"86",
		X"07",X"20",X"29",X"4F",X"D6",X"84",X"C4",X"0F",X"CB",X"F8",X"EB",X"04",X"DB",X"5E",X"89",X"00",
		X"44",X"56",X"96",X"86",X"84",X"07",X"27",X"0A",X"96",X"5F",X"81",X"81",X"25",X"0A",X"86",X"EA",
		X"20",X"08",X"96",X"5F",X"81",X"81",X"23",X"F6",X"86",X"18",X"1E",X"89",X"97",X"2B",X"4F",X"E0",
		X"05",X"82",X"00",X"ED",X"88",X"10",X"D6",X"2B",X"4F",X"E0",X"04",X"82",X"00",X"ED",X"0E",X"F6",
		X"BE",X"65",X"86",X"40",X"3D",X"1F",X"89",X"4F",X"58",X"49",X"58",X"49",X"34",X"06",X"43",X"53",
		X"34",X"06",X"58",X"49",X"34",X"06",X"43",X"53",X"34",X"06",X"EC",X"0E",X"10",X"A3",X"64",X"2F",
		X"1F",X"10",X"A3",X"66",X"2C",X"1A",X"EC",X"88",X"10",X"10",X"A3",X"62",X"2F",X"12",X"10",X"A3",
		X"E4",X"2C",X"0D",X"58",X"49",X"ED",X"88",X"10",X"EC",X"0E",X"58",X"49",X"ED",X"0E",X"20",X"DC",
		X"32",X"68",X"9F",X"17",X"96",X"85",X"84",X"1F",X"8B",X"30",X"A7",X"4E",X"CC",X"4B",X"11",X"BD",
		X"D0",X"4B",X"35",X"D0",X"AE",X"47",X"EC",X"0A",X"E3",X"0E",X"81",X"07",X"25",X"23",X"81",X"8B",
		X"22",X"1F",X"EC",X"0C",X"E3",X"88",X"10",X"81",X"18",X"25",X"1C",X"81",X"E3",X"22",X"18",X"6A",
		X"4E",X"27",X"08",X"86",X"02",X"8E",X"4F",X"94",X"7E",X"D0",X"66",X"BD",X"D0",X"75",X"7E",X"D0",
		X"63",X"63",X"0E",X"63",X"0F",X"20",X"06",X"63",X"88",X"10",X"63",X"88",X"11",X"CC",X"4B",X"16",
		X"BD",X"D0",X"4B",X"20",X"DE",X"96",X"48",X"26",X"14",X"0A",X"F1",X"BD",X"5B",X"43",X"BD",X"D0",
		X"78",X"CC",X"00",X"25",X"BD",X"D0",X"0C",X"CC",X"4B",X"1E",X"7E",X"D0",X"4B",X"39",X"04",X"07",
		X"4F",X"F2",X"00",X"0A",X"00",X"00",X"0A",X"CC",X"CA",X"00",X"0C",X"0B",X"0C",X"A0",X"AC",X"BB",
		X"BC",X"A0",X"0C",X"0B",X"0C",X"A0",X"0A",X"CC",X"CA",X"00",X"00",X"0A",X"00",X"00",X"02",X"04",
		X"50",X"36",X"FF",X"FF",X"04",X"07",X"50",X"3E",X"00",X"FF",X"04",X"08",X"50",X"5A",X"FF",X"FE",
		X"06",X"0C",X"50",X"7A",X"00",X"FE",X"07",X"10",X"55",X"1E",X"07",X"10",X"55",X"8E",X"07",X"10",
		X"55",X"FE",X"07",X"10",X"56",X"6E",X"01",X"00",X"11",X"10",X"11",X"10",X"97",X"90",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"11",X"00",X"16",X"66",X"61",X"00",X"11",X"11",
		X"11",X"00",X"79",X"79",X"79",X"00",X"07",X"97",X"90",X"00",X"00",X"11",X"10",X"00",X"00",X"19",
		X"10",X"00",X"11",X"11",X"11",X"10",X"16",X"60",X"66",X"10",X"16",X"06",X"06",X"10",X"11",X"11",
		X"11",X"10",X"97",X"79",X"77",X"90",X"07",X"97",X"79",X"00",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"00",X"19",X"91",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"00",X"10",X"60",X"06",X"01",X"00",X"00",X"16",
		X"06",X"60",X"61",X"00",X"00",X"10",X"60",X"06",X"01",X"00",X"00",X"11",X"11",X"11",X"11",X"00",
		X"00",X"97",X"79",X"77",X"97",X"00",X"07",X"00",X"00",X"00",X"00",X"70",X"00",X"79",X"77",X"97",
		X"79",X"00",X"08",X"0F",X"50",X"E6",X"08",X"0F",X"51",X"5E",X"08",X"0F",X"51",X"D6",X"08",X"0F",
		X"52",X"4E",X"08",X"0F",X"52",X"C6",X"08",X"0F",X"53",X"3E",X"08",X"0F",X"53",X"B6",X"08",X"0F",
		X"54",X"2E",X"08",X"0F",X"54",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EA",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"0E",X"A0",X"AE",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0A",X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"A0",X"AE",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"EA",X"00",X"0A",X"E0",X"00",X"00",X"00",X"00",
		X"E0",X"A0",X"A0",X"E0",X"00",X"00",X"00",X"00",X"E0",X"0A",X"00",X"E0",X"00",X"00",X"00",X"00",
		X"E0",X"A0",X"A0",X"E0",X"00",X"00",X"00",X"00",X"EA",X"00",X"0A",X"E0",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"0E",X"A0",X"00",X"00",X"AE",X"00",X"00",X"00",X"0E",
		X"0A",X"00",X"0A",X"0E",X"00",X"00",X"00",X"0E",X"00",X"A0",X"A0",X"0E",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"A0",X"A0",X"0E",X"00",X"00",X"00",X"0E",
		X"0A",X"00",X"0A",X"0E",X"00",X"00",X"00",X"0E",X"A0",X"00",X"00",X"AE",X"00",X"00",X"00",X"0E",
		X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"00",X"EE",X"E0",X"0E",X"E0",X"00",X"00",X"EA",X"00",X"00",X"00",X"0A",X"E0",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"E0",X"E0",X"00",X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"E0",
		X"00",X"E0",X"E0",X"00",X"E0",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"0A",X"E0",X"00",X"00",X"EE",
		X"00",X"EE",X"E0",X"0E",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",
		X"00",X"EE",X"E0",X"00",X"EE",X"00",X"0E",X"A0",X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"0E",X"A0",X"00",X"00",X"00",X"00",X"AE",X"00",X"0E",X"E0",
		X"00",X"EE",X"E0",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E0",X"0A",X"00",X"00",X"0E",X"00",X"00",X"0A",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"0E",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"E0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"0E",X"00",X"00",X"0A",X"00",X"E0",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"19",X"09",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"06",X"60",X"00",X"66",X"01",X"00",X"01",X"06",X"06",X"06",X"06",X"01",X"00",X"01",X"00",X"66",
		X"66",X"60",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"00",X"09",X"77",X"79",X"77",X"79",X"77",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"70",
		X"07",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"79",X"77",X"79",X"77",X"70",X"00",X"00",X"00",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"19",X"09",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"06",X"06",X"06",X"66",X"01",X"00",X"01",X"06",X"06",X"00",X"00",X"01",X"00",X"01",X"06",X"06",
		X"66",X"66",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"00",X"07",X"97",X"77",X"97",X"77",X"97",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"70",
		X"07",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"97",X"77",X"97",X"77",X"90",X"00",X"00",X"00",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"00",X"66",X"06",X"60",X"01",X"00",X"01",X"06",X"06",X"06",X"06",X"01",X"00",X"01",X"06",X"60",
		X"60",X"66",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"00",X"07",X"79",X"77",X"79",X"77",X"79",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"70",
		X"09",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"77",X"79",X"77",X"79",X"70",X"00",X"00",X"00",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"01",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",
		X"06",X"66",X"06",X"06",X"01",X"00",X"01",X"00",X"00",X"06",X"06",X"01",X"00",X"01",X"06",X"66",
		X"66",X"06",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"11",X"11",X"11",
		X"11",X"00",X"07",X"77",X"97",X"77",X"97",X"77",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"90",
		X"07",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"77",X"97",X"77",X"97",X"70",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"57",X"03",X"35",X"06",X"DE",X"15",X"ED",X"47",X"BD",X"D0",X"54",X"59",X"B0",X"86",X"EF",
		X"8E",X"3B",X"80",X"10",X"8E",X"5A",X"82",X"AF",X"49",X"10",X"AF",X"4B",X"A7",X"4D",X"86",X"01",
		X"8E",X"57",X"26",X"7E",X"D0",X"66",X"AE",X"49",X"10",X"AE",X"4B",X"A6",X"4D",X"C6",X"02",X"E7",
		X"4E",X"BD",X"5A",X"11",X"4D",X"27",X"1A",X"81",X"12",X"26",X"04",X"86",X"EF",X"20",X"12",X"81",
		X"F1",X"26",X"04",X"86",X"DE",X"20",X"0A",X"81",X"23",X"26",X"04",X"86",X"F1",X"20",X"02",X"80",
		X"22",X"8C",X"06",X"16",X"27",X"0E",X"30",X"89",X"FE",X"FE",X"31",X"A9",X"01",X"02",X"6A",X"4E",
		X"26",X"CF",X"20",X"B3",X"4D",X"27",X"03",X"4F",X"20",X"A6",X"6E",X"D8",X"07",X"59",X"84",X"1F",
		X"00",X"59",X"00",X"3F",X"00",X"58",X"A8",X"3F",X"00",X"57",X"9D",X"0F",X"00",X"57",X"B5",X"0F",
		X"00",X"57",X"CD",X"0F",X"00",X"57",X"E9",X"0F",X"00",X"58",X"39",X"1F",X"00",X"58",X"6B",X"1F",
		X"00",X"58",X"91",X"0F",X"00",X"58",X"07",X"1F",X"00",X"59",X"58",X"1F",X"00",X"01",X"02",X"03",
		X"04",X"05",X"06",X"07",X"0F",X"17",X"1F",X"2D",X"34",X"3A",X"7A",X"BA",X"FA",X"F8",X"F0",X"E0",
		X"D0",X"C0",X"C0",X"00",X"00",X"C0",X"C0",X"D0",X"E0",X"F0",X"F8",X"FA",X"BA",X"7A",X"3A",X"34",
		X"2D",X"1F",X"17",X"0F",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"00",X"C0",X"C1",X"C2",
		X"C3",X"C4",X"C5",X"C6",X"C7",X"87",X"87",X"47",X"47",X"07",X"07",X"47",X"47",X"87",X"87",X"C7",
		X"C7",X"C6",X"C5",X"C4",X"C3",X"C2",X"C1",X"00",X"00",X"38",X"38",X"31",X"3A",X"3B",X"3C",X"2D",
		X"2E",X"2F",X"27",X"1F",X"17",X"17",X"0F",X"07",X"07",X"0F",X"17",X"17",X"1F",X"27",X"2F",X"2E",
		X"2D",X"2C",X"3B",X"3A",X"39",X"00",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"37",
		X"2F",X"27",X"17",X"0F",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"01",X"01",X"49",X"CA",X"DA",
		X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"C0",X"C0",X"C0",X"07",X"07",X"38",
		X"38",X"38",X"07",X"C0",X"38",X"FF",X"FF",X"00",X"00",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",
		X"CA",X"DA",X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"C0",X"C0",X"C0",X"07",
		X"07",X"38",X"38",X"38",X"07",X"C0",X"38",X"FF",X"FF",X"00",X"00",X"38",X"39",X"3A",X"3B",X"3C",
		X"3D",X"3E",X"3F",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",
		X"CC",X"CB",X"CA",X"DA",X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"3C",X"00",
		X"00",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",
		X"CA",X"C0",X"D0",X"98",X"38",X"33",X"00",X"00",X"07",X"0F",X"17",X"1F",X"27",X"2F",X"37",X"3F",
		X"3F",X"7F",X"7F",X"BF",X"BF",X"FF",X"FF",X"FF",X"BF",X"BF",X"7F",X"7F",X"3F",X"3F",X"3E",X"3D",
		X"3C",X"3B",X"3A",X"39",X"38",X"38",X"30",X"28",X"20",X"08",X"08",X"49",X"52",X"A5",X"FB",X"FC",
		X"FD",X"FE",X"FF",X"FF",X"FE",X"FD",X"FC",X"FB",X"FA",X"F9",X"F8",X"F0",X"E8",X"E0",X"D8",X"D0",
		X"C8",X"C0",X"80",X"40",X"01",X"01",X"01",X"01",X"02",X"03",X"04",X"05",X"06",X"4F",X"EF",X"F7",
		X"FF",X"FF",X"F7",X"EF",X"E7",X"DF",X"D7",X"CF",X"C7",X"87",X"87",X"47",X"47",X"07",X"00",X"00",
		X"07",X"0F",X"17",X"1F",X"27",X"2F",X"37",X"3F",X"3F",X"7F",X"7F",X"BF",X"BF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"7F",X"7F",X"3F",X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"38",X"78",X"78",
		X"B8",X"B8",X"F8",X"F8",X"F9",X"FA",X"FB",X"FC",X"FD",X"FE",X"FF",X"FF",X"FE",X"FD",X"FC",X"FB",
		X"FA",X"F9",X"F8",X"F0",X"E8",X"E0",X"D8",X"D0",X"C8",X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",
		X"C7",X"C7",X"CF",X"D7",X"DF",X"E7",X"EF",X"F7",X"FF",X"FF",X"F7",X"EF",X"E7",X"DF",X"D7",X"CF",
		X"C7",X"87",X"87",X"47",X"47",X"07",X"00",X"00",X"07",X"0F",X"17",X"1F",X"27",X"2F",X"37",X"3F",
		X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",X"38",X"78",X"78",X"B8",X"B8",X"F8",X"F8",X"F0",X"E8",
		X"E0",X"D8",X"D0",X"C8",X"C0",X"80",X"41",X"01",X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"07",
		X"07",X"07",X"00",X"00",X"07",X"0F",X"17",X"1F",X"27",X"2F",X"37",X"3F",X"3E",X"3D",X"3C",X"3B",
		X"3A",X"39",X"38",X"38",X"78",X"78",X"B8",X"B8",X"F8",X"F8",X"F0",X"E8",X"E0",X"D8",X"D0",X"C8",
		X"C0",X"C1",X"C2",X"C3",X"C4",X"C5",X"C6",X"C7",X"C7",X"87",X"87",X"47",X"47",X"07",X"00",X"00",
		X"10",X"8E",X"57",X"6D",X"BD",X"D0",X"39",X"84",X"0F",X"81",X"0C",X"24",X"F7",X"48",X"48",X"1F",
		X"89",X"AE",X"A5",X"CB",X"02",X"BD",X"D0",X"39",X"A4",X"A5",X"AF",X"47",X"30",X"86",X"AF",X"49",
		X"AE",X"49",X"30",X"01",X"6D",X"84",X"26",X"02",X"AE",X"47",X"AF",X"49",X"10",X"8E",X"98",X"01",
		X"A6",X"80",X"26",X"04",X"AE",X"47",X"20",X"F8",X"A7",X"A0",X"10",X"8C",X"98",X"10",X"25",X"F0",
		X"C6",X"00",X"A6",X"4B",X"4A",X"81",X"05",X"25",X"02",X"86",X"04",X"A7",X"4B",X"8E",X"98",X"01",
		X"E7",X"86",X"30",X"05",X"8C",X"98",X"10",X"25",X"F7",X"86",X"01",X"8E",X"59",X"D0",X"7E",X"D0",
		X"66",X"34",X"76",X"84",X"F0",X"97",X"CC",X"A6",X"E4",X"84",X"0F",X"97",X"CD",X"1F",X"10",X"97",
		X"CA",X"D7",X"C8",X"1F",X"20",X"97",X"CB",X"D7",X"C9",X"D0",X"C8",X"56",X"24",X"02",X"0A",X"C9",
		X"BD",X"5A",X"C3",X"96",X"C8",X"BD",X"5A",X"89",X"4C",X"BD",X"5A",X"CC",X"8D",X"6C",X"96",X"C9",
		X"BD",X"5A",X"C3",X"8D",X"44",X"4A",X"BD",X"5A",X"CC",X"8D",X"5F",X"96",X"CA",X"BD",X"5A",X"D5",
		X"8D",X"09",X"96",X"CB",X"BD",X"5A",X"DA",X"8D",X"02",X"35",X"F6",X"34",X"17",X"8D",X"1C",X"1A",
		X"10",X"B7",X"CA",X"01",X"86",X"05",X"C8",X"04",X"FD",X"CA",X"06",X"CC",X"00",X"00",X"FD",X"CA",
		X"02",X"BF",X"CA",X"04",X"86",X"12",X"B7",X"CA",X"00",X"35",X"97",X"34",X"04",X"D6",X"C8",X"5C",
		X"1F",X"01",X"D6",X"C9",X"D0",X"C8",X"5A",X"35",X"82",X"34",X"17",X"8D",X"28",X"5C",X"1A",X"10",
		X"B7",X"CA",X"01",X"C8",X"04",X"F7",X"CA",X"06",X"86",X"05",X"B7",X"CA",X"07",X"FD",X"CA",X"02",
		X"BF",X"CA",X"04",X"86",X"12",X"B7",X"CA",X"00",X"35",X"97",X"34",X"17",X"8D",X"07",X"5A",X"30",
		X"89",X"01",X"00",X"20",X"D9",X"34",X"04",X"1F",X"89",X"96",X"CA",X"1F",X"01",X"D6",X"CB",X"D0",
		X"CA",X"35",X"82",X"D6",X"CC",X"54",X"54",X"54",X"54",X"DA",X"CC",X"39",X"D6",X"CD",X"58",X"58",
		X"58",X"58",X"DA",X"CD",X"39",X"D6",X"CC",X"DA",X"CD",X"39",X"D6",X"CC",X"54",X"54",X"54",X"54",
		X"34",X"04",X"D6",X"CD",X"58",X"58",X"58",X"58",X"EA",X"E0",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"5B",X"5E",X"7E",X"5C",X"1F",X"7E",X"5B",X"C6",X"7E",X"5E",X"15",X"7E",X"5E",X"38",X"7E",
		X"5C",X"0A",X"7E",X"5C",X"14",X"7E",X"5B",X"98",X"7E",X"5B",X"B1",X"7E",X"5B",X"BB",X"0F",X"96",
		X"0F",X"97",X"0F",X"98",X"0F",X"99",X"BD",X"F0",X"09",X"7E",X"46",X"80",X"34",X"10",X"DE",X"1B",
		X"27",X"0E",X"AE",X"C4",X"9F",X"1B",X"9E",X"96",X"AF",X"C4",X"DF",X"96",X"1C",X"FE",X"35",X"90",
		X"1A",X"01",X"35",X"90",X"34",X"10",X"DE",X"1B",X"27",X"F6",X"AE",X"C4",X"9F",X"1B",X"9E",X"98",
		X"AF",X"C4",X"DF",X"98",X"1C",X"FE",X"35",X"90",X"34",X"76",X"8D",X"E8",X"25",X"6A",X"ED",X"49",
		X"CC",X"0E",X"0E",X"ED",X"C8",X"10",X"20",X"30",X"34",X"02",X"B6",X"CC",X"13",X"84",X"0F",X"35",
		X"82",X"8D",X"F5",X"10",X"26",X"94",X"58",X"34",X"76",X"20",X"0D",X"8D",X"EB",X"10",X"26",X"94",
		X"4B",X"34",X"76",X"7E",X"5C",X"3A",X"34",X"76",X"8D",X"BA",X"25",X"3C",X"CC",X"0A",X"0A",X"ED",
		X"C8",X"10",X"EC",X"04",X"ED",X"49",X"AE",X"02",X"D6",X"A7",X"E7",X"44",X"E0",X"4A",X"25",X"04",
		X"E1",X"01",X"25",X"0B",X"E6",X"84",X"54",X"E7",X"45",X"EB",X"4A",X"E7",X"44",X"20",X"02",X"E7",
		X"45",X"EC",X"84",X"ED",X"4B",X"C6",X"01",X"E7",X"4F",X"88",X"04",X"C8",X"04",X"ED",X"4D",X"AE",
		X"02",X"AF",X"42",X"CC",X"10",X"00",X"ED",X"46",X"35",X"F6",X"CC",X"01",X"00",X"DD",X"88",X"8D",
		X"0E",X"7E",X"5B",X"5B",X"CC",X"01",X"01",X"DD",X"88",X"8D",X"04",X"86",X"FF",X"97",X"88",X"34",
		X"76",X"96",X"88",X"26",X"07",X"BD",X"5B",X"5B",X"24",X"7D",X"20",X"13",X"D6",X"89",X"27",X"0A",
		X"98",X"89",X"43",X"BD",X"46",X"83",X"24",X"6F",X"20",X"05",X"BD",X"5B",X"6C",X"24",X"0A",X"10",
		X"AE",X"02",X"EC",X"04",X"BD",X"D0",X"1E",X"20",X"5E",X"EC",X"04",X"AE",X"02",X"ED",X"49",X"CC",
		X"0A",X"0A",X"ED",X"C8",X"10",X"D6",X"A7",X"E7",X"44",X"E0",X"4A",X"25",X"04",X"E1",X"01",X"25",
		X"0B",X"E6",X"01",X"54",X"E7",X"45",X"EB",X"4A",X"E7",X"44",X"20",X"02",X"E7",X"45",X"10",X"8E",
		X"C3",X"A5",X"EC",X"84",X"ED",X"4B",X"E7",X"4F",X"C6",X"01",X"88",X"04",X"C8",X"04",X"ED",X"4D",
		X"96",X"59",X"2B",X"16",X"A6",X"A9",X"FA",X"CD",X"81",X"4A",X"27",X"0E",X"96",X"86",X"26",X"0A",
		X"D6",X"85",X"86",X"98",X"34",X"06",X"EF",X"F4",X"35",X"06",X"AE",X"02",X"AF",X"42",X"CC",X"01",
		X"00",X"ED",X"46",X"86",X"10",X"A7",X"48",X"35",X"F6",X"E6",X"2F",X"C0",X"10",X"50",X"86",X"06",
		X"3D",X"BE",X"F0",X"17",X"3A",X"34",X"10",X"A6",X"26",X"97",X"A8",X"A6",X"29",X"C6",X"12",X"1A",
		X"10",X"B7",X"CA",X"04",X"A6",X"2A",X"CE",X"00",X"00",X"FF",X"CA",X"01",X"B7",X"CA",X"03",X"EE",
		X"2D",X"FF",X"CA",X"06",X"CE",X"CA",X"05",X"8E",X"CA",X"00",X"39",X"CE",X"98",X"96",X"10",X"AC",
		X"C4",X"27",X"08",X"EE",X"C4",X"26",X"F7",X"1A",X"10",X"20",X"FE",X"EC",X"A4",X"ED",X"C4",X"DC",
		X"1B",X"ED",X"A4",X"10",X"9F",X"1B",X"31",X"C4",X"39",X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",
		X"4F",X"4E",X"3A",X"20",X"32",X"30",X"38",X"34",X"20",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",
		X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",
		X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",
		X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",
		X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"EC",X"26",X"83",X"00",X"80",X"A1",X"26",X"26",
		X"03",X"E7",X"27",X"39",X"BD",X"5C",X"A9",X"96",X"59",X"26",X"08",X"DC",X"5E",X"A7",X"29",X"EB",
		X"25",X"E7",X"24",X"A6",X"2C",X"97",X"9C",X"EC",X"26",X"81",X"01",X"22",X"08",X"8D",X"27",X"CE",
		X"98",X"98",X"7E",X"5C",X"DE",X"83",X"00",X"80",X"81",X"01",X"22",X"1A",X"A6",X"A8",X"10",X"81",
		X"0E",X"26",X"EC",X"86",X"01",X"20",X"0F",X"6A",X"28",X"10",X"27",X"FF",X"4E",X"A6",X"2C",X"97",
		X"9C",X"EC",X"26",X"C3",X"01",X"00",X"97",X"A8",X"ED",X"26",X"44",X"E6",X"25",X"26",X"01",X"4F",
		X"97",X"9F",X"AE",X"22",X"96",X"A8",X"E6",X"25",X"3D",X"DD",X"9D",X"E6",X"24",X"4F",X"93",X"9D",
		X"DB",X"9F",X"89",X"00",X"26",X"04",X"C1",X"18",X"22",X"16",X"0A",X"9C",X"DB",X"A8",X"89",X"00",
		X"26",X"F8",X"C1",X"18",X"23",X"F4",X"E7",X"2A",X"EC",X"2B",X"D0",X"9C",X"3D",X"3A",X"20",X"02",
		X"E7",X"2A",X"96",X"9C",X"4A",X"D6",X"A8",X"3D",X"EB",X"2A",X"89",X"00",X"27",X"08",X"0A",X"9C",
		X"D0",X"A8",X"82",X"00",X"26",X"F8",X"C1",X"EA",X"24",X"F4",X"96",X"9C",X"10",X"27",X"FE",X"EB",
		X"A7",X"2F",X"80",X"10",X"40",X"C6",X"0B",X"3D",X"F3",X"F0",X"15",X"34",X"26",X"EE",X"A8",X"10",
		X"EC",X"2D",X"1A",X"10",X"FD",X"CA",X"06",X"A6",X"29",X"B7",X"CA",X"04",X"E6",X"2B",X"A6",X"2A",
		X"10",X"8E",X"CA",X"05",X"39",X"10",X"9E",X"96",X"27",X"0B",X"BD",X"5C",X"A9",X"BD",X"5D",X"87",
		X"10",X"AE",X"A4",X"26",X"F5",X"10",X"9E",X"98",X"27",X"08",X"BD",X"5D",X"48",X"10",X"AE",X"A4",
		X"26",X"F8",X"BD",X"F0",X"12",X"7E",X"46",X"89",X"DE",X"15",X"35",X"06",X"ED",X"4D",X"86",X"0A",
		X"A7",X"47",X"8E",X"98",X"5A",X"BD",X"D0",X"15",X"8E",X"98",X"5A",X"86",X"99",X"BD",X"38",X"88",
		X"86",X"02",X"8E",X"5E",X"58",X"7E",X"D0",X"66",X"96",X"84",X"84",X"03",X"8E",X"5E",X"AE",X"A6",
		X"86",X"8E",X"98",X"5A",X"BD",X"38",X"88",X"6A",X"47",X"27",X"08",X"86",X"06",X"8E",X"5E",X"48",
		X"7E",X"D0",X"66",X"BD",X"D0",X"60",X"BD",X"D0",X"24",X"BD",X"D0",X"5D",X"DE",X"15",X"8E",X"5E",
		X"B2",X"AF",X"47",X"8E",X"98",X"5A",X"86",X"CC",X"BD",X"38",X"88",X"AE",X"47",X"A6",X"80",X"97",
		X"0C",X"27",X"0A",X"AF",X"47",X"86",X"04",X"8E",X"5E",X"8B",X"7E",X"D0",X"66",X"8E",X"98",X"5A",
		X"6F",X"88",X"12",X"BD",X"D0",X"15",X"BD",X"D0",X"24",X"DE",X"15",X"6E",X"D8",X"0D",X"00",X"11",
		X"33",X"77",X"FF",X"F6",X"AD",X"A4",X"5B",X"52",X"09",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"5F",X"BE",X"7E",X"60",X"23",X"7E",X"61",X"3F",X"7E",X"61",X"47",X"7E",X"5F",X"A2",X"7E",
		X"60",X"96",X"34",X"02",X"86",X"11",X"97",X"CF",X"35",X"02",X"34",X"02",X"86",X"07",X"97",X"D2",
		X"0F",X"D0",X"0F",X"D5",X"0F",X"D7",X"86",X"01",X"97",X"D1",X"9F",X"D3",X"35",X"82",X"34",X"66",
		X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"05",X"D7",X"D2",X"81",X"20",X"26",X"02",X"86",X"3A",X"10",
		X"BE",X"E9",X"C8",X"81",X"5E",X"22",X"4A",X"80",X"30",X"25",X"46",X"48",X"10",X"AE",X"A6",X"A6",
		X"A4",X"44",X"4C",X"88",X"04",X"C6",X"01",X"34",X"21",X"1A",X"10",X"FD",X"CA",X"06",X"31",X"21",
		X"10",X"BF",X"CA",X"02",X"96",X"CF",X"B7",X"CA",X"01",X"BF",X"CA",X"04",X"86",X"1A",X"D6",X"D0",
		X"27",X"02",X"86",X"3A",X"B7",X"CA",X"00",X"35",X"21",X"A6",X"A4",X"4C",X"5F",X"44",X"30",X"8B",
		X"24",X"0F",X"96",X"D0",X"27",X"07",X"30",X"89",X"01",X"00",X"5F",X"20",X"02",X"C6",X"FF",X"D7",
		X"D0",X"35",X"E6",X"34",X"66",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"07",X"D7",X"D2",X"81",X"20",
		X"26",X"02",X"86",X"3A",X"10",X"BE",X"E9",X"CA",X"81",X"5E",X"22",X"E5",X"80",X"30",X"25",X"E1",
		X"48",X"10",X"AE",X"A6",X"A6",X"A4",X"44",X"4C",X"88",X"04",X"D6",X"D7",X"2F",X"01",X"50",X"CB",
		X"06",X"C8",X"04",X"34",X"21",X"1A",X"10",X"FD",X"CA",X"06",X"31",X"21",X"D6",X"D7",X"2F",X"05",
		X"88",X"04",X"3D",X"31",X"A5",X"10",X"BF",X"CA",X"02",X"96",X"CF",X"B7",X"CA",X"01",X"BF",X"CA",
		X"04",X"86",X"1A",X"D6",X"D0",X"27",X"8D",X"20",X"89",X"0F",X"D0",X"34",X"66",X"86",X"05",X"5F",
		X"20",X"2F",X"0F",X"D0",X"34",X"66",X"86",X"05",X"C6",X"01",X"20",X"25",X"0F",X"D0",X"34",X"66",
		X"86",X"07",X"C6",X"01",X"20",X"1B",X"0F",X"D0",X"34",X"66",X"C6",X"07",X"D7",X"D2",X"C6",X"02",
		X"D7",X"D1",X"8D",X"65",X"A6",X"E4",X"8D",X"65",X"35",X"E6",X"0F",X"D0",X"34",X"66",X"86",X"07",
		X"5F",X"97",X"D2",X"D7",X"D1",X"A6",X"E4",X"20",X"02",X"34",X"66",X"0F",X"D6",X"8D",X"4A",X"0C",
		X"D6",X"A6",X"E4",X"8D",X"48",X"35",X"E6",X"0F",X"D0",X"34",X"66",X"86",X"05",X"5F",X"20",X"1B",
		X"0F",X"D0",X"34",X"66",X"86",X"05",X"C6",X"01",X"20",X"11",X"0F",X"D0",X"34",X"66",X"86",X"07",
		X"C6",X"01",X"20",X"07",X"0F",X"D0",X"34",X"66",X"86",X"07",X"5F",X"97",X"D2",X"D7",X"D1",X"A6",
		X"E4",X"20",X"02",X"34",X"66",X"0F",X"D6",X"8D",X"10",X"A6",X"E4",X"8D",X"10",X"A6",X"61",X"8D",
		X"08",X"0C",X"D6",X"A6",X"61",X"8D",X"06",X"35",X"E6",X"44",X"44",X"44",X"44",X"84",X"0F",X"26",
		X"08",X"D6",X"D6",X"26",X"04",X"D6",X"D1",X"26",X"0F",X"0C",X"D6",X"8B",X"30",X"D6",X"D2",X"C1",
		X"07",X"10",X"27",X"FE",X"FE",X"7E",X"5F",X"BE",X"C1",X"02",X"26",X"0E",X"30",X"89",X"02",X"00",
		X"D6",X"D2",X"C1",X"05",X"27",X"04",X"30",X"89",X"01",X"00",X"39",X"34",X"66",X"20",X"12",X"0F",
		X"D0",X"34",X"66",X"C6",X"05",X"20",X"06",X"0F",X"D0",X"34",X"66",X"C6",X"07",X"D7",X"D2",X"0F",
		X"D7",X"34",X"42",X"CE",X"99",X"4B",X"C6",X"37",X"0D",X"59",X"2B",X"13",X"E1",X"C8",X"A8",X"27",
		X"0E",X"96",X"85",X"81",X"30",X"22",X"08",X"D6",X"84",X"86",X"98",X"1F",X"03",X"63",X"C4",X"35",
		X"42",X"1F",X"89",X"4F",X"58",X"49",X"10",X"8E",X"62",X"91",X"10",X"AE",X"AB",X"A6",X"A0",X"27",
		X"1F",X"81",X"17",X"24",X"0B",X"4A",X"48",X"CE",X"61",X"A2",X"EE",X"C6",X"AD",X"C4",X"20",X"ED",
		X"D6",X"D2",X"C1",X"07",X"26",X"05",X"BD",X"60",X"23",X"20",X"E2",X"BD",X"5F",X"BE",X"20",X"DD",
		X"35",X"E6",X"61",X"D8",X"61",X"D8",X"61",X"D8",X"61",X"D9",X"61",X"DE",X"62",X"16",X"62",X"1D",
		X"62",X"2A",X"62",X"37",X"62",X"3C",X"62",X"44",X"62",X"49",X"62",X"4E",X"62",X"53",X"62",X"75",
		X"62",X"58",X"62",X"6B",X"62",X"0F",X"62",X"70",X"61",X"CE",X"62",X"3F",X"62",X"5D",X"B6",X"C8",
		X"06",X"10",X"2B",X"00",X"A0",X"EC",X"A1",X"39",X"39",X"A6",X"A0",X"97",X"CF",X"39",X"1F",X"10",
		X"AB",X"A4",X"EB",X"21",X"1F",X"01",X"6D",X"22",X"27",X"22",X"6D",X"A4",X"2B",X"0F",X"96",X"D0",
		X"27",X"06",X"30",X"89",X"01",X"00",X"86",X"FF",X"4C",X"97",X"D0",X"20",X"0F",X"96",X"D0",X"81",
		X"01",X"27",X"06",X"30",X"89",X"FF",X"00",X"86",X"02",X"4A",X"97",X"D0",X"31",X"23",X"39",X"AE",
		X"A1",X"A6",X"A0",X"97",X"D0",X"39",X"D6",X"D0",X"D7",X"D5",X"9F",X"D3",X"39",X"96",X"D2",X"81",
		X"07",X"27",X"06",X"86",X"07",X"97",X"D2",X"30",X"1F",X"39",X"96",X"D2",X"81",X"05",X"27",X"F9",
		X"86",X"05",X"97",X"D2",X"30",X"01",X"39",X"86",X"01",X"97",X"D1",X"39",X"0F",X"D1",X"39",X"86",
		X"02",X"97",X"D1",X"39",X"EC",X"A1",X"7E",X"60",X"F3",X"EC",X"B1",X"7E",X"60",X"F3",X"A6",X"A0",
		X"7E",X"60",X"B9",X"A6",X"B1",X"7E",X"60",X"B9",X"A6",X"63",X"7E",X"60",X"B9",X"A6",X"63",X"81",
		X"05",X"23",X"05",X"81",X"FB",X"24",X"01",X"4F",X"97",X"D7",X"39",X"EC",X"64",X"7E",X"60",X"F3",
		X"A6",X"B1",X"97",X"CF",X"39",X"32",X"78",X"E6",X"6B",X"E7",X"61",X"EC",X"6C",X"ED",X"62",X"CC",
		X"62",X"8E",X"ED",X"66",X"EC",X"A1",X"10",X"AF",X"64",X"1F",X"02",X"7E",X"61",X"7D",X"1F",X"32",
		X"39",X"6D",X"1B",X"6C",X"D1",X"6D",X"58",X"6D",X"4D",X"6B",X"B4",X"6B",X"FC",X"6C",X"08",X"6C",
		X"25",X"6C",X"2F",X"6C",X"8A",X"6D",X"37",X"6D",X"42",X"6B",X"A2",X"6A",X"D0",X"6A",X"D8",X"6A",
		X"E0",X"6A",X"EB",X"6A",X"FC",X"6B",X"06",X"6B",X"12",X"6B",X"1E",X"6B",X"29",X"6B",X"36",X"6B",
		X"43",X"6B",X"51",X"6B",X"56",X"6B",X"65",X"6B",X"70",X"6B",X"7D",X"6B",X"8A",X"6A",X"9B",X"69",
		X"62",X"6A",X"5C",X"6A",X"6C",X"6A",X"7E",X"69",X"9E",X"69",X"B3",X"69",X"CC",X"69",X"E9",X"69",
		X"FC",X"6D",X"E4",X"69",X"55",X"69",X"58",X"69",X"5B",X"67",X"90",X"67",X"96",X"68",X"14",X"68",
		X"24",X"68",X"32",X"68",X"44",X"68",X"4C",X"68",X"56",X"68",X"6B",X"68",X"75",X"68",X"85",X"68",
		X"B6",X"68",X"C9",X"68",X"DC",X"68",X"FF",X"69",X"0A",X"69",X"13",X"69",X"2A",X"69",X"35",X"69",
		X"4E",X"65",X"4C",X"65",X"5B",X"65",X"9F",X"65",X"A2",X"65",X"B9",X"65",X"BF",X"65",X"D5",X"66",
		X"14",X"66",X"18",X"66",X"1B",X"66",X"2C",X"6D",X"F2",X"66",X"33",X"66",X"3A",X"65",X"6E",X"66",
		X"EB",X"67",X"49",X"65",X"F0",X"66",X"51",X"66",X"73",X"66",X"85",X"66",X"9C",X"66",X"AC",X"66",
		X"C1",X"66",X"D0",X"66",X"E1",X"66",X"41",X"69",X"6E",X"64",X"28",X"69",X"7F",X"64",X"A6",X"64",
		X"FD",X"65",X"29",X"65",X"3C",X"65",X"42",X"65",X"45",X"64",X"35",X"63",X"CF",X"65",X"82",X"6E",
		X"01",X"6E",X"0B",X"6C",X"C4",X"6A",X"13",X"6A",X"33",X"6A",X"37",X"6A",X"58",X"63",X"95",X"63",
		X"CA",X"6D",X"6C",X"6D",X"B7",X"6E",X"1F",X"6E",X"28",X"6E",X"3B",X"6E",X"41",X"6E",X"2E",X"6E",
		X"47",X"6E",X"5B",X"6E",X"7D",X"6E",X"99",X"66",X"66",X"6E",X"BD",X"68",X"05",X"63",X"BB",X"6D",
		X"AD",X"6E",X"C8",X"6E",X"DD",X"04",X"77",X"12",X"35",X"25",X"00",X"0F",X"63",X"BC",X"45",X"53",
		X"12",X"35",X"6E",X"00",X"41",X"4C",X"4C",X"20",X"05",X"00",X"00",X"01",X"54",X"49",X"4D",X"45",
		X"20",X"05",X"01",X"00",X"00",X"48",X"45",X"52",X"4F",X"45",X"53",X"00",X"52",X"4F",X"42",X"4F",
		X"54",X"52",X"4F",X"4E",X"20",X"48",X"45",X"52",X"4F",X"00",X"15",X"10",X"5C",X"3A",X"00",X"04",
		X"99",X"12",X"25",X"70",X"01",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"54",X"48",X"45",X"20",
		X"4C",X"49",X"4E",X"45",X"20",X"55",X"53",X"49",X"4E",X"47",X"20",X"40",X"46",X"49",X"52",X"45",
		X"40",X"12",X"24",X"7E",X"01",X"0F",X"64",X"0E",X"57",X"48",X"45",X"4E",X"20",X"43",X"45",X"4E",
		X"54",X"45",X"52",X"45",X"44",X"04",X"BB",X"08",X"12",X"49",X"50",X"01",X"3E",X"00",X"50",X"52",
		X"45",X"53",X"53",X"20",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"00",X"0F",X"64",X"0E",
		X"54",X"4F",X"20",X"45",X"58",X"49",X"54",X"00",X"04",X"BB",X"12",X"2E",X"16",X"00",X"0F",X"69",
		X"39",X"0F",X"64",X"69",X"00",X"04",X"BB",X"12",X"20",X"70",X"00",X"35",X"20",X"45",X"4E",X"54",
		X"52",X"49",X"45",X"53",X"20",X"4D",X"41",X"58",X"49",X"4D",X"55",X"4D",X"0F",X"68",X"29",X"12",
		X"28",X"90",X"01",X"4C",X"4F",X"57",X"45",X"53",X"54",X"20",X"45",X"4E",X"54",X"52",X"59",X"20",
		X"52",X"45",X"50",X"4C",X"41",X"43",X"45",X"44",X"00",X"08",X"04",X"99",X"12",X"2F",X"C0",X"01",
		X"0F",X"67",X"EF",X"4C",X"45",X"54",X"54",X"45",X"52",X"12",X"32",X"CC",X"00",X"40",X"46",X"49",
		X"52",X"45",X"20",X"55",X"50",X"40",X"20",X"54",X"4F",X"20",X"45",X"4E",X"54",X"45",X"52",X"20",
		X"4C",X"45",X"54",X"54",X"45",X"52",X"04",X"44",X"00",X"00",X"12",X"40",X"10",X"00",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"00",X"04",X"BB",X"0F",X"64",X"9A",X"09",X"11",X"12",X"2C",X"28",
		X"00",X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",X"54",X"48",X"45",X"20",X"47",X"52",X"45",
		X"41",X"54",X"45",X"53",X"54",X"12",X"36",X"38",X"00",X"0F",X"63",X"BC",X"12",X"34",X"58",X"00",
		X"0F",X"64",X"F1",X"4E",X"41",X"4D",X"45",X"12",X"31",X"68",X"00",X"5B",X"55",X"50",X"20",X"54",
		X"4F",X"20",X"09",X"10",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"53",X"5C",X"0F",X"64",X"69",
		X"00",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"00",X"04",X"44",X"0F",
		X"64",X"9A",X"09",X"10",X"12",X"29",X"30",X"00",X"59",X"4F",X"55",X"20",X"41",X"52",X"45",X"20",
		X"41",X"20",X"0F",X"63",X"BC",X"12",X"2D",X"58",X"01",X"0F",X"64",X"F1",X"49",X"4E",X"49",X"54",
		X"49",X"41",X"4C",X"53",X"3F",X"0F",X"64",X"69",X"00",X"04",X"99",X"0F",X"64",X"9A",X"09",X"10",
		X"12",X"43",X"67",X"00",X"41",X"4C",X"53",X"4F",X"0F",X"65",X"15",X"00",X"15",X"10",X"5C",X"3A",
		X"3A",X"00",X"15",X"11",X"00",X"05",X"08",X"00",X"00",X"15",X"11",X"00",X"15",X"10",X"30",X"30",
		X"30",X"20",X"20",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"00",X"15",X"10",X"30",X"30",X"30",
		X"20",X"20",X"52",X"45",X"43",X"4F",X"4D",X"4D",X"45",X"4E",X"44",X"45",X"44",X"00",X"15",X"10",
		X"30",X"30",X"30",X"20",X"20",X"43",X"4F",X"4E",X"53",X"45",X"52",X"56",X"41",X"54",X"49",X"56",
		X"45",X"00",X"15",X"10",X"30",X"30",X"30",X"20",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"0F",
		X"65",X"75",X"00",X"05",X"08",X"00",X"00",X"00",X"0F",X"65",X"93",X"0F",X"65",X"62",X"00",X"15",
		X"10",X"00",X"0F",X"66",X"0E",X"48",X"49",X"47",X"48",X"20",X"56",X"4F",X"4C",X"55",X"4D",X"45",
		X"20",X"41",X"52",X"43",X"41",X"44",X"45",X"53",X"00",X"15",X"10",X"0F",X"65",X"98",X"00",X"0F",
		X"66",X"0E",X"46",X"4F",X"52",X"20",X"57",X"45",X"41",X"4B",X"45",X"52",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"53",X"00",X"0F",X"66",X"0E",X"43",X"55",X"53",X"54",X"4F",X"4D",X"20",X"40",
		X"3A",X"5B",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"42",X"45",X"4C",X"4F",X"57",X"5C",X"00",
		X"59",X"45",X"53",X"0F",X"65",X"93",X"05",X"FE",X"00",X"00",X"41",X"44",X"56",X"41",X"4E",X"43",
		X"45",X"20",X"54",X"4F",X"20",X"41",X"43",X"54",X"49",X"56",X"41",X"54",X"45",X"00",X"15",X"10",
		X"0F",X"65",X"93",X"00",X"59",X"45",X"53",X"00",X"4E",X"4F",X"00",X"0F",X"66",X"22",X"0F",X"65",
		X"53",X"00",X"0F",X"66",X"0E",X"45",X"58",X"54",X"52",X"41",X"20",X"00",X"0F",X"66",X"0E",X"0F",
		X"65",X"53",X"00",X"0F",X"66",X"0E",X"0F",X"65",X"75",X"00",X"0F",X"66",X"22",X"0F",X"65",X"75",
		X"00",X"0F",X"66",X"0E",X"4E",X"4F",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",X"45",X"4E",
		X"00",X"0F",X"66",X"0E",X"31",X"5E",X"46",X"49",X"46",X"54",X"59",X"20",X"20",X"33",X"5E",X"44",
		X"4F",X"4C",X"4C",X"41",X"52",X"00",X"0F",X"66",X"0E",X"46",X"52",X"45",X"45",X"20",X"50",X"4C",
		X"41",X"59",X"00",X"0F",X"66",X"0E",X"31",X"5E",X"31",X"20",X"44",X"4D",X"20",X"20",X"36",X"5E",
		X"35",X"20",X"44",X"4D",X"00",X"0F",X"66",X"0E",X"31",X"5E",X"51",X"55",X"41",X"52",X"54",X"45",
		X"52",X"20",X"20",X"34",X"5E",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"00",X"0F",X"66",X"0E",X"31",
		X"5E",X"32",X"20",X"46",X"20",X"20",X"33",X"5E",X"35",X"20",X"46",X"00",X"0F",X"66",X"0E",X"31",
		X"5E",X"46",X"49",X"46",X"54",X"59",X"20",X"20",X"32",X"5E",X"44",X"4F",X"4C",X"4C",X"41",X"52",
		X"00",X"0F",X"66",X"0E",X"31",X"5E",X"32",X"35",X"20",X"20",X"34",X"5E",X"31",X"20",X"47",X"00",
		X"0F",X"66",X"0E",X"31",X"5E",X"35",X"20",X"46",X"20",X"20",X"32",X"5E",X"31",X"30",X"20",X"46",
		X"00",X"0F",X"66",X"0E",X"31",X"5E",X"31",X"30",X"20",X"46",X"00",X"04",X"11",X"12",X"30",X"80",
		X"00",X"0F",X"67",X"E4",X"20",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",X"12",X"20",X"A0",X"00",
		X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"0F",X"67",X"36",X"42",X"59",X"12",X"20",X"B0",X"00",
		X"0F",X"67",X"5C",X"14",X"67",X"6F",X"12",X"20",X"C0",X"00",X"41",X"4E",X"44",X"20",X"54",X"55",
		X"52",X"4E",X"49",X"4E",X"47",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"46",X"46",X"20",X"41",
		X"4E",X"44",X"20",X"4F",X"4E",X"00",X"20",X"46",X"41",X"43",X"54",X"4F",X"52",X"59",X"20",X"53",
		X"45",X"54",X"54",X"49",X"4E",X"47",X"53",X"20",X"00",X"04",X"99",X"12",X"21",X"80",X"00",X"0F",
		X"67",X"36",X"20",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"44",X"00",X"4F",X"50",X"45",X"4E",
		X"49",X"4E",X"47",X"20",X"46",X"52",X"4F",X"4E",X"54",X"20",X"44",X"4F",X"4F",X"52",X"00",X"12",
		X"20",X"B0",X"00",X"04",X"00",X"0F",X"67",X"5C",X"12",X"20",X"B0",X"00",X"04",X"11",X"52",X"41",
		X"49",X"53",X"49",X"4E",X"47",X"20",X"54",X"41",X"42",X"4C",X"45",X"20",X"54",X"4F",X"50",X"00",
		X"04",X"99",X"5D",X"04",X"66",X"00",X"07",X"04",X"99",X"12",X"37",X"0F",X"00",X"47",X"41",X"4D",
		X"45",X"20",X"0F",X"67",X"E4",X"08",X"12",X"2E",X"CD",X"00",X"04",X"99",X"0F",X"67",X"EF",X"0F",
		X"67",X"E4",X"12",X"2B",X"D5",X"00",X"55",X"53",X"45",X"20",X"40",X"46",X"49",X"52",X"45",X"40",
		X"20",X"4C",X"45",X"56",X"45",X"52",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",
		X"20",X"54",X"48",X"45",X"20",X"56",X"41",X"4C",X"55",X"45",X"12",X"39",X"E2",X"00",X"04",X"55",
		X"0F",X"64",X"1D",X"00",X"41",X"44",X"4A",X"55",X"53",X"54",X"4D",X"45",X"4E",X"54",X"00",X"55",
		X"53",X"45",X"20",X"40",X"4D",X"4F",X"56",X"45",X"40",X"20",X"54",X"4F",X"20",X"53",X"45",X"4C",
		X"45",X"43",X"54",X"20",X"00",X"04",X"66",X"12",X"36",X"EE",X"00",X"0F",X"68",X"14",X"3A",X"10",
		X"30",X"30",X"30",X"00",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",X"41",X"4E",X"20",X"45",X"56",
		X"45",X"52",X"59",X"00",X"54",X"55",X"52",X"4E",X"53",X"20",X"50",X"45",X"52",X"20",X"0F",X"64",
		X"9E",X"00",X"50",X"52",X"49",X"43",X"49",X"4E",X"47",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",
		X"49",X"4F",X"4E",X"00",X"4C",X"45",X"46",X"54",X"0F",X"68",X"5F",X"00",X"43",X"45",X"4E",X"54",
		X"45",X"52",X"0F",X"68",X"5F",X"00",X"52",X"49",X"47",X"48",X"54",X"0F",X"68",X"5F",X"00",X"20",
		X"53",X"4C",X"4F",X"54",X"20",X"55",X"4E",X"49",X"54",X"53",X"00",X"0F",X"68",X"A2",X"43",X"52",
		X"45",X"44",X"49",X"54",X"00",X"0F",X"68",X"A2",X"42",X"4F",X"4E",X"55",X"53",X"20",X"43",X"52",
		X"45",X"44",X"49",X"54",X"00",X"4D",X"49",X"4E",X"49",X"4D",X"55",X"4D",X"20",X"55",X"4E",X"49",
		X"54",X"53",X"20",X"46",X"4F",X"52",X"20",X"41",X"4E",X"59",X"20",X"43",X"52",X"45",X"44",X"49",
		X"54",X"00",X"55",X"4E",X"49",X"54",X"53",X"20",X"52",X"45",X"51",X"55",X"49",X"52",X"45",X"44",
		X"20",X"46",X"4F",X"52",X"20",X"00",X"46",X"41",X"4E",X"43",X"59",X"20",X"41",X"54",X"54",X"52",
		X"41",X"43",X"54",X"20",X"4D",X"4F",X"44",X"45",X"00",X"44",X"49",X"46",X"46",X"49",X"43",X"55",
		X"4C",X"54",X"59",X"20",X"4F",X"46",X"20",X"50",X"4C",X"41",X"59",X"00",X"4C",X"45",X"54",X"54",
		X"45",X"52",X"53",X"20",X"46",X"4F",X"52",X"0F",X"68",X"EB",X"00",X"20",X"48",X"49",X"47",X"48",
		X"45",X"53",X"54",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"4E",X"41",X"4D",X"45",X"00",X"52",
		X"45",X"53",X"54",X"4F",X"52",X"45",X"0F",X"67",X"36",X"00",X"43",X"4C",X"45",X"41",X"52",X"0F",
		X"69",X"89",X"00",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"54",X"41",
		X"42",X"4C",X"45",X"20",X"52",X"45",X"53",X"45",X"54",X"00",X"41",X"55",X"54",X"4F",X"20",X"43",
		X"59",X"43",X"4C",X"45",X"00",X"53",X"45",X"54",X"20",X"41",X"54",X"54",X"52",X"41",X"43",X"54",
		X"20",X"4D",X"4F",X"44",X"45",X"20",X"4D",X"45",X"53",X"53",X"41",X"47",X"45",X"00",X"53",X"45",
		X"54",X"0F",X"68",X"EB",X"00",X"15",X"10",X"00",X"0A",X"11",X"00",X"05",X"06",X"00",X"00",X"15",
		X"11",X"00",X"12",X"2F",X"10",X"00",X"04",X"99",X"0F",X"69",X"89",X"04",X"11",X"00",X"12",X"20",
		X"60",X"00",X"04",X"33",X"0F",X"69",X"89",X"43",X"4C",X"45",X"41",X"52",X"45",X"44",X"00",X"12",
		X"2A",X"40",X"00",X"04",X"88",X"0F",X"69",X"13",X"00",X"20",X"42",X"4F",X"4F",X"4B",X"4B",X"45",
		X"45",X"50",X"49",X"4E",X"47",X"20",X"54",X"4F",X"54",X"41",X"4C",X"53",X"20",X"00",X"12",X"1C",
		X"60",X"00",X"50",X"41",X"49",X"44",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"12",X"6C",
		X"60",X"00",X"00",X"12",X"1C",X"70",X"00",X"45",X"58",X"54",X"52",X"41",X"20",X"4D",X"45",X"4E",
		X"20",X"45",X"41",X"52",X"4E",X"45",X"44",X"12",X"6C",X"70",X"00",X"00",X"12",X"1C",X"80",X"00",
		X"50",X"4C",X"41",X"59",X"20",X"54",X"49",X"4D",X"45",X"20",X"49",X"4E",X"20",X"4D",X"49",X"4E",
		X"55",X"54",X"45",X"53",X"12",X"6C",X"80",X"00",X"00",X"12",X"1C",X"90",X"00",X"4D",X"45",X"4E",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"44",X"12",X"6C",X"90",X"00",X"00",X"12",X"1C",X"A0",X"00",
		X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"44",X"12",X"6C",
		X"A0",X"00",X"00",X"12",X"1C",X"C0",X"00",X"41",X"56",X"45",X"52",X"41",X"47",X"45",X"20",X"54",
		X"49",X"4D",X"45",X"20",X"50",X"45",X"52",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"12",X"64",
		X"C0",X"00",X"00",X"3F",X"0A",X"10",X"00",X"12",X"1C",X"D0",X"00",X"41",X"56",X"45",X"52",X"41",
		X"47",X"45",X"20",X"54",X"55",X"52",X"4E",X"53",X"20",X"50",X"45",X"52",X"20",X"43",X"52",X"45",
		X"44",X"49",X"54",X"12",X"64",X"D0",X"00",X"00",X"3D",X"0A",X"10",X"00",X"12",X"1C",X"30",X"00",
		X"4C",X"45",X"46",X"54",X"0F",X"6A",X"8F",X"12",X"6C",X"30",X"00",X"00",X"12",X"1C",X"40",X"00",
		X"43",X"45",X"4E",X"54",X"45",X"52",X"0F",X"6A",X"8F",X"12",X"6C",X"40",X"00",X"00",X"12",X"1C",
		X"50",X"00",X"52",X"49",X"47",X"48",X"54",X"0F",X"6A",X"8F",X"12",X"6C",X"50",X"00",X"00",X"20",
		X"53",X"4C",X"4F",X"54",X"20",X"43",X"4F",X"49",X"4E",X"53",X"00",X"04",X"33",X"12",X"3A",X"80",
		X"00",X"43",X"4F",X"4C",X"4F",X"52",X"20",X"52",X"41",X"4D",X"20",X"54",X"45",X"53",X"54",X"12",
		X"27",X"B0",X"00",X"56",X"45",X"52",X"54",X"49",X"43",X"41",X"4C",X"20",X"42",X"41",X"52",X"53",
		X"20",X"49",X"4E",X"44",X"49",X"43",X"41",X"54",X"45",X"20",X"45",X"52",X"52",X"4F",X"52",X"00",
		X"41",X"55",X"54",X"4F",X"20",X"55",X"50",X"00",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"00",
		X"52",X"49",X"47",X"48",X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",X"48",X"49",X"47",X"48",X"20",
		X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"45",X"53",X"45",X"54",X"00",X"4C",X"45",X"46",X"54",
		X"20",X"43",X"4F",X"49",X"4E",X"00",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"43",X"4F",X"49",
		X"4E",X"00",X"53",X"4C",X"41",X"4D",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"00",X"4D",X"4F",
		X"56",X"45",X"20",X"55",X"50",X"14",X"6B",X"98",X"00",X"4D",X"4F",X"56",X"45",X"20",X"44",X"4F",
		X"57",X"4E",X"14",X"6B",X"98",X"00",X"4D",X"4F",X"56",X"45",X"20",X"4C",X"45",X"46",X"54",X"14",
		X"6B",X"98",X"00",X"4D",X"4F",X"56",X"45",X"20",X"52",X"49",X"47",X"48",X"54",X"14",X"6B",X"98",
		X"00",X"31",X"0F",X"6B",X"5B",X"00",X"32",X"0F",X"6B",X"5B",X"00",X"3A",X"0F",X"64",X"9E",X"53",
		X"54",X"41",X"52",X"54",X"00",X"46",X"49",X"52",X"45",X"20",X"55",X"50",X"14",X"6B",X"98",X"00",
		X"46",X"49",X"52",X"45",X"20",X"44",X"4F",X"57",X"4E",X"14",X"6B",X"98",X"00",X"46",X"49",X"52",
		X"45",X"20",X"4C",X"45",X"46",X"54",X"14",X"6B",X"98",X"00",X"46",X"49",X"52",X"45",X"20",X"52",
		X"49",X"47",X"48",X"54",X"14",X"6B",X"98",X"00",X"20",X"20",X"5B",X"0F",X"64",X"9E",X"09",X"10",
		X"5C",X"00",X"04",X"88",X"12",X"3A",X"1A",X"00",X"53",X"57",X"49",X"54",X"43",X"48",X"20",X"54",
		X"45",X"53",X"54",X"00",X"04",X"99",X"12",X"3E",X"50",X"00",X"41",X"4C",X"4C",X"20",X"52",X"4F",
		X"4D",X"53",X"20",X"4F",X"4B",X"12",X"36",X"90",X"00",X"04",X"33",X"52",X"41",X"4D",X"20",X"54",
		X"45",X"53",X"54",X"20",X"46",X"4F",X"4C",X"4C",X"4F",X"57",X"53",X"0F",X"6B",X"DF",X"00",X"12",
		X"2F",X"A0",X"00",X"0F",X"64",X"1D",X"00",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",
		X"52",X"53",X"20",X"44",X"45",X"54",X"45",X"43",X"54",X"45",X"44",X"00",X"04",X"99",X"12",X"2A",
		X"80",X"00",X"4E",X"4F",X"0F",X"6B",X"E7",X"00",X"04",X"99",X"12",X"23",X"80",X"00",X"4E",X"4F",
		X"20",X"43",X"4D",X"4F",X"53",X"0F",X"6B",X"E7",X"00",X"43",X"4D",X"4F",X"53",X"20",X"52",X"41",
		X"4D",X"0F",X"6D",X"63",X"00",X"04",X"11",X"12",X"36",X"80",X"00",X"0F",X"6C",X"19",X"00",X"0F",
		X"6C",X"25",X"12",X"28",X"90",X"00",X"4F",X"52",X"20",X"57",X"52",X"49",X"54",X"45",X"20",X"50",
		X"52",X"4F",X"54",X"45",X"43",X"54",X"20",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",X"04",X"99",
		X"0F",X"6C",X"7E",X"14",X"6C",X"57",X"00",X"04",X"00",X"0F",X"6C",X"7E",X"04",X"99",X"12",X"17",
		X"B0",X"00",X"40",X"0F",X"67",X"86",X"20",X"4D",X"55",X"53",X"54",X"20",X"42",X"45",X"20",X"4F",
		X"50",X"45",X"4E",X"20",X"46",X"4F",X"52",X"20",X"54",X"45",X"53",X"54",X"40",X"00",X"12",X"1B",
		X"B0",X"00",X"40",X"0F",X"67",X"64",X"0F",X"6C",X"66",X"00",X"04",X"00",X"12",X"57",X"80",X"00",
		X"3E",X"04",X"99",X"12",X"3A",X"80",X"00",X"53",X"4F",X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",
		X"45",X"20",X"09",X"10",X"00",X"3D",X"3A",X"3A",X"12",X"30",X"70",X"00",X"49",X"4E",X"49",X"54",
		X"49",X"41",X"4C",X"20",X"54",X"45",X"53",X"54",X"53",X"20",X"49",X"4E",X"44",X"49",X"43",X"41",
		X"54",X"45",X"3F",X"00",X"04",X"11",X"0F",X"6C",X"A8",X"12",X"3C",X"90",X"00",X"0F",X"6D",X"1B",
		X"00",X"04",X"99",X"0F",X"6C",X"A8",X"12",X"3F",X"90",X"01",X"4F",X"50",X"45",X"52",X"41",X"54",
		X"49",X"4F",X"4E",X"41",X"4C",X"00",X"04",X"11",X"0F",X"6C",X"A8",X"12",X"40",X"90",X"00",X"00",
		X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"2E",X"20",X"12",X"40",X"80",X"00",X"04",X"11",X"00",X"0F",X"6D",X"14",X"05",X"E2",
		X"00",X"00",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"43",X"48",X"49",X"50",X"20",X"46",
		X"41",X"49",X"4C",X"55",X"52",X"45",X"00",X"0F",X"6D",X"14",X"52",X"4F",X"4D",X"0F",X"6D",X"63",
		X"10",X"00",X"0F",X"6D",X"14",X"52",X"41",X"4D",X"0F",X"6D",X"63",X"10",X"00",X"0F",X"6C",X"E6",
		X"52",X"4F",X"4D",X"0F",X"6D",X"63",X"10",X"00",X"0F",X"6C",X"E6",X"52",X"41",X"4D",X"0F",X"6D",
		X"63",X"10",X"00",X"20",X"45",X"52",X"52",X"4F",X"52",X"20",X"09",X"00",X"04",X"AA",X"12",X"24",
		X"C8",X"00",X"0F",X"6D",X"BB",X"04",X"66",X"12",X"38",X"B5",X"00",X"44",X"45",X"53",X"49",X"47",
		X"4E",X"45",X"44",X"20",X"42",X"59",X"20",X"56",X"49",X"44",X"20",X"4B",X"49",X"44",X"5A",X"12",
		X"2E",X"BC",X"00",X"46",X"4F",X"52",X"20",X"0F",X"6D",X"CA",X"04",X"22",X"12",X"3D",X"A8",X"00",
		X"07",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"3F",X"3A",X"09",X"10",X"00",X"04",X"AA",X"12",
		X"41",X"EE",X"00",X"0F",X"6D",X"A1",X"00",X"12",X"24",X"EE",X"00",X"43",X"4F",X"50",X"59",X"52",
		X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"3D",X"00",X"12",X"3E",X"80",X"00",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",
		X"52",X"00",X"12",X"3F",X"79",X"01",X"0F",X"6E",X"05",X"12",X"3E",X"86",X"00",X"0F",X"6D",X"E8",
		X"00",X"12",X"3F",X"7A",X"01",X"0F",X"64",X"9E",X"09",X"10",X"00",X"12",X"3E",X"EE",X"00",X"15",
		X"04",X"AA",X"10",X"05",X"03",X"00",X"00",X"04",X"BB",X"20",X"57",X"41",X"56",X"45",X"00",X"05",
		X"04",X"00",X"00",X"09",X"04",X"AA",X"10",X"00",X"4D",X"4F",X"4D",X"4D",X"59",X"00",X"47",X"52",
		X"55",X"4E",X"54",X"20",X"40",X"20",X"31",X"30",X"30",X"00",X"00",X"44",X"41",X"44",X"44",X"59",
		X"00",X"4D",X"49",X"4B",X"45",X"59",X"00",X"49",X"4E",X"44",X"45",X"53",X"54",X"52",X"55",X"43",
		X"54",X"41",X"42",X"4C",X"45",X"20",X"48",X"55",X"4C",X"4B",X"00",X"53",X"50",X"48",X"45",X"52",
		X"45",X"4F",X"49",X"44",X"20",X"40",X"20",X"31",X"30",X"30",X"30",X"20",X"20",X"20",X"20",X"20",
		X"51",X"55",X"41",X"52",X"4B",X"20",X"40",X"20",X"31",X"30",X"30",X"30",X"00",X"45",X"4E",X"46",
		X"4F",X"52",X"43",X"45",X"52",X"20",X"40",X"20",X"31",X"35",X"30",X"20",X"20",X"20",X"54",X"41",
		X"4E",X"4B",X"20",X"40",X"20",X"32",X"30",X"30",X"00",X"42",X"52",X"41",X"49",X"4E",X"20",X"40",
		X"20",X"35",X"30",X"30",X"20",X"20",X"20",X"20",X"20",X"43",X"52",X"55",X"49",X"53",X"45",X"20",
		X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"20",X"40",X"20",X"32",X"35",X"00",X"50",X"52",X"4F",
		X"47",X"20",X"40",X"20",X"31",X"30",X"30",X"00",X"04",X"AA",X"12",X"36",X"24",X"00",X"52",X"4F",
		X"42",X"4F",X"54",X"52",X"4F",X"4E",X"3F",X"3A",X"32",X"30",X"38",X"34",X"00",X"04",X"AA",X"12",
		X"25",X"84",X"00",X"53",X"41",X"56",X"45",X"20",X"54",X"48",X"45",X"20",X"4C",X"41",X"53",X"54",
		X"20",X"48",X"55",X"4D",X"41",X"4E",X"20",X"46",X"41",X"4D",X"49",X"4C",X"59",X"00",X"FF",X"FF",
		X"7E",X"70",X"FD",X"7E",X"74",X"B8",X"7E",X"75",X"2C",X"7E",X"75",X"3A",X"7E",X"6F",X"11",X"6F",
		X"65",X"34",X"02",X"A6",X"80",X"1E",X"12",X"BD",X"D0",X"AB",X"1E",X"12",X"5A",X"26",X"F4",X"35",
		X"82",X"8E",X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",X"36",X"8E",X"6F",
		X"53",X"10",X"8E",X"CC",X"00",X"C6",X"12",X"8D",X"D8",X"35",X"B6",X"34",X"36",X"8E",X"6F",X"65",
		X"10",X"8E",X"CC",X"24",X"C6",X"34",X"8D",X"C9",X"BD",X"74",X"91",X"8E",X"CC",X"8E",X"BD",X"D0",
		X"AB",X"35",X"B6",X"25",X"03",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"03",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"50",X"52",X"45",X"53",X"45",X"4E",
		X"54",X"45",X"44",X"20",X"42",X"59",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"3D",X"2F",X"28",X"01",X"04",X"01",X"01",X"00",X"00",X"01",
		X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"01",X"00",
		X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",X"01",X"02",X"00",X"00",X"01",X"00",X"04",
		X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"01",X"00",X"02",X"02",X"00",X"00",X"01",
		X"04",X"01",X"01",X"00",X"00",X"00",X"50",X"70",X"41",X"00",X"1E",X"01",X"20",X"70",X"4C",X"00",
		X"27",X"00",X"09",X"70",X"5A",X"00",X"32",X"00",X"99",X"70",X"57",X"01",X"3B",X"00",X"99",X"70",
		X"57",X"01",X"44",X"00",X"99",X"70",X"57",X"01",X"4D",X"01",X"99",X"70",X"57",X"01",X"56",X"00",
		X"99",X"70",X"57",X"01",X"5F",X"00",X"99",X"70",X"57",X"01",X"68",X"00",X"01",X"70",X"6F",X"00",
		X"73",X"00",X"10",X"70",X"79",X"00",X"7C",X"03",X"20",X"70",X"84",X"00",X"85",X"00",X"01",X"70",
		X"74",X"00",X"90",X"00",X"01",X"70",X"74",X"00",X"99",X"00",X"01",X"70",X"74",X"00",X"A2",X"00",
		X"01",X"70",X"74",X"00",X"AB",X"00",X"01",X"70",X"74",X"00",X"B4",X"00",X"01",X"70",X"74",X"00",
		X"BD",X"00",X"5A",X"20",X"40",X"25",X"41",X"30",X"4E",X"50",X"66",X"FF",X"00",X"42",X"02",X"43",
		X"03",X"44",X"04",X"45",X"05",X"42",X"FF",X"00",X"42",X"FF",X"00",X"46",X"01",X"52",X"02",X"53",
		X"03",X"54",X"04",X"55",X"05",X"56",X"06",X"57",X"07",X"58",X"08",X"59",X"09",X"7B",X"FF",X"00",
		X"48",X"01",X"47",X"FF",X"00",X"48",X"01",X"51",X"FF",X"00",X"49",X"03",X"4A",X"05",X"44",X"06",
		X"4C",X"08",X"4D",X"FF",X"00",X"44",X"04",X"42",X"FF",X"34",X"22",X"86",X"11",X"6D",X"44",X"27",
		X"02",X"86",X"16",X"E6",X"45",X"1F",X"01",X"A6",X"E4",X"BD",X"5F",X"96",X"8D",X"02",X"35",X"A2",
		X"34",X"36",X"1E",X"12",X"BD",X"D0",X"A5",X"C1",X"FF",X"26",X"02",X"C6",X"EE",X"1E",X"12",X"1E",
		X"10",X"86",X"59",X"E6",X"45",X"1E",X"10",X"34",X"06",X"CC",X"3C",X"05",X"BD",X"D0",X"1B",X"35",
		X"06",X"8D",X"05",X"BD",X"5F",X"96",X"35",X"B6",X"34",X"20",X"10",X"AE",X"42",X"E1",X"A1",X"24",
		X"FC",X"A6",X"3D",X"35",X"A0",X"BD",X"D0",X"12",X"86",X"66",X"97",X"CF",X"CE",X"6F",X"D5",X"10",
		X"8E",X"CC",X"00",X"86",X"2E",X"8E",X"CC",X"24",X"34",X"10",X"8D",X"9D",X"33",X"46",X"31",X"22",
		X"4C",X"10",X"AC",X"E4",X"26",X"F4",X"86",X"2D",X"BD",X"5F",X"96",X"35",X"90",X"BD",X"74",X"AB",
		X"27",X"03",X"BD",X"6F",X"2C",X"8E",X"CC",X"18",X"6F",X"80",X"8C",X"CC",X"24",X"25",X"F9",X"BD",
		X"74",X"78",X"8D",X"C1",X"CE",X"6F",X"D5",X"10",X"8E",X"CC",X"00",X"86",X"2E",X"BD",X"74",X"33",
		X"BD",X"71",X"FE",X"BD",X"D0",X"54",X"72",X"9F",X"BD",X"72",X"1D",X"8D",X"08",X"86",X"01",X"8E",
		X"71",X"28",X"7E",X"D0",X"66",X"35",X"06",X"DE",X"15",X"ED",X"4D",X"86",X"20",X"A7",X"47",X"B6",
		X"C8",X"04",X"2B",X"22",X"85",X"40",X"26",X"03",X"6E",X"D8",X"0D",X"8D",X"32",X"86",X"01",X"8E",
		X"71",X"55",X"7E",X"D0",X"66",X"B6",X"C8",X"04",X"85",X"40",X"27",X"EC",X"6A",X"47",X"26",X"ED",
		X"86",X"05",X"A7",X"47",X"20",X"E5",X"8D",X"3D",X"86",X"01",X"8E",X"71",X"70",X"7E",X"D0",X"66",
		X"B6",X"C8",X"04",X"2A",X"D3",X"6A",X"47",X"26",X"EF",X"86",X"05",X"A7",X"47",X"20",X"E7",X"BD",
		X"74",X"3E",X"1F",X"21",X"BD",X"D0",X"A2",X"10",X"8C",X"CC",X"00",X"27",X"32",X"8B",X"01",X"19",
		X"25",X"12",X"A1",X"41",X"22",X"0E",X"1F",X"21",X"BD",X"D0",X"AB",X"BD",X"74",X"78",X"BD",X"70",
		X"A0",X"BD",X"74",X"49",X"39",X"BD",X"74",X"3E",X"1F",X"21",X"BD",X"D0",X"A2",X"4D",X"27",X"F4",
		X"10",X"8C",X"CC",X"00",X"27",X"0F",X"8B",X"99",X"19",X"A1",X"C4",X"25",X"E7",X"20",X"D7",X"8D",
		X"0A",X"A6",X"01",X"20",X"D1",X"8D",X"04",X"A6",X"1F",X"20",X"CB",X"8E",X"71",X"DB",X"A1",X"84",
		X"23",X"07",X"30",X"01",X"8C",X"71",X"DF",X"25",X"F5",X"39",X"00",X"00",X"20",X"25",X"30",X"50",
		X"50",X"34",X"12",X"A6",X"44",X"27",X"13",X"8E",X"CC",X"04",X"4A",X"27",X"03",X"8E",X"CC",X"14",
		X"BD",X"D0",X"A2",X"4D",X"27",X"04",X"1A",X"01",X"35",X"92",X"1C",X"FE",X"35",X"92",X"34",X"16",
		X"E6",X"45",X"86",X"0C",X"1F",X"01",X"86",X"2C",X"BD",X"5F",X"96",X"35",X"96",X"34",X"16",X"E6",
		X"45",X"86",X"0C",X"1F",X"01",X"CC",X"03",X"05",X"BD",X"D0",X"1B",X"35",X"96",X"35",X"06",X"DE",
		X"15",X"ED",X"4D",X"86",X"30",X"A7",X"47",X"B6",X"C8",X"04",X"46",X"25",X"21",X"46",X"25",X"03",
		X"6E",X"D8",X"0D",X"8D",X"33",X"86",X"01",X"8E",X"72",X"3D",X"7E",X"D0",X"66",X"B6",X"C8",X"04",
		X"85",X"02",X"27",X"EC",X"6A",X"47",X"26",X"ED",X"86",X"08",X"A7",X"47",X"20",X"E5",X"8D",X"34",
		X"86",X"01",X"8E",X"72",X"58",X"7E",X"D0",X"66",X"B6",X"C8",X"04",X"46",X"24",X"D2",X"6A",X"47",
		X"26",X"EE",X"86",X"08",X"A7",X"47",X"20",X"E6",X"BD",X"74",X"3E",X"8D",X"A0",X"10",X"8C",X"CC",
		X"22",X"27",X"0D",X"31",X"22",X"4C",X"33",X"46",X"BD",X"71",X"E1",X"25",X"F0",X"BD",X"74",X"33",
		X"BD",X"71",X"FE",X"39",X"BD",X"74",X"3E",X"8D",X"84",X"10",X"8C",X"CC",X"00",X"27",X"F1",X"31",
		X"3E",X"4A",X"33",X"5A",X"BD",X"71",X"E1",X"25",X"F0",X"BD",X"74",X"33",X"7E",X"71",X"FE",X"86",
		X"01",X"8E",X"72",X"A7",X"7E",X"D0",X"66",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F1",X"BD",X"D0",
		X"60",X"BD",X"D0",X"12",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1B",X"84",X"0F",
		X"27",X"14",X"7F",X"CC",X"1B",X"BD",X"74",X"78",X"BD",X"D0",X"12",X"BD",X"75",X"15",X"86",X"40",
		X"8E",X"72",X"D6",X"7E",X"D0",X"66",X"B6",X"CC",X"1D",X"84",X"0F",X"27",X"11",X"7F",X"CC",X"1D",
		X"BD",X"74",X"78",X"BD",X"E3",X"D9",X"86",X"40",X"8E",X"72",X"EE",X"7E",X"D0",X"66",X"B6",X"CC",
		X"21",X"84",X"0F",X"27",X"5D",X"7F",X"CC",X"21",X"BD",X"74",X"78",X"86",X"3A",X"8E",X"CC",X"24",
		X"C6",X"32",X"BD",X"D0",X"AB",X"5A",X"26",X"FA",X"BD",X"D0",X"12",X"86",X"5C",X"BD",X"5F",X"99",
		X"10",X"8E",X"CC",X"24",X"8E",X"25",X"30",X"CC",X"19",X"80",X"BD",X"75",X"3A",X"C6",X"30",X"8E",
		X"CC",X"88",X"10",X"8E",X"CC",X"24",X"BD",X"73",X"8A",X"86",X"5C",X"BD",X"5F",X"99",X"BD",X"74",
		X"0D",X"10",X"8E",X"CC",X"56",X"8E",X"25",X"40",X"CC",X"19",X"80",X"BD",X"75",X"3A",X"C6",X"40",
		X"8E",X"CC",X"8A",X"10",X"8E",X"CC",X"56",X"8D",X"41",X"BD",X"74",X"91",X"8E",X"CC",X"8E",X"BD",
		X"D0",X"AB",X"B6",X"CC",X"23",X"84",X"0F",X"27",X"09",X"7F",X"CC",X"23",X"BD",X"74",X"78",X"BD",
		X"E3",X"D6",X"B6",X"CC",X"1F",X"84",X"0F",X"27",X"0B",X"7F",X"CC",X"1F",X"BD",X"74",X"78",X"8D",
		X"08",X"7E",X"F0",X"06",X"8D",X"03",X"7E",X"D0",X"00",X"B6",X"CC",X"19",X"84",X"0F",X"27",X"09",
		X"7C",X"CC",X"8C",X"7C",X"CC",X"8C",X"7F",X"CC",X"19",X"39",X"DE",X"15",X"86",X"25",X"ED",X"47",
		X"35",X"06",X"ED",X"4D",X"AF",X"4B",X"10",X"AF",X"49",X"86",X"25",X"BD",X"D0",X"AB",X"86",X"65",
		X"BD",X"5F",X"99",X"86",X"04",X"8E",X"73",X"AB",X"7E",X"D0",X"66",X"B6",X"C8",X"0C",X"85",X"02",
		X"26",X"F1",X"B6",X"C8",X"06",X"85",X"02",X"27",X"10",X"AE",X"4B",X"BD",X"D0",X"A2",X"AE",X"4B",
		X"4C",X"81",X"3A",X"23",X"15",X"86",X"3A",X"20",X"11",X"46",X"24",X"1D",X"AE",X"4B",X"BD",X"D0",
		X"A2",X"AE",X"4B",X"4A",X"81",X"13",X"24",X"02",X"86",X"13",X"BD",X"D0",X"AB",X"A7",X"47",X"8D",
		X"2C",X"86",X"10",X"8E",X"73",X"B2",X"7E",X"D0",X"66",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"08",
		X"86",X"04",X"8E",X"73",X"B2",X"7E",X"D0",X"66",X"BD",X"D0",X"12",X"86",X"04",X"8E",X"74",X"03",
		X"7E",X"D0",X"66",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F1",X"6E",X"D8",X"0D",X"0F",X"D0",X"AE",
		X"47",X"30",X"89",X"FF",X"00",X"86",X"5A",X"C6",X"09",X"BD",X"D0",X"1B",X"AE",X"47",X"0F",X"D0",
		X"10",X"AE",X"49",X"C6",X"19",X"1E",X"12",X"BD",X"D0",X"A2",X"1E",X"12",X"BD",X"5F",X"93",X"5A",
		X"26",X"F3",X"39",X"10",X"BF",X"B3",X"EC",X"FF",X"B3",X"EF",X"B7",X"B3",X"EE",X"39",X"10",X"BE",
		X"B3",X"EC",X"FE",X"B3",X"EF",X"B6",X"B3",X"EE",X"39",X"10",X"8C",X"CC",X"04",X"27",X"01",X"39",
		X"1F",X"21",X"BD",X"D0",X"A2",X"48",X"34",X"02",X"48",X"AB",X"E0",X"8E",X"6F",X"99",X"30",X"86",
		X"33",X"46",X"31",X"22",X"A6",X"80",X"34",X"10",X"1F",X"21",X"BD",X"D0",X"AB",X"35",X"10",X"BD",
		X"70",X"A0",X"10",X"8C",X"CC",X"10",X"25",X"E8",X"34",X"12",X"8D",X"08",X"8E",X"CC",X"8C",X"BD",
		X"D0",X"AB",X"35",X"92",X"34",X"34",X"8E",X"CC",X"00",X"10",X"8E",X"CC",X"24",X"8D",X"09",X"35",
		X"B4",X"8E",X"CC",X"24",X"10",X"8E",X"CC",X"8C",X"10",X"9F",X"2B",X"4F",X"E6",X"80",X"C4",X"0F",
		X"34",X"04",X"AB",X"E0",X"9C",X"2B",X"26",X"F4",X"8B",X"37",X"39",X"8D",X"D7",X"34",X"02",X"8E",
		X"CC",X"8C",X"BD",X"D0",X"A2",X"A1",X"E0",X"39",X"8D",X"6B",X"8D",X"EF",X"27",X"3A",X"86",X"39",
		X"B7",X"CB",X"FF",X"BD",X"6F",X"2C",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"AB",X"86",X"39",X"B7",
		X"CB",X"FF",X"BD",X"D0",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"23",X"BD",X"E3",X"DC",X"BD",
		X"E3",X"D0",X"8D",X"C7",X"27",X"15",X"86",X"4F",X"BD",X"5F",X"99",X"86",X"39",X"B7",X"CB",X"FF",
		X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F4",X"39",X"7E",X"E3",X"D0",X"86",X"50",X"20",X"E9",X"8E",
		X"CD",X"02",X"C6",X"04",X"A6",X"80",X"84",X"0F",X"81",X"09",X"23",X"03",X"5A",X"27",X"06",X"8C",
		X"CD",X"32",X"26",X"F0",X"39",X"86",X"5B",X"BD",X"5F",X"99",X"8E",X"CD",X"02",X"6F",X"80",X"8C",
		X"CD",X"32",X"26",X"F9",X"39",X"8D",X"05",X"27",X"FB",X"7E",X"6F",X"3B",X"BD",X"74",X"91",X"34",
		X"02",X"8E",X"CC",X"8E",X"BD",X"D0",X"A2",X"A1",X"E0",X"39",X"DE",X"15",X"ED",X"47",X"AF",X"49",
		X"10",X"AF",X"4B",X"35",X"06",X"ED",X"4D",X"86",X"04",X"8E",X"75",X"4F",X"7E",X"D0",X"66",X"8D",
		X"34",X"26",X"F4",X"BD",X"D0",X"54",X"77",X"49",X"EC",X"4D",X"ED",X"0D",X"EC",X"47",X"ED",X"07",
		X"EF",X"09",X"9F",X"D8",X"86",X"99",X"97",X"CF",X"0F",X"D0",X"0F",X"DA",X"0F",X"DB",X"0F",X"DC",
		X"8D",X"08",X"86",X"02",X"8E",X"75",X"8B",X"7E",X"D0",X"66",X"BD",X"76",X"2A",X"BD",X"76",X"36",
		X"86",X"3A",X"7E",X"76",X"5D",X"B6",X"C8",X"04",X"85",X"40",X"39",X"B6",X"C8",X"04",X"46",X"10",
		X"25",X"01",X"16",X"46",X"10",X"25",X"00",X"F3",X"8D",X"EB",X"27",X"D6",X"A6",X"48",X"84",X"80",
		X"8B",X"20",X"A7",X"48",X"BD",X"76",X"48",X"81",X"5E",X"27",X"4D",X"96",X"D0",X"97",X"DC",X"BD",
		X"76",X"45",X"BD",X"76",X"48",X"AE",X"49",X"9F",X"DA",X"BD",X"5F",X"93",X"AF",X"49",X"BD",X"76",
		X"72",X"6A",X"47",X"27",X"2B",X"BD",X"75",X"7A",X"86",X"02",X"8E",X"75",X"D0",X"7E",X"D0",X"66",
		X"8D",X"B3",X"27",X"0F",X"A6",X"47",X"4A",X"27",X"EF",X"6A",X"48",X"27",X"06",X"A6",X"48",X"81",
		X"80",X"26",X"E5",X"BD",X"75",X"85",X"27",X"8A",X"A6",X"48",X"84",X"80",X"8B",X"04",X"20",X"B2",
		X"9E",X"D8",X"BD",X"D0",X"5D",X"6E",X"D8",X"0D",X"8D",X"4B",X"8D",X"2E",X"86",X"3A",X"8D",X"5D",
		X"9E",X"DA",X"AF",X"49",X"D6",X"DC",X"D7",X"D0",X"6C",X"47",X"10",X"AE",X"4B",X"31",X"3F",X"10",
		X"8C",X"C0",X"00",X"25",X"02",X"31",X"3F",X"10",X"AF",X"4B",X"86",X"01",X"8E",X"76",X"22",X"7E",
		X"D0",X"66",X"BD",X"75",X"85",X"26",X"F3",X"7E",X"75",X"6A",X"34",X"06",X"AE",X"49",X"CC",X"04",
		X"07",X"BD",X"D0",X"1B",X"35",X"86",X"86",X"99",X"AE",X"49",X"A7",X"08",X"A7",X"89",X"01",X"08",
		X"A7",X"89",X"02",X"08",X"39",X"4F",X"20",X"F0",X"10",X"AE",X"4B",X"10",X"8C",X"C0",X"00",X"24",
		X"03",X"A6",X"A4",X"39",X"34",X"10",X"AE",X"4B",X"BD",X"D0",X"A2",X"35",X"90",X"10",X"AE",X"4B",
		X"10",X"8C",X"C0",X"00",X"24",X"03",X"A7",X"A4",X"39",X"34",X"10",X"AE",X"4B",X"BD",X"D0",X"AB",
		X"35",X"90",X"10",X"AE",X"4B",X"31",X"21",X"10",X"8C",X"C0",X"00",X"25",X"02",X"31",X"21",X"10",
		X"AF",X"4B",X"39",X"8E",X"20",X"00",X"30",X"1F",X"26",X"FC",X"39",X"86",X"0A",X"8D",X"7F",X"8D",
		X"F2",X"F6",X"C8",X"04",X"C5",X"02",X"10",X"27",X"FE",X"FE",X"4A",X"26",X"F2",X"86",X"01",X"8E",
		X"76",X"A5",X"7E",X"D0",X"66",X"86",X"01",X"20",X"E4",X"86",X"0A",X"8D",X"19",X"8D",X"D4",X"F6",
		X"C8",X"04",X"56",X"10",X"24",X"FE",X"E1",X"4A",X"26",X"F3",X"86",X"01",X"8E",X"76",X"C2",X"7E",
		X"D0",X"66",X"86",X"01",X"20",X"E5",X"34",X"02",X"BD",X"76",X"48",X"4C",X"6D",X"48",X"2A",X"15",
		X"0D",X"DA",X"27",X"04",X"81",X"5E",X"23",X"06",X"81",X"5D",X"23",X"02",X"86",X"30",X"81",X"3E",
		X"26",X"1B",X"4C",X"20",X"18",X"81",X"5A",X"23",X"0E",X"0D",X"DA",X"27",X"08",X"81",X"5E",X"22",
		X"04",X"86",X"5E",X"20",X"02",X"86",X"3A",X"81",X"3B",X"26",X"02",X"86",X"41",X"BD",X"76",X"5D",
		X"BD",X"76",X"2A",X"D6",X"D0",X"AE",X"49",X"BD",X"5F",X"93",X"D7",X"D0",X"35",X"82",X"34",X"02",
		X"BD",X"76",X"48",X"4A",X"6D",X"48",X"2A",X"15",X"81",X"30",X"24",X"0A",X"0D",X"DA",X"27",X"04",
		X"86",X"5E",X"20",X"02",X"86",X"5D",X"81",X"3E",X"26",X"1D",X"4A",X"20",X"1A",X"81",X"39",X"26",
		X"0A",X"0D",X"DA",X"27",X"04",X"86",X"5E",X"20",X"02",X"86",X"5A",X"81",X"40",X"26",X"02",X"86",
		X"3A",X"81",X"5D",X"26",X"02",X"86",X"5A",X"20",X"B4",X"6D",X"48",X"2B",X"34",X"86",X"FF",X"8E",
		X"77",X"55",X"7E",X"D0",X"66",X"86",X"FF",X"8E",X"77",X"5D",X"7E",X"D0",X"66",X"86",X"82",X"8E",
		X"77",X"65",X"7E",X"D0",X"66",X"6A",X"47",X"26",X"E4",X"AE",X"49",X"33",X"84",X"BD",X"76",X"48",
		X"81",X"5E",X"26",X"05",X"86",X"3A",X"BD",X"76",X"5D",X"DE",X"15",X"BD",X"D0",X"5D",X"6E",X"D8",
		X"0D",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"E1",X"86",X"01",X"8E",X"77",X"81",X"7E",X"D0",X"66",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"77",X"A5",X"79",X"2D",X"BD",X"D0",X"60",X"0F",X"F4",X"BD",X"D0",X"54",X"77",X"B9",X"8E",
		X"77",X"E4",X"4F",X"BD",X"D0",X"5A",X"7E",X"D0",X"63",X"96",X"51",X"A7",X"47",X"96",X"51",X"A1",
		X"47",X"27",X"05",X"0C",X"F4",X"7E",X"79",X"9D",X"86",X"08",X"8E",X"77",X"BD",X"7E",X"D0",X"66",
		X"8A",X"77",X"8A",X"CA",X"8B",X"16",X"8A",X"CA",X"8B",X"95",X"8A",X"77",X"8A",X"CA",X"8B",X"CB",
		X"8C",X"07",X"00",X"00",X"BD",X"D0",X"12",X"BD",X"DF",X"40",X"0F",X"F4",X"7E",X"79",X"9D",X"0F",
		X"F4",X"BD",X"D0",X"60",X"BD",X"D0",X"30",X"BD",X"D0",X"12",X"BD",X"D0",X"54",X"77",X"B9",X"0F",
		X"0C",X"0F",X"0E",X"86",X"03",X"8E",X"78",X"0B",X"7E",X"D0",X"66",X"8E",X"18",X"3A",X"AF",X"49",
		X"8E",X"9A",X"B0",X"10",X"8E",X"77",X"D0",X"10",X"AF",X"47",X"AF",X"4B",X"86",X"01",X"8E",X"78",
		X"24",X"7E",X"D0",X"66",X"10",X"AE",X"4B",X"CC",X"0B",X"0E",X"ED",X"A4",X"C6",X"0D",X"ED",X"24",
		X"30",X"2A",X"AF",X"22",X"30",X"A9",X"00",X"A4",X"AF",X"26",X"AE",X"49",X"AF",X"28",X"10",X"AE",
		X"47",X"EE",X"A4",X"27",X"33",X"5F",X"86",X"CE",X"34",X"10",X"BD",X"8D",X"69",X"DE",X"15",X"30",
		X"89",X"02",X"00",X"AF",X"49",X"35",X"10",X"10",X"AE",X"4B",X"31",X"2A",X"CC",X"0B",X"1B",X"BD",
		X"D0",X"B7",X"AE",X"4B",X"30",X"89",X"01",X"33",X"10",X"AE",X"47",X"31",X"22",X"20",X"A8",X"34",
		X"02",X"B6",X"CC",X"13",X"84",X"0F",X"35",X"82",X"8D",X"F5",X"27",X"03",X"BD",X"D0",X"12",X"86",
		X"07",X"97",X"0C",X"86",X"3F",X"97",X"0E",X"8D",X"E6",X"10",X"27",X"0F",X"19",X"96",X"59",X"84",
		X"FB",X"97",X"59",X"DE",X"15",X"10",X"8E",X"9A",X"B0",X"10",X"AF",X"47",X"86",X"09",X"A7",X"49",
		X"20",X"08",X"86",X"08",X"8E",X"78",X"AA",X"7E",X"D0",X"66",X"10",X"AE",X"47",X"EC",X"28",X"CB",
		X"0D",X"D7",X"A7",X"C0",X"0D",X"30",X"A4",X"BD",X"5B",X"55",X"CB",X"0E",X"D7",X"A7",X"30",X"24",
		X"BD",X"5B",X"55",X"31",X"A9",X"01",X"33",X"10",X"AF",X"47",X"6A",X"49",X"26",X"D4",X"86",X"20",
		X"8E",X"87",X"A6",X"7E",X"D0",X"66",X"86",X"3F",X"97",X"0F",X"86",X"07",X"97",X"0D",X"BD",X"D0",
		X"54",X"D0",X"C3",X"10",X"8E",X"8C",X"E8",X"5F",X"8E",X"39",X"5C",X"86",X"FD",X"EE",X"B1",X"27",
		X"05",X"BD",X"8D",X"69",X"20",X"F7",X"EE",X"A1",X"27",X"05",X"BD",X"8D",X"69",X"20",X"F7",X"BD",
		X"D0",X"54",X"79",X"2D",X"8E",X"79",X"75",X"10",X"8E",X"98",X"0E",X"86",X"01",X"DE",X"15",X"AF",
		X"49",X"10",X"AF",X"4B",X"A7",X"4D",X"AE",X"49",X"AF",X"47",X"AE",X"47",X"A6",X"80",X"27",X"F6",
		X"A7",X"D8",X"0B",X"AF",X"47",X"A6",X"4D",X"8E",X"79",X"1A",X"7E",X"D0",X"66",X"96",X"86",X"2A",
		X"10",X"86",X"07",X"97",X"0C",X"BD",X"D0",X"39",X"84",X"07",X"4C",X"8E",X"79",X"41",X"7E",X"D0",
		X"66",X"96",X"84",X"84",X"03",X"27",X"0A",X"0F",X"0C",X"86",X"03",X"8E",X"79",X"51",X"7E",X"D0",
		X"66",X"8E",X"79",X"8B",X"BD",X"D0",X"39",X"84",X"0F",X"A6",X"86",X"97",X"0C",X"86",X"07",X"8E",
		X"79",X"65",X"7E",X"D0",X"66",X"96",X"86",X"84",X"03",X"27",X"C2",X"0F",X"0C",X"86",X"04",X"8E",
		X"79",X"2D",X"7E",X"D0",X"66",X"3F",X"3F",X"3F",X"37",X"2F",X"27",X"1F",X"17",X"0F",X"07",X"07",
		X"07",X"0F",X"17",X"1F",X"27",X"2F",X"37",X"3F",X"3F",X"3F",X"00",X"FF",X"C0",X"C7",X"1F",X"07",
		X"07",X"C0",X"C7",X"FF",X"C0",X"C7",X"16",X"07",X"FF",X"C0",X"C7",X"20",X"37",X"96",X"F4",X"8A",
		X"80",X"97",X"F4",X"8D",X"0A",X"86",X"81",X"BD",X"5F",X"99",X"8E",X"83",X"B2",X"20",X"2A",X"BD",
		X"D0",X"60",X"BD",X"D0",X"C0",X"BD",X"D0",X"12",X"BD",X"D0",X"24",X"BD",X"D0",X"54",X"7E",X"C8",
		X"96",X"59",X"84",X"F3",X"97",X"59",X"0F",X"3F",X"86",X"CC",X"97",X"8F",X"BD",X"26",X"D2",X"86",
		X"80",X"7E",X"5F",X"99",X"8D",X"D9",X"8E",X"7F",X"A3",X"DE",X"15",X"AF",X"47",X"AE",X"47",X"A6",
		X"80",X"AF",X"47",X"81",X"09",X"22",X"08",X"8E",X"7A",X"08",X"48",X"AD",X"96",X"20",X"EE",X"81",
		X"5F",X"25",X"06",X"8E",X"79",X"DD",X"7E",X"D0",X"66",X"AE",X"49",X"BD",X"5F",X"93",X"AF",X"49",
		X"86",X"03",X"8E",X"79",X"DD",X"7E",X"D0",X"66",X"7A",X"93",X"7A",X"9C",X"7A",X"B6",X"7A",X"C1",
		X"7A",X"C7",X"7A",X"60",X"7A",X"84",X"7A",X"5A",X"7A",X"29",X"7A",X"1C",X"96",X"F4",X"84",X"7F",
		X"97",X"F4",X"10",X"27",X"FD",X"C9",X"7E",X"79",X"9B",X"8E",X"7A",X"31",X"86",X"00",X"7E",X"D0",
		X"57",X"86",X"0E",X"A7",X"47",X"86",X"10",X"8E",X"7A",X"3D",X"7E",X"D0",X"66",X"BD",X"D0",X"39",
		X"84",X"06",X"8E",X"7A",X"52",X"10",X"AE",X"86",X"BD",X"7B",X"0F",X"6A",X"47",X"26",X"E6",X"7E",
		X"D0",X"63",X"84",X"F5",X"85",X"17",X"85",X"40",X"85",X"67",X"BD",X"7D",X"6E",X"97",X"CF",X"39",
		X"86",X"14",X"C6",X"D8",X"1F",X"01",X"CC",X"74",X"06",X"BD",X"D0",X"1B",X"96",X"D0",X"34",X"02",
		X"BD",X"7D",X"6E",X"C6",X"D8",X"0F",X"D0",X"1F",X"01",X"BD",X"7D",X"6E",X"BD",X"5F",X"96",X"35",
		X"02",X"97",X"D0",X"39",X"96",X"59",X"8A",X"0C",X"97",X"59",X"BD",X"D0",X"30",X"BD",X"D0",X"60",
		X"7E",X"77",X"A0",X"BD",X"7D",X"5E",X"10",X"AF",X"49",X"0F",X"D0",X"39",X"BD",X"7D",X"6E",X"1F",
		X"89",X"86",X"14",X"ED",X"49",X"8E",X"14",X"30",X"0F",X"D0",X"BD",X"7D",X"6E",X"1F",X"89",X"C0",
		X"10",X"86",X"74",X"7E",X"D0",X"1B",X"E6",X"4A",X"86",X"14",X"CB",X"0B",X"ED",X"49",X"0F",X"D0",
		X"39",X"BD",X"7D",X"5E",X"7E",X"7B",X"0F",X"BD",X"7D",X"6E",X"8E",X"79",X"DD",X"7E",X"D0",X"66",
		X"10",X"8E",X"FD",X"80",X"CC",X"FF",X"06",X"20",X"07",X"10",X"8E",X"02",X"80",X"CC",X"02",X"06",
		X"BD",X"D0",X"6F",X"10",X"AF",X"0E",X"10",X"AE",X"47",X"EB",X"2C",X"E7",X"0C",X"AB",X"2A",X"A7",
		X"0A",X"ED",X"04",X"FC",X"26",X"D7",X"ED",X"02",X"ED",X"88",X"14",X"9F",X"17",X"AF",X"47",X"A6",
		X"49",X"8E",X"7B",X"07",X"7E",X"D0",X"66",X"AE",X"47",X"BD",X"D0",X"75",X"7E",X"D0",X"63",X"34",
		X"12",X"86",X"00",X"8E",X"7B",X"1E",X"BD",X"D0",X"5A",X"10",X"AF",X"07",X"35",X"92",X"BD",X"D0",
		X"6F",X"AF",X"4B",X"6F",X"C8",X"12",X"8D",X"11",X"8D",X"0F",X"DE",X"15",X"AE",X"4B",X"EC",X"02",
		X"ED",X"88",X"14",X"9F",X"17",X"8D",X"02",X"20",X"FC",X"35",X"06",X"DE",X"15",X"ED",X"4E",X"BD",
		X"7D",X"6E",X"48",X"8E",X"7B",X"58",X"AE",X"86",X"9F",X"2B",X"AE",X"4B",X"10",X"AE",X"49",X"AD",
		X"9F",X"98",X"2B",X"DE",X"15",X"6E",X"D8",X"0E",X"8D",X"A0",X"7D",X"31",X"7D",X"4B",X"7D",X"19",
		X"7D",X"1F",X"7D",X"25",X"7D",X"2B",X"7C",X"C1",X"7C",X"B2",X"7C",X"B9",X"7C",X"8F",X"7C",X"87",
		X"7C",X"81",X"7C",X"6F",X"7C",X"68",X"7C",X"54",X"7C",X"5C",X"7C",X"4E",X"7C",X"1F",X"7C",X"26",
		X"7C",X"37",X"7C",X"05",X"7C",X"CB",X"D0",X"63",X"7D",X"41",X"7B",X"90",X"7C",X"D9",X"7B",X"FD",
		X"35",X"06",X"ED",X"C8",X"10",X"BD",X"7C",X"54",X"6F",X"88",X"12",X"BD",X"7D",X"5E",X"10",X"AF",
		X"C8",X"15",X"BD",X"7D",X"5E",X"10",X"AF",X"C8",X"17",X"A6",X"0A",X"E6",X"0C",X"ED",X"04",X"ED",
		X"06",X"86",X"03",X"8E",X"7B",X"B9",X"7E",X"D0",X"66",X"AE",X"4B",X"8D",X"2F",X"EC",X"04",X"AB",
		X"0E",X"EB",X"88",X"10",X"ED",X"04",X"EC",X"C8",X"15",X"10",X"AE",X"02",X"BD",X"1A",X"C8",X"EC",
		X"04",X"ED",X"06",X"A6",X"C8",X"18",X"27",X"05",X"8D",X"1A",X"BD",X"D0",X"18",X"6A",X"C8",X"17",
		X"26",X"CF",X"8D",X"10",X"8D",X"06",X"BD",X"7C",X"5C",X"6E",X"D8",X"10",X"EC",X"06",X"10",X"AE",
		X"02",X"7E",X"D0",X"1E",X"EC",X"04",X"A7",X"0A",X"E7",X"0C",X"6F",X"0B",X"39",X"AF",X"47",X"BD",
		X"7C",X"54",X"7E",X"38",X"95",X"BD",X"7D",X"5E",X"8E",X"7B",X"35",X"86",X"00",X"BD",X"D0",X"5A",
		X"10",X"AF",X"07",X"EC",X"4B",X"ED",X"0B",X"EC",X"49",X"ED",X"09",X"6F",X"88",X"12",X"39",X"BD",
		X"D0",X"54",X"7A",X"D0",X"20",X"05",X"BD",X"D0",X"54",X"7A",X"D9",X"EC",X"4B",X"ED",X"07",X"BD",
		X"7D",X"6E",X"A7",X"09",X"7E",X"7C",X"87",X"BD",X"7D",X"6E",X"BD",X"7D",X"5E",X"E6",X"C8",X"12",
		X"26",X"03",X"A7",X"C8",X"12",X"6A",X"C8",X"12",X"27",X"03",X"10",X"AF",X"47",X"39",X"BD",X"7D",
		X"5E",X"7E",X"7B",X"0F",X"BD",X"D0",X"75",X"EC",X"84",X"DD",X"1B",X"39",X"EC",X"02",X"ED",X"88",
		X"14",X"DC",X"17",X"ED",X"84",X"9F",X"17",X"39",X"BD",X"7D",X"5E",X"10",X"AF",X"47",X"39",X"BD",
		X"D0",X"75",X"86",X"A6",X"97",X"A7",X"CC",X"FF",X"00",X"DD",X"88",X"BD",X"5B",X"43",X"7E",X"D0",
		X"63",X"BD",X"D0",X"75",X"7E",X"D0",X"63",X"35",X"10",X"BD",X"7D",X"6E",X"7E",X"D0",X"66",X"35",
		X"06",X"ED",X"C8",X"10",X"BD",X"7D",X"5E",X"10",X"AF",X"C8",X"13",X"10",X"AE",X"49",X"BD",X"7D",
		X"41",X"A6",X"C8",X"13",X"8E",X"7C",X"AA",X"7E",X"D0",X"66",X"6A",X"C8",X"14",X"26",X"EC",X"6E",
		X"D8",X"10",X"BD",X"7D",X"5E",X"10",X"AF",X"0E",X"39",X"BD",X"7D",X"5E",X"10",X"AF",X"88",X"10",
		X"39",X"BD",X"7D",X"5E",X"1F",X"20",X"E7",X"0C",X"A7",X"0A",X"39",X"BD",X"7D",X"5E",X"1F",X"20",
		X"AB",X"0A",X"A7",X"0A",X"EB",X"0C",X"E7",X"0C",X"39",X"A6",X"05",X"A7",X"C8",X"13",X"86",X"40",
		X"A7",X"C8",X"15",X"BD",X"D0",X"39",X"84",X"07",X"AB",X"C8",X"13",X"A7",X"05",X"86",X"01",X"8E",
		X"7C",X"F5",X"7E",X"D0",X"66",X"AE",X"4B",X"BD",X"D0",X"39",X"84",X"07",X"40",X"AB",X"C8",X"13",
		X"A7",X"05",X"86",X"01",X"8E",X"7D",X"0A",X"7E",X"D0",X"66",X"AE",X"4B",X"6A",X"C8",X"15",X"26",
		X"D2",X"A6",X"C8",X"13",X"A7",X"05",X"7E",X"D0",X"63",X"BD",X"7D",X"6E",X"6E",X"B8",X"04",X"BD",
		X"7D",X"6E",X"6E",X"B8",X"06",X"BD",X"7D",X"6E",X"6E",X"B8",X"08",X"BD",X"7D",X"6E",X"6E",X"B8",
		X"0A",X"BD",X"7D",X"5E",X"10",X"AF",X"49",X"4F",X"A7",X"4D",X"8D",X"14",X"AE",X"4B",X"ED",X"02",
		X"39",X"A6",X"4D",X"4C",X"A1",X"22",X"25",X"F0",X"4F",X"20",X"ED",X"BD",X"7D",X"6E",X"20",X"EA",
		X"34",X"60",X"DE",X"15",X"10",X"AE",X"49",X"E6",X"23",X"3D",X"E3",X"B4",X"35",X"E0",X"34",X"50",
		X"8D",X"07",X"10",X"AE",X"81",X"AF",X"47",X"35",X"D0",X"DE",X"15",X"AE",X"47",X"39",X"34",X"50",
		X"8D",X"F7",X"A6",X"80",X"20",X"EF",X"5F",X"ED",X"C8",X"13",X"A6",X"2C",X"40",X"20",X"1C",X"C6",
		X"03",X"ED",X"C8",X"13",X"A6",X"2C",X"5F",X"20",X"12",X"C6",X"06",X"ED",X"C8",X"13",X"E6",X"2C",
		X"20",X"08",X"C6",X"09",X"ED",X"C8",X"13",X"E6",X"2C",X"50",X"4F",X"ED",X"C8",X"15",X"35",X"06",
		X"ED",X"C8",X"10",X"CC",X"7D",X"F2",X"ED",X"C8",X"17",X"10",X"AE",X"49",X"8E",X"7D",X"B4",X"A6",
		X"2D",X"7E",X"D0",X"66",X"AE",X"4B",X"EC",X"C8",X"15",X"8D",X"24",X"10",X"AE",X"C8",X"17",X"31",
		X"21",X"10",X"8C",X"7D",X"F3",X"25",X"04",X"10",X"8E",X"7D",X"EF",X"A6",X"A4",X"10",X"AF",X"C8",
		X"17",X"AB",X"C8",X"14",X"BD",X"7D",X"38",X"6A",X"C8",X"13",X"26",X"CD",X"6E",X"D8",X"10",X"34",
		X"04",X"5F",X"47",X"56",X"E3",X"0A",X"ED",X"0A",X"35",X"04",X"EB",X"0C",X"E7",X"0C",X"39",X"00",
		X"01",X"00",X"02",X"5F",X"20",X"0A",X"C6",X"0D",X"20",X"06",X"C6",X"1A",X"20",X"02",X"C6",X"27",
		X"AE",X"B8",X"0C",X"3A",X"AF",X"C8",X"13",X"A7",X"C8",X"15",X"35",X"06",X"ED",X"C8",X"10",X"86",
		X"08",X"8E",X"7E",X"17",X"7E",X"D0",X"66",X"8D",X"08",X"6A",X"C8",X"15",X"26",X"F1",X"6E",X"D8",
		X"10",X"AE",X"4B",X"10",X"AE",X"C8",X"13",X"EC",X"21",X"8D",X"B4",X"A6",X"A4",X"44",X"44",X"BD",
		X"7D",X"38",X"31",X"23",X"E6",X"A4",X"C1",X"FF",X"26",X"02",X"31",X"34",X"10",X"AF",X"C8",X"13",
		X"39",X"00",X"0E",X"0C",X"04",X"7D",X"F3",X"7D",X"F6",X"7D",X"FA",X"7D",X"FE",X"00",X"18",X"1A",
		X"CB",X"01",X"04",X"00",X"10",X"0C",X"04",X"7D",X"F3",X"7D",X"F6",X"7D",X"FA",X"7D",X"FE",X"00",
		X"18",X"00",X"12",X"0C",X"04",X"7D",X"F3",X"7D",X"F6",X"7D",X"FA",X"7D",X"FE",X"00",X"18",X"00",
		X"14",X"0C",X"04",X"7D",X"F3",X"7D",X"F6",X"7D",X"FA",X"7D",X"FE",X"00",X"16",X"1A",X"C3",X"0C",
		X"04",X"7D",X"76",X"7D",X"7F",X"7D",X"89",X"7D",X"92",X"02",X"08",X"38",X"91",X"03",X"04",X"38",
		X"93",X"24",X"04",X"11",X"48",X"06",X"04",X"26",X"D5",X"0C",X"04",X"7D",X"76",X"7D",X"7F",X"7D",
		X"89",X"7D",X"92",X"01",X"02",X"4B",X"06",X"09",X"04",X"11",X"46",X"08",X"04",X"4B",X"08",X"05",
		X"06",X"4B",X"0A",X"04",X"04",X"00",X"0C",X"05",X"04",X"00",X"1A",X"01",X"04",X"0D",X"F4",X"26",
		X"05",X"0C",X"F4",X"7E",X"79",X"9D",X"0C",X"F4",X"CC",X"10",X"05",X"8E",X"50",X"EE",X"BD",X"D0",
		X"1B",X"D6",X"51",X"E7",X"47",X"86",X"7F",X"8D",X"55",X"86",X"20",X"A7",X"4A",X"86",X"08",X"8E",
		X"7E",X"E5",X"7E",X"D0",X"66",X"8D",X"39",X"96",X"51",X"A1",X"47",X"26",X"D0",X"6A",X"4A",X"26",
		X"EC",X"8E",X"CC",X"00",X"BD",X"D0",X"A5",X"5D",X"27",X"DF",X"8D",X"47",X"86",X"7D",X"8D",X"2E",
		X"86",X"0A",X"A7",X"4A",X"96",X"51",X"A1",X"47",X"27",X"04",X"8D",X"37",X"20",X"AF",X"86",X"08",
		X"8E",X"7F",X"16",X"7E",X"D0",X"66",X"8D",X"08",X"6A",X"4A",X"26",X"E8",X"8D",X"25",X"20",X"A8",
		X"96",X"F4",X"2B",X"09",X"B6",X"C8",X"04",X"81",X"41",X"10",X"27",X"FB",X"57",X"39",X"34",X"06",
		X"96",X"D0",X"D6",X"CF",X"34",X"06",X"EC",X"62",X"BD",X"5F",X"96",X"35",X"06",X"97",X"D0",X"D7",
		X"CF",X"35",X"86",X"34",X"16",X"8E",X"20",X"EE",X"CC",X"50",X"05",X"BD",X"D0",X"1B",X"35",X"96",
		X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",
		X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"2E",X"20",
		X"20",X"22",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",X"3A",X"20",X"32",X"30",X"38",X"34",
		X"22",X"20",X"20",X"01",X"38",X"80",X"07",X"DD",X"49",X"4E",X"53",X"50",X"49",X"52",X"45",X"44",
		X"20",X"42",X"59",X"20",X"48",X"49",X"53",X"20",X"4E",X"45",X"56",X"45",X"52",X"20",X"45",X"4E",
		X"44",X"49",X"4E",X"47",X"02",X"51",X"55",X"45",X"53",X"54",X"20",X"46",X"4F",X"52",X"20",X"50",
		X"52",X"4F",X"47",X"52",X"45",X"53",X"53",X"3C",X"02",X"49",X"4E",X"20",X"07",X"AA",X"32",X"30",
		X"38",X"34",X"07",X"DD",X"20",X"4D",X"41",X"4E",X"20",X"50",X"45",X"52",X"46",X"45",X"43",X"54",
		X"53",X"20",X"54",X"48",X"45",X"20",X"07",X"AA",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",
		X"53",X"3F",X"04",X"20",X"02",X"02",X"07",X"FF",X"41",X"20",X"52",X"4F",X"42",X"4F",X"54",X"20",
		X"53",X"50",X"45",X"43",X"49",X"45",X"53",X"20",X"53",X"4F",X"20",X"41",X"44",X"56",X"41",X"4E",
		X"43",X"45",X"44",X"20",X"54",X"48",X"41",X"54",X"02",X"4D",X"41",X"4E",X"20",X"49",X"53",X"20",
		X"49",X"4E",X"46",X"45",X"52",X"49",X"4F",X"52",X"20",X"54",X"4F",X"20",X"48",X"49",X"53",X"20",
		X"4F",X"57",X"4E",X"20",X"43",X"52",X"45",X"41",X"54",X"49",X"4F",X"4E",X"3D",X"02",X"02",X"04",
		X"20",X"07",X"DD",X"47",X"55",X"49",X"44",X"45",X"44",X"20",X"42",X"59",X"20",X"54",X"48",X"45",
		X"49",X"52",X"20",X"49",X"4E",X"46",X"41",X"4C",X"4C",X"49",X"42",X"4C",X"45",X"20",X"4C",X"4F",
		X"47",X"49",X"43",X"3C",X"02",X"54",X"48",X"45",X"20",X"07",X"AA",X"52",X"4F",X"42",X"4F",X"54",
		X"52",X"4F",X"4E",X"53",X"07",X"DD",X"20",X"43",X"4F",X"4E",X"43",X"4C",X"55",X"44",X"45",X"3F",
		X"02",X"02",X"04",X"30",X"07",X"AA",X"54",X"48",X"45",X"20",X"48",X"55",X"4D",X"41",X"4E",X"20",
		X"52",X"41",X"43",X"45",X"20",X"49",X"53",X"20",X"49",X"4E",X"45",X"46",X"46",X"49",X"43",X"49",
		X"45",X"4E",X"54",X"3C",X"02",X"41",X"4E",X"44",X"20",X"54",X"48",X"45",X"52",X"45",X"46",X"4F",
		X"52",X"45",X"20",X"4D",X"55",X"53",X"54",X"20",X"42",X"45",X"20",X"44",X"45",X"53",X"54",X"52",
		X"4F",X"59",X"45",X"44",X"3D",X"70",X"01",X"36",X"C0",X"07",X"DD",X"03",X"83",X"B7",X"59",X"4F",
		X"55",X"20",X"41",X"52",X"45",X"20",X"54",X"48",X"45",X"20",X"4C",X"41",X"53",X"54",X"20",X"48",
		X"4F",X"50",X"45",X"20",X"4F",X"46",X"20",X"4D",X"41",X"4E",X"4B",X"49",X"4E",X"44",X"3D",X"02",
		X"02",X"60",X"07",X"FF",X"44",X"55",X"45",X"20",X"54",X"4F",X"20",X"41",X"20",X"47",X"45",X"4E",
		X"45",X"54",X"49",X"43",X"20",X"45",X"4E",X"47",X"49",X"4E",X"45",X"45",X"52",X"49",X"4E",X"47",
		X"20",X"45",X"52",X"52",X"4F",X"52",X"3C",X"02",X"59",X"4F",X"55",X"20",X"50",X"4F",X"53",X"53",
		X"45",X"53",X"53",X"20",X"53",X"55",X"50",X"45",X"52",X"48",X"55",X"4D",X"41",X"4E",X"20",X"50",
		X"4F",X"57",X"45",X"52",X"53",X"3D",X"07",X"DD",X"02",X"02",X"59",X"4F",X"55",X"52",X"20",X"4D",
		X"49",X"53",X"53",X"49",X"4F",X"4E",X"20",X"49",X"53",X"20",X"54",X"4F",X"07",X"AA",X"20",X"53",
		X"54",X"4F",X"50",X"20",X"54",X"48",X"45",X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",
		X"53",X"3C",X"02",X"07",X"DD",X"41",X"4E",X"44",X"20",X"07",X"AA",X"53",X"41",X"56",X"45",X"20",
		X"54",X"48",X"45",X"20",X"4C",X"41",X"53",X"54",X"20",X"48",X"55",X"4D",X"41",X"4E",X"20",X"46",
		X"41",X"4D",X"49",X"4C",X"59",X"3F",X"03",X"84",X"77",X"04",X"20",X"05",X"1C",X"73",X"04",X"58",
		X"05",X"18",X"74",X"04",X"58",X"05",X"14",X"75",X"70",X"05",X"10",X"7E",X"70",X"01",X"58",X"80",
		X"07",X"33",X"08",X"54",X"48",X"45",X"20",X"46",X"4F",X"52",X"43",X"45",X"20",X"4F",X"46",X"20",
		X"47",X"52",X"4F",X"55",X"4E",X"44",X"20",X"52",X"4F",X"56",X"49",X"4E",X"47",X"02",X"55",X"4E",
		X"49",X"54",X"20",X"4E",X"45",X"54",X"57",X"4F",X"52",X"4B",X"20",X"54",X"45",X"52",X"4D",X"49",
		X"4E",X"41",X"54",X"4F",X"52",X"20",X"02",X"07",X"AA",X"05",X"74",X"76",X"5B",X"47",X"52",X"55",
		X"4E",X"54",X"5C",X"3A",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",X"53",X"07",X"33",X"20",
		X"53",X"45",X"45",X"4B",X"20",X"54",X"4F",X"02",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"20",
		X"59",X"4F",X"55",X"3D",X"FF",X"01",X"58",X"80",X"07",X"55",X"03",X"85",X"A1",X"54",X"48",X"45",
		X"07",X"AA",X"05",X"14",X"77",X"20",X"48",X"55",X"4C",X"4B",X"20",X"52",X"4F",X"42",X"4F",X"54",
		X"52",X"4F",X"4E",X"53",X"20",X"07",X"55",X"53",X"45",X"45",X"4B",X"20",X"4F",X"55",X"54",X"02",
		X"41",X"4E",X"44",X"20",X"45",X"4C",X"49",X"4D",X"49",X"4E",X"41",X"54",X"45",X"20",X"54",X"48",
		X"45",X"20",X"4C",X"41",X"53",X"54",X"20",X"48",X"55",X"4D",X"41",X"4E",X"20",X"46",X"41",X"4D",
		X"49",X"4C",X"59",X"3D",X"F9",X"05",X"14",X"7E",X"80",X"01",X"70",X"80",X"07",X"DD",X"03",X"85",
		X"BD",X"54",X"48",X"45",X"07",X"AA",X"05",X"2C",X"78",X"20",X"53",X"50",X"48",X"45",X"52",X"45",
		X"4F",X"49",X"44",X"53",X"20",X"41",X"4E",X"44",X"20",X"51",X"55",X"41",X"52",X"4B",X"53",X"20",
		X"20",X"07",X"DD",X"02",X"41",X"52",X"45",X"20",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"4D",
		X"45",X"44",X"20",X"54",X"4F",X"20",X"4D",X"41",X"4E",X"55",X"46",X"41",X"43",X"54",X"55",X"52",
		X"45",X"02",X"07",X"AA",X"05",X"33",X"79",X"45",X"4E",X"46",X"4F",X"52",X"43",X"45",X"52",X"20",
		X"41",X"4E",X"44",X"20",X"54",X"41",X"4E",X"4B",X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",
		X"4E",X"53",X"3D",X"A0",X"05",X"10",X"7E",X"01",X"58",X"80",X"07",X"FF",X"42",X"45",X"57",X"41",
		X"52",X"45",X"20",X"4F",X"46",X"20",X"54",X"48",X"45",X"20",X"49",X"4E",X"47",X"45",X"4E",X"49",
		X"4F",X"55",X"53",X"02",X"07",X"AA",X"05",X"20",X"7A",X"42",X"52",X"41",X"49",X"4E",X"20",X"52",
		X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",X"53",X"07",X"FF",X"20",X"54",X"48",X"41",X"54",X"20",
		X"50",X"4F",X"53",X"53",X"45",X"53",X"53",X"02",X"54",X"48",X"45",X"20",X"50",X"4F",X"57",X"45",
		X"52",X"20",X"54",X"4F",X"20",X"52",X"45",X"50",X"52",X"4F",X"47",X"52",X"41",X"4D",X"02",X"48",
		X"55",X"4D",X"41",X"4E",X"53",X"20",X"49",X"4E",X"54",X"4F",X"20",X"53",X"49",X"4E",X"49",X"53",
		X"54",X"45",X"52",X"20",X"07",X"AA",X"50",X"52",X"4F",X"47",X"53",X"3D",X"73",X"05",X"2C",X"7C",
		X"80",X"03",X"86",X"CC",X"01",X"64",X"80",X"04",X"20",X"05",X"10",X"7E",X"04",X"40",X"07",X"DD",
		X"41",X"53",X"20",X"59",X"4F",X"55",X"20",X"53",X"54",X"52",X"55",X"47",X"47",X"4C",X"45",X"20",
		X"54",X"4F",X"20",X"53",X"41",X"56",X"45",X"02",X"48",X"55",X"4D",X"41",X"4E",X"49",X"54",X"59",
		X"3C",X"20",X"42",X"45",X"20",X"53",X"55",X"52",X"45",X"20",X"54",X"4F",X"20",X"41",X"56",X"4F",
		X"49",X"44",X"02",X"07",X"AA",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"44",X"45",X"53",X"07",
		X"DD",X"20",X"49",X"4E",X"20",X"59",X"4F",X"55",X"52",X"20",X"50",X"41",X"54",X"48",X"3D",X"D0",
		X"AD",X"06",X"03",X"87",X"15",X"FF",X"09",X"01",X"7E",X"97",X"07",X"18",X"A0",X"15",X"84",X"0F",
		X"04",X"60",X"02",X"06",X"0B",X"90",X"0B",X"FF",X"0B",X"FF",X"03",X"50",X"04",X"68",X"02",X"03",
		X"0B",X"80",X"0B",X"80",X"02",X"06",X"0B",X"40",X"03",X"18",X"05",X"23",X"02",X"00",X"0B",X"FF",
		X"02",X"06",X"0B",X"E0",X"06",X"3C",X"02",X"03",X"0B",X"38",X"05",X"38",X"02",X"03",X"0B",X"20",
		X"02",X"06",X"0B",X"E3",X"06",X"20",X"02",X"00",X"0B",X"3C",X"02",X"06",X"0B",X"F1",X"0B",X"30",
		X"05",X"20",X"02",X"00",X"0B",X"20",X"02",X"06",X"0B",X"90",X"0B",X"90",X"04",X"80",X"0D",X"0B",
		X"FF",X"0B",X"60",X"13",X"1D",X"05",X"14",X"0A",X"84",X"13",X"12",X"1B",X"05",X"14",X"08",X"84",
		X"1A",X"13",X"1D",X"05",X"14",X"14",X"84",X"21",X"12",X"1B",X"05",X"14",X"05",X"84",X"28",X"13",
		X"1D",X"05",X"14",X"0A",X"84",X"2F",X"0B",X"FF",X"0B",X"FF",X"0B",X"50",X"13",X"0B",X"10",X"14",
		X"0E",X"84",X"3C",X"0B",X"E0",X"12",X"0B",X"0B",X"14",X"0A",X"84",X"45",X"0B",X"FF",X"0B",X"E3",
		X"0B",X"10",X"13",X"0E",X"80",X"13",X"18",X"08",X"13",X"20",X"08",X"14",X"03",X"84",X"58",X"0B",
		X"FF",X"0B",X"44",X"12",X"09",X"C0",X"0B",X"E0",X"12",X"08",X"FF",X"0B",X"90",X"13",X"04",X"10",
		X"13",X"06",X"10",X"13",X"08",X"01",X"17",X"01",X"7E",X"41",X"07",X"18",X"A0",X"11",X"84",X"AD",
		X"11",X"84",X"C6",X"04",X"28",X"0F",X"01",X"7E",X"B5",X"02",X"00",X"16",X"00",X"04",X"10",X"0B",
		X"30",X"0F",X"01",X"7E",X"53",X"07",X"18",X"A0",X"0B",X"40",X"10",X"04",X"30",X"06",X"10",X"04",
		X"10",X"05",X"13",X"03",X"12",X"0F",X"01",X"7E",X"B9",X"10",X"0B",X"80",X"0C",X"01",X"7E",X"53",
		X"07",X"18",X"A0",X"0F",X"0B",X"70",X"10",X"04",X"1E",X"0F",X"01",X"7E",X"B5",X"02",X"01",X"16",
		X"00",X"04",X"10",X"0B",X"30",X"0C",X"01",X"7E",X"61",X"07",X"18",X"A0",X"0F",X"0B",X"D8",X"10",
		X"04",X"15",X"0F",X"01",X"7E",X"B5",X"02",X"02",X"16",X"00",X"04",X"10",X"0B",X"30",X"0F",X"01",
		X"7E",X"61",X"07",X"18",X"A0",X"0B",X"C0",X"10",X"04",X"04",X"05",X"08",X"04",X"10",X"05",X"18",
		X"03",X"01",X"0E",X"84",X"A5",X"01",X"7E",X"8B",X"07",X"86",X"85",X"0B",X"10",X"16",X"FE",X"04",
		X"02",X"01",X"0B",X"08",X"16",X"FD",X"04",X"02",X"00",X"0B",X"20",X"16",X"FE",X"04",X"02",X"02",
		X"14",X"02",X"84",X"FB",X"0E",X"85",X"8B",X"01",X"7E",X"8B",X"07",X"88",X"90",X"0B",X"09",X"16",
		X"FE",X"02",X"02",X"02",X"0B",X"12",X"16",X"FE",X"02",X"02",X"00",X"0B",X"12",X"16",X"FE",X"02",
		X"02",X"01",X"0B",X"0B",X"16",X"FE",X"02",X"02",X"00",X"14",X"02",X"85",X"1D",X"0E",X"85",X"8B",
		X"01",X"7E",X"8B",X"07",X"88",X"BC",X"0B",X"10",X"16",X"FE",X"FD",X"02",X"01",X"0B",X"06",X"16",
		X"FE",X"FD",X"02",X"00",X"0B",X"1A",X"16",X"FE",X"FD",X"02",X"02",X"0B",X"08",X"16",X"FE",X"FD",
		X"14",X"02",X"85",X"46",X"0E",X"85",X"8B",X"01",X"7E",X"8B",X"07",X"88",X"B1",X"0B",X"04",X"16",
		X"FE",X"FE",X"02",X"01",X"0B",X"09",X"16",X"FD",X"FE",X"02",X"00",X"0B",X"18",X"16",X"FE",X"FE",
		X"02",X"02",X"0B",X"15",X"16",X"FE",X"FE",X"14",X"02",X"85",X"74",X"02",X"00",X"16",X"FC",X"02",
		X"0B",X"04",X"02",X"02",X"16",X"FE",X"FE",X"0B",X"20",X"02",X"00",X"16",X"FC",X"02",X"0B",X"12",
		X"0D",X"01",X"7E",X"6F",X"07",X"10",X"C0",X"15",X"85",X"B1",X"04",X"1C",X"06",X"10",X"04",X"36",
		X"0C",X"0B",X"7C",X"16",X"FE",X"00",X"0B",X"0B",X"14",X"0A",X"85",X"B3",X"17",X"01",X"7E",X"A9",
		X"07",X"88",X"87",X"11",X"85",X"D6",X"11",X"85",X"E3",X"11",X"86",X"03",X"11",X"86",X"1A",X"08",
		X"FF",X"40",X"0A",X"02",X"60",X"0C",X"01",X"7E",X"A5",X"07",X"0A",X"B4",X"08",X"00",X"C0",X"0A",
		X"02",X"60",X"0C",X"01",X"7E",X"AD",X"07",X"10",X"B4",X"0F",X"0B",X"10",X"10",X"0B",X"14",X"16",
		X"00",X"FF",X"18",X"14",X"03",X"85",X"ED",X"0F",X"01",X"7E",X"B1",X"10",X"08",X"00",X"80",X"0A",
		X"02",X"70",X"0D",X"01",X"7E",X"93",X"07",X"80",X"87",X"0F",X"0B",X"10",X"10",X"0B",X"14",X"18",
		X"14",X"05",X"86",X"0D",X"08",X"FF",X"A0",X"0B",X"30",X"0D",X"01",X"7E",X"41",X"07",X"0A",X"B4",
		X"0F",X"0B",X"C0",X"10",X"04",X"20",X"11",X"86",X"8D",X"05",X"0A",X"03",X"08",X"04",X"1A",X"16",
		X"03",X"FE",X"0B",X"02",X"15",X"86",X"8C",X"19",X"AA",X"BB",X"28",X"00",X"11",X"86",X"48",X"08",
		X"02",X"00",X"19",X"00",X"AA",X"2C",X"00",X"0C",X"01",X"7E",X"41",X"07",X"31",X"BC",X"02",X"03",
		X"0F",X"0B",X"03",X"11",X"86",X"66",X"11",X"86",X"7B",X"0B",X"04",X"10",X"08",X"02",X"00",X"19",
		X"EE",X"00",X"2C",X"00",X"00",X"0C",X"01",X"7E",X"41",X"07",X"31",X"BC",X"0F",X"0B",X"04",X"02",
		X"03",X"10",X"08",X"02",X"00",X"19",X"EE",X"00",X"2C",X"00",X"0C",X"01",X"7E",X"41",X"07",X"31",
		X"BC",X"02",X"03",X"08",X"02",X"00",X"19",X"EE",X"00",X"2C",X"00",X"0C",X"1A",X"01",X"7E",X"7D",
		X"07",X"0A",X"A0",X"04",X"10",X"11",X"86",X"A4",X"05",X"0C",X"04",X"10",X"19",X"BB",X"BB",X"38",
		X"01",X"04",X"0B",X"0D",X"01",X"86",X"B0",X"07",X"1A",X"A4",X"08",X"00",X"60",X"0B",X"40",X"0C",
		X"86",X"B4",X"01",X"04",X"86",X"B6",X"09",X"02",X"86",X"BA",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DA",X"A0",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DA",X"A0",X"01",X"7E",X"8F",X"07",
		X"86",X"C1",X"02",X"0C",X"0F",X"0B",X"48",X"11",X"86",X"ED",X"0B",X"0A",X"11",X"86",X"F9",X"0B",
		X"0A",X"11",X"87",X"07",X"0B",X"10",X"10",X"19",X"00",X"DD",X"B8",X"00",X"1B",X"01",X"7E",X"8F",
		X"07",X"68",X"C1",X"19",X"00",X"FF",X"8D",X"00",X"1B",X"01",X"7E",X"8F",X"07",X"72",X"C1",X"02",
		X"04",X"19",X"00",X"AA",X"91",X"00",X"1B",X"01",X"7E",X"8F",X"07",X"7C",X"C1",X"02",X"08",X"19",
		X"00",X"CC",X"92",X"00",X"1B",X"01",X"7E",X"41",X"07",X"50",X"68",X"11",X"87",X"39",X"11",X"87",
		X"42",X"11",X"87",X"5B",X"11",X"87",X"74",X"11",X"87",X"8D",X"04",X"09",X"0F",X"01",X"7E",X"B5",
		X"02",X"00",X"16",X"00",X"05",X"10",X"0B",X"50",X"0C",X"01",X"7E",X"97",X"07",X"68",X"6A",X"03",
		X"80",X"0C",X"01",X"7E",X"53",X"07",X"48",X"69",X"0F",X"0B",X"10",X"10",X"04",X"0A",X"0F",X"01",
		X"7E",X"B5",X"02",X"01",X"16",X"00",X"04",X"10",X"0B",X"50",X"0C",X"01",X"7E",X"61",X"07",X"40",
		X"6B",X"0F",X"0B",X"20",X"10",X"04",X"0C",X"0F",X"01",X"7E",X"B5",X"02",X"02",X"16",X"00",X"02",
		X"10",X"0B",X"50",X"0C",X"01",X"7E",X"41",X"07",X"38",X"68",X"0F",X"0B",X"30",X"10",X"04",X"0D",
		X"0F",X"01",X"7E",X"B5",X"02",X"03",X"16",X"00",X"05",X"10",X"0B",X"50",X"0C",X"01",X"7E",X"61",
		X"07",X"30",X"6B",X"0F",X"0B",X"40",X"10",X"04",X"0F",X"0F",X"01",X"7E",X"B5",X"02",X"04",X"16",
		X"00",X"02",X"10",X"0B",X"50",X"0C",X"BD",X"D0",X"30",X"96",X"59",X"8A",X"04",X"97",X"59",X"BD",
		X"D0",X"54",X"78",X"D6",X"BD",X"8A",X"3A",X"BD",X"D0",X"54",X"87",X"F8",X"BD",X"78",X"6F",X"26",
		X"15",X"BD",X"D0",X"54",X"8A",X"4F",X"86",X"FF",X"8E",X"87",X"CE",X"7E",X"D0",X"66",X"86",X"FF",
		X"8E",X"79",X"9B",X"7E",X"D0",X"66",X"BD",X"88",X"BF",X"86",X"1C",X"DE",X"15",X"A7",X"47",X"9E",
		X"E6",X"96",X"E9",X"BD",X"8A",X"19",X"BD",X"89",X"6C",X"86",X"04",X"8E",X"87",X"F1",X"7E",X"D0",
		X"66",X"6A",X"47",X"26",X"EA",X"7E",X"88",X"CD",X"BD",X"6F",X"06",X"27",X"13",X"BE",X"6F",X"0F",
		X"10",X"8E",X"B3",X"EA",X"EC",X"81",X"ED",X"A1",X"10",X"8C",X"B4",X"1E",X"25",X"F6",X"20",X"12",
		X"8E",X"CC",X"24",X"10",X"8E",X"B3",X"EA",X"BD",X"D0",X"A8",X"ED",X"A1",X"10",X"8C",X"B4",X"1E",
		X"25",X"F5",X"B6",X"B4",X"1C",X"C6",X"86",X"10",X"8E",X"B3",X"EA",X"8D",X"15",X"B6",X"B4",X"1D",
		X"C6",X"96",X"10",X"8E",X"B4",X"03",X"8D",X"0A",X"D6",X"51",X"86",X"70",X"BD",X"5F",X"96",X"7E",
		X"D0",X"63",X"35",X"10",X"DE",X"15",X"AF",X"47",X"1F",X"01",X"86",X"19",X"A7",X"49",X"86",X"66",
		X"97",X"CF",X"A6",X"A0",X"BD",X"5F",X"93",X"AF",X"4A",X"10",X"AF",X"4C",X"86",X"02",X"8E",X"88",
		X"64",X"7E",X"D0",X"66",X"AE",X"4A",X"10",X"AE",X"4C",X"6A",X"49",X"26",X"E5",X"6E",X"D8",X"07",
		X"20",X"52",X"4F",X"42",X"4F",X"54",X"52",X"4F",X"4E",X"3A",X"20",X"32",X"30",X"38",X"34",X"20",
		X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",
		X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"BD",
		X"89",X"4B",X"10",X"8E",X"B4",X"26",X"86",X"10",X"8D",X"6A",X"7E",X"89",X"4B",X"8D",X"F0",X"BD",
		X"D0",X"54",X"8A",X"4F",X"DE",X"15",X"8E",X"02",X"C0",X"AF",X"4D",X"86",X"06",X"A7",X"4B",X"9E",
		X"E6",X"96",X"E9",X"20",X"0A",X"86",X"06",X"A7",X"4B",X"BD",X"89",X"6C",X"BD",X"89",X"E6",X"10",
		X"9E",X"EB",X"F6",X"CB",X"00",X"D7",X"2B",X"E1",X"21",X"25",X"0E",X"E0",X"21",X"C1",X"14",X"23",
		X"EE",X"D6",X"2B",X"C1",X"EC",X"24",X"E8",X"20",X"0D",X"E6",X"21",X"C1",X"1E",X"23",X"E0",X"F0",
		X"CB",X"00",X"C1",X"1E",X"23",X"D9",X"BD",X"89",X"F8",X"BD",X"8A",X"19",X"DE",X"15",X"6A",X"4B",
		X"26",X"C7",X"AE",X"4D",X"30",X"1F",X"10",X"27",X"F0",X"71",X"AF",X"4D",X"86",X"01",X"8E",X"88",
		X"E5",X"7E",X"D0",X"66",X"34",X"22",X"9E",X"E6",X"35",X"02",X"34",X"10",X"5F",X"CE",X"8C",X"F4",
		X"BD",X"8D",X"69",X"35",X"30",X"CC",X"0E",X"1B",X"7E",X"D0",X"B7",X"34",X"16",X"86",X"05",X"C6",
		X"0F",X"DD",X"E6",X"0F",X"E8",X"0F",X"EA",X"86",X"77",X"97",X"E9",X"8E",X"B5",X"AE",X"9F",X"EB",
		X"CC",X"13",X"AF",X"ED",X"81",X"8C",X"B5",X"E6",X"25",X"F9",X"35",X"96",X"34",X"04",X"96",X"E8",
		X"84",X"03",X"4A",X"2B",X"4E",X"4A",X"2B",X"3B",X"4A",X"2B",X"24",X"DC",X"E6",X"C0",X"20",X"25",
		X"04",X"C1",X"0F",X"22",X"4F",X"96",X"EA",X"8B",X"02",X"81",X"10",X"25",X"08",X"0F",X"EA",X"86",
		X"15",X"C6",X"0F",X"20",X"3D",X"97",X"EA",X"C6",X"0F",X"86",X"05",X"9B",X"EA",X"20",X"33",X"DC",
		X"E6",X"80",X"10",X"25",X"04",X"81",X"05",X"22",X"2B",X"86",X"05",X"D6",X"EA",X"50",X"58",X"CB",
		X"CF",X"20",X"1F",X"DC",X"E6",X"CB",X"20",X"C1",X"CF",X"25",X"19",X"C6",X"CF",X"86",X"85",X"90",
		X"EA",X"20",X"0F",X"DC",X"E6",X"8B",X"10",X"81",X"85",X"25",X"09",X"86",X"85",X"D6",X"EA",X"58",
		X"CB",X"0F",X"0C",X"E8",X"DD",X"E6",X"1F",X"01",X"96",X"E9",X"80",X"11",X"25",X"02",X"26",X"02",
		X"86",X"77",X"97",X"E9",X"35",X"84",X"34",X"10",X"9E",X"EB",X"30",X"02",X"8C",X"B5",X"E6",X"25",
		X"03",X"8E",X"B5",X"AE",X"9F",X"EB",X"35",X"90",X"34",X"17",X"AE",X"9F",X"98",X"EB",X"1A",X"10",
		X"BF",X"CA",X"04",X"CC",X"0A",X"1F",X"FD",X"CA",X"06",X"7F",X"CA",X"01",X"CC",X"B4",X"26",X"FD",
		X"CA",X"02",X"86",X"1E",X"B7",X"CA",X"00",X"35",X"97",X"34",X"03",X"AF",X"9F",X"98",X"EB",X"1A",
		X"10",X"B7",X"CA",X"01",X"BF",X"CA",X"04",X"CC",X"0A",X"1F",X"FD",X"CA",X"06",X"CC",X"B4",X"26",
		X"FD",X"CA",X"02",X"86",X"1E",X"B7",X"CA",X"00",X"35",X"83",X"34",X"32",X"8E",X"8A",X"70",X"10",
		X"8E",X"98",X"01",X"A6",X"80",X"A7",X"A0",X"10",X"8C",X"98",X"08",X"25",X"F6",X"35",X"B2",X"8E",
		X"98",X"01",X"AF",X"49",X"8D",X"E4",X"AE",X"49",X"30",X"01",X"8C",X"98",X"08",X"25",X"03",X"8E",
		X"98",X"01",X"AF",X"49",X"86",X"FF",X"A7",X"84",X"86",X"03",X"8E",X"8A",X"54",X"7E",X"D0",X"66",
		X"07",X"C0",X"17",X"30",X"C7",X"1F",X"3F",X"01",X"39",X"90",X"22",X"57",X"22",X"90",X"21",X"59",
		X"21",X"90",X"21",X"43",X"27",X"4F",X"21",X"90",X"21",X"43",X"21",X"05",X"22",X"4D",X"22",X"90",
		X"21",X"43",X"21",X"06",X"21",X"42",X"2C",X"90",X"21",X"43",X"21",X"06",X"21",X"42",X"21",X"90",
		X"C6",X"21",X"43",X"22",X"05",X"21",X"42",X"21",X"90",X"21",X"44",X"27",X"42",X"21",X"90",X"21",
		X"4D",X"21",X"90",X"23",X"4B",X"22",X"90",X"02",X"2A",X"43",X"2B",X"90",X"0A",X"22",X"4D",X"22",
		X"90",X"0B",X"22",X"4C",X"22",X"90",X"0C",X"2E",X"90",X"A0",X"01",X"39",X"90",X"22",X"57",X"22",
		X"90",X"21",X"59",X"21",X"90",X"21",X"43",X"33",X"43",X"21",X"90",X"21",X"42",X"22",X"11",X"22",
		X"42",X"21",X"90",X"21",X"42",X"21",X"13",X"21",X"42",X"21",X"90",X"C8",X"21",X"42",X"24",X"10",
		X"21",X"42",X"21",X"90",X"21",X"45",X"22",X"0F",X"21",X"42",X"21",X"90",X"21",X"46",X"22",X"0D",
		X"22",X"42",X"21",X"90",X"21",X"47",X"2F",X"43",X"21",X"90",X"21",X"59",X"21",X"90",X"22",X"57",
		X"22",X"90",X"01",X"39",X"90",X"A0",X"01",X"39",X"90",X"22",X"57",X"21",X"90",X"21",X"58",X"22",
		X"90",X"21",X"42",X"27",X"50",X"21",X"90",X"21",X"42",X"21",X"05",X"22",X"4F",X"21",X"90",X"21",
		X"42",X"21",X"06",X"21",X"4F",X"21",X"90",X"21",X"42",X"21",X"06",X"21",X"43",X"29",X"43",X"21",
		X"90",X"21",X"42",X"21",X"06",X"21",X"42",X"22",X"07",X"22",X"42",X"21",X"90",X"21",X"42",X"21",
		X"06",X"21",X"42",X"21",X"09",X"21",X"42",X"21",X"90",X"C5",X"21",X"42",X"22",X"05",X"21",X"42",
		X"21",X"09",X"21",X"42",X"21",X"90",X"21",X"43",X"27",X"42",X"21",X"09",X"21",X"42",X"21",X"90",
		X"21",X"4C",X"21",X"09",X"21",X"42",X"21",X"90",X"22",X"4B",X"22",X"07",X"22",X"42",X"21",X"90",
		X"01",X"2A",X"43",X"29",X"43",X"21",X"90",X"0A",X"21",X"4E",X"22",X"90",X"0A",X"22",X"4B",X"23",
		X"90",X"0B",X"2D",X"90",X"A0",X"01",X"23",X"90",X"22",X"41",X"22",X"90",X"21",X"43",X"21",X"90",
		X"C4",X"21",X"43",X"22",X"90",X"21",X"44",X"35",X"90",X"21",X"58",X"22",X"90",X"21",X"59",X"21",
		X"90",X"C1",X"21",X"44",X"27",X"4D",X"22",X"90",X"21",X"43",X"22",X"05",X"2F",X"90",X"21",X"43",
		X"21",X"90",X"C4",X"22",X"41",X"22",X"90",X"01",X"23",X"90",X"A0",X"01",X"39",X"90",X"22",X"57",
		X"22",X"90",X"21",X"59",X"21",X"90",X"21",X"42",X"28",X"4F",X"21",X"90",X"21",X"42",X"21",X"06",
		X"21",X"4F",X"21",X"90",X"21",X"42",X"21",X"06",X"22",X"4C",X"22",X"90",X"21",X"42",X"21",X"07",
		X"2E",X"90",X"21",X"42",X"21",X"90",X"C8",X"21",X"42",X"37",X"90",X"21",X"58",X"22",X"90",X"22",
		X"57",X"22",X"90",X"01",X"39",X"90",X"A0",X"03",X"24",X"0E",X"24",X"90",X"02",X"22",X"42",X"22",
		X"0C",X"22",X"42",X"22",X"90",X"02",X"21",X"44",X"21",X"0C",X"21",X"44",X"21",X"90",X"C5",X"02",
		X"22",X"42",X"22",X"0C",X"22",X"42",X"22",X"90",X"03",X"24",X"0E",X"24",X"90",X"A0",X"01",X"21",
		X"4C",X"23",X"4C",X"21",X"90",X"02",X"21",X"4C",X"21",X"4C",X"21",X"90",X"03",X"21",X"57",X"21",
		X"90",X"04",X"21",X"55",X"21",X"90",X"05",X"21",X"43",X"26",X"41",X"26",X"43",X"21",X"90",X"06",
		X"21",X"43",X"21",X"04",X"21",X"04",X"21",X"43",X"21",X"90",X"07",X"21",X"43",X"21",X"03",X"21",
		X"03",X"21",X"43",X"21",X"90",X"08",X"21",X"43",X"23",X"41",X"23",X"43",X"21",X"90",X"09",X"21",
		X"4B",X"21",X"90",X"0A",X"21",X"49",X"21",X"90",X"0B",X"21",X"43",X"21",X"43",X"21",X"90",X"0C",
		X"28",X"90",X"A0",X"0D",X"21",X"45",X"21",X"90",X"0C",X"21",X"46",X"21",X"90",X"0B",X"21",X"47",
		X"21",X"90",X"0A",X"21",X"48",X"21",X"90",X"09",X"21",X"45",X"21",X"43",X"21",X"90",X"08",X"21",
		X"45",X"22",X"43",X"21",X"90",X"08",X"21",X"44",X"21",X"01",X"21",X"43",X"21",X"90",X"08",X"21",
		X"43",X"21",X"02",X"21",X"43",X"21",X"90",X"08",X"21",X"43",X"24",X"43",X"25",X"90",X"08",X"21",
		X"4E",X"21",X"90",X"C3",X"08",X"28",X"43",X"25",X"90",X"0F",X"21",X"43",X"21",X"90",X"C3",X"0E",
		X"21",X"44",X"21",X"90",X"C4",X"0F",X"21",X"43",X"21",X"90",X"10",X"21",X"42",X"21",X"90",X"11",
		X"21",X"41",X"21",X"90",X"12",X"22",X"90",X"A0",X"F0",X"19",X"F0",X"1B",X"8C",X"F2",X"8C",X"2E",
		X"8C",X"83",X"00",X"00",X"0A",X"47",X"90",X"08",X"4B",X"90",X"06",X"4F",X"90",X"05",X"51",X"90",
		X"04",X"44",X"22",X"4D",X"90",X"03",X"47",X"22",X"4C",X"90",X"02",X"49",X"24",X"4A",X"90",X"02",
		X"4A",X"25",X"48",X"90",X"01",X"4C",X"27",X"46",X"90",X"01",X"4D",X"28",X"44",X"90",X"4D",X"27",
		X"47",X"90",X"48",X"22",X"42",X"26",X"49",X"90",X"49",X"27",X"4B",X"90",X"4A",X"24",X"4D",X"90",
		X"49",X"27",X"4B",X"90",X"48",X"22",X"42",X"26",X"49",X"90",X"4D",X"27",X"47",X"90",X"01",X"4D",
		X"28",X"44",X"90",X"01",X"4C",X"27",X"46",X"90",X"02",X"4A",X"25",X"48",X"90",X"02",X"49",X"24",
		X"4A",X"90",X"03",X"47",X"22",X"4C",X"90",X"04",X"44",X"22",X"4D",X"90",X"05",X"51",X"90",X"06",
		X"4F",X"90",X"08",X"4B",X"90",X"0A",X"47",X"90",X"A0",X"34",X"62",X"84",X"F0",X"34",X"02",X"44",
		X"44",X"44",X"44",X"AA",X"E0",X"97",X"DF",X"A6",X"E4",X"84",X"0F",X"34",X"02",X"48",X"48",X"48",
		X"48",X"AA",X"E0",X"97",X"E0",X"8D",X"04",X"24",X"FC",X"35",X"E2",X"A6",X"C4",X"43",X"85",X"C0",
		X"27",X"02",X"DF",X"E4",X"9F",X"DD",X"A6",X"C0",X"2A",X"27",X"85",X"20",X"27",X"03",X"1A",X"01",
		X"39",X"85",X"10",X"27",X"05",X"8D",X"5B",X"1C",X"FE",X"39",X"85",X"40",X"27",X"E8",X"84",X"0F",
		X"97",X"E1",X"DF",X"E2",X"DE",X"E4",X"8D",X"DC",X"0A",X"E1",X"26",X"F8",X"DE",X"E2",X"1C",X"FE",
		X"39",X"85",X"60",X"26",X"04",X"30",X"86",X"20",X"CD",X"34",X"03",X"84",X"1F",X"1A",X"10",X"BF",
		X"CA",X"04",X"30",X"86",X"88",X"04",X"B7",X"CA",X"07",X"86",X"05",X"B7",X"CA",X"06",X"FD",X"CA",
		X"02",X"A6",X"61",X"85",X"40",X"27",X"04",X"96",X"DF",X"20",X"02",X"96",X"E0",X"B7",X"CA",X"01",
		X"86",X"12",X"5D",X"27",X"04",X"8A",X"80",X"20",X"02",X"8A",X"40",X"B7",X"CA",X"00",X"35",X"03",
		X"20",X"94",X"9E",X"DD",X"5D",X"27",X"06",X"C6",X"FF",X"30",X"89",X"01",X"00",X"53",X"39",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
