-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "243C003C3C183C000606FFFFFFFF3C3C00000000FFFFFFFF0000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000004921FFFFB6DE00006969AAAAB6FE0000B6DE0000";
    attribute INIT_02 of inst : label is "D99BD99BC003C00303C003C0FFFF0000B49980080000000000000000B6DE0000";
    attribute INIT_03 of inst : label is "FFFFFFFF3FFC2AA8000000005B94A46803000300A768632413101B905BE58C32";
    attribute INIT_04 of inst : label is "33CC33CC2A2A2A2AD5D5D5D5BEBEBEBEFFFFFFFF2A2A2A2AC963E00BD5D5D5D5";
    attribute INIT_05 of inst : label is "C963E00BFFFFFFFFD557D557FFFFFFFF30EB7AD5999999990B9F600B318C0CCC";
    attribute INIT_06 of inst : label is "00000000000000006CDEDC7F9321238093212380932123809321238000000000";
    attribute INIT_07 of inst : label is "FFFFFFFF4146064203E000C003E000C0DEB707D0FC1FFF3F36F800C03FF800C0";
    attribute INIT_08 of inst : label is "9006003C90063C00C1800098C180009871C7F7DFC71CDF7DF7DFBAEBDF7DEBAE";
    attribute INIT_09 of inst : label is "BE140000BC160000B41E0000943E000014BE000016BC00001EB400003E940000";
    attribute INIT_0A of inst : label is "AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "FFFFAAAAFFFF0410FFFF1964FFFF73CDAAAAE6DB0410D9F71964F7BF73CDFF7F";
    attribute INIT_0E of inst : label is "000055500000FFF50000FFFF0000EABF5550D57FFFF5AAEAFFFF00C0EABF0080";
    attribute INIT_0F of inst : label is "000055500000FFF50000EABF0000807A555000E0FFF500C0EABF00C0807A0080";
    attribute INIT_10 of inst : label is "000055550000FBEF0000E69B00008C3255551924FBEF2608E69B08408C320080";
    attribute INIT_11 of inst : label is "000055550000FBEF0000E69B00008C3255551924FBEF2608E69B08408C320080";
    attribute INIT_12 of inst : label is "000055550000EEEE000099990000666655559999EEEE66669999999966666666";
    attribute INIT_13 of inst : label is "000055550000FFFF0000BEBE0000696955559286FFFF2148BEBE56C46969A888";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2FB007D0FFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F3DBDFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "03DB007D02FB003DC000000000000000FF6F07D02FB03DBD0000000000000000";
    attribute INIT_21 of inst : label is "003E00000002000FFFBC7D00FB0040B800FF0007002F003D6F00D000B000BD00";
    attribute INIT_22 of inst : label is "0CCC0C4CC4CC0CCC33303130331333301ED7AFFF17AF0A83AAA4F825FD75AAA0";
    attribute INIT_23 of inst : label is "C2DA6CFE03FF005CA783BF39FFC03500194103000AEB75758E90C000A000555D";
    attribute INIT_24 of inst : label is "000F0BBF042D02B4C000FF007AB07A0001FDBBFE02D709010000A000AC008000";
    attribute INIT_25 of inst : label is "0000000A0000000005C0BFE02D7B207A000000BB000200005C00FEA0D7AC1D00";
    attribute INIT_26 of inst : label is "036800FB003D00773000D000E50060003C830FD903DE01D40000000050000000";
    attribute INIT_27 of inst : label is "0003000000000000C230FD903DE57760003C000F0003001D8300D900DE507600";
    attribute INIT_28 of inst : label is "02660DEA00020022E000DE00FA0000002FFEDEAD002F01900000E000A0000000";
    attribute INIT_29 of inst : label is "0002000D00000000FFE0629E06FA2200002F004E00000000FE00ADE02FA00000";
    attribute INIT_2A of inst : label is "0003000200332BFFF400B000F3008B00003F002B030FAFF840000000F000B000";
    attribute INIT_2B of inst : label is "00000000000000AF03F402B03C0FFF8B0000000000032AFF7F402B00FC30F8B0";
    attribute INIT_2C of inst : label is "002F0F1A0F000F3FFE0000000000F00002FFF155F000F3FFE000500000000000";
    attribute INIT_2D of inst : label is "0000000F000F000F2FFE1A0000003FF0000200F100F000F3FFE080001800FF00";
    attribute INIT_2E of inst : label is "002E0FFF07FC0000E000FFC03F40000002EEFFFD7F0F01DD00004000E8000000";
    attribute INIT_2F of inst : label is "0000000F000700002EE0FF50F5F80000000300FF007F0000FF00FD400FE80000";
    attribute INIT_30 of inst : label is "00FF001F003D1A0A40008000000050001EFC03F900DD800200000000C0000000";
    attribute INIT_31 of inst : label is "000000000000001AFF401F803D0000A0000300000000057EF900DDC00000FD40";
    attribute INIT_32 of inst : label is "D01F015F00BE05C0F407F540BE000350381E007F00BE005CB42CFD00BE003500";
    attribute INIT_33 of inst : label is "00192D3F00B400A76400FC781E00DA0000190B7F14B400E76400FDE01E14DB00";
    attribute INIT_34 of inst : label is "0C19005A018900A5830050002400A000C09025A504910A5A3000000080000000";
    attribute INIT_35 of inst : label is "000C00080009000006035A502424A5A000CA00050024000A6530A58024905A00";
    attribute INIT_36 of inst : label is "058E0ABF050B0288EE58FDB03510F280858EEABF0543071CEE52FDA93604C340";
    attribute INIT_37 of inst : label is "058E0ABF050B0288EE58FDB03510F28001AE02BF00490000EE40FD401C00A000";
    attribute INIT_38 of inst : label is "0AAF000F000F0BE0AA0000000000B600AAFA00F000F09E0BA000000000006000";
    attribute INIT_39 of inst : label is "000A00000000000BAFAA0F000F00E0B600AA0000000000B6FAA0F000F00009E0";
    attribute INIT_3A of inst : label is "03DB007D02FB003DC000000000000000FF6F07D02FB03DBD0000000000000000";
    attribute INIT_3B of inst : label is "003E00000002000FFFBC7D00FB0040B800FF0007002F003D6F00D000B000BD00";
    attribute INIT_3C of inst : label is "03DA00BF3EAF0FFFA7C0FE2AFA94FFF003DA00BF1EAF0FFFA7C0FE00FAB4FFF0";
    attribute INIT_3D of inst : label is "03DAA8BF16AF0FFFA7C0FE00FABCFFF003DA00BF1EAF0FFFA7C0FE00FAB4FFF0";
    attribute INIT_3E of inst : label is "00AD003B00370215A400C000C00018001A7A24F118F224540000800040008000";
    attribute INIT_3F of inst : label is "00010000000000028F84CF30CF3051500012000000000005F240F000F0004580";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "FFFF02FCFFFF3F80FFFF60603C3C3C3C00000000FFFFFFFF0000000000000000";
    attribute INIT_01 of inst : label is "00000000000000000000000000004FDDFFFFB022FFFF6969FFFFB022FFFFB022";
    attribute INIT_02 of inst : label is "D99BD99BEAABC003FFFF03C0FFFF8888FFFF86480000000000000000FFFFB022";
    attribute INIT_03 of inst : label is "FFFFFFFF15543FFC0000000053141A90030003000300A76803005B9498261FF4";
    attribute INIT_04 of inst : label is "33CC33CCA2A2A2A25D5D5D5DEBEBEBEBFFFFFFFFA2A2A2A2D007C6935D5D5D5D";
    attribute INIT_05 of inst : label is "D007C693FFFFFFFFEAABEAABFFFFFFFF75C3BAEA99999999BFF906BF30CC3264";
    attribute INIT_06 of inst : label is "0000000000000000DB9FA4C924605B3624605B3624605B3624605B3600000000";
    attribute INIT_07 of inst : label is "FFFFFFFF8EE262862FF802C02FF802C00BE0ED7BD007FD3FFFFE30F0FFFE30F0";
    attribute INIT_08 of inst : label is "EAAB0AE0EAAB0BA01A4028901A402890F7DFBAEBDF7DEBAEBAEB71C7EBAEC71C";
    attribute INIT_09 of inst : label is "EE4428286EC428284EE4282846EE282844EE2828C46E2828E44E2828EC462828";
    attribute INIT_0A of inst : label is "BEBC0000AFAD0000EBE90000FAF80000BEBC0000AFAD0000EBE90000FAF80000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFAAAAFFFF0410FFFF1964FFFF73CDAAAAE6DB0410D9F7";
    attribute INIT_0E of inst : label is "0000000000000000000055500000FFF50000FFFF0000EABF5550D57FFFF5AAEA";
    attribute INIT_0F of inst : label is "0000000000000000000055500000FFF50000EABF0000807A555000E0FFF500C0";
    attribute INIT_10 of inst : label is "0000000000000000000055550000FBEF0000E69B00008C3255551924FBEF2608";
    attribute INIT_11 of inst : label is "0000000000000000000055550000FBEF0000E69B00008C3255551924FBEF2608";
    attribute INIT_12 of inst : label is "0000000000000000000055550000EEEE000099990000666655559999EEEE6666";
    attribute INIT_13 of inst : label is "0000000000000000000055550000FFFF0000BEBE0000696955559286FFFF2148";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF057C0FF8FFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFC1FB4FFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "03CF00FF005700BEC0008000C00000003FFC0FF8057C1FB40000000000000000";
    attribute INIT_21 of inst : label is "0007000000000001FFD0FF8057C0FBC4003F000F0005001FFC00F8007C00B400";
    attribute INIT_22 of inst : label is "0CCC218CBFAE0CCC33303248BAFE33300001AB5D001937570000AFD598055556";
    attribute INIT_23 of inst : label is "CB570A56005F202ED5E395A0F500B808060601D70D99303090004000B000200C";
    attribute INIT_24 of inst : label is "063F033F007E003CFE00F400B570F00083FF93FF07EB9F8BE00040005C00D800";
    attribute INIT_25 of inst : label is "00000000000000001BF53FF57EB710F00081009300070000BFE0FF40EB5C2C00";
    attribute INIT_26 of inst : label is "03CF00F8001F06F530006000400060003CE30F8601F46F560000000000000000";
    attribute INIT_27 of inst : label is "0003000000000006CB30F8601F40F560003C000F0001006FE3008600F4005640";
    attribute INIT_28 of inst : label is "0780000000010226F0002D00E400000064470002001E00C00000D00040000000";
    attribute INIT_29 of inst : label is "000700000000000055F0666D01E40C000064000000000001470002D01E409000";
    attribute INIT_2A of inst : label is "0003002600060C5FB000F600F400FD00003B024F006F31FF0000E0004000D000";
    attribute INIT_2B of inst : label is "000000000000003003B02D1E07B45FFD0000000200000C173B00FC607E40FFD0";
    attribute INIT_2C of inst : label is "0F7F0F000F0007F7FF0058000000F800F7FFF000F0007F7FF000000000008000";
    attribute INIT_2D of inst : label is "000F000F000F00077FFF00580000F7F800F700F000F0007FFFF0600000007F80";
    attribute INIT_2E of inst : label is "03FF0FFE017F001DFF00AA80F500D0003FFFFFE817FF00CCF800000050000000";
    attribute INIT_2F of inst : label is "0003000F00010000FFFDFE007AF51DD0003F00FF00170000FFF8E800FF500000";
    attribute INIT_30 of inst : label is "003F000D000001EF9000DC000000C0000FF401F003D030240000000000000000";
    attribute INIT_31 of inst : label is "00000000000000033F900DDC0000EF80000100030000000FF800D0000000F400";
    attribute INIT_32 of inst : label is "7EBF002600DB0078FEBD9800E7002D0007AF0026035B08B4FAD09800E5C01E20";
    attribute INIT_33 of inst : label is "02FF2C1F2B40027DFF80F43801E87D8000BF1C1F02B4007DFE00F4341E807D00";
    attribute INIT_34 of inst : label is "03000188010903801C00240004000C0030302481009130C0C00080000000C000";
    attribute INIT_35 of inst : label is "0003000900010003240C20242424024C003000240004003000C02090240000C0";
    attribute INIT_36 of inst : label is "1EBF02A700110865FD50F1A00400C9207A3F2827019C3861FD75F1A81C40CC2C";
    attribute INIT_37 of inst : label is "1EBF02A700110865FD50F1A00400C92003BF002700000066FD40F1800000CD00";
    attribute INIT_38 of inst : label is "000F000F000F0690000000000000790000F000F000F07906000000000000D000";
    attribute INIT_39 of inst : label is "00000000000000060F000F000F009079000000000000006DF000F000F0000790";
    attribute INIT_3A of inst : label is "03CF00FF03B000BEC000C000000000003FFC0FFC3B001FB40000000000000000";
    attribute INIT_3B of inst : label is "0007000000030001FFD0FFC0B000FBC4003F000F003B001FFC00FC000000B400";
    attribute INIT_3C of inst : label is "00E500C01FF50FFF5B00233F5000FFF000E5FCCA00000FFF5B00A33F0000FFF0";
    attribute INIT_3D of inst : label is "00E5FCC800050FFF5B0003005FF4FFF000E5FCCA00000FFF5B00A33F0000FFF0";
    attribute INIT_3E of inst : label is "000F00CF000F0FFF000030000000FD000278C0F001B47FFF000030000000F000";
    attribute INIT_3F of inst : label is "000000030000000B2D800F0C1E40FFFF00000000000000FFF000C000F000FFE0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFF0606FFFF0000C3C3FFFFFFFFFFFFFFFFFFFFFFFF00000000";
    attribute INIT_01 of inst : label is "B6DE0000A9FE00C0C3C32828B6DE0000B6DE00006969AAAA4901FFFFB6DE0000";
    attribute INIT_02 of inst : label is "26642664C003C00303C003C0FFFF0000B49980084921FFFFB6DE0000FFFFFFFF";
    attribute INIT_03 of inst : label is "FD00FFFD00000000030003005B94A46803000300A768632413101B90FFFFFFFF";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD5D7D5D5FFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0B9F600BFFFFFFFF";
    attribute INIT_06 of inst : label is "23A698973030FDFD9321238093212380FFFFFFFF93212380FFFFFFFF93212380";
    attribute INIT_07 of inst : label is "007F7FFFFFFFFFFFFFFFFFFF03E000C0DEB707D0FFFFFFFFFFFFFFFF3FF800C0";
    attribute INIT_08 of inst : label is "9006003C90063C00C1800098FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_09 of inst : label is "BE140000BC160000B41E0000943E000014BE000016BC00001EB400003E940000";
    attribute INIT_0A of inst : label is "AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000AAA80000";
    attribute INIT_0B of inst : label is "BC16AAAAB41EAAAA943EAAAA14BEAAAA16BCAAAA1EB4AAAA3E94AAAABE14AAAA";
    attribute INIT_0C of inst : label is "0000FFFF0003FFFF000FFFFF003FFFFF00FFFFFF03FFFFFF0FFFFFFF3FFFFFFF";
    attribute INIT_0D of inst : label is "000055550000FBEF0000E69B00008C3255551924FBEF2608E69B08408C320080";
    attribute INIT_0E of inst : label is "000055500000FFF50000FFFF0000EABF5550D57FFFF5AAEAFFFF00C0EABF0080";
    attribute INIT_0F of inst : label is "000055500000FFF50000EABF0000807A555000E0FFF500C0EABF00C0807A0080";
    attribute INIT_10 of inst : label is "000055550000FBEF0000E69B00008C3255551924FBEF2608E69B08408C320080";
    attribute INIT_11 of inst : label is "FFFFAAAAFFFF0410FFFF1964FFFF73CDAAAAE6DB0410D9F71964F7BF73CDFF7F";
    attribute INIT_12 of inst : label is "000055550000EEEE000099990000666655559999EEEE66669999999966666666";
    attribute INIT_13 of inst : label is "000055550000FFFF0000BEBE0000696955559286FFFF2148BEBE56C46969A888";
    attribute INIT_14 of inst : label is "FDFFFFFFF67FF577D79FDFD7F117F517D147F7DFF7DFFFFFFCFFFDFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFE7F7FFFFFFFD7FFFFFFFFFFFFFFE7FFF3FFF7FFD9FFDDFFCFFF7FFFF3FFFDF";
    attribute INIT_16 of inst : label is "FFE7FDFFCAAFF55FCAAFF55FF93FFF7FDFA7F55FDFF3D557F73FF557CF93F55F";
    attribute INIT_17 of inst : label is "DFE7FF7FFDBFFDFFFAABFFFFFF9FFFDFFDFFF9FFFEFFFDFFCFF3F55FDAA7F55F";
    attribute INIT_18 of inst : label is "CFF7F55FCAAFDFFFCAAFD557CFDBD57FCFF7F55FCAA7D55FCFF3DFF7CE63F55F";
    attribute INIT_19 of inst : label is "CFF3F55FC6F3DFF7C693DFF7CFFFD557CA7FDFF7FFF3F55FFF3FF557CAA3DFF7";
    attribute INIT_1A of inst : label is "CFF3F7DFCFF3FD7FCFF3F55FFCFFFDFFDAAFF55FCFF3DFF7CFF3F55FCFF3DFFF";
    attribute INIT_1B of inst : label is "F7DFBAEBDF7DEBAEFCFFD5FFDBFFFFDF00000000FF9FD557DB9FFDFFF69FDFF7";
    attribute INIT_1C of inst : label is "E54FFA9FFCBFFDFFE56FF55FFA8FF55FF95FFD5FF2AFF55FF56FF55FE2B7D557";
    attribute INIT_1D of inst : label is "E56FF57FC56FDFDFC66FDDDFFCFFFF5FF27FF7DFFFEFF69FFAFFF57FCABFDFDF";
    attribute INIT_1E of inst : label is "CECFF77FCFCFFDFFCFCFF57FF47FFF5FE57FD57FF95FF7FFE54FFFCBC56FCFFF";
    attribute INIT_1F of inst : label is "71C7F7DFC71CDF7D397CDAA7FF3FFF7F00000000D51FD55FCFCFFA9FDB9FDFDF";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000006BE00FF00140A8A714000000000AAA0";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFFFFF6060C3C3C3C3FFFFFFFFFFFFFFFFFFFFFFFF00000000";
    attribute INIT_01 of inst : label is "FFFFB0227FF500E0FFFFEBEBFFFFB022FFFFB022FFFF696900004FDDFFFFB022";
    attribute INIT_02 of inst : label is "26642664EAABC003FFFF03C0FFFF8888FFFF864800004FDDFFFFB022FFFFFFFF";
    attribute INIT_03 of inst : label is "D000FFD0000000000300030053141A90030003000300A76803005B94FFFFFFFF";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5D5D5D5DFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF906BFFFFFFFFF";
    attribute INIT_06 of inst : label is "65846E5430307C7C24605B3624605B36FFFFFFFF24605B36FFFFFFFF24605B36";
    attribute INIT_07 of inst : label is "000707FFFFFFFFFFFFFFFFFF2FF802C00BE0ED7BFFFFFFFFFFFFFFFFFFFE30F0";
    attribute INIT_08 of inst : label is "EAAB0AE0EAAB0BA01A402890FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_09 of inst : label is "EE4428286EC428284EE4282846EE282844EE2828C46E2828E44E2828EC462828";
    attribute INIT_0A of inst : label is "BEBC0000AFAD0000EBE90000FAF80000BEBC0000AFAD0000EBE90000FAF80000";
    attribute INIT_0B of inst : label is "3E9441411EB4414116BC414114BE4141943E4141B41E4141BC164141BE144141";
    attribute INIT_0C of inst : label is "FFFF0000FFFF0003FFFF000FFFFF003FFFFF00FFFFFF03FFFFFF0FFFFFFF3FFF";
    attribute INIT_0D of inst : label is "0000000000000000000055550000FBEF0000E69B00008C3255551924FBEF2608";
    attribute INIT_0E of inst : label is "0000000000000000000055500000FFF50000FFFF0000EABF5550D57FFFF5AAEA";
    attribute INIT_0F of inst : label is "0000000000000000000055500000FFF50000EABF0000807A555000E0FFF500C0";
    attribute INIT_10 of inst : label is "0000000000000000000055550000FBEF0000E69B00008C3255551924FBEF2608";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFFFFFFFFFFAAAAFFFF0410FFFF1964FFFF73CDAAAAE6DB0410D9F7";
    attribute INIT_12 of inst : label is "0000000000000000000055550000EEEE000099990000666655559999EEEE6666";
    attribute INIT_13 of inst : label is "0000000000000000000055550000FFFF0000BEBE0000696955559286FFFF2148";
    attribute INIT_14 of inst : label is "FFBFFFFFFEFFE767EBFBF9EBFFBFF513FBEFE28BFBEFFFFFFEFFFDFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFE7FFFFFFEBFFFFFF557FFFFFFBFFFFFF517FFFFF517FBFFFCFFFFEFFF3F";
    attribute INIT_16 of inst : label is "EAABFE7FFAAFCFF3EAABEFF3FFBFCA2BFAAFEFF3FAAFE55FFEBFFF3FFAAFC9F3";
    attribute INIT_17 of inst : label is "FAAFFF7FFFFFFF9FFFFFFAABFFFFFDBFFFFFFEFFFFFFFFFFFAAFF553FAAFCFF3";
    attribute INIT_18 of inst : label is "FAAFCF53EAABCFFFEAABCFFFEABFCFE7FAAFCFFBEAAFCFF3FAAFC553FAAFCD57";
    attribute INIT_19 of inst : label is "FAAFCFF3EFFBCF63EFFBCFF3EFFFCFFFEFEFCF6FFFFBCFF3FAABFF3FEFFBCFF3";
    attribute INIT_1A of inst : label is "EFFBCEB3EFFBDBE7EFFBCFF3AAABFCFFFAAFEFF3EAAFC54FFAAFCDB3EAAFC55F";
    attribute INIT_1B of inst : label is "BAEB71C7EBAEC71CEAFFFCFFFFFFFDBF00000000EAABF9FFBFFBFCFFEFFBF96F";
    attribute INIT_1C of inst : label is "FFFFDA8FFFAFFCFFFFFFC57FFFEFCFCFFFFFF3FFFBFFF3F3FFFFE54FFEAFF3FF";
    attribute INIT_1D of inst : label is "FFFFCFCFFFFFCFCFFFFFCCCFFEFFFCFFFBFFF1BFFFEFFFCFFEFFFCFFEFFFCFCF";
    attribute INIT_1E of inst : label is "FFFFCCCFFFFFF33FFFFFCFCFFEFFFCFFFFFFF56FFFFFF3FFFFFFDA8FFFFFCA9F";
    attribute INIT_1F of inst : label is "F7DFBAEBDF7DEBAEE55B36BCFFBFFF3F00000000FFFFF9FFFFFFDA8FFFFFF9BF";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000001F9002802660FCF400000004000DFF0";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
