-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "1800117FE0C19B4215612C583156C790D440D440000000000000000000000035";
    attribute INIT_01 of inst : label is "084F3A6E5B00148822A6360200B44454D44301B5501217E7B50A3BB44AF325D9";
    attribute INIT_02 of inst : label is "BDEAA50000000031FFAEA5AC46BE0EA5FFAD80054AA020E94A1081812C21600B";
    attribute INIT_03 of inst : label is "5A6A92825554E1A8A860A20255400000000000000000084A05050001E585FF9A";
    attribute INIT_04 of inst : label is "4541555154A212AA520885100552143013450201AA10544540E0C42500AAA103";
    attribute INIT_05 of inst : label is "FDFE00002EE36E7565C97DF0F81414141410419FE0419FF06A22C440A9014545";
    attribute INIT_06 of inst : label is "04FFE21A5B6C9280047A9EFE000015500864902268E232800005555555552FFF";
    attribute INIT_07 of inst : label is "8AAAA3426B52C82C26F845051441544446FE96AAA8AAAACC4C4C494889028000";
    attribute INIT_08 of inst : label is "DD553852926280A4290A4101523806080000000155544B848AEFEEAAAAA4EFEE";
    attribute INIT_09 of inst : label is "1E4739BFDFFC1C8FF65D9328F239CDFE0000227D214C49BA543894DD1140000C";
    attribute INIT_0A of inst : label is "019410016C43F531BD54C9508845020D48B2D55849584BE3BBCEE269B72AE4D5";
    attribute INIT_0B of inst : label is "BAB515BAA5102054272A451444434350B448104A95A8854552818DB6305E2050";
    attribute INIT_0C of inst : label is "EAFB2AE1B4D242140A0845294243667646DCD22E80A43667646DCCB888420905";
    attribute INIT_0D of inst : label is "65766AC9492B21242C8690480E002C70FC0450586DB54AAF5ACBEB9B003EFBED";
    attribute INIT_0E of inst : label is "23133236D34AC36A366469AEB0FA9CC6F4FBAD01007DD952D110141472923604";
    attribute INIT_0F of inst : label is "0000000000000000000000000681A2415A82D0CB423DA51E92D92FF644AD0DB2";
    attribute INIT_10 of inst : label is "95949F00000000000000000000000006F42EAC32D51728A084A1421292820480";
    attribute INIT_11 of inst : label is "AA807159BE9A69BEFA66666666AEE8D3BEA3767DDD493B0B3F55D50DA8CC2AB7";
    attribute INIT_12 of inst : label is "3788F457D65DE726977E42DBBF206CAA89110B655448881B77E42D2A02842A80";
    attribute INIT_13 of inst : label is "72A92ADA440168557C989A04F6C24008088080081011000000880155AEC8374F";
    attribute INIT_14 of inst : label is "63801770C516DD000BA0084202B92488DF74F36BA03C9891014B6BA829EFA129";
    attribute INIT_15 of inst : label is "5BFD82FA408817881834026E8440BF9AE9D65FA59B102F25662CF23C9F23C9FC";
    attribute INIT_16 of inst : label is "11A336120E8AA8B2255439558957AA91110AB7642D92AA2499035A802100E491";
    attribute INIT_17 of inst : label is "4854042C7A3B55500C2A245215010B1DE6BA7544446CDA3A3371FA5FAC97CDC5";
    attribute INIT_18 of inst : label is "70C074264C08E4D081CA10420500DAB3EB3EB3E8A12A214A0CFBE9E6DC572091";
    attribute INIT_19 of inst : label is "CE5B36F2DB9ED5556AD5AAFBABFCACF2CE0CE4CFB40F58956B89080824A458C0";
    attribute INIT_1A of inst : label is "6E8113DA7B349409111191D1F2816B528A23EE8102AA71CF2FB7795A9CE5B369";
    attribute INIT_1B of inst : label is "00000000000000000000000000000000005D3CD76B32D4B17DF7D8603F01BDDA";
    attribute INIT_1C of inst : label is "4D4D4D4D3F3F3F3F0C0C3C3C0C0C3C3C0D0D3D3D0C0C3C3C0D0D3C3C1B1B3F3F";
    attribute INIT_1D of inst : label is "3D3D3D3D2D2D2D2D1D1D1D1D0D0D0D0D3D3D3D3D2D2D2D2D3D3D3D3D4D4D4D4D";
    attribute INIT_1E of inst : label is "1D0D1D0D2D3D3D2D3F3D3F3F08083F3F4D4D4D4D3D3D1D1D4D4D4D4D2D2D3D3D";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "1071474C5E8DAF5595595145105485A8FAF55955951451054C5A8D92A54B9E04";
    attribute INIT_21 of inst : label is "9D65D65C51C41D3A3E0000000000000000000C404294A6B5A529622AF7597597";
    attribute INIT_22 of inst : label is "D8415F43626AEACAA6890AA1B7E1116111AA25145694A9655955951051454A8D";
    attribute INIT_23 of inst : label is "009126CF995954DE42634A48556DBB082BEA4A434C434ACA8AB4AAD4B242AA6F";
    attribute INIT_24 of inst : label is "2A88A40B8E74A92CB849249A8520531415451060215473B9C8A0B4101090404A";
    attribute INIT_25 of inst : label is "B3B504100A4C9142890B98C016F258AF4B2CA2C298632302F4BACB2C29863230";
    attribute INIT_26 of inst : label is "FEF95089240041486499D142851164398C318C63762D70C0C54775D7598E5460";
    attribute INIT_27 of inst : label is "598DA4E58F584F947AC9FA3D613F4799354794E4AC5E9A6DA77CFF9B0DECE830";
    attribute INIT_28 of inst : label is "C739738011111A68347FC689362FA100469069251F591B933A3591851F42F555";
    attribute INIT_29 of inst : label is "5C289B571C4F00543407D5065094B4C618C6D5A3CC2688DDDD127E5FF2B70B70";
    attribute INIT_2A of inst : label is "FDB6A00FBD6064F7C9837A99988FF6559228F2F839CDFE91ABF201205A012466";
    attribute INIT_2B of inst : label is "0A92208A5A580012AAAAAAAAAAAAAA5B102BD692B9F402EA2BE040400E240AFF";
    attribute INIT_2C of inst : label is "CC6BFA9E17EAFB219C42FAFB3537188FFFE7F55281E41C64257B2A2F52444218";
    attribute INIT_2D of inst : label is "EEBAF6745FBAEBD9D97EEBAF6745FBAEB9305A0E6233A6063187EFB21EE766BE";
    attribute INIT_2E of inst : label is "889719961098942581B6DA6BA431C31C3756575657544085AF6745FBAEBD9D97";
    attribute INIT_2F of inst : label is "939CCC000FFC013248EFCF9F91E44001010080510828000208822225E8888D88";
    attribute INIT_30 of inst : label is "A0140451200BE2A22204000044008020228054502A8A0002FE84ED2075952122";
    attribute INIT_31 of inst : label is "0911C065B751FD581F03EA49910570ACA1AC0F891BF4AAA8257C655752B0BAB0";
    attribute INIT_32 of inst : label is "2D31FA993402231A01950D022B27EE90BFBA427FE92F224C60A460B470A14296";
    attribute INIT_33 of inst : label is "FA6F2B0EB4DF2B0EB4FF2B3AD37E82EEDD24F800020824A1A544949684051A35";
    attribute INIT_34 of inst : label is "4EFE8EB09FA2AC9FFD9564EC547AD5445113EBFAA14739332ED7F45B71107289";
    attribute INIT_35 of inst : label is "F593F5273C3E0CFFB0BECBFB2BFFA887B9421EE5085F96FF333FFF67584FD956";
    attribute INIT_36 of inst : label is "7E02A96ADB495F659CC9D65115F8EDF72E3FCCBBCE64EB18C487B6CB6A42A7D1";
    attribute INIT_37 of inst : label is "9E4D88511412221C0A004B8F9569B3F46FB77019D3B7F2B0E8DF2B0E8FF2B3A3";
    attribute INIT_38 of inst : label is "6A8EAF15944A680A1A792CAAA8290931557A1090249CA8A20C14575A85108026";
    attribute INIT_39 of inst : label is "F73672324EC6CC447C6E99D9A2BB3315DCC8C2CC0B3D9C09D9500C651407D50A";
    attribute INIT_3A of inst : label is "0BF0056C3B618EDD178465AF2F27793BC9416AA621A1825B52802408481297A4";
    attribute INIT_3B of inst : label is "04ACBE8081164508140B2131ADD34D14B518BAD694A6FA8D4950AB894F49D58A";
    attribute INIT_3C of inst : label is "12242097BD40F5FFFB6D4019BC84BD195AF788AA4280814244A8ADB4210842F0";
    attribute INIT_3D of inst : label is "618C61564FD448079271A482A0DA9FF581506E516838890CFF1FE00980480240";
    attribute INIT_3E of inst : label is "800E002AAAB9EE23D1D77D2D00A4C9FFF8A12243B8CF710CAD0D24E7121B48CC";
    attribute INIT_3F of inst : label is "000000000000000000000000000000000000000000000000000000000000757B";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "81B58280095438B587E8152A833A8D028CA58C80000000000000000000000013";
    attribute INIT_01 of inst : label is "7520DFB3C2C0064D6698E95942722CD30DCED67137252FC2062CF549AD047397";
    attribute INIT_02 of inst : label is "20745300000000B2001853F1CBC8505300F01AC8ED3DD620A63D92BA9DF4EFA7";
    attribute INIT_03 of inst : label is "7B2CD9AB7D37FCBBBBFA795B55500000000000000000012D01970002F8130077";
    attribute INIT_04 of inst : label is "DCCD9D9E66DB594CDED3365ACE66F3CAD95C9ECCBB6B3223266E48B7525AE729";
    attribute INIT_05 of inst : label is "FFFE00016C637EA9E5337CAAA3500550B420419FE0419FFE6611976B26565CCD";
    attribute INIT_06 of inst : label is "247FE2937BEC920024CC299600009AAEEA65D212E8EB1680040398E663986FFF";
    attribute INIT_07 of inst : label is "8BAAB24AE6D7F57FB6B951514511555446FEB4CCCD9AB244CC44C95203018000";
    attribute INIT_08 of inst : label is "888841DE66F4F6529CE52DADC9E224A0000000059998CA3D98FFEF6FFEF4FFEF";
    attribute INIT_09 of inst : label is "E4880B40007149D550A6006F24405A0000004440E7799BC1CBE05C119DD5D5D9";
    attribute INIT_0A of inst : label is "DFAA7F96FAAD57DED0F3066894B89EDB6734029A029A001C2FFEBDF25055003D";
    attribute INIT_0B of inst : label is "9E6DC3BE6DA2D26AB166DC724A8E6F5B6CD928D9B76D1679C05A5468EB7AEB6F";
    attribute INIT_0C of inst : label is "410241284B27FECCED64DCBCFE10830010110B6859810830010111A3996D2C97";
    attribute INIT_0D of inst : label is "80CDB1322646CCD99B3164A81604B6D86A0C600002012B02A5505E29B7010010";
    attribute INIT_0E of inst : label is "3C51A4030C33431BC348061865D5971E83041BAD55F30DD684996412CF324F28";
    attribute INIT_0F of inst : label is "000000000000000000000000079C07928CF31AE3CBC9E1E4646644F2CD9F6C72";
    attribute INIT_10 of inst : label is "392EA4000000000000000000000000022AD57AB49AAA5AFEDE7DEB7B4B6B56DE";
    attribute INIT_11 of inst : label is "31129B8030C30A38C39898989D313F74C1D0808FC718FD5040663E42591563CB";
    attribute INIT_12 of inst : label is "D877198B6D92C86F4C90BDE6485EF213106AFF90988357FCC90BDEBFFD6F8CFB";
    attribute INIT_13 of inst : label is "88F0DFFC5EF6DF1A82043DEB3F77FC8888888881089888899889986A315F4596";
    attribute INIT_14 of inst : label is "94B5B9995F79E6D2ACB7B5F8DF440371E0596D8D5DC2043E6FAF8D469A2035B6";
    attribute INIT_15 of inst : label is "BC52F7F9BC7FF5F5F65FDDF17BB9436CB26CFFB63CEE5080D1D437CDE378DF32";
    attribute INIT_16 of inst : label is "EECD7ABFE33133274FAB73E11FFC352E2AAC4CCBDE404C41F2F7ADFF5FE0203E";
    attribute INIT_17 of inst : label is "BFDA96558CD786A255F0796FF6A595E6DB2C99B9BBB7EFECDF9E6CFFC93FD0EA";
    attribute INIT_18 of inst : label is "BB6B9BF481B58DEBF81D6DFD7A6FA06C925B6C9535B4B5EDE91FFBE020BAEE65";
    attribute INIT_19 of inst : label is "0C0924659438198CF333CC047419C92573F30DC0B8FDB57ADD3BB2FACB4FAD6B";
    attribute INIT_1A of inst : label is "2FFFEB9D40A05ADFFEBEBEBE4D5F94EFF7FC411AD5359732445592BC0C252129";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000165B6CAE5FBFEA82152AD5C2AEA050";
    attribute INIT_1C of inst : label is "4C464C464C444E461B112B213B310A000A003A303B310A003A300B012C243A32";
    attribute INIT_1D of inst : label is "282228222822282238323832383238301C161C161C161C160C060C064C464C46";
    attribute INIT_1E of inst : label is "26360616360626360C3806303B3102027C765C566C666C666C667C765C564C46";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "A28A68D6A352304E38E38A68A68D6A350304E38E38A68A68D2A3500090FD08DE";
    attribute INIT_21 of inst : label is "778E78E69A69A74D4000000000000000000000FDB67959DA4ED38C5304E38E38";
    attribute INIT_22 of inst : label is "27FAD094B496942CCEF85DDF001FFF6EEE6FDDE9E9AB5EDEE3AE3AA2AA2AD552";
    attribute INIT_23 of inst : label is "7BA34110468599D195B4B6C2EEF804FF5A3FD494B694B6B46CC9B3E9BE1776C0";
    attribute INIT_24 of inst : label is "41529587DF79248222C30C30F2B7844FDA9A7E9FDCE8940A1BCBD9A5A5369693";
    attribute INIT_25 of inst : label is "4A5A4BD01A5CC3FECEDEF3B00404E144BCF3DB3526A4D4F44BC73DB3526A4D4F";
    attribute INIT_26 of inst : label is "4206F231E608434C348363B7FD9C0FEF3BDEF7BD89F7E7BFFEE8C30C22CBAB5D";
    attribute INIT_27 of inst : label is "06F7D9CEB2D2833996906CCB4A0D9952030B383B52012D970094028250577258";
    attribute INIT_28 of inst : label is "4A53A5252666600500868F1A0897683EA96586726D92203708D2A5206ED00F0F";
    attribute INIT_29 of inst : label is "15A4411C71C1B61B025C0DDD3B12877B6F7BD2E415085522226CECE6C7245245";
    attribute INIT_2A of inst : label is "104156B1038A0C002EF8F76C2DD550AE016F24BDC05A006652AB6ED6A56A4A80";
    attribute INIT_2B of inst : label is "1930725FF6FF795A000000000000004033C5B53EE0762BEC6FF7D7F79E6C9B80";
    attribute INIT_2C of inst : label is "960D51A6D821525824DB01525E4479BE00440B2E5CDD3B99C815D5412608C949";
    attribute INIT_2D of inst : label is "1060298A806182A6A241060298880618426723AC7C7C4DBBDECD15258109C0D4";
    attribute INIT_2E of inst : label is "A0A6F7ACB7C34A5AB810418411455045444455455447C18E02988806182A6AA4";
    attribute INIT_2F of inst : label is "8301460AAAA99756D577D5A8B79A0009B0B2D10B24B4C28859A28281AA0A0BA0";
    attribute INIT_30 of inst : label is "DBEDF2AB97DFEAFD4F7ADEDEFADE5F6F955CEAEB9D5B797A64DF30456127F3FC";
    attribute INIT_31 of inst : label is "D5AB2F08266EF6ADACB59DB52ADECBDBDE53D672A4CE5576FBFD4FA9EF5BDF5B";
    attribute INIT_32 of inst : label is "8BAFB5227EF5D4BF7A6E5FF4D598012D4444BD8012D6FF3ACD5BDD4ACD4DFF7D";
    attribute INIT_33 of inst : label is "05167257FD267257FD06725FF409E917ABF5200001D76BDECFEEFFFFFB8F3E7C";
    attribute INIT_34 of inst : label is "811B312506CD490036E2480199873A08E235B1DCE5CA4370101C20804222E71A";
    attribute INIT_35 of inst : label is "49204ED5954AA5804747141CD0005F3846BDE80A738069004C400D9A92836624";
    attribute INIT_36 of inst : label is "09E95F97A07CAA4FA01FEEEA8A850B1061D4A9DFD00FF16B5B7A79E7D7FD4B6E";
    attribute INIT_37 of inst : label is "0C904C2A0A7C401D0500F305A0D20CD9BA5CABD22003672575267257506725D4";
    attribute INIT_38 of inst : label is "09D958A21E14B5F738E38C4C5DE7337EABFBFBFEF9F6D394FBA9E845FD99D2F4";
    attribute INIT_39 of inst : label is "0989998C31111110FFFFC22B750CD7A8295610154052BD4000001C46D185E1D2";
    attribute INIT_3A of inst : label is "365FDA97A4BD6927EA7A8AD2F2F497A4BD9F85594A4AD5A4BF7B7EDEBDFF6C3E";
    attribute INIT_3B of inst : label is "F7C7C75E809D0FFC9AADDBDED025B32BFAF767A93D4865D2322DD5DAF87C6FF3";
    attribute INIT_3C of inst : label is "72022B4000DF9A080000AD76EBFF62AEE0003B15B76BFAFF667672069CA72986";
    attribute INIT_3D of inst : label is "DEF7B28890AEBD7375EE3E5775216C0A6BBA81A48EB0F187D5DAA55DA9CD4F6A";
    attribute INIT_3E of inst : label is "EEEC0043D2C0EA4A0D79400D01A5CC0801FFB3B66D34DA535252DF4DA4A4F739";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000002400006509";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "D00C407FCA9D0A53C00C0113A510D4C085210440000000000000000000000021";
    attribute INIT_01 of inst : label is "6148A30AD24000290AAA284040310155444210A5010100000708002421BA94E5";
    attribute INIT_02 of inst : label is "C8A4110000000015FF0C115001441C110A5004C040C9A6A0221AA0B0A5852D29";
    attribute INIT_03 of inst : label is "4282120888410620AA833C5A0008000000000000000002090121000079010280";
    attribute INIT_04 of inst : label is "55540036540654C015B2A032B200A8E2C0060422228818110307152415308ADC";
    attribute INIT_05 of inst : label is "A855E00060477EF5F4033DD4D015544030107F9FE07F9FF0CA2AA1CBCB178445";
    attribute INIT_06 of inst : label is "2401E09B7FFEDA002400940800009FF0025DD826EEEE26000C041FF87FE06552";
    attribute INIT_07 of inst : label is "E6FE6C8A2BB7CAFF6FF14FBFFFEBFFFFF6FF30F0F27AA24444CCC8C445408000";
    attribute INIT_08 of inst : label is "9919009427E410108C63086050FA202000000005E1E0C2D59A2AA2E6FE666FE6";
    attribute INIT_09 of inst : label is "B6CD1B6FC00868DAB0B500A5B668DB7E000044014A129F905078109959919111";
    attribute INIT_0A of inst : label is "404A028514238539FF55794925252A15000400020007000ABFE8FA1FF15AA044";
    attribute INIT_0B of inst : label is "AA15150A0570950A8A28571493C14A12440A0C08142B85444E177E9A28502848";
    attribute INIT_0C of inst : label is "C6AB66AA08414A95210065244BD43F03D015428A149D43F03D01572C82490921";
    attribute INIT_0D of inst : label is "B638738A614C298530A6152FF7FDB61879F98FE48C314A23C998DED6754E3CF1";
    attribute INIT_0E of inst : label is "D2A56D461C72DF752ADA8C38E0FB5CBAC71E3361333C7BF5DBB72C9D2EEE4473";
    attribute INIT_0F of inst : label is "00000000000000000000000005B80A549CE5547AD52D6A9614C14C9246A94DCF";
    attribute INIT_10 of inst : label is "AFF0B10000000000000000000000000091821D22D4410A90942952C250505030";
    attribute INIT_11 of inst : label is "BFB7D2C11C71C50C10C5544557BFAA16288430DF0E18F7F82A731BD0A98B4365";
    attribute INIT_12 of inst : label is "6D879DEDB6FB6D7E066240F3312078D9B9410BC6CDCA081E66242F4148440641";
    attribute INIT_13 of inst : label is "32D95A1FB39C881DCC94A90A17AD20000000019899899888888998773B887EFB";
    attribute INIT_14 of inst : label is "C7462F33D146F8ACA218C6418A992544F3EFB6CEEA8C94B8C55BCEED6B73E464";
    attribute INIT_15 of inst : label is "DF9B17FB28AF5F2F58F0AB7C4153EDB7DF77BF839E54FB25147CED5956759C48";
    attribute INIT_16 of inst : label is "54EF3F7903BD99F7EEF29BB39D40BB90354EE6A44F1366E5511BE6731D00C4BA";
    attribute INIT_17 of inst : label is "2942A096EEFBC7F6FE58A50A50A8253D6DF7DCCDD53EFCAEFBD3B6FF7FBFFB9B";
    attribute INIT_18 of inst : label is "FA4AD237C5612FC0409B18210F18B03EFBFDF7D984040C210DB7EBF2213EEE14";
    attribute INIT_19 of inst : label is "F15EDE36F6BC5E03FC0FF0269FAD6DB59A59AFC7AD86D84F69ABA58A9214294B";
    attribute INIT_1A of inst : label is "C2D7B5FE9B4DA1853B5F1F4FEAF5FF18D87EF3B4A7B8E9DB6761DB5EA3F05E83";
    attribute INIT_1B of inst : label is "00000000000000000000000000000000003BEDB6D36B5AD7DF61F0A56D2B0D86";
    attribute INIT_1C of inst : label is "3C363C360C040E062A200A000A000B013A300A000A000B010A000A000C040A02";
    attribute INIT_1D of inst : label is "1C161C161C161C160C060C060C060C044C464C464C464C464C464C467C767C76";
    attribute INIT_1E of inst : label is "46466666464646460C0C0600080202026C666C664C464C465C564C464C464C46";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "73D77D5A8858AA832C32C73C73C5A8A5A8A932D32D77D77D5A8858E425209630";
    attribute INIT_21 of inst : label is "A4CB4DB5CF5DF5696A00000000000000000001520208424282916690A932D32D";
    attribute INIT_22 of inst : label is "8ABAAEA4042527AA850F5771A2ABAE92029242480A482D4932D36D73D73D5A58";
    attribute INIT_23 of inst : label is "C6BD6851C0F550AEA505057ABBAD115D55D4A42420850507AA90AA4843D5DC6A";
    attribute INIT_24 of inst : label is "624AA50BD73828B41B0410411CE403620CF3D070AA3DCAA5767E6F777FCDDDFE";
    attribute INIT_25 of inst : label is "5762121FF961E54A2009CA7000E3D264C7DC7DCE79CF17164E75E7DEE7DCF979";
    attribute INIT_26 of inst : label is "4F1ED04A2FF6FF2B7DB045029445AC1CA739CE73B8327080C7438718715DC8EC";
    attribute INIT_27 of inst : label is "01CF256B5B9BD5AEDCF8B76E6F56EDDF178DAC628A4A01052A39570F78ECEA58";
    attribute INIT_28 of inst : label is "CF5BF5A53FBFB223105395AB42A848615195595BB6DF32BF18256C2050900FF0";
    attribute INIT_29 of inst : label is "A73B1B33CCD51DF75D8B21E39C4ED8E71CE7D8C4090E2A737312B6B7E5F67F67";
    attribute INIT_2A of inst : label is "E1C60437805A0C7001530A95A8DAB0B500A5B6FB68DB7E352D50936136136E22";
    attribute INIT_2B of inst : label is "AA3114B4A529CEC7FFFFDFFFFFFFFF1B9066E73E00A198432105050D041428B8";
    attribute INIT_2C of inst : label is "DA32AE8EA566AB6AADD4AEAB6C51DBA4E399C1CD98D99B05295E676B461652E2";
    attribute INIT_2D of inst : label is "78C2BCCCD5E30AF3B3570C23CECC5C30CD950E1FFB5132E739C7CAB68EAA4B2A";
    attribute INIT_2E of inst : label is "FF5FDB932ED0421D6830C30C395C30D71F7F6E6E7E7F7F3223CEEC5C308F3331";
    attribute INIT_2F of inst : label is "0203AA66799831A49C486ABDD52E8001208C508B0B14A394589D57FD955FF7D5";
    attribute INIT_30 of inst : label is "1284A021A42FEE20A28290948290342501045061AA0850D0B6B1492304B0A086";
    attribute INIT_31 of inst : label is "25454A16F3B01B0141282C23F0100202D6108414B18A043085FDC41550420042";
    attribute INIT_32 of inst : label is "1D74DA3324AD2D1252120925240D44A1315284C44A1429804240525142420844";
    attribute INIT_33 of inst : label is "173B5F78458B5F7845AB5FE1162F0DDAB4A5A8CD3492D20A0D74D24051020205";
    attribute INIT_34 of inst : label is "D44DD9B78B766FAA9B337C47765B951CB3DEDC772253EBF14AB4726AB73DBDCB";
    attribute INIT_35 of inst : label is "6DF558A533399002FD1DF5775102AEEE188AB8722EE5CAFFBB3FC6ECDBC5BBB7";
    attribute INIT_36 of inst : label is "2F8DE55EB520956DF45FBCBC8D54AEF145AAEDBEFA2FDBE1FAAAEDA6939EC1BB";
    attribute INIT_37 of inst : label is "F14A9C65191220064CA04851D66ED26EF378F29FB152B5F7E58B5F7C5AB5FF96";
    attribute INIT_38 of inst : label is "12E8A9415690A45202082822A04213F093F850A189FE02A4291555169442A586";
    attribute INIT_39 of inst : label is "1110000002220000FD7E8512540A24A012B6100940256340000004314003545D";
    attribute INIT_3A of inst : label is "422A109AA8D50A150950869151550AA854818A50528212921AC615AD6B0A45B4";
    attribute INIT_3B of inst : label is "A6AAD854FBA5952D42A10139C9402148420E294A0840A0CE4A40A4348B684ED0";
    attribute INIT_3C of inst : label is "F7BF9DEC32509271E30C084EA546259C63876A290292024B1111142CC77B9EB2";
    attribute INIT_3D of inst : label is "39CE749877073663666C14258789197292C3C720283DED6EB376733F67FB3ED9";
    attribute INIT_3E of inst : label is "145C0056A8430042191D8B15FF961E71E2A58802A15142159490830421213145";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000004041";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "80258A5420850F5B80C00810A114C58084350680000000000000000000000021";
    attribute INIT_01 of inst : label is "202A82A1D0801021021A004A56256043440C92C620203123AF22122504B602C0";
    attribute INIT_02 of inst : label is "6010110000000042500A119CCE7044110B9D1644524882A0221A1B1410A08504";
    attribute INIT_03 of inst : label is "434251691A012D22CC96FAEB089810000000000000000C0104C100012D118282";
    attribute INIT_04 of inst : label is "4445D1C7568958E8143AB44AC740A5C25A85C82523031712729684A2D234021A";
    attribute INIT_05 of inst : label is "CA32A0AAE9CA77EFC6977D454504450074601E1FE01E1FF50BAB19495212A664";
    attribute INIT_06 of inst : label is "2C3CE3BFFAC813C02C322B030000BAAEEEE1F63BE07BBED55C021FFF8000ECCC";
    attribute INIT_07 of inst : label is "09AA92AAA28FF55FFB2551504130411045807700FFFA954444444D5001114000";
    attribute INIT_08 of inst : label is "88082094B31D877BD6B5AF0F8FC225A000000005FE00AA3BBADFED4DFED09AA9";
    attribute INIT_09 of inst : label is "92C79868108F77DAB23D814C963CC3400000C8914A50CC628D41098008880088";
    attribute INIT_0A of inst : label is "4CA97A559E27C539FDC37F4804345C4C2C600630223002119BF86D59331EE069";
    attribute INIT_0B of inst : label is "F079D59069F295403BCF1F22034F030070D304D1A747913C5E1F7EFA1158114D";
    attribute INIT_0C of inst : label is "CE796C500A0102952949618503E03E03E005438A1E3E03E03E00572E00010801";
    attribute INIT_0D of inst : label is "AD627B0B616E2FC5F8BE142802002040340FC0706EB223A34888EBC6361F79F5";
    attribute INIT_0E of inst : label is "75182F365D6232FB505E6EB2E05BD55EB77CBAAD0FD154D8E58D87247FF9B73E";
    attribute INIT_0F of inst : label is "00000000000000000000000007D52250DCD3692BE355F1AA96C96CD30C3C6BF2";
    attribute INIT_10 of inst : label is "CC973100000000000000000000000004B4368DA2515B2C56D2059B5A095B4656";
    attribute INIT_11 of inst : label is "88BACED70C30410430DCDDCDC9889326B930247D884CB61A9F115B00A8800564";
    attribute INIT_12 of inst : label is "ACB1C446BACB2F30D76B5A3BB5AC1E88CD1D60F4466CEB0776B5A30D2959A258";
    attribute INIT_13 of inst : label is "9BDD09068AD6934466D7A96801B5AC0404404010110100EE88CD991188931359";
    attribute INIT_14 of inst : label is "9425AC4DC61836B68D56B59A6CCDBD0039359AE22AE6D7A03668E22593F2B1B1";
    attribute INIT_15 of inst : label is "460A10FC06802C002666241B5D5964D66B1A1FB5475659B6185BAC0902609820";
    attribute INIT_16 of inst : label is "56220DA56888AA9264D2C934889A88D715623735A3DA233F0560C35AD66017E0";
    attribute INIT_17 of inst : label is "205026192228D117595A2508140986C9359AC554558A34A228EC935F64D7D96B";
    attribute INIT_18 of inst : label is "CDC8F2D2E7CF661D5CCE9E2CAB8B3C965975D75AC1D4D6B575E3FC129FBE8294";
    attribute INIT_19 of inst : label is "555FFED777975FE0000000B356A465998E58E625CCB2C9CB2C9418B2E8E1DFED";
    attribute INIT_1A of inst : label is "657B3D7F89C4EAF7B3D787C7AEF97DCF9E4F389EF58CB0DDEBF86F86AAA00001";
    attribute INIT_1B of inst : label is "00000000000000000000000000000000004D66B2E17CA729FF38FED4672384C2";
    attribute INIT_1C of inst : label is "0E040E040C040E060C060C060C060C060C060C060C060C060C060C060C040E06";
    attribute INIT_1D of inst : label is "0E040E040E040E040E040E040E040E060E040E040E040E040E040E040E040E04";
    attribute INIT_1E of inst : label is "0404040404040404080A02020E0406060E040E040E040E040E040E040E040E04";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "B0D34D9B085AA61B0D34DB4D34D9B0A58A60B0C34CB4C34C9B0A5880252D9656";
    attribute INIT_21 of inst : label is "86C34C36D34C3669620000000000000000000C534A4A58524292E21861B0D30D";
    attribute INIT_22 of inst : label is "AE622289898504A245036C64223D989ADA535A29696BAD60B0C30CB0C30C985A";
    attribute INIT_23 of inst : label is "5B326075149448A28981A59A630115CC445094893121A524A240894948D19808";
    attribute INIT_24 of inst : label is "6A6A31AC59C5456C7600000056958EDAD5514746AC2C6181D2736D39B1A4C6D9";
    attribute INIT_25 of inst : label is "49524210368F3102AD2D6F5012ABB04E9698719630C61616EB61A71B634C6969";
    attribute INIT_26 of inst : label is "3C7A0284360B46C1C651914A055B68D6F539CE73F0281808C88F555555C50B2A";
    attribute INIT_27 of inst : label is "C9CE85234988F48E4C5E97262392E4CB9084CE5AEB6A4125BAAA4549989B9882";
    attribute INIT_28 of inst : label is "DD29108E1DD99B3D9639E1D30360942D5C9E09C992CB1B989B8D1C018128FCCC";
    attribute INIT_29 of inst : label is "A3DF4B37DCFE1D767D8FB171DFBC60E71CE72FD26080ABDD9983D33529DA9929";
    attribute INIT_2A of inst : label is "E5D6043FA220240421798E14D5DAB23D814C96433CC340F5E55969729729682A";
    attribute INIT_2B of inst : label is "B39136B94AFDADDD5555755555555509A2226398F4C5BB8B4E41E9E15C70AAFD";
    attribute INIT_2C of inst : label is "58B8AD0CE3F4A97AA89E7EA96E55E13DF793E18D180CC1052D5B222A72169A62";
    attribute INIT_2D of inst : label is "FAEAB46457CB2AD1115F2EA344447EB2C8D90C37B26B9AC739E7CA978CEBA38A";
    attribute INIT_2E of inst : label is "AAA3A15F3508421C10B2EB2EB079E78A2E9E9E9E8E8E81F9AB46457CB2AD1915";
    attribute INIT_2F of inst : label is "0580DA01E87C178000404A3DA338000C00AC4A88AB122255618802AA8AA00080";
    attribute INIT_30 of inst : label is "58D695359083E68624405266005246B4A9A51D7583AA9A1892D6592D45B410B6";
    attribute INIT_31 of inst : label is "843103539916896D68AD3CAC963612C1CE52B456B5C8A6B6107CC0C4881A501A";
    attribute INIT_32 of inst : label is "A49249112101819004C0C80880A556A1B15A86556A142D94985D984C98482948";
    attribute INIT_33 of inst : label is "5459199949A919994989196526251D883019AB32CABA48EB4556895B4D282058";
    attribute INIT_34 of inst : label is "F5658891E96225C8CB112E44DCCF2647B1465836C5997989AE19543871149193";
    attribute INIT_35 of inst : label is "2CB954B9B3066042B454D0534182ADA054B680425A21495066EA12C448E4B112";
    attribute INIT_36 of inst : label is "255DA088312D0526BE4DB534D052E633040A64DB5F26DBDE05A2A0824D2B4CB1";
    attribute INIT_37 of inst : label is "0ADC0C130450701642304292F120872E516A40CB1D149199A5A9199858919616";
    attribute INIT_38 of inst : label is "2E43AD5CFA20A6014B2CB9F7EC421987917B50A42CCCF61D80969D1A055C3ABA";
    attribute INIT_39 of inst : label is "C74D65AAB8E98C9400AE5C901831A0C1848A80C0238D03000000010000500000";
    attribute INIT_3A of inst : label is "6BA894EA075271F54D44C29D4D40EA475095FA5246923BFBFD7BDED7BDAF6B82";
    attribute INIT_3B of inst : label is "107DFC6285DFC40D500D2539FD48250A62EEA1C90C4EEAEFCB52A75EF7054C82";
    attribute INIT_3C of inst : label is "C6EEEA79B20AD3FBCB2C086EB516B0DD7B3641E94A06030357D7D3BEF7FDED73";
    attribute INIT_3D of inst : label is "A9CE70DD7F873660320402A1A1A9707254D4C72430DFC8388FF1E0F32F1978CB";
    attribute INIT_3E of inst : label is "BAEC0064CC99283AB2F32F050368F3FBC881AB4AA07144871224D3144C4C3937";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000600004293";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "C1A59A954A95249495C90112A2A00810AAB56AC000000000000000000000000A";
    attribute INIT_01 of inst : label is "60289488980002ED44B0C3DB56C76896198CF62960202A21170400480D0482A1";
    attribute INIT_02 of inst : label is "C0975A000000001355D55A5C0566135A4B58804E9008AA82B4389AB015A0AC05";
    attribute INIT_03 of inst : label is "004EC24B1A472D031186BAE80A095000000000000000016D019200006D8A52AA";
    attribute INIT_04 of inst : label is "888D1106768058C81C33B402D640E5D75099D8ED0003677676969D8496B48E5A";
    attribute INIT_05 of inst : label is "0B0E6A66EB0C34A992577D35351050007410EFDFE0EFDFF50DBB131D061A0888";
    attribute INIT_06 of inst : label is "2C1C61B36C9249402CDC98650000B00AA6D871C3861A4EB33C53E0000000EC3F";
    attribute INIT_07 of inst : label is "4DFED6AA222AC78C6B656101041044455DD57400FFFA95444444456465414000";
    attribute INIT_08 of inst : label is "08880B8CF7100694A5295C0C5872B6A000000005FFFEAA8FBA9AA929AA96DFED";
    attribute INIT_09 of inst : label is "96CD906D4A0BEADAB01108BCB66C836A00000005CE71DC405870008080000080";
    attribute INIT_0A of inst : label is "5A485212082C065AC016106915A1C2C562C4006221622142B028CA097108A257";
    attribute INIT_0B of inst : label is "4255864255A2D773302C58568A88B4AD44AB24A9562D1769845A5000D360D36B";
    attribute INIT_0C of inst : label is "606B6063092524D9AD6D85B42406202202154B4A588042002021542891B52DB6";
    attribute INIT_0D of inst : label is "6DE0B0D20A4148690521A4A8120430002806B060030D6B0ED99A81403048A298";
    attribute INIT_0E of inst : label is "6318BE80820AEBF2317D010C115C94C48193052DFF5FC98AF151943662D3C606";
    attribute INIT_0F of inst : label is "00000000000000000000000006CA849282AAF1C36231B118241243044AB56FCA";
    attribute INIT_10 of inst : label is "8D92B5000000000000000000000000014638C5E921DC3117D3275F5E0C5FE716";
    attribute INIT_11 of inst : label is "99FEFAC49269A492493766677599E997BCB620FCCADC86191E37DF1891E12771";
    attribute INIT_12 of inst : label is "2DE18ECDB6DB6F70C8D29EB4694E5A19DC9A72D0CEE0D3968D29EB918C658659";
    attribute INIT_13 of inst : label is "C8FC01D7A318CB0CD242516035E72C4400044052516142EE88CDDC3319CB365B";
    attribute INIT_14 of inst : label is "F677AEED824CBCBACF1CE759ECE49206B465B2C66ED24240F672C675CBEAE9E1";
    attribute INIT_15 of inst : label is "973BD007061B2B1B2B62675E59D97196CB360033D6765C930C5A48100401006E";
    attribute INIT_16 of inst : label is "32672E3961D999BA74F2D931988C99A637666889CB487772027AE46399609240";
    attribute INIT_17 of inst : label is "A49B3654667AC33FDD58496926CD951E65B2CCCCCC9CB84672D1B2806CA01B8B";
    attribute INIT_18 of inst : label is "E19CE2F6F74F6E1E5CDFFF2DAB8BB837DF6DB6D9C9C4C6316DF01C32372CA225";
    attribute INIT_19 of inst : label is "555FFE36E7B640000000002716AE6DB59E59EE253CB6D98B6D993CB860E5B38C";
    attribute INIT_1A of inst : label is "F47238E73F9FC8E62383C3C36EFC5BAC1C467198C59E73FB6778DBD6AAA00001";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000196CBFE7FDEF7AE379BCEE6F33DFEF";
    attribute INIT_1C of inst : label is "0C060C0608000C044A404A404A404A404A404A404A404A404A404A400C040800";
    attribute INIT_1D of inst : label is "0C060C060C060C060C060C060C060C040C060C060C060C060C060C060C060C06";
    attribute INIT_1E of inst : label is "4646464646464646080C00060A00000008020802080208020802080208020802";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "B8DB2D580858860BCCB2CBCCB2C580858A61BCDB2DB8DB2D580A5886492C04D6";
    attribute INIT_21 of inst : label is "86F36C36F36C356962000000000000000000008B242A49424A92265061BCDB6D";
    attribute INIT_22 of inst : label is "886820909495142EC92A85850220B09242504A4909491C80BCCB2CB8CB0C5858";
    attribute INIT_23 of inst : label is "5AB16C450285D920909C95542C0811050414A490929C95142EC93B0942A36040";
    attribute INIT_24 of inst : label is "6356B5AD14A52C002A10010090858552DDD15686EC2CC194C36B6DB5B586F6DA";
    attribute INIT_25 of inst : label is "4C524AD03CCF0224EC90C210081489609719699732E616160B79B69B736E6969";
    attribute INIT_26 of inst : label is "089352184400479E84DF422449D8018C215AD6B5A2C81B1B195A60860A514988";
    attribute INIT_27 of inst : label is "F2D689731B9CF5CCDCDEB66E73D6CDDBD08DAF42528125B2522A454B58A8A8C2";
    attribute INIT_28 of inst : label is "AB5B3594333335A5903757AB6200442DD9A41A4B36DB35B89000389040880FFF";
    attribute INIT_29 of inst : label is "639F493EF8B01F3B4FCE79F3FE18616B2D6BCEC021803B333304B6BB61B75B61";
    attribute INIT_2A of inst : label is "8861BDA809286E2292534A259ADAB415083CB6C76C836A2301509B61B61B602A";
    attribute INIT_2B of inst : label is "99B05250006F18CDDDDD88888F77761B1266E7B844A31946250880A094549122";
    attribute INIT_2C of inst : label is "D8A0AA8843E82B60AA8A7A2B671155108A21164C9A9B534B5876766B360C4941";
    attribute INIT_2D of inst : label is "44106ECCC51043BB3354430EECCD530C14891454AEA810CB5AE802B60A656A8A";
    attribute INIT_2E of inst : label is "000A55F7D2A14A54200410C10C00000004C4C4C4C4C540D006ECCC530C3BB335";
    attribute INIT_2F of inst : label is "9A05201FE7F99685902002B516A08006D0BC4B882F12E25C458002AA8AAAAAAA";
    attribute INIT_30 of inst : label is "644A90A3C0900D44704B938389930254851748E3C9140E0969D7A6959A6818BC";
    attribute INIT_31 of inst : label is "B566D131CB13993F3AE76F2593733A64E79C9D98B1E014781201B88E09727132";
    attribute INIT_32 of inst : label is "8DB6DB336730B0B3985859B0B490452D4154B59552DCD5BA0C4A1C4B1C4CCC75";
    attribute INIT_33 of inst : label is "50339B1E758B9B1E758B9B79D62FDDDCBC15895554517A46C0920C5D488E3871";
    attribute INIT_34 of inst : label is "E44D9DB9CB676DC89B3B6E477673930FB3D6DE67265B7B89EE755219933EB5CB";
    attribute INIT_35 of inst : label is "6DBD18948CC00012E01D807601529E06189810726041C955B3AAA6CEDCF5B3B6";
    attribute INIT_36 of inst : label is "2FDDE0DCB52C85633E5C3838C8546E37650AEC599F2E1BDEF200C924D39ED9B3";
    attribute INIT_37 of inst : label is "640450280A6C00000500B10002D4086CF378F45BBD5339B1C58B9B1E58B9B796";
    attribute INIT_38 of inst : label is "16E3147CB6C0174169B699BB2CC63087180362E6B848F4BDA08F4C2C49DCBAB8";
    attribute INIT_39 of inst : label is "0F48F48691E91E9200A04C8260110500C618C841210822200000000000000000";
    attribute INIT_3A of inst : label is "648052A0250129622C029E540404A0250093A149CE4A54E8CC7319C7318C6602";
    attribute INIT_3B of inst : label is "1067E76281D0089DDB4C925AF224B629624245892C4851D3128915B8CC042EC3";
    attribute INIT_3C of inst : label is "AB4D650A16590A5D71C57BC2500E47A4E143EB85244A4A2777131248CE398CCB";
    attribute INIT_3D of inst : label is "0AD6B28A95DB366A6E4D02199989386248C8C7244110BBD08010000116A8B545";
    attribute INIT_3E of inst : label is "BFAC0108110B00BA30F0660D03CCF05D7113BB2447308A7392424B08A484B121";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000600000573";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "C9A59ABA48F4AC9095A82B5A93B40D12EEB46EC000000000000000000000002B";
    attribute INIT_01 of inst : label is "61240B2AC3000AED46B4E25B56E768D69DCC962961A1AFE687244A482C041231";
    attribute INIT_02 of inst : label is "F9835B0000000053E9DF5BA0CE90575B37A410CED0218E42B63A9AB49D84EC27";
    attribute INIT_03 of inst : label is "7B4EDB4B1A778D3B55C6BAFB2AAD1000000000000000056D01DB0001781B4DAA";
    attribute INIT_04 of inst : label is "AAAD9D9676CA5ACCDE33B652D666F1C7D89D5AED3B4B757676969DB696B4EF1A";
    attribute INIT_05 of inst : label is "F201E61EE95AE72B4E177D050515000074E1F7FAA1F7FAA54EBB1B4B5696AAAA";
    attribute INIT_06 of inst : label is "2C0C25B6DA4937402C402F190000B55446E3B40B71728E80FC9A00000000EBFF";
    attribute INIT_07 of inst : label is "89AA94AAAA0AF80CFB2555451441544445E677FF000695444444455001114000";
    attribute INIT_08 of inst : label is "008813DEE196961084210D2D584A24A000000005FFFEAA2BBADFEDA9AA94DFED";
    attribute INIT_09 of inst : label is "868D3052491068D5580522A43469829200000009EF7986595848088888080880";
    attribute INIT_0A of inst : label is "580B52D0412F275AF216906815A9C2C562D4116A086E0928B42ADA121900A8C4";
    attribute INIT_0B of inst : label is "4A55C30A4582533A14A548560A0AB62D448B2C8916A41321C4584524E374E368";
    attribute INIT_0C of inst : label is "02A3422029256E4CA524C4946E906906900D89445A89049049009D1A91B52DB7";
    attribute INIT_0D of inst : label is "1200B01202424C09813124AFE3F8200225F04F9400016B029111050970200010";
    attribute INIT_0E of inst : label is "88A420000413020488400008211006200100012DFF1022208A2247C9820404C1";
    attribute INIT_0F of inst : label is "000000000000000000000000042006928084060214810A40242240414A912803";
    attribute INIT_10 of inst : label is "0902A6000000000000000000000000002634D5A081DA3896B62D5A5A4A587296";
    attribute INIT_11 of inst : label is "11369280410412410404444555110954A0B040D2BB81C4108A735B0199079B41";
    attribute INIT_12 of inst : label is "092508A934D34D08C44E1AA2230D51515218628A8A90C35444E1AA4148558459";
    attribute INIT_13 of inst : label is "A4D213549294AB088924096055252C0440404412170366CCAAEFFE22112B2412";
    attribute INIT_14 of inst : label is "8D2D28452698A0B0E414A5582CD24008A24120844EC9244116628445AB770C85";
    attribute INIT_15 of inst : label is "1412910525152C152046655259D94904822420125476524A1850202A0A828080";
    attribute INIT_16 of inst : label is "32442829611511234692D1A12D9B910627644441AA2545400862825215600801";
    attribute INIT_17 of inst : label is "ADCB925244428226D050696B72E49412412088888C92A4644A8120214808521A";
    attribute INIT_18 of inst : label is "890E82D68C6C231859844D2C4A4B26269A69A6992CA4A52969A416063428F225";
    attribute INIT_19 of inst : label is "555FFE26B685C0000000004497E869A19259030AA8B6990A6DD1B4B2D2D5C10A";
    attribute INIT_1A of inst : label is "8052A4B4924924842A4A0A0A4850120850545114A512495245489254AAA00001";
    attribute INIT_1B of inst : label is "000000000000000000000000000000000010482492400000824925A7487A0904";
    attribute INIT_1C of inst : label is "0C040C044C444840080008000800080008000800080008000800080008000800";
    attribute INIT_1D of inst : label is "080008000800080008000800080008000C040C040C040C040C040C0408000800";
    attribute INIT_1E of inst : label is "0000000000000000080800004840000008000800080008000800080008000800";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "34A30A5A9E514BA30A30A30A30A5A9C516BB30B30B30B30B5A9E5100122F6916";
    attribute INIT_21 of inst : label is "4CC2CC2CC2CC2D794400000000000000000000CB6E2C49624B932656BA30A30A";
    attribute INIT_22 of inst : label is "92844C90909616264E4E500D864A013262664CC9C9893CD230A30A34A30A5C51";
    attribute INIT_23 of inst : label is "5EB940D242C4C9CC90909672804C3250899CE49092109616264999C993940361";
    attribute INIT_24 of inst : label is "414294AD9EF4ACD0631450419CE58C72CCF3D606EF2C9A0D66666B33316CCCD4";
    attribute INIT_25 of inst : label is "4C724ADFC130036E65BC63101840C964C614614628C517144E61661662CC5979";
    attribute INIT_26 of inst : label is "0206D21047FC78200720036EDCCE81C6315AD6B58CF23B9B9A58820C3051898C";
    attribute INIT_27 of inst : label is "F2D78B629BD88D88DED1B46F62368DDA31C908F253336C938658CB1A116EC800";
    attribute INIT_28 of inst : label is "8A53A544322228512302F56A0447612DD927124224D33804219CE0448EC20FFF";
    attribute INIT_29 of inst : label is "2BB7FE7CF0915FBAEFCC7B7FFF31F96B2D6B9ED545723B2222C4A43241A41A41";
    attribute INIT_2A of inst : label is "308235F3061C80C2727394258ED5580D232434C1098292474FF9B15315314A64";
    attribute INIT_2B of inst : label is "BB0716FC63318C5DF5F5DF5F5A8283129254B50CE9478B8F2E45C5E5D964BB8C";
    attribute INIT_2C of inst : label is "D059FE98E1347341B09C24734632913830D067CF9BCD996B4814444560DE5BF3";
    attribute INIT_2D of inst : label is "1060A888984180A222210402888886104CC110462101188B5ACF67343422679C";
    attribute INIT_2E of inst : label is "5543010008056B5CE3184186100000000606060606043E0002888884182A2226";
    attribute INIT_2F of inst : label is "8F0B647FFFF99796D0C7E5AAD7404002D0BD5BAAAF56E2DD55FFFD50F55550D5";
    attribute INIT_30 of inst : label is "E2DCB1A7E5B4076CF2D99797999796E58D3759E7EB3E5C586D973499D36CBCBC";
    attribute INIT_31 of inst : label is "B567CB204A271073726E6F2D0797A6F4E718B91CA2C034F8B680FD9F5B22E322";
    attribute INIT_32 of inst : label is "8DA6D3324630B0A3185851B0B091D92D6724B50C92DCF1BA5C4B4C4A4C4CCE65";
    attribute INIT_33 of inst : label is "25221A1E759A1A1C659A1A79D6698D14A8B5100000D360CEA1B65C5E59ACB265";
    attribute INIT_34 of inst : label is "8C8D19B11B466D191A3368CB777B9309B2D4D675A75B48C7E8349260D228A16A";
    attribute INIT_35 of inst : label is "69A328948000000DC02D00B4024D9E05289814B2605289E9BB3D268CD88DA336";
    attribute INIT_36 of inst : label is "69CD6596A22C8F66A4C62C2CC8F42F791D9EECC55263100002016BAEF9CC49A3";
    attribute INIT_37 of inst : label is "FE07FEF83EFF103FDFF1FFFF87FFF068F358F2DA332221A1C59A1A1E59A1A716";
    attribute INIT_38 of inst : label is "1EEE1C782602175B6DA699BBAEF7B0C7D88172F6386A6CBF2D9F5E08DCCEBCBC";
    attribute INIT_39 of inst : label is "0F48F48691C91C938190C8CB40911604CE7022658918FC880000000000000000";
    attribute INIT_3A of inst : label is "2E80D6B0258129436C068A540404A0250097B149CE4A50C8DEE73CE6318E6716";
    attribute INIT_3B of inst : label is "B2F6F676FE200DBCCA64B75AE46D93296262E5C92E4843C3931B9518EE2C2FD9";
    attribute INIT_3C of inst : label is "0210100C1B5B8A1041046BE2701EE285E1836BC56EDADA6F33131288CE79CEE3";
    attribute INIT_3D of inst : label is "8AD6B288111F3E6F36659631311130A258988B2441188400FF1FFFF1400A0050";
    attribute INIT_3E of inst : label is "BFFC0000000FE56933B13621FC13001041B7996E6438C84312424B8C8484B931";
    attribute INIT_3F of inst : label is "00000000000000000000000000000000000000000000000000000002000042DB";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "A236487FF3023242428084204882E0C8A211E240000000000000000000000018";
    attribute INIT_01 of inst : label is "E592C33324001910714709E429188E28E212F8468D8D9B024F93016CB1B65842";
    attribute INIT_02 of inst : label is "5897080000000069FFC708D267410F08FFD242E60B0FB702109349F2C7963CB1";
    attribute INIT_03 of inst : label is "C679B66E3BCD3DE6449E79FE776800000000000000000C9006480000FA48FFBB";
    attribute INIT_04 of inst : label is "2227735FCDA373FA34FE6D1B8FD1A3CFF2F1B599E66EC6CDD2DEF36CDC779A3B";
    attribute INIT_05 of inst : label is "02001E00EEA05288C1D77DF5F54000007413FBF543FBF5457966C96B32566222";
    attribute INIT_06 of inst : label is "2C040DB136C800402D3AF0B90000B00006E14BD4A02D4E8FFDE200000000E800";
    attribute INIT_07 of inst : label is "EDFED8AA220AC00C26F541010401544555FF77FFFFFFD5555555554005414000";
    attribute INIT_08 of inst : label is "0808BEB5A394DCD6B5AD6DB9A37A24A0000000040000AA8BBA9AA929AA96DFED";
    attribute INIT_09 of inst : label is "36C5987FDF6BEBDAB8320C41B62CC3FE0000001F5AD48E51A378800808088088";
    attribute INIT_0A of inst : label is "632B1AC365B198319968DB80C20645028B4065A0B1A023E4B424D9DB79192348";
    attribute INIT_0B of inst : label is "6D9A182D8A1D089AC2D1A16860F390640B14CB162850E88E17A108B70C830C83";
    attribute INIT_0C of inst : label is "4B2B6B2086D8912210921A4190C12C1AC0267473A32C12C1AC0264C91C90D248";
    attribute INIT_0D of inst : label is "000262885188330660CD1A0802004184200000004822943A588ED520B0CC30D1";
    attribute INIT_0E of inst : label is "000020241452020000404A2082100400255821B1001000008000040002000400";
    attribute INIT_0F of inst : label is "00000000000000000000000004003048108000020001000090A90A28B1428802";
    attribute INIT_10 of inst : label is "AD9D3D00000000000000000000000004B8C71232DA2340D8D8D1A3636161F858";
    attribute INIT_11 of inst : label is "88FEDAD96DB6596D9659999889889666C941345AE88C475A4B113B04E090376D";
    attribute INIT_12 of inst : label is "2CB5C445B6DB6D29172A613B95309C88C96184E4464B0C67722613256B4A2360";
    attribute INIT_13 of inst : label is "33D95466DA52B4446C94C5818994B04000440056732500EEAAEFFF118894965B";
    attribute INIT_14 of inst : label is "9CB5AC89D96332C7F1D294A2D31926313B65B2E2312C9486698CE23613779E16";
    attribute INIT_15 of inst : label is "26D8D505B8EFD1EFD679999B66256D96CB16A04167895B26DB5C90C4310C6312";
    attribute INIT_16 of inst : label is "CC324DA5888888BD6ACB1EB5966288991882372633923324318CCB4AD28064C6";
    attribute INIT_17 of inst : label is "1223C90B222CD11FDB5B068488F2424965B2C444730B37822CE4B2A06CA8192B";
    attribute INIT_18 of inst : label is "EB3ECB36F5F1A723668C2CB02B2CB0B6DB6DB6D8BE3735AD8DB41E22BCAEE69A";
    attribute INIT_19 of inst : label is "555FFEB6C691401FC000FEE257ED6DB58B58A7374EC6DE6B71BBF2CBCB0A452A";
    attribute INIT_1A of inst : label is "495AB6C6C964B6B5AB6B2B2B61425929595768D6B58B2D9B76645B26AAA00001";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000596CB6DB6D6B5ADB25B29764BB2492";
    attribute INIT_1C of inst : label is "0800080008000800080008000800080008000800080008000800080008000800";
    attribute INIT_1D of inst : label is "080008000800080008000800080008000C040C040C040C040C040C0408000800";
    attribute INIT_1E of inst : label is "4040404040404040080800004840000008000800080008000800080008000800";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "92C92C98495E92592D92D92D92D984B5E92592D92D92D92D984B5E802CB19658";
    attribute INIT_21 of inst : label is "B64B64B64B64B66D7A0000000000000000000E3490C3761BB05C630B2492C92C";
    attribute INIT_22 of inst : label is "E80036676761E09131B300027BA000DB8B9B736E6E6ECB2D92D92D92D92D9B5E";
    attribute INIT_23 of inst : label is "6136624D1C122636676761980033DD0006C637676CE761E09136442E6CC0009E";
    attribute INIT_24 of inst : label is "6C094A5304A6516C10C34D305296020B045B685911AC6C8659292C9495925259";
    attribute INIT_25 of inst : label is "711BA11000001891124318C00CA21C2A1259299232465656A125929923246565";
    attribute INIT_26 of inst : label is "2C5A6CA08400400004001891222366318C318C63350DCC2465A3451041042E21";
    attribute INIT_27 of inst : label is "098CC46B0B9AF5AC5CDEB62E6BD6C5DBD085AF5B884EDB6C7BA774EB5E911104";
    attribute INIT_28 of inst : label is "C3DABDA0111117ADD49B4993121006B22091890116DB1694DA420011200C0000";
    attribute INIT_29 of inst : label is "044048830E8E0040102BC1C3108404C618C6218FB0C6C411116236B365B65B65";
    attribute INIT_2A of inst : label is "D1454245BD800677C909291089DAB8360C41B6C06CC3FEBD9156496C96C961B2";
    attribute INIT_2B of inst : label is "6E1CDD86B5AD297200AA200AA002A8C96C22E71D86BC6E78D9B63616430B6634";
    attribute INIT_2C of inst : label is "D92CAB6F99732B64EC71292B66DD68E2D345A86CDC98738431D2223BC3B1B60E";
    attribute INIT_2D of inst : label is "60A3A44475828E9111D60A3A44475A28A63020842002C60631B192B66920BACA";
    attribute INIT_2E of inst : label is "00020100000C21020620828A28C30C30C4040404040400013244465828E9111D";
    attribute INIT_2F of inst : label is "810CD80000065841031012B528A1800240401C07900700E01C80000080000080";
    attribute INIT_30 of inst : label is "0B22C619364418D30D2278586278591630C1A65934C36360B658DB652DB2C2C6";
    attribute INIT_31 of inst : label is "42986C589B38D98D8DF19CB198784B09CE52C6D6BDC0C326C8830A60A44F0C4F";
    attribute INIT_32 of inst : label is "2E38DC1138C7471C63A38E47472F74989DD2627749878D64B375B375B373294B";
    attribute INIT_33 of inst : label is "D05B5B5B59EB5B5B59EB5B6527AC298932C9E800030C1B32462963616621858A";
    attribute INIT_34 of inst : label is "F76D88B5EB622DEEDB116F7588A76D47B166DB66D9A369CD920B64883112B593";
    attribute INIT_35 of inst : label is "6DBDD2EB3FDFEF7F90D243490DFFE982D2E60B5B982D6EFE445FF6C45AF5B116";
    attribute INIT_36 of inst : label is "AC69B60B3DB1656B364A32B2D2792EF936CAED759B251BDEF5869451052975B1";
    attribute INIT_37 of inst : label is "FF07DC7C1F3E101F0F90FBDFC7DF796C5B6C5B1B1DD5B5B5B5EB5B595EB5B657";
    attribute INIT_38 of inst : label is "2351E1961A0861A436CB2444525291C822848D28C8E303445220A313222142C2";
    attribute INIT_39 of inst : label is "F5B75B3B6EB6EB658251122002244011630008B032C600200000000000000000";
    attribute INIT_3A of inst : label is "916108585AC2D6BC8308718B0B0B585AC2E95E36B5B182376B5AD294A52B58D8";
    attribute INIT_3B of inst : label is "CB0B4B788000624A22F348319BDB6C860B99186EC374AC88C8E462D691B1C4A4";
    attribute INIT_3C of inst : label is "0200001521A47169A28A84198C251C1252A434789121219288DCDD77B4AD291B";
    attribute INIT_3D of inst : label is "618C681046A1B37261CE58C5C5EDC74BA2E2F5B882108000FF1FEFF100080040";
    attribute INIT_3E of inst : label is "155C00000019C850F056490900000169AC49449199CF339CDD9DB0F33B3B05CC";
    attribute INIT_3F of inst : label is "00000000000000000000000000000000000000000000000000000000000002A9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "0034007FE3001246070004600112C4808401C440000000000000000000000031";
    attribute INIT_01 of inst : label is "4502C333C000100023820B4030200470442050E7050D11020E02116DA19250C3";
    attribute INIT_02 of inst : label is "9896010000000071FF8E018046042601FF8007804907140002118122811408A0";
    attribute INIT_03 of inst : label is "4228926A3B443CA2001E71F220A000000000000000000800040100009001FFBB";
    attribute INIT_04 of inst : label is "0001515F448353E810FA241A9F40878F92D4D088A22A5344405E5124D4768839";
    attribute INIT_05 of inst : label is "020001FEEFFF88083FD77DF5F500000075E7FDE007FDE0056BA2007E207C4000";
    attribute INIT_06 of inst : label is "2C03FDB00137FF402D3B9FC10000BFFFF6DEABD55FD54E8003FBFFFFFFFEE800";
    attribute INIT_07 of inst : label is "09AA90AAAAAFFFFFFFF555545154411045F877FFFFFFD5555555555551014000";
    attribute INIT_08 of inst : label is "08803A108184D4D6B5AD69A9C35AF6F8000000040000AAABBADFEDCDFED89AA9";
    attribute INIT_09 of inst : label is "1245113FDF6B43CAB81600F0922889FE0000445D08400600C158000880088800";
    attribute INIT_0A of inst : label is "432A1A836DA091738B705901800C0E03098104C000C003E4940451493909204E";
    attribute INIT_0B of inst : label is "261C15661C10845AA6E9D130C04102C01C38083870E8844456110D9218121803";
    attribute INIT_0C of inst : label is "0B292B004000029508495D2102C0AC02C015422A11AC0AC02C0154A988000001";
    attribute INIT_0D of inst : label is "0002E61CC318610C2185300802002002200000005A6B186248889420A00D34C3";
    attribute INIT_0E of inst : label is "0000202C34D2020000405A69A01004002C5A68A1001000008000040002000400";
    attribute INIT_0F of inst : label is "000000000000000000000000040022E03480000200010000B98B9820C1A34802";
    attribute INIT_10 of inst : label is "A4B1910000000000000000000000000490821016C80108505060C14141417450";
    attribute INIT_11 of inst : label is "88FE5A5B6DB65B6DB65999999C88B8724B80B6522800424A4B11390288901724";
    attribute INIT_12 of inst : label is "64B4C444924925081762C39BB161CC8C89430E64644A1833762C196D294C2340";
    attribute INIT_13 of inst : label is "33C950724A52B8446C948D001CB5A0444400003415414088CC899911889892C9";
    attribute INIT_14 of inst : label is "94BDE4CC90419687E8D6B5C2601924039B2C9662202C94803006623419779D14";
    attribute INIT_15 of inst : label is "3248D501A0850185072001CB44052CB25912A02133014B245148900401004013";
    attribute INIT_16 of inst : label is "002264A5088888952A5A0A94D40088B11002376C199222240306594A53002480";
    attribute INIT_17 of inst : label is "0053A40B232E511FCB4A2C0014E902CB2C96444640099223266C96A025A80929";
    attribute INIT_18 of inst : label is "4A2E4A0245E1A303408069A069681492492492489D1414A504A40602A8A5D4B0";
    attribute INIT_19 of inst : label is "555FFE9242894000007FFEE2D3E524948948A3076682482920A3A2868A0C452A";
    attribute INIT_1A of inst : label is "495A9642C964B6B5A96929292346C96B4B5328D29489248932244932AAA00001";
    attribute INIT_1B of inst : label is "00000000000000000000000000000000004B25924925294A5924929724B92492";
    attribute INIT_1C of inst : label is "0800080008000800080008000800080008000800080008000800080008000800";
    attribute INIT_1D of inst : label is "0800080008000800080008000800080008000800080008000800080008000800";
    attribute INIT_1E of inst : label is "0000000000000000080800000800000008000800080008000800080008000800";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "BA4BA4C82948B25BA5BA5BA5BA5C82B48924BA4BA4BA4BA4C829488024A09650";
    attribute INIT_21 of inst : label is "96E96E96E96E972D220000000000000000000C400201400A0050420B24BA4BA4";
    attribute INIT_22 of inst : label is "880036040401818885BB0007222000CA1A1B432828688864BA4BA4BA4BA4C948";
    attribute INIT_23 of inst : label is "41932141103110B6040401D80039110006C21404008401818880A22866C000C8";
    attribute INIT_24 of inst : label is "2A19AD604109616C38C30C30D6B4031A044A30D000A46C86496964B4B492D2C9";
    attribute INIT_25 of inst : label is "431A001000001102880B18C005A6182E374B6CB796F2D2D2E17496C9792F2525";
    attribute INIT_26 of inst : label is "2C5A70800400400004001102051360318C739CE73424804080C34D34D30C2861";
    attribute INIT_27 of inst : label is "0B9C4C29090A44A448489224291244891084A44A084800012224448948911082";
    attribute INIT_28 of inst : label is "A1CE94B01111122D15991CB90A3000A000B08B01124912841242000120000000";
    attribute INIT_29 of inst : label is "227A482596970960592DE1A2949CCDCE39CE7987900680111166129934934934";
    attribute INIT_2A of inst : label is "C30C000CBD800077DB196B3083CAB81200F0927C2889FEB491524B24B24B202A";
    attribute INIT_2B of inst : label is "22045486B5AD2B57FF557FF557FD54493022420C90942A2868B41414020C2AB0";
    attribute INIT_2C of inst : label is "48ACAB88997329228A132B2926117422C30D81285010220C6352222A4090D20A";
    attribute INIT_2D of inst : label is "6986244445A618911116986244445861823000042002460E738492922920C2CA";
    attribute INIT_2E of inst : label is "00020100000800060261869A6800000004040404040400016A44455A61891111";
    attribute INIT_2F of inst : label is "2B2FF800000450C00030321570A00000000030020004008010E00000E0000080";
    attribute INIT_30 of inst : label is "0A0684113C0408E20E02D0D0C2F0D0342080C45118894140B650C92525928286";
    attribute INIT_31 of inst : label is "03116848B190CB0D0DE1BDA0B0F0DA1BDED686D291C0822380810C40C04A084E";
    attribute INIT_32 of inst : label is "241048113084041842020C04042C4480B11202C44806250DC144C144C141294C";
    attribute INIT_33 of inst : label is "1059494B5C89494B5C89492D7224688B968C880002080E20002141414401060C";
    attribute INIT_34 of inst : label is "4464889489222488C911244599A731479132492260C128C1120C448821129499";
    attribute INIT_35 of inst : label is "2491128C0000007FB016C05B01FF88821682084A082128FECCDFF2444A449112";
    attribute INIT_36 of inst : label is "2468B40B91A1652814421696967B24F9164A45240A2108000480904105294491";
    attribute INIT_37 of inst : label is "0000000000000240000200000000012449244A09111494949489494948949252";
    attribute INIT_38 of inst : label is "23808B061C0401C036CB2CCCC00000C00282100080628184E000C11605118282";
    attribute INIT_39 of inst : label is "C1C41C218838838780101660012CC00921000090024200000000000000000000";
    attribute INIT_3A of inst : label is "4360005862C318910300400B0B0C5862C2814800000006136B5AD6B5AD694DD0";
    attribute INIT_3B of inst : label is "8A1B5B708000440912E80173890001001A1820280145A8985C4082529BA10482";
    attribute INIT_3C of inst : label is "0200001561C0C161861800182C04303056AC18200200050244505136B5A529BB";
    attribute INIT_3D of inst : label is "639CE034C604A14041885084848D0C5A024244A0001080008010000100080040";
    attribute INIT_3E of inst : label is "BFFC0000001AC060C1876D0D000001618881220221044210501000442020050C";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000400004552";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
