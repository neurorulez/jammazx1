-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "5EED595E58E5E5DE58CCB9C488EE9B14E5AA7DCEA236071C8868C6B2E384045C";
    attribute INIT_01 of inst : label is "044101049550465559F5B9E0ACC966A5A69761BF2DEB619EDDC56565656DA269";
    attribute INIT_02 of inst : label is "D62DBA09C6995AB6F78271A456DBDE996FE11ED005C5C05B65975DE551A46955";
    attribute INIT_03 of inst : label is "558B73720573B435EDFB61AB52FEADEDC8177B4041815E54185597B70C80B55B";
    attribute INIT_04 of inst : label is "6502514D59CDE5A86D962E2FF2945927189757805275D74DB6E1B6D965C5D559";
    attribute INIT_05 of inst : label is "615B58775156D45DD415B50459E48792484BDE1206E141D859D8BA07585E5A85";
    attribute INIT_06 of inst : label is "105794A0106779C05796DE105ED81C65C11E50574BC9C19676150575956D65DD";
    attribute INIT_07 of inst : label is "36361281265D4952657809C1814575EDDED745D67765A49C0794105795E00794";
    attribute INIT_08 of inst : label is "3C87ADACA1B558149A2580D9F576367D5D84A818569E5295D6A1894357C5E968";
    attribute INIT_09 of inst : label is "85B657965C85F67FC1607008A0107F9B655B5B56805A23F23D16C90A575AB682";
    attribute INIT_0A of inst : label is "7F97ED6874E169400C87657D57D965D686595D786B67EA84A5949DB490AAAC04";
    attribute INIT_0B of inst : label is "03A275E89D682AAC4961EB1849DA4909499D69D7BD7974996D26D95566650752";
    attribute INIT_0C of inst : label is "EBDD596D70BFFEABAAAAAB0E8DC498D0D890D8D000159D6D7B657AA0AAA0AAAC";
    attribute INIT_0D of inst : label is "06596397A8B5B4E927D6AD7DEDD57B4EDB4ED0AAAF0E8DC7A375EBC5EBCD5B45";
    attribute INIT_0E of inst : label is "9DED7F222389A0FAE02000C9ADC9ADC9A95D7AA0017165BF94927C1F65419595";
    attribute INIT_0F of inst : label is "659FA4B66DA7B630046D9F92D9B69ED8C074659F5A4B69ED80061C510730C3C1";
    attribute INIT_10 of inst : label is "7B899B67FF2300F7D967E92D9B69ED8C1472D9B6359967E4B69ED8C05810A69A";
    attribute INIT_11 of inst : label is "9E7BA1D12866E6569867C99967F8434104D0C0101878574D6251967B21E19196";
    attribute INIT_12 of inst : label is "6AAD99D111199001122236E666D223EFB8396662766A86960934765BC117B255";
    attribute INIT_13 of inst : label is "15D5D5151501044659FE000574A59B4C357D65759967FA996519FE84115AD56B";
    attribute INIT_14 of inst : label is "FFFCEE1BCFCEE3BFDFCE6FBFFFD595D7D5959F97D517555D5DD5151515555715";
    attribute INIT_15 of inst : label is "FF38EFBFFFFCCE3B3823BFFFFC3B7B61BFFFFCDE3B78EFFFFF378EFFFF37BE1B";
    attribute INIT_16 of inst : label is "B8EF8E3AFB8E3BEFAFFFFFFFFFFCFE3BFFF86DBFFFFCFE3BFFFB6DBFFFFCCE3B";
    attribute INIT_17 of inst : label is "FFECCE3BEC6FB28E3FFFF338ECE3BEFFFFF378EDEF7FF7FF378EDEF7FFFFF3FF";
    attribute INIT_18 of inst : label is "FFFF3B8EEEF7FF7FF3B8EEEF7FFBFFE3BFFF86FBFFFFCFEB8EFFFFF3FBEFE3BF";
    attribute INIT_19 of inst : label is "5C555554554555554557555557554554557408A2378EDEE7EF7FFF378EDADBEF";
    attribute INIT_1A of inst : label is "5555555555555575555555555555555D75D75545575575575555555555555555";
    attribute INIT_1B of inst : label is "65555557165965575565575565575555555555575D7554554556555554554556";
    attribute INIT_1C of inst : label is "155955155155355B55355F5555555515575D3559555551555555655755755755";
    attribute INIT_1D of inst : label is "5555555555155555355D55955155555755555D5557D55DD55D55555D55D55155";
    attribute INIT_1E of inst : label is "57D57D57F57D57D57D55D55D55D551D55C55C55C55C55C55C55C557595556D95";
    attribute INIT_1F of inst : label is "555545545555545765745775765745775765745775765745775B55D55D55D57D";
    attribute INIT_20 of inst : label is "2355D9EADDC6A116D7E8E6DBFFFDD55155D55D55155D55555155155555155145";
    attribute INIT_21 of inst : label is "AAB3A83AAEAAAEAABA0CAACEB3ACEAAABAAC0AAAAAB14A5F0457A5F205DC8557";
    attribute INIT_22 of inst : label is "AFFC2AABFF0AAAFFC2AAAAAFFC2AABFF0ABAAAFFC2AAABAAABFFC0EABAAABACE";
    attribute INIT_23 of inst : label is "56984A5BCEF3B4EC3BA6499C606011A3BDE17D61F626285076975C70AAFFC2AA";
    attribute INIT_24 of inst : label is "154496072355C85772055E8567A355C8D6765BDEE82AF2AABCAEAB0098041E8D";
    attribute INIT_25 of inst : label is "0FFFC0AAAAAAB1805807FAFB57EBE117C5315AFEE05666253291567F06E141C9";
    attribute INIT_26 of inst : label is "7BA0AABAAAB03AABAABC0A83A0AABAAEAAA0AAFFFFFAA0AABAAAAA0AAAEAEAAC";
    attribute INIT_27 of inst : label is "32AEAAB004BA3559D1432F549F6C861CBD5E7DB2AD417B7665D9976B45C8D476";
    attribute INIT_28 of inst : label is "79C9556CAD57237DD9EE89AC9C140B3AA9DC33AEAC0CFFEB03B0EC3B0EC3B0EC";
    attribute INIT_29 of inst : label is "F79D6FCAD97A3E257CA3DD7D1CA0797C3EC0F832AAEAAC012E8D57205D79C85F";
    attribute INIT_2A of inst : label is "675ED9E563605D8D20105A3123643A355C89C7217DC8DF767AB9E5965E980492";
    attribute INIT_2B of inst : label is "40DBA1858041E85E7A355CB2AB6D87B6DB7A7D5A57BFEE16D59A6A5D7E7DF679";
    attribute INIT_2C of inst : label is "B03AEAAC0EAAEAAEB3AACEA0EAABAABAAAE832AB3ACEB3AAAAEAB02AAEAAC603";
    attribute INIT_2D of inst : label is "958D8176360105A3123643A355C89D7217DC8DF6A65965D9EB7EA82AF2ABCAEA";
    attribute INIT_2E of inst : label is "B3A83AAAEAAEAABA0CAACEB3ACEAAABAAC0AABAAB180E952957BF5B6716D5B67";
    attribute INIT_2F of inst : label is "0BB85BB81159251F07E8D572151C81772059C8D6767BA0EBAAB03AABAAABACEA";
    attribute INIT_30 of inst : label is "3AAAAABABF0AAABAAAABFC0AABAAAC55603AD805E947A1010757405005005005";
    attribute INIT_31 of inst : label is "AAF00AAF00AAB00AAF00AFFC0AAA00AA00AA00AA802A802B03EAABFFFFEAAB00";
    attribute INIT_32 of inst : label is "DEA5A56856D6B7607269E632315DD91E8DB9AEEAEB409051EBE175FAFE0AAA00";
    attribute INIT_33 of inst : label is "21A61A69A6597B65ADCCBCE096D696DD2DA566615595BFB8524A49595ADEDD4E";
    attribute INIT_34 of inst : label is "C2AA00AAB17A95D7B94112FB6D2DB50D695C204C8557581668C8D6767B6A17AD";
    attribute INIT_35 of inst : label is "DA9A25F5A51D956DF86D7B355686D15BFEE16DA7A9A75A98617B0AAAFEBC2AAB";
    attribute INIT_36 of inst : label is "AB02AA82ABAAC164BD271761F732259895F5A5E548584BC5D5DA322517AE4BE5";
    attribute INIT_37 of inst : label is "B676556116AA2298716D075B807569E50496BA5540843892256599A50AAA0AAB";
    attribute INIT_38 of inst : label is "6191E0A5556A4290A66DB4426519FF9045585A59B619769527353B449D6661A7";
    attribute INIT_39 of inst : label is "7B4697E56B6DA95D75DD75D656EE59D6EE51204656D5B56D5B569A16D59615B5";
    attribute INIT_3A of inst : label is "97BB6215FEF5FEF5567F9E7F9E6611ED8750D00DD8DE817B43634361F2DBAD69";
    attribute INIT_3B of inst : label is "B7B56E05B5E5DB56FBB85B7B85E70437986384BF69A4D7B94B795A1DB5F495B7";
    attribute INIT_3C of inst : label is "885E21E225E1B87D1ADE18C2D75E54BF6F99866D6698CD85ED95A53AE0D8D05D";
    attribute INIT_3D of inst : label is "AD58967BB8C689856844581D556944574BF837A61AF3F90E035952A59A699863";
    attribute INIT_3E of inst : label is "8C11B479D8598DEDD8505E5D7DB95BA97B6663607198589C5E8BD8DF5850B77B";
    attribute INIT_3F of inst : label is "ABE778795B59595661356EAA5358ED31DA5869D69E2D0445A667DA26559F9A64";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A80AAAACB8EF36B365EC662861712E383A55EA894B0FD9EBFFC6CB490F98DBE0";
    attribute INIT_01 of inst : label is "CCCA875E6FBCCDFEF1EB2BA0D88AACAA6A7FDB6EEE2BA3F323DAAAAAAAAFD4CA";
    attribute INIT_02 of inst : label is "AE3E2557DC33AB49AA54F70DEA26A977AE2373247EFE15C6996FBAFF371DF6FB";
    attribute INIT_03 of inst : label is "6ADEBE863EE7FDEBBEAAC52EF9A97EFA18FBCE95F33EF36F33EC7CDA9855F994";
    attribute INIT_04 of inst : label is "F2576EBFF3BB369E9FC9686AA460979A28D8FE8FB5EBAEAAABBFEBACB2FA0AAB";
    attribute INIT_05 of inst : label is "E3B7F8FFFEEDFFBBFE3B7F8DA6D85B6195A6A57CFA8F9593E9B3A2FAF3B369EA";
    attribute INIT_06 of inst : label is "63EEFB557D9FE743EEEBE275B3A53DFAF673A3EEB793F67A7FFBFEFFEEDFFBFF";
    attribute INIT_07 of inst : label is "7DFDE9561BE286A1BEE557368FBEEF3EB3EBDFF6AFF75A695CEB63EEEB955CFB";
    attribute INIT_08 of inst : label is "5B4A7A7E477FF57D995F95E4ABE8F92AFA3A5571EC3326EBFD972FA6BE2F2FA5";
    attribute INIT_09 of inst : label is "73EBEEEBAE63FD68F5FD8E7B9BEFBA04FA3EAEBC15B0166D3A3FE65BAFF5BC11";
    attribute INIT_0A of inst : label is "AD6F1FCEB924AC955E4ACAA2AA2CF3BCEB7DFDF8CFAE95597ADE7BCE7AD58658";
    attribute INIT_0B of inst : label is "57D9EBF67BD6965586C7F77FE7BFE7539ABFDBAEAAE3CA3DDB8F37DDEEFFDEB9";
    attribute INIT_0C of inst : label is "E7ABFEF26A5FE5C90B27409F7FADB53535B57575553AABE7ECBAE55AAFAA50F6";
    attribute INIT_0D of inst : label is "FFF7AEFC55DAD98B9AF8A6EFF3FFFD93EA9EBA46359F7BDFDEE3E7BBE7BBFDBB";
    attribute INIT_0E of inst : label is "B8A8EA48AECA8905B77155B72FB72FB72DFFE5555FBF9E8EDFAFBBAE5FFFFD7F";
    attribute INIT_0F of inst : label is "FFBA59B5AD5A35687BF7BA66D6B568D5A1EBFFBAF59B568D555D34D38F209207";
    attribute INIT_10 of inst : label is "E65ABDEEAA4E85EC3FEE966D6B568D5A29C2D6B57DBFEE99B568D5A1F5EDFEA9";
    attribute INIT_11 of inst : label is "796B7E835FAA2AFCBDEEBABDEEAF960A9981A1A93FBFAEBFDEA7FEE6FE8EA7FE";
    attribute INIT_12 of inst : label is "955FFBBFBFBFB55EE9ECE8C888BECECF314AAACA2ED558387AE0EF7A9ABEA7FF";
    attribute INIT_13 of inst : label is "FA7A7EBABA9A9BBF7BA9557EED6AAAD14FEF6BEDBDEEA5AA9F3BAAE9B6F3EBCF";
    attribute INIT_14 of inst : label is "155134936410595164129551543A7A6F7A7A3FBFBE7BBA3E7E3EFAFA7AFAFFFF";
    attribute INIT_15 of inst : label is "5082510D1741379C86595515C19C85595454C1179C065545304DE73110450590";
    attribute INIT_16 of inst : label is "DE7575D6C9E7D1556C5401551541279F50B2551D1751279F50B1551D0751279F";
    attribute INIT_17 of inst : label is "1165279D505D4755D074541E7179D5F75D041A60649A89404DA63649B8540550";
    attribute INIT_18 of inst : label is "457055A6574DD855051A64649B850779F51F2510D0751775677045D5014479DC";
    attribute INIT_19 of inst : label is "EFBEBBEDBEDBEFBEDBECBEDBE9BEBBEEBEC962B155E7570DFDC25555E7495551";
    attribute INIT_1A of inst : label is "BEFBEFBEFBEFBEEBEFBEFBEFBEFBEFB6DB6DBEDBEDBEDBEDBEFBEFBEFBEFBEFB";
    attribute INIT_1B of inst : label is "EBEFBEFBEBA69BEBBE9BEBBE9BEBBEBAEBBE9BEBAEBBECBEDBEEBEFBECBEDBEE";
    attribute INIT_1C of inst : label is "2FFEFFEFFAFF7FFFFFFFFFFFEFFAFBAFB7FBAFFEFF2FF6FBEFBEEBEDBEDBEDBE";
    attribute INIT_1D of inst : label is "BAFBAFBAFBAFB2FBBFB3FB6FA2FBEFA7FE6FEA9BEFFEDFEFBAFBAFBAFBEFBEFF";
    attribute INIT_1E of inst : label is "FFAFEAFEBFEAFFAFFAFEAFEAFFAFF6FBF9FF9FF9FF9FF9FF9FF9FF8AEABFEBFF";
    attribute INIT_1F of inst : label is "EDFEFFEEFEDFEFFFFFFDFFCFFFFFDFFCFFBFF9FF8FFBFF9FF8FFFFAFEAFEAFFA";
    attribute INIT_20 of inst : label is "98F7A657E38A7AFB6E95F9551543BFFFFFFFFBFFFFFFFBBFBFFBBFBBFBFFBBEF";
    attribute INIT_21 of inst : label is "2449D68E7566571593A2216609F641EC1612A878055B0FFBD8EE8FB99FBE63DF";
    attribute INIT_22 of inst : label is "C59AA4C966A9655DA9049805DAA4B566A591DE59AA07D9C6B1762A39D7C75327";
    attribute INIT_23 of inst : label is "AD7CC4F2089238CD3398A62CCCE3E6DE6A27EFCEEE0E3FEDBE3EB3BADD5DAA0F";
    attribute INIT_24 of inst : label is "FBBE74FB99EBE63BF9BEFF678FDEEBE639E9A6A516974918D2C5DC9538DBEF7B";
    attribute INIT_25 of inst : label is "ABEB6A076C401BC578FAB9AADEE687AEABFCB2ACCE6888CE796BBAEABE8DB6E6";
    attribute INIT_26 of inst : label is "945A545D1BCA954551D2A0290A4C95171BDA6555555E5A595F7105AD58676042";
    attribute INIT_27 of inst : label is "896477995C7DEEB7E6979FED2EDE5CFE7FB8BB795FEFADFDBFF6FFDDFFE639E9";
    attribute INIT_28 of inst : label is "E3D7FFDD4BFF98F7A651570D3D39C80A57F2890706A25540A9BA5E9FA5E93A4E";
    attribute INIT_29 of inst : label is "AB6A9AD72E857D7AAE5FFF7B6E55F7829B2A6E881452D6571F7BAF163CE3C67D";
    attribute INIT_2A of inst : label is "AEBCB2DFE2E3EF8B23EDADE61DD97DEEBE67BF98EFE63AE9954AF3CFE17C5C69";
    attribute INIT_2B of inst : label is "8596938B8FB6F7FBFDEEBD615EBEEBFBA98EAAF1DEBACCDAFF3FAFA3BAEF2CB3";
    attribute INIT_2C of inst : label is "CAA05652A1657F64C954275A2471595C564E88859827D907B0584A8145656F17";
    attribute INIT_2D of inst : label is "7F8B8FBE2E3EDADE61DD97DEEBE679F98EFE63BD6B3CFEA65F89569748552C75";
    attribute INIT_2E of inst : label is "09D6891C53271593A2216609F641EC1612A0514C9BC594F99EAABD2CB7A2E2CB";
    attribute INIT_2F of inst : label is "8A2BEA2BE3AAEFFEE8F7BAF9FF7E6FCF9AFFE63FE9945A814C8A84C97C753255";
    attribute INIT_30 of inst : label is "85D1515655A83F15A6D552A0510FC6FEF16538FBDFFF6FF6E8FA74B84B84B84B";
    attribute INIT_31 of inst : label is "545AA215AAD19AAC55AAF556A110AA54AA21AAD1AAB16ABDAA675D5557675DAA";
    attribute INIT_32 of inst : label is "AA4F3A94E5FC9A5DA187173331777FD5DACF58A695F535F3E687EBE5A9AC91AA";
    attribute INIT_33 of inst : label is "7EEBEFBAFB2DBE9EB30609B0DAFCFBA932BF888DBECA2B3367A7E7F7B7EFE203";
    attribute INIT_34 of inst : label is "EB9EAAA6C9F5EAAE3EB679AEBAE9BBCB8AFB2F9E679EF2FAD9E6BBE994A7AE7B";
    attribute INIT_35 of inst : label is "29A27A3E3EF2DEF33EE6947ABCEB362BACCDAB2BBFEEF3BFFA94A9D7661EA75D";
    attribute INIT_36 of inst : label is "D0AA75EA6154665A5B9EDBB28E79AEB5EB9F3EFEB595A5B6FEA279AEB951E7BA";
    attribute INIT_37 of inst : label is "BBCAFBE705980084EFEE5EA7C4FF4B9A5D71A3D7D13D23E97EFE6ABAA9D7AD59";
    attribute INIT_38 of inst : label is "C3A6D12AAE9490240AAF6AA6AEBBABA7BAA5D5AA8C366ABB9A7A4B9D7AAAC36C";
    attribute INIT_39 of inst : label is "CBAEFBDFCFAA94FABA72BA3CAA8EA72A8EA756A9AA2A8AA2A8AAF0F82AAE2F0A";
    attribute INIT_3A of inst : label is "AC03E22F21EF25EAABC86BC96AAC3B2E56B4BC4BB8B893E3D3E3D3E1AFE2BEF6";
    attribute INIT_3B of inst : label is "7CBB9B1DAA9FB6BCE803FA803F2BC96CB1D6CE6B9B1DAC03D3CBD22B9BAD2D2C";
    attribute INIT_3C of inst : label is "C8AB22B22E812C6FD2AB13C26EFE3E6B9AAB1EA31C350B8B2EBB1A65B1F8FCFB";
    attribute INIT_3D of inst : label is "2AF8BAC02C0C5B1E8EAAA53FEB1ABAAEE7AC7CAC7D83865B17DAB56AA6C7B0D6";
    attribute INIT_3E of inst : label is "7F25A963F8FB3F2EF8FCB4FEDB23F227CB9ECFE3C3B3F8B2E956B8BEF8FCBAC0";
    attribute INIT_3F of inst : label is "258FF3F2E2E2F3EEC3BFC89AA7A93E779DB826F22E1A6A986AEEADEAE3BAB1DB";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "7BE8787FED2A32A3A05D065D8A7D355B3214C75C633CFED7DB505456D8CDFBE4";
    attribute INIT_01 of inst : label is "54480515756545F5984E27C4C1180660731D461F9A56BCA32201E1E1E1E7CBF8";
    attribute INIT_02 of inst : label is "F876345A5493133DFF569524C4F7FDFB0F58E3243EBE545597583834B1247756";
    attribute INIT_03 of inst : label is "FF9DAD9C7E6CF1D9BE607DAE19EC76B671FA8D90DFBEE3ADFBE458E94D11DAD4";
    attribute INIT_04 of inst : label is "FE472DAD9BE63A558FF856155A05459601E9661FA9E18E3861BCDB6CB6B67FFB";
    attribute INIT_05 of inst : label is "5867570F5E19D7CBD586757175DC5579D567F1BAF96F947BE47A59FB9A63A559";
    attribute INIT_06 of inst : label is "E3E6DA45BF89F553E6CBE584E3A126FEBE23E3E656DA7EB0F7C7F1F5E19D7CFD";
    attribute INIT_07 of inst : label is "7535B5551FE54751FE654A3E8DBE6E36E3E1CD637F70167D08FBE3E6F98448DB";
    attribute INIT_08 of inst : label is "1F0B7E3D097F55B41C6D15F73EBE3DCFAFAD5552581320F9F416CFAF6E061F95";
    attribute INIT_09 of inst : label is "58EBE6FB6C7C741387CFFD43DBFDE146FE3F8F9A946231FC3D77D143E7D11893";
    attribute INIT_0A of inst : label is "E55DD665A32EDF91444CFDCF4CFE75E65B9F571F6F9F45157ED50FF540DDD444";
    attribute INIT_0B of inst : label is "53143DC54F4437794741C51750F5544B001F41867B998D8C4773535FCEDFDE19";
    attribute INIT_0C of inst : label is "D6FB5F3AA0E089D65F775D1C78D6BAFAFEBE7E7D14B13C7CFCB261408880888C";
    attribute INIT_0D of inst : label is "F5CB0F7111E8EB69966AB266389E6EB3EEB380775B1C70471D31D5F8D5EB5EBC";
    attribute INIT_0E of inst : label is "7D5715A0579CC405A165145FAD5FAD5FAE3DF1444DADAC1FE36D9BEE8F7D723D";
    attribute INIT_0F of inst : label is "5C7D00791E41B91960787D01E47906E465E25C7D6407906E454D79E7DF5175D1";
    attribute INIT_10 of inst : label is "F50CDE1F55A9943A571F401E47906E4655E5E4791A971F407906E46564087488";
    attribute INIT_11 of inst : label is "7CD61675D58071EE9D1F4CDE1F5581D805746508A7878E2D917571F51E693571";
    attribute INIT_12 of inst : label is "8141DD1DD5DDD448358FEFFF7FF8FEF9DC534DF956513E26769DE785489F51C6";
    attribute INIT_13 of inst : label is "7FD7D73F7F58102787D545366760CF81176E219A9E1F518C0507D578719B6E6F";
    attribute INIT_14 of inst : label is "D7D6CE3F4DEC63DD4D6D27DD5D775737F775DFF73537D5BDBDF57F3F3D3D77B7";
    attribute INIT_15 of inst : label is "F730DF7FD7F6DE3F78D3EFF5D6373BD3EF7D5EEE3FB8FBFD75BF0DD577B73F37";
    attribute INIT_16 of inst : label is "38FFEDB4D78F37FFCD7D5F7FF7D64E3FF530DF5FE7F65E3FF573DF5FF7F6CE3F";
    attribute INIT_17 of inst : label is "7F4E7E3DD4AFDBAFB57FD9F2D7EBFFFD5F7938F4CF76D6FD978F5CF75D6FDB7D";
    attribute INIT_18 of inst : label is "FDFDB30DCEEFE70DFB78FDCF75DEDCE3FF730DF5FF7F6FEBCFF5FDFBF1DDE3DD";
    attribute INIT_19 of inst : label is "D77DE7D67D77DF7D77D67D77DE7DE7D67D7541E5B38FCC776F25F5BF8FFEF5FF";
    attribute INIT_1A of inst : label is "7D67DF5D75D77D77D77D77D77DF7DF71C71C7DF7DC7DC7DC7DF7DF7DF7DF7DF7";
    attribute INIT_1B of inst : label is "77D67DF5D77DF7D67DF7D67DF7D67D75D77D77D65967DD7DF7D77D67DD7DF7D7";
    attribute INIT_1C of inst : label is "7F75F79F55F7DF75F79F79F5DF51FFBFF7FFBF57F57F5BFBD67D77DC7DC7DC7D";
    attribute INIT_1D of inst : label is "F9FF1FF9FFDF75FF9F71F77F73FDFFD3F53F5FEFD6FDDF9FF3FFBFF3FF9FF7F7";
    attribute INIT_1E of inst : label is "F5FF7FF5DF7FF5FF7FF5FF7FF5FF7977DF7DF7DF7DF7DF7DF7DF7DFFBEFD47BF";
    attribute INIT_1F of inst : label is "DE7DE7D57D67D67FE7FF7FF7F67F77F77FE7FF7FF7F67F77F779F5FF7FF5FF7F";
    attribute INIT_20 of inst : label is "1F31F797E5CF56FBA6C6D2FFF5D7DF7DF79F5DF5DF59FF9FF9FFDFD9FD9FDDD7";
    attribute INIT_21 of inst : label is "7752DE2D7B757B5D678CD7CB72D495D5E75C0575D5D1177DD0CEC3F1E1DC5CE7";
    attribute INIT_22 of inst : label is "7A2A1F56AA8777A2A175DF5AAA15F68A85E5DDAAA177D6F7D68A40B5E75767C9";
    attribute INIT_23 of inst : label is "D53146B9B6DF976EFB766FB36B87E51B7B787668D94977EFBF0F2210DDAAA1DF";
    attribute INIT_24 of inst : label is "1677CEFB1C19C78771E1DC5CE71D35C78C7D77B95037B1DD64D9DF11A1FBEC74";
    attribute INIT_25 of inst : label is "0888C0D7757D531161F9B5679ED789D3B07F8D5EE3A3660C3115675F712FBEC5";
    attribute INIT_26 of inst : label is "E540DD6F5F702DD67DEC0F42D0F5675B5FD0F7AAAAA558DDE7D5F70DDDB79DDC";
    attribute INIT_27 of inst : label is "317977511471D35E10071E5ABD5C54DC7966F5710D586C717CC5F31C7CC7C47D";
    attribute INIT_28 of inst : label is "49D79F0D65B31F39F7951AA0A530022313D4325B740CAA9702E0982E0B82E098";
    attribute INIT_29 of inst : label is "F559DE472C94713E6C4B9EB57C449B3421C0A4315D97D4451C74D7D34E41F7CC";
    attribute INIT_2A of inst : label is "C6621FAD9797EA1DC7EF91B1150D31D35C74E71735C7CF7DE453B8C7E5311459";
    attribute INIT_2B of inst : label is "D4A79A1E1FBEC78C71D354451CBA5AFBEC979BB8D665EEF939B7A5B3E8E607C7";
    attribute INIT_2C of inst : label is "7027B7740B77B759F2F5CB78B75EDDED759E335F2DCB5257579D7015DB774C45";
    attribute INIT_2D of inst : label is "3E5E5FA8687EF91B1150D31D35C74571719C7C444F8C7EF79F9C5037B17ECDBD";
    attribute INIT_2E of inst : label is "72DE2DD7BD5B5D678CD7CB72D495D5E75C0576F55311C6D9AFA39987C7C7887E";
    attribute INIT_2F of inst : label is "1587E587EB13F3DFF9C74D7173DC5CD7173DC7CF7DE5409EF5502F5675767CBD";
    attribute INIT_30 of inst : label is "2DF5F5E76A877DED57DEAC0576DF74F7C471A1F9D7075CBEF96E21E91E19E99E";
    attribute INIT_31 of inst : label is "F5A88D7A88F5E88F7A88DAAC0DD588F588D788F5E23DE23702B57EAAA8B57D22";
    attribute INIT_32 of inst : label is "A079BAF4FD66CA9F85F5D0202140006CFFC0BF8FBD15317DD7C9EEE47D05DD88";
    attribute INIT_33 of inst : label is "5679E5967BAEAFAC3C4551A4CAE6CB227638766F92FBD7BBE7D3D3DFF76BE473";
    attribute INIT_34 of inst : label is "03DD8857F2F9D9BBADBE59EDB201BE9EEB9E5F8C78D79B8C48C70C7DC5F56638";
    attribute INIT_35 of inst : label is "7D1A7A5BB263C5B5A532C540E65B47F65EEF81E29C77994556C50D5FAB60357E";
    attribute INIT_36 of inst : label is "D70357E3765545166D96785EA631C191E989B232554466DE1ABA31C11C4465BA";
    attribute INIT_37 of inst : label is "6982757C203D55203F1A4E035046E38D1A5D0A61AF8ADAF47E7E0CFE0D5F875E";
    attribute INIT_38 of inst : label is "4103CFA07B427E972F3F242334C7D480200014001490A0C996C0C48878334118";
    attribute INIT_39 of inst : label is "869DEA166F9A84D800B4203FC06207406A06120005F17C4F43D0E2EEF4084BBD";
    attribute INIT_3A of inst : label is "9BBB872A197A197003865E865F34921A0FF5ED5FE5EE5599D784C787C3627664";
    attribute INIT_3B of inst : label is "1868D6786A575BE6F79866BB8A231D38924196791907FBBBBB8A9B23C99B9A98";
    attribute INIT_3C of inst : label is "B906E46E5ACF997639A6F857A6E346591E01240414909A9A1A68501D64E9E175";
    attribute INIT_3D of inst : label is "9A6969BB99914123F6A0001F4016A006679938949CEBB0164586895A8249D041";
    attribute INIT_3E of inst : label is "4CF468FBEDF58E1AEDE5EEFDBF98A890869D63B58B586DE1E50BEDFF6DE56ABB";
    attribute INIT_3F of inst : label is "93EE9BB899BB99D64136E247AC0F3E6FACE176FFEF49020B734E69336C7D904B";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "551909055FA77E77E0322EFED2D71D937A444557F70F18B3F7ED65DC25261040";
    attribute INIT_01 of inst : label is "76313246D47760515737A92F7FFBC7EF06651035B01CBDD769856564242E7889";
    attribute INIT_02 of inst : label is "54FE94DDCA40C1C85777729230615DE84D31976E0484117D38D4513D42815D45";
    attribute INIT_03 of inst : label is "55BF210FC644F711BCE15EAC7B27F0BC1F1BDFB12C46D7E2C464E5FACA31F15E";
    attribute INIT_04 of inst : label is "BEC7C125D96F7E5F86F8FD1FF1215FBEA9F076B193451451C73DC3CD30841559";
    attribute INIT_05 of inst : label is "555E557A5557955A9555E5576D74F4D74F4E5B251BD1B4D46C46F518DAB7E5F9";
    attribute INIT_06 of inst : label is "4846F24D8127765846E3030C57235F3C8417E8467E71C484555657A5557955A9";
    attribute INIT_07 of inst : label is "57979F713BC04E13BC631544A1046372772EA27B553144D705F84846F18C45F8";
    attribute INIT_08 of inst : label is "ADC37535E55957881CE2346D060E9B4183A7C7291E8764DA51006F22566F4FA3";
    attribute INIT_09 of inst : label is "D9CBC6D367D9515920F18A2388E3A590B4AD5DF6B45A99B70CAF7C536D550E99";
    attribute INIT_0A of inst : label is "24D9B76F8F6ACCB115F57F5FF57D3976FB4E675B6CA45136F4E196C19A3052D4";
    attribute INIT_0B of inst : label is "C5775C5DD512A0274FA85D4C556F55DCD12513B4599ADD1D564795674545347B";
    attribute INIT_0C of inst : label is "4E494574EA57D4656594E8B5D54337773A3A72331184243D9D38644A500AAA5E";
    attribute INIT_0D of inst : label is "03D845F453D5DD5BB642B46535250DD72D135A2137B5D151745C4C554C594D55";
    attribute INIT_0E of inst : label is "9165555BE361BC5B701B1165A665A665AC54544C5121210DC4C118C63444F4D1";
    attribute INIT_0F of inst : label is "BD9114737CC6735D04B99151CDF319CD7444BD91DD47319CDD1D79E75C55559E";
    attribute INIT_10 of inst : label is "4141AE645559D01E2F64453CD7319CD740E4CDB37EAF64547319CD74DC11DDD9";
    attribute INIT_11 of inst : label is "D4563E67BF842C36AF646D6C645F959110657431DF2F944F7922F641BC9822F6";
    attribute INIT_12 of inst : label is "844BFFB337733C511FB1155555231159570E187A5D050E3ACC994B19412493DD";
    attribute INIT_13 of inst : label is "D797D7D797F1044B1914C4446EE51BD54667A75AAC6455955BD917F061DB2D6C";
    attribute INIT_14 of inst : label is "6575D491221D1955645D95554457D71717D71797579717975757D797D7D7D794";
    attribute INIT_15 of inst : label is "477655554755C597365D75754597B149313161C597375D515171651088755597";
    attribute INIT_16 of inst : label is "5651F4967965904D64DE01017545D597775655557775D597775555555775D597";
    attribute INIT_17 of inst : label is "5565E5955C5575555D1557565C4904414487D24F55572D5D7524D5554215D5D3";
    attribute INIT_18 of inst : label is "551D6D24B4111214C6924A555621D9597765655557775A5D65995596F5595945";
    attribute INIT_19 of inst : label is "5655555555755555755755555755555755472F9865E794113ED77765659D545D";
    attribute INIT_1A of inst : label is "5545555145145565545545545555555145145555545545545555555555555555";
    attribute INIT_1B of inst : label is "45545555965145575545575545575555555545575D7557555554554557555554";
    attribute INIT_1C of inst : label is "555155955D55D55155955955555551B55155955555555D515455455455455455";
    attribute INIT_1D of inst : label is "5155D55155155155D55155D55155555D55555D45545555D55D55155155955555";
    attribute INIT_1E of inst : label is "5595595595595595595595595595515557557557557557557557554554556575";
    attribute INIT_1F of inst : label is "5555655755555655555755455555755455555755455555755455559559559559";
    attribute INIT_20 of inst : label is "F54C4D370166FC13C67D59555445955155955955155955155955955155955975";
    attribute INIT_21 of inst : label is "12393EA1041D044858A288E5894A771ED0A2A5C6873898929634475F4407DD21";
    attribute INIT_22 of inst : label is "151A922546A60251A86042951A9A5156A9571155A92C052145566A8410131827";
    attribute INIT_23 of inst : label is "010D2EF8760D8F63D8362D8F684C6571701155E946DDC861291D56DA3C5DA9A0";
    attribute INIT_24 of inst : label is "C721D519F4487D101F4445D10175407D51136D9312BC4884DE24F0B1131065D5";
    attribute INIT_25 of inst : label is "A0152AAC50CA78D1131A1325CE4CA446117407FB990175B15F4043354791847C";
    attribute INIT_26 of inst : label is "4C4A8293352A9829251AA0A9AA2250A4541A1755555D4A809C870CA305515682";
    attribute INIT_27 of inst : label is "8A55C47B12D7540D9151F31C7207CA47CC7DC81F41116F4B352C54BF157D5013";
    attribute INIT_28 of inst : label is "291D5541E955F5444D3135A9DD0430F3155289E4AAA2557AA94A6294A6298A72";
    attribute INIT_29 of inst : label is "94C9B67F4E04D334E7C8C78877CE7852942A528B4D694EC4B5D500F112293D10";
    attribute INIT_2A of inst : label is "06565618EDDC6FF1CC6117153458575407D101F7407D51134D00BDF3C10D12D3";
    attribute INIT_2B of inst : label is "91CDF1FF31845DD2175407D74C38F2C30D0F398A16EFB919AD9F2F2218A55486";
    attribute INIT_2C of inst : label is "CABA6022AA02501609A5A4FA9189809121628A23962529DC7B428AB4D602E344";
    attribute INIT_2D of inst : label is "63B771BFCCC6117153458575407D121F7487D53103DF3C4D3C07D2BC4969A259";
    attribute INIT_2E of inst : label is "693EA46248944858A288E5894A771ED0A2AD352278D17CBBA86096948E015958";
    attribute INIT_2F of inst : label is "F7706F7868420645205D501F4607D1A1F7607D59134C4AE9224AA22501318269";
    attribute INIT_30 of inst : label is "A033B3D155A68050514152AD35A01E55345F131AF46BD184205E2F5B757F5F75";
    attribute INIT_31 of inst : label is "A55AA885AA335AA025AA455AABB9AAA5AA88AA336A80AA92A9536555555366AA";
    attribute INIT_32 of inst : label is "21E5BA8FAB76DB31179EB666650CCC4E5DFC3E8E3F0D41944D64E4E4D5AC48AA";
    attribute INIT_33 of inst : label is "F0F30F3CF34D2C2131272AD8D276E3247839575190C17EE46F0F0D469F0B0237";
    attribute INIT_34 of inst : label is "6851AA514897D19BAD84FB6C3084B1326BDFD197D1B1D91A197DDB136C6FC671";
    attribute INIT_35 of inst : label is "1B1EF81DBA76D1F8AF746CC576FB9D72FB918564BDF55BDC7E6CA4D955969365";
    attribute INIT_36 of inst : label is "02A936690924AD74C7B24284A65F7647E1ADB8BA9F5C4C509C9A5F7686D0EDB8";
    attribute INIT_37 of inst : label is "FA5E9CB9B23AEE1C757ED45697975D58C4E366B846A47AC771F355F3A4D9AC45";
    attribute INIT_38 of inst : label is "E93695A5BE1A9EA3AAC6A8C46BD916B445556DF30A874CFBB2455C96D175A84D";
    attribute INIT_39 of inst : label is "5F9BCABD6CBC90B94FA14F2194DAF614DAFDB44553645B0611847A7E6126CC98";
    attribute INIT_3A of inst : label is "8D965F676F5F635556DBF5D8F46A837E576777F6F3754EF6ADFD9DCDFBCAFE4E";
    attribute INIT_3B of inst : label is "4DF9384EF9F949555D165F996F66985DAA161EF97A81CD96DAD96B66D19DBDBD";
    attribute INIT_3C of inst : label is "13584F8DF3B7A1B58BE8CA9746D3DEF9761290C13A05FFF17EC5BF6785735394";
    attribute INIT_3D of inst : label is "7ED3CE596136D2944D8455E53D3EC454EDA15DAA87B18518455C9379B2A86A16";
    attribute INIT_3E of inst : label is "CAE2F97E77EDEF7E3F3796EE9FB79A6CDF8B7BEDDEDEB3F49F5933653BF7F859";
    attribute INIT_3F of inst : label is "6DEADBD9D8D8DA72A02429BBE45D72E1A77B3A63AA6A4CD4C6B55F869991A815";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
