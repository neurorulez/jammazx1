-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "4BFFD0783552C0EA031A9A75E6E9AD86B7DFD4FFFFA9FD693DFCC581FDE7E7DD";
    attribute INIT_01 of inst : label is "122218EBAA9724E0B09FFFFE585E76517DBD5B895A92EB013445FB7B96A1E59D";
    attribute INIT_02 of inst : label is "7AC115F5095A243B320ACC06E96074A3E64A228060029211310CA70809C85DF7";
    attribute INIT_03 of inst : label is "05827AA9F4637D9F1A6619987CBEB9FB9D7F9FFE7F351881FFFFEDFF759FFF11";
    attribute INIT_04 of inst : label is "A6A82D563436C75C7B9ED0DD2E1F4FE3AACCFA89FCD27A78D84DD8D37423FC2F";
    attribute INIT_05 of inst : label is "A9FFDE19FF99B9FB6F9819142DEEC335569DBA772EB1EC7BA6BD5177FF3C0F22";
    attribute INIT_06 of inst : label is "882800020A0A08AA2A80001F5DD74AAA7D6AFD054B8D9AAAA81EAC2FFECB979E";
    attribute INIT_07 of inst : label is "5695A5695A5695A5695A5695AF3815A5695A5695A5695A5695A5695774BAF888";
    attribute INIT_08 of inst : label is "8CDEF3C8D65D1DCFC2CB13CF2279E44F3C8A4211405B1777582220A5D3FBA95A";
    attribute INIT_09 of inst : label is "920A41ACBA1E786B2E87FD963CF1ACBA359746B2E8B2C4F3C8CDEF3C89E79165";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFE8200000C0000112444431002AAC200001089090100900";
    attribute INIT_0B of inst : label is "FFFFF0778B3C971B49E8AFFC455B7B1D03FC455B79D08010697392A23A3AE709";
    attribute INIT_0C of inst : label is "066D6E046AE39085524CCDB30028A348815980855276CCCDB30332944A669101";
    attribute INIT_0D of inst : label is "B4F53B24BC1C200433824B4859A4DA5B512D3873F99C6616A4B40709FFFF8000";
    attribute INIT_0E of inst : label is "E01041041041055567D8025242B3CF789D14D3F5FF0DC78A67939839EF5B5871";
    attribute INIT_0F of inst : label is "8C28838C201BE3BE21851041C4510514180101040E4EFFFFFE30410020805FB2";
    attribute INIT_10 of inst : label is "8200208009A28808A088698EF9024545501810011041171040B4C34CEA26B2C8";
    attribute INIT_11 of inst : label is "08218608A38E28A21441C61C66B9699C11431C41410C7104490412417D71DF38";
    attribute INIT_12 of inst : label is "67B6700010416FA4BA4BA4BA4B26BA6FB4FB4FB6F34BB77C75C830830830E58E";
    attribute INIT_13 of inst : label is "B04608C11823056C15B29B39B39B39B39B3C4CF533865B3839B392DB3DC4CF5A";
    attribute INIT_14 of inst : label is "E22CFFFFECF664BD0CED6DA19FAF1A3330BC46613708CC33B119E2321555460B";
    attribute INIT_15 of inst : label is "974026019CF7873B7CBC9F3EF3E8F9CEEFEDEED977F1CFF52CADCAD90AF212EF";
    attribute INIT_16 of inst : label is "FE4F9FF27FFF81C27C9FF3E4F9FE23C7F9327EC5CE07FC1FF07F88888A6069A2";
    attribute INIT_17 of inst : label is "3E7299729D659205A65C92465E55E9F7299B473CF5BE92647198727886D1FFFF";
    attribute INIT_18 of inst : label is "739E7BD7CA646B76E838EAD5E306F54844CBE5A82DCFE8FC88199FC853F902FC";
    attribute INIT_19 of inst : label is "116424584998842390CD6511D153B9534BC9A7493CCC1C1B79C8B9DCF9A739CE";
    attribute INIT_1A of inst : label is "B724FAA3B54AEE000004437CEE848A47E4321EEA5A89D51511ECAA2E6EAA0111";
    attribute INIT_1B of inst : label is "8952093D65C725016854133092848C23960A4E84265E45224E0421365A4D3650";
    attribute INIT_1C of inst : label is "DA485469282C81B56D3A473089352C21C808721CBEF6C8A230CCB93B64CDE9BD";
    attribute INIT_1D of inst : label is "6DCBBC8817E9EFF621C085F8CCFCDF4E1ECDE8EE20495D757CDFCA4E9A92C841";
    attribute INIT_1E of inst : label is "28E035B4E9B54D010E3CA9526A95655BB565084A5084389E1802020204521ADA";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE5767621C38EBEC3800001";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "187CD56BA4EB2CA409274AE7BE6C9CE4B1FCB8E265CF30033A4EEC0674AA33FF";
    attribute INIT_23 of inst : label is "157AD69B2883656DFF0946320BF3E3E71EC91FCEF4726B9EAC90D2D559E770B6";
    attribute INIT_24 of inst : label is "ECD3FF0D8FFBFD4FE7E9F9276F753F336CE52E0344AB90A89DC31C5AC4D86F4F";
    attribute INIT_25 of inst : label is "820000005D6FBF6793F551CBAE7A0020800C108208300108008556F8C2029278";
    attribute INIT_26 of inst : label is "34110EE438C07454ECB6F8D5FF86DF6028044337900FBED679299CC104100820";
    attribute INIT_27 of inst : label is "B06669002930D0D441E4C4D8631E59F69DED0ECFF33738FB2FA0C868325831F6";
    attribute INIT_28 of inst : label is "2031882081BB063401768B4AA406340610BB462AA176C338BDB5FE79CE549851";
    attribute INIT_29 of inst : label is "1341B158C1A8B4AA4063406EC02063F79F68B35480C6208206ED18D547DA2CD5";
    attribute INIT_2A of inst : label is "47D1B4A99823C8A8D2B90EC85643B9D09D29E69F889041FB986E61A083BFE644";
    attribute INIT_2B of inst : label is "CEAD255ED53F36C04A6D93DBDD6C74AC7FA4C5E6B49B54FCDB01306D9274AC7E";
    attribute INIT_2C of inst : label is "6963311CF28162579F5555D9248541E3A1256507C75CDA8A4840840855A36769";
    attribute INIT_2D of inst : label is "3900329E296824D5D1ADAED7E80CFFFFFECF364097B3B812D998910220F8AC18";
    attribute INIT_2E of inst : label is "5DB4FFFFF5602EF75408A230910A11468D80E6AABD95D20167929D6ED4E0CC64";
    attribute INIT_2F of inst : label is "05F1B6CCC6AF9E36CC6AF91B7034EB980DDBB23D2E35EFE4986CF2BCBA4B4962";
    attribute INIT_30 of inst : label is "59A2649324A493B5FE426F4DF09A9180DA957C6D84CC6AFDC6DB31ABE06DDAB6";
    attribute INIT_31 of inst : label is "843231AF0CA68C1BE6BE94E6DE5795FBF6AFCB5DB7E9274247D8CF91F5F29652";
    attribute INIT_32 of inst : label is "072AB528C1BE6BE9CD22F272E771824C93289BE9DB02CABCAF95A94327EFEF2C";
    attribute INIT_33 of inst : label is "5211F49290CC1213E549A92534A4D4929A536A6D4DAB3D5BAF97A6AFB7CBDD37";
    attribute INIT_34 of inst : label is "FB81567850050C817E53ED48817F9D9604A6D910B3129F6A442CC73B2C094DBE";
    attribute INIT_35 of inst : label is "E9EF256DF90B2172902D908F902F908D908DE1204D42684E5FF35E0C9A7B699C";
    attribute INIT_36 of inst : label is "20595508E704431423DEEF38124348690D218D2CDBD473F8E9B2930E343DC4B2";
    attribute INIT_37 of inst : label is "B857EE15E6B0EB389597029C48E270100804221531A3987181223000000804E5";
    attribute INIT_38 of inst : label is "109190104D04DA82ACD1251112F629092058D23318AE152275DEEC3F0C34C658";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFF090901211929191139193918043C041C340C24340C0C1019010";
    attribute INIT_3A of inst : label is "D980927958D9811B2B79DBFF9DCE739FFF87B4915C63F19E86DFD56400F3C835";
    attribute INIT_3B of inst : label is "FC136ED3ACE7EB673EE63D03363826629158844EF59FF5111D153B9653E2D916";
    attribute INIT_3C of inst : label is "10186AB57E7CD4DE76BEDDA9594DA65B4D948ECB47D21B64C2330F6EBB4ED367";
    attribute INIT_3D of inst : label is "28889E0D781A3C051820DA309E9D3D0E46089685122900D28458EF23B34D5CFB";
    attribute INIT_3E of inst : label is "FFFFF7EFDFFFFF9FFFFFF6FFFFFFFCFBFF7FE7EDFCF8DB5402B4AD2B4ACD42E2";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFF7C58DCFE98FEE4FC63369779938F58DFFFFFFFDFFFFFFF9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "D48009907FF7F968B386397F8460B569980090BFFEF3C783FAFC8B13FC0EC79C";
    attribute INIT_01 of inst : label is "A50E5BD515038DE4340008FECCBCA46FE9A28D19AB8FB189EABC876CA79E8A97";
    attribute INIT_02 of inst : label is "D6B43D7F53FB6D081CDE17E9266D80DA3AC70B5F6D3375CF141569363D5979D7";
    attribute INIT_03 of inst : label is "20162114188415C1E54055015B20221853D0070080331B31FFFFED5414AAAA43";
    attribute INIT_04 of inst : label is "08028603091014D4ADED7AB2DBA091CB9CC02914116D458290A9692A5A6C8460";
    attribute INIT_05 of inst : label is "73FFB6297F9951C1E8C9C8A043604A000320408387C2E4B819E0054C0516E594";
    attribute INIT_06 of inst : label is "82088888200A02882A88AA2088001F5FFF40027D6AFD87FFFA23D1281061D52F";
    attribute INIT_07 of inst : label is "2008020080200802008020080810000200802008020080200802008160C8FA82";
    attribute INIT_08 of inst : label is "684B4996A932DA22FB06DC22DB845B708B697AC86F42C8A20008A2864143C080";
    attribute INIT_09 of inst : label is "004979C22D9936708B602E0DB26DC22DAA4CB708B6C1B708B684B4996E116D83";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFE8600444800440061011240077F8000024400002400000";
    attribute INIT_0B of inst : label is "FFFFF4AB90816550B0F659576A63B82A9D576A63B8A99133AA48FB5C4CD49164";
    attribute INIT_0C of inst : label is "023E41DB5E299D5BA1B9B25132D2F6F457C39D5BA18B25B250133D269B0DE8AC";
    attribute INIT_0D of inst : label is "485340615B5100000F643413A48951F528D237ED263B0CA2466EB6F4FFFF8000";
    attribute INIT_0E of inst : label is "3000000000000BBBAD3691AC9D49B50F0BC12198FF025C6596000DC210289BCE";
    attribute INIT_0F of inst : label is "C31430C71C628E0858E08A3861CF6CB18648268A210FFFFFFE00000020827F56";
    attribute INIT_10 of inst : label is "71CF1C33C30E30E39C3B8A3800C59A18278418E78E38718638451C2050CF0C73";
    attribute INIT_11 of inst : label is "E71E71F75F75E71DB7CF3DB6D8A2060668A48218209A28E14D3CD1450106000C";
    attribute INIT_12 of inst : label is "8A181F3DEF8E9861A69863AEB861A69861A698E3A69C7841C207DF3CF7DF3775";
    attribute INIT_13 of inst : label is "A0C4188310620DC83722B23B23B23B23B23FE8FFA3AB7239EB238EF238D88E22";
    attribute INIT_14 of inst : label is "C649FFFFE8E4661EE8FD73511DAE6E2325F4C4619E988C27D311FF23FFFF841C";
    attribute INIT_15 of inst : label is "8F462A390C7B4A0190492802007E8200B1A33260808BB12BE5F25F227C012E13";
    attribute INIT_16 of inst : label is "FE4F9FF27FFF81C27C9FF3E4F9FE23C7F9327EC5CE07FC1FF07FDF5F5AA2D171";
    attribute INIT_17 of inst : label is "4017079703998466C285606282F8324E628B297C012208198005818462CAFFFF";
    attribute INIT_18 of inst : label is "A52480715F793D9B27E5B6CCE591F09804A7C42004063627D3A24013E0027603";
    attribute INIT_19 of inst : label is "EAAC4DEB06A45D4CF9673EE266A00A0194609B3C5851090B7290B2D9608A5294";
    attribute INIT_1A of inst : label is "58CB0FF09326335AD6AA6DC000C153B02D56E724893E2BABE2558150A6542BAB";
    attribute INIT_1B of inst : label is "BFCCA0C008717C44DCAA2D4B3F8B124CFF4EBDCB1EBDCB128D085A006D5A0064";
    attribute INIT_1C of inst : label is "A8DC88A3D449726F3A08F17888CA4997A445E9B96F70926FAAA93A8097183A07";
    attribute INIT_1D of inst : label is "321035D3A0360014423D2B0100022150A200D47A6602C121912DF58237F65AF2";
    attribute INIT_1E of inst : label is "8EF9DCE83B9904D5B3533A7C114EA2241696358521484701860220022156B773";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC510014402086201063860";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "730E0BC00B76C9C1F65AFE0C4050630B576153BE4298A2D810B1B2F95117A8FF";
    attribute INIT_23 of inst : label is "66A018EBBAD67603FED67AA4E62D4C9AA90E2A40F8E8A045FFC9C622625EA764";
    attribute INIT_24 of inst : label is "2CCA6011F7C321D81A3D2618A473C16C943A5C052878B9510059C26E5778CD15";
    attribute INIT_25 of inst : label is "8008008016D080102C9FF8D695500400000000010400400400008A7F0D2D2436";
    attribute INIT_26 of inst : label is "C2EAC03FD59499A815082CCCFE1BEE583000ADADA660816102DD4D4804800800";
    attribute INIT_27 of inst : label is "B363E52B42DD7F6A8DC338771D2CB649750EB802AAB35E8054255AADD6E35C06";
    attribute INIT_28 of inst : label is "9942E1475E413840AD48B4C45338D83AA94128422D4BD9412FF7FEAFFFE16EF8";
    attribute INIT_29 of inst : label is "AC2B42A166CB4D55338DD3904952842A549B528A650B851D3904E1209426D422";
    attribute INIT_2A of inst : label is "000A9114234E1711444B955C8AE55C4DEBFA022026EEA208208022273E005DDD";
    attribute INIT_2B of inst : label is "AA785A8A2260291E35982CA91CF3511540CB1AD5E1688980A478CF982D511140";
    attribute INIT_2C of inst : label is "90848A75A62011842289EEEB8DC8A250B087AE4962E04E3E8000020044150193";
    attribute INIT_2D of inst : label is "BEFFCFD19680032C22571209840000000776EABB608D076D0C256A334B83CD8F";
    attribute INIT_2E of inst : label is "04F2FFFFD9C441089CAD1C4F4FB7FF6BC598764C0B292CCC102DD2924B9BB9DB";
    attribute INIT_2F of inst : label is "68ED400CCDF41DAC2CDF60AD9F98302FD26CB689407282123B0A286228800005";
    attribute INIT_30 of inst : label is "059D006803000CDFFEC80600D559BAFD27AF1B5928ECDF41B500B37D92B657D9";
    attribute INIT_31 of inst : label is "6357337145F1BDAD0672711202F8BE0D16665B220CA3753AE81392B841280100";
    attribute INIT_32 of inst : label is "B0E1F37BDAD06722240037B7D896E5A00CF621B62002DF05C2B99E2568C955C3";
    attribute INIT_33 of inst : label is "84F821010C05A1846800000000020048010000000007BCFAE2BC11E4F15E023A";
    attribute INIT_34 of inst : label is "385CE4CB1A22E93A0380227D3A03630C631A2BA749BD251BE9D26ED65AC6B44B";
    attribute INIT_35 of inst : label is "B0D04B06C2749CEC27C027C1274027432751280A01903202E4C330E938806500";
    attribute INIT_36 of inst : label is "86036622403C982CB3F11411641C8380760ED4E03439DFF96400DD777C801BA6";
    attribute INIT_37 of inst : label is "C0B0B02C240166118858160CC50030389C06030309722C00D383002000000461";
    attribute INIT_38 of inst : label is "5050D0505F31EBAA849586559BE74D2508CD92B25AE0C7B4808A064004135041";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE0000080818180810000010012101390901013921010125250D2";
    attribute INIT_3A of inst : label is "9E5424A2D81109A9F272067FBF94A524FF06B14C876C1DA2FA347F9199A8FD8C";
    attribute INIT_3B of inst : label is "4ADEA5E1C0065400317A8B535680589102A332802FF52662266A00A2C5174F90";
    attribute INIT_3C of inst : label is "DC5E03FF0BDEE3057D6D5B5E4B3892C50CB3C058A05E815D8AA7E7AF317D9AFD";
    attribute INIT_3D of inst : label is "B5F5E5C1E9C2C628E25482461A3035A4102E1250038F7A1AF21C3F20F37FC7BF";
    attribute INIT_3E of inst : label is "5D555B854CCD4E19CCD55AD7335559A9CDB542A524A85AEEEAB5A52B5A510280";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFF8C2AC02A8A607031786C950585462FE0F66666A5AEAAAAA3";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "32280482CAA518219A84280A6A6510690A9F917FFE539293F9FE8301F80FD3AC";
    attribute INIT_01 of inst : label is "A50210C545018CA00407F4028C0000AE8D064195910D219DC4B8142EB506C180";
    attribute INIT_02 of inst : label is "9CD789EF50A8E91918D41EAA0F4104AA0A855A5649008247A00B4B292C585DA6";
    attribute INIT_03 of inst : label is "3596592FEC85DD7EFF264C993DB88827CAAB880BFF211031FFFFC4AA45155378";
    attribute INIT_04 of inst : label is "A8FAFE7F1D129281C6B5A2677FB6DBACEC86419FF7B72EB26CA5E1597A4B7A4F";
    attribute INIT_05 of inst : label is "520024A9555174CFEC0484B46A43C91FFDA7EADD7A73ECFAFD77F431E0826096";
    attribute INIT_06 of inst : label is "2A028282088288A02A82882A80AA208A281F5FFF4002FD5552815903ABDE8237";
    attribute INIT_07 of inst : label is "0040100401004010040100401817E9500401004010040100401004AA8203FA80";
    attribute INIT_08 of inst : label is "0A020090C0161802C32611064220C8441908430458C20880222228A018410401";
    attribute INIT_09 of inst : label is "00084110641830441900A64C306110643005844190C9844190A0200908832193";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFEC311110911110030000201120A9080000060400024024";
    attribute INIT_0B of inst : label is "FFFFF4CC1F6FB4480802060A3BBAC333960A3BBAC3311B42CB11AD80E66623C4";
    attribute INIT_0C of inst : label is "231A3E88942E2080063959B0328B22A00686B080061FA159B192A8A404C5400C";
    attribute INIT_0D of inst : label is "3442E04BBA4520000A44759BAA3CC0A539D424FC4F925166B22BA4BCFFFF8002";
    attribute INIT_0E of inst : label is "0000000000000FAFAF3413ACDF55F0E31AF52B84FF0259CC4040351F90A2D2EB";
    attribute INIT_0F of inst : label is "A59258001024104924820C20028210424B34D249550FFFFFFE20000020820056";
    attribute INIT_10 of inst : label is "41400000009838C01E3090412412C92490491493410C60002149249269208209";
    attribute INIT_11 of inst : label is "C30D34C30D34D34C75D71D31E924924020800020000000828808800852492480";
    attribute INIT_12 of inst : label is "104906D96DB69A6B8E38E3AE9AEB8E38E3AE9AEB8638F4820920D34C34C32430";
    attribute INIT_13 of inst : label is "E0EC1D83B0760FD83F633623623623623627D89F626B3E27BBE27BFE278F88A4";
    attribute INIT_14 of inst : label is "8E2AFFFFE88C43EA9897D8FB12FB1F621F54EC40EA9D881D53B13E62FFFFEC1F";
    attribute INIT_15 of inst : label is "14721A982E388699769AD10A90D45B66DF1E70B8711BF483C56CD6EB7C3B69C6";
    attribute INIT_16 of inst : label is "FE4F9FF27FFF81C27C9FF3E4F9FE23C7F9327EC5CE07FC1FF07FFDD779A0B4E0";
    attribute INIT_17 of inst : label is "4D150AD50EE85C32A000A1300AB56AC20A22097E67660A19C20883F66882FFFF";
    attribute INIT_18 of inst : label is "D6BADF12D7A18BB74E208E84EF06916C414A02790440AA855AAA0E9BE1D35C7D";
    attribute INIT_19 of inst : label is "B4F8E8EABFAB40EDA9E27BB733B11A143E081A1CD05C5454AB580BD5A8056B5A";
    attribute INIT_1A of inst : label is "C07DF55A468D0294A53C2C662B3788F5EFF7B547D1E9B5F5B775428F057665F5";
    attribute INIT_1B of inst : label is "0A9428C15975E96554CE3F59B50FD6EDAD1E3CC30E3CC3020C000A153D1A1534";
    attribute INIT_1C of inst : label is "B3D4CDCFD47FB7EA5B12F5E8A31B7F3E6CEF9127B9A6DEAB9A65338A65D5CB19";
    attribute INIT_1D of inst : label is "8954055BE2AE89A273DDAEB981C1F35EE058C414E701DB2164A1F444BDBE5AD3";
    attribute INIT_1E of inst : label is "1771C1CADB010060F151BF7719CEE3B5B6C0802008020088400222200AB6BD13";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC5455451A1921A21482000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "985E0EBF7D9F6D6DC3EFB40E675981FDD735DB3D31E182D107DEF0BB27A891FF";
    attribute INIT_23 of inst : label is "B79FCE73E39646CB54BB6C9F3F55D759A4EB2596CC90DA8D554094B573ABB7CE";
    attribute INIT_24 of inst : label is "0A8075AD65D21E50FF97CF61CF21F0566C7FF204D650E9D988D1507783F4C85B";
    attribute INIT_25 of inst : label is "000000001BF3EDEDF6EAAD9E1C730020810800820820010810C5F2EFCF2FFB3E";
    attribute INIT_26 of inst : label is "0A16846A00ADCCEC7D1CE884FE5FFD563801E6F93423EDFEDF77E9C924920000";
    attribute INIT_27 of inst : label is "204242AE5F73F1EA219F8441043FFBEFCDEF2444003272510983DBE076B168E4";
    attribute INIT_28 of inst : label is "19F7E9F1CB5B2C60890D0687632E782EF95B3C68810E5141BA8354B94A6FB8F8";
    attribute INIT_29 of inst : label is "F6A163B3E3D0686632E782D6CCF3C62A14D070CC67DFA7D72D6CB18805341C33";
    attribute INIT_2A of inst : label is "017507A8A17AFB9D9EAA9DD4CEA775171ED038A50652C650A9AA4F11BAAFFEFE";
    attribute INIT_2B of inst : label is "E2D3EEE0B573AD56C0D3F7F3C87127AD22FD8BF14FB2D5CEB55B0AD3F727A922";
    attribute INIT_2C of inst : label is "11ED574DA4A0138C9FFF00FB0D4CC36494A6BBCDB2A714B400400408EB6AF381";
    attribute INIT_2D of inst : label is "37FFC17F31BB0C23E68E0F870944453FF5DF9AD1193AFA2308A5F3996EB8E83E";
    attribute INIT_2E of inst : label is "7C92FFFFD86A998CC52BA688801B0043C1005400CE2FBC84EDF77B9C975B75FD";
    attribute INIT_2F of inst : label is "2D7566CA856CAEA8E856CCBB33B468BD5459D48D6A21FD33AB14DE265A824449";
    attribute INIT_30 of inst : label is "050A205101A0069354C284509D50EBD5450A1D59EC8856C9D59BA15B36EC95B3";
    attribute INIT_31 of inst : label is "48F5A55F4561B58B3434E5324AB5ADF93426D2067F4B5E52BFD5FDADFEDEA010";
    attribute INIT_32 of inst : label is "20B4215B58B3434A64001515E802854406B4A12A0703568F6DAD0E2769D6DFC0";
    attribute INIT_33 of inst : label is "86F8A5011C50A3A428400801002004008014028050022842ADA9E0E596D4F122";
    attribute INIT_34 of inst : label is "28552CC9CA3209BE2B868A55BE2BE9342700EAB755DD105AADD577C2284E81DF";
    attribute INIT_35 of inst : label is "A3C22A95D37549CBB54537C537C537D537D5286B05592B02A7DA1AA8B4B04000";
    attribute INIT_36 of inst : label is "A6C97880242CD82CD2B8EE8974D01E03C26857640029DEA8400005644C0188AA";
    attribute INIT_37 of inst : label is "2476891DA2894B11F4C4820CF89030100804022C08E1F8608102000000080465";
    attribute INIT_38 of inst : label is "81818000000004555322588A440892925722294C2511284875D4D98C86290040";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE080808280838181020103000101000100808183000003000002";
    attribute INIT_3A of inst : label is "2B540222D848CDB15CAB3AD52F5AD6BDFF26A258A60A183A680DAAA31BC3553C";
    attribute INIT_3B of inst : label is "B0E122000813A8409E0AC018341C7EA1B3B1B2C46A22C333733B11A383144AC3";
    attribute INIT_3C of inst : label is "20E2334AF001165940C0D0111E70979521E706F2A3D44CB89C55316ADF089C08";
    attribute INIT_3D of inst : label is "3D77DDE85410D814FC088058808505B82A0C8A5E042E4282FC6066819A62B802";
    attribute INIT_3E of inst : label is "A2AAAC5EB112B176222AA56888AAA6D6224AAB598AD5BABEAF39CE718C79B34D";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFF96CDC4456BC756C3EE565C115D7C6BC4F888895BD155555F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "07A82AF862218C9313AA3987BFEE4C628AB5737FFF9964C1BBFFC281FAA4F184";
    attribute INIT_01 of inst : label is "E01A4DD4555588E6600C17564AC630B5450AD0FEB4CEF2EEEDDD330887265340";
    attribute INIT_02 of inst : label is "8C4158871DB7EE19989F1E328E7663E4A0158073FC009A174008782D160908FB";
    attribute INIT_03 of inst : label is "3B13B1592CC6E992976BD9AE658EBA2158AACA8AD4FABDB0FFFFD4AB0F655115";
    attribute INIT_04 of inst : label is "6E8E8F45049E1600463194F18D345F621BE652A924B77318DCEED993B6524E52";
    attribute INIT_05 of inst : label is "98FFD69F2ADE7C6266B8E8BB34989E44463186858B8B164423B115CA0D5C7D17";
    attribute INIT_06 of inst : label is "00AA802A02808288A208A02A82882A8282208A281F5F7888889660B958E2DD8E";
    attribute INIT_07 of inst : label is "08421084210842108421084212C7CA108421084210842108421084184283FA80";
    attribute INIT_08 of inst : label is "68100097C016D802DA02D8025E004B400B785A20CB42DDFFFF7FD7641934C421";
    attribute INIT_09 of inst : label is "082CDB8025D016E00B6F5405A02D802DA004B6009780B6009781000978012D01";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFF924400184400442010060447F4A1136D2A50848292492";
    attribute INIT_0B of inst : label is "FFFFF4470925941898D1D38AAB10F111978AAB10F119D7B2E39988CD22233324";
    attribute INIT_0C of inst : label is "071BAFBFCB2C2EFCE61E5BAD31F55E3B65663EFCE604305BAC1BBF5BED7C76CC";
    attribute INIT_0D of inst : label is "77178A6A2D23000033A44D1A6A3A875829369AF2479D62D3A1636F7CFFFF8000";
    attribute INIT_0E of inst : label is "7000000000000BEEAF355268D1D5C97F48F463BCFFFEC957A650370452439DE3";
    attribute INIT_0F of inst : label is "050810040000820020820000000830C08A000104151BFFFFFE000008000000B3";
    attribute INIT_10 of inst : label is "00041000040441001000020800A20408430A20200C0000080001041040461440";
    attribute INIT_11 of inst : label is "C30D34D34C30C30C75D75C30E020800000020820000000000220800000410000";
    attribute INIT_12 of inst : label is "0200061A698638E38E38E3AE9A69A69A698618E3863870004000D34D30C30430";
    attribute INIT_13 of inst : label is "70DE1BC3786F0CDC33737737737737737733DCCF732AB733AF733AB733ADCD80";
    attribute INIT_14 of inst : label is "DA45FFFFECDE67FFDCFFFAFB9FFF5F733FFCEE61FF9DCC3FF3B99E73FFFFEE1E";
    attribute INIT_15 of inst : label is "84410E00A80C030BD5154308B0C651C2542D30E3A583CD232478C7AB452336C7";
    attribute INIT_16 of inst : label is "FE4F9FF27FFF81C27C9FF3E4F9FE23C7F9327EC5CE07FC1FF07FA0A288E10C61";
    attribute INIT_17 of inst : label is "0B1998119817B1CE7A4550F2023F7EB9E8C7BB064F41A69FBAA6820651EEFFFF";
    attribute INIT_18 of inst : label is "D6B253F1C440FF3F4F34E6ECE50882088002732188D6B9A45A38829A3053464A";
    attribute INIT_19 of inst : label is "3EC97CB98DBE3E6D88E25119119999110EEA9B18744B37724B5DE9A5888D2B4A";
    attribute INIT_1A of inst : label is "7C6C8112CB3779DEF7AF6794616DDEC9546A39D6F5BAB838313C939408323C3C";
    attribute INIT_1B of inst : label is "D89E2AD11A696946C4451F7DB146DF7D8DFE3CC30E3CC3020C00051D0FB10D07";
    attribute INIT_1C of inst : label is "12E4444B3224BBE25992E969A3196432F50CB76D9DC24F33B2ED1B9839A4D39B";
    attribute INIT_1D of inst : label is "F8C4765A3AB9A0A22371A8A8C182E498825ED4DC56004C33E5A5CD64B1B658D1";
    attribute INIT_1E of inst : label is "ACB179E08980C77293718B078CA8F19FE0E318C6318C69863A200000001639D5";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7401404C10008A08618E0";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "4D9D87C96C89646D43662B0A329D818CF115F88FA9111A49D6CA4F1F6578B9FF";
    attribute INIT_23 of inst : label is "11B265BC3AD3EEE8AB594D36D994E2538E53ECAC6DBC4CCC54649CAF1129F1A3";
    attribute INIT_24 of inst : label is "9FEC7C7B9C8720802F24AB6052DB6816EB0976009D2C88C8CCE9A334E58C4E73";
    attribute INIT_25 of inst : label is "000000006B352424B24289DA5190000000000000000000000000AEB1A224BEB9";
    attribute INIT_26 of inst : label is "71EF666324EC44666C9497ECFF63D2AD3806F691B42D27924B248D8210210000";
    attribute INIT_27 of inst : label is "13E0F6B75B20E0F55646CC08E812CB2EBB575E66F7CB6EDB513DC4CF713964AB";
    attribute INIT_28 of inst : label is "9D61D578ABFE2E35FECF76A333AC3FAF93FEAE3FFECC69A09F03FE518CED90D8";
    attribute INIT_29 of inst : label is "B3FF7198E1F76A333AC3AAFF8A2EE37F6CF77466758755F26FFAB8DD5B3DDD19";
    attribute INIT_2A of inst : label is "05678579A56488889DF888C44723321758FC30A5556ADB59A6E1DBBDA4CAC9C9";
    attribute INIT_2B of inst : label is "92FB6650AF594FE2C4DB3214B6CF657973ECC9C9ED92BD653F8B0EDB33657972";
    attribute INIT_2C of inst : label is "17566D3DA4A0526C9601008B4C44713C9E46A204BA2614BF00000000AECF7A79";
    attribute INIT_2D of inst : label is "1FFFF24D5F96AC2DE36B48A45404557FFCCD7E77F92CBEFE79A7F195692E0FBA";
    attribute INIT_2E of inst : label is "4C91FFFFFA5348C46671C7DD48958A2EC09C6F7FE62CBC8524B24B94BFD7FDB5";
    attribute INIT_2F of inst : label is "2D720247CC788E404CC7A8BE3D3F7CBC6575D044727AD928818E93253A3644D2";
    attribute INIT_30 of inst : label is "A1D73B39D8A363A1FE4A22465B3D8BC657C59C808C7CC78BC809331EA2F8F1E3";
    attribute INIT_31 of inst : label is "4F313F17A47158CEAF44A52A2A3DCF10AF40D3AC36CB92562DEADB896D92A911";
    attribute INIT_32 of inst : label is "59287B158CEAF44A54001151E61364E7632AACB9830347CE4989D9956B0DD736";
    attribute INIT_33 of inst : label is "668EA4691322E24C244688D9132244488911223444D37EC1C989395C84C4909C";
    attribute INIT_34 of inst : label is "40443454ABCFFDA3AA678BC5A3AB983124C0F8B4D57318562D355F20224981EE";
    attribute INIT_35 of inst : label is "5BD26A975B4D4AB5B4753475347534653475746B07502A062757AA89B08EF600";
    attribute INIT_36 of inst : label is "0041800124A0CCA0C599A90522D09E034278574400641159F4038702E4C92F15";
    attribute INIT_37 of inst : label is "941225048801C3198082820CC05030100804021010612858810200000000066C";
    attribute INIT_38 of inst : label is "00000080000000000000000000000000000000000000000000A2800680050C00";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE001000000000000808080818002000003000000818380000001";
    attribute INIT_3A of inst : label is "90650602D86AABB9124B9C7F955AD2B9FF049198ECE43383763C08D8DBEAC5BC";
    attribute INIT_3B of inst : label is "237665914C105060805E6B192ACA3EE89191AAE6630489911119999346140896";
    attribute INIT_3C of inst : label is "BF7C65A37BEDFF7C3E76AFBEA243889B1A24AD12972BA4FEAFF6325508CCAEC1";
    attribute INIT_3D of inst : label is "15D77F808081E001810201E0808101F1600400F880020000F8C4D3D34BF8DFDB";
    attribute INIT_3E of inst : label is "0000080C00000030000008C0000005800000160101800AABFEB5AD6B5AC18604";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFD24575457325C2C08C96DF31CA6263A4F000000180000003";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "94AAA8DC40A519DE5291168A0C990C6442854DBFFE5B1AD380FFAA5AFE6DDAA3";
    attribute INIT_01 of inst : label is "A58D41D050114896C4069502A0AA0036885A8531AD4D7E89CBD804B315069A6A";
    attribute INIT_02 of inst : label is "9CD8099700AB089514943422034409410A74055A4D008A36A00948293C45B1A6";
    attribute INIT_03 of inst : label is "781881D360841936922608982D981929482A884A1562B110FFFFC6AB38055380";
    attribute INIT_04 of inst : label is "02921549001A12AA52B5A26008344F2A2087519B6C9320125585930164D6D074";
    attribute INIT_05 of inst : label is "DA5552DA001566840F20A09B71B10C488802010A950912C44122208A02405813";
    attribute INIT_06 of inst : label is "AAAA8000AA802A82A08288A208A02A80882A8282208A2A828200081511254880";
    attribute INIT_07 of inst : label is "0842108421084210842108421087C2108421084210842108421084000201F82A";
    attribute INIT_08 of inst : label is "180000B08016380242023802C70058E0090CC20048E60A88A208888008000421";
    attribute INIT_09 of inst : label is "4108C1002C3831400B108C047063002C60048C00B0808C00B180000B0C016301";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFEAA8A888A82208A20A28AAA88A28148002844200000000";
    attribute INIT_0B of inst : label is "FFFFF4EC1B7094085109261E7B3AC33B361E7B32C3B1D526EB1589A167762A11";
    attribute INIT_0C of inst : label is "2A1EDAA9542853B4483234D3B0A0AE283E80C3B44C185A34D3522A05A2D45079";
    attribute INIT_0D of inst : label is "98DE0F445B570000042702300A194A012C0802818A4151651063E051FFFF8002";
    attribute INIT_0E of inst : label is "10000000000004056E3D1815811406C558A81C09FF03D554C832650019A09346";
    attribute INIT_0F of inst : label is "2082080010A000000000002002000000000000006FF5FFFFFE00000000000074";
    attribute INIT_10 of inst : label is "4000004100000004004280000000000000010410402080002140000001000000";
    attribute INIT_11 of inst : label is "5144104104104105104104516800000000000000820820808208228A50000000";
    attribute INIT_12 of inst : label is "8000020820A28A28A28A288228A28A28A28A28208A0834100004C30C30C32514";
    attribute INIT_13 of inst : label is "F0DE1BC3786F0DDC37737737737737737737DCDF737FF737FF737FF737FDCDA0";
    attribute INIT_14 of inst : label is "A149FFFFECDE67FFBCFEBFF79FD7FEF33AFCDE61FF9BCC3BF3799EF3FFFFDE1E";
    attribute INIT_15 of inst : label is "0920310100436D102499CF2A32C553CAD41B2471B120004A0644E46E0D2DA5A6";
    attribute INIT_16 of inst : label is "FE4F9FF27FFF81C27C9FF3E4F9FE23C7F9327EC5CE07FC1FF07FDD75D3115181";
    attribute INIT_17 of inst : label is "4991F319F30615ABC84837A00F2346CA503024007883023DE40098404C09FFFF";
    attribute INIT_18 of inst : label is "56B25E2B47AA91A246311489E28932908D84C7118240918C702802B060560448";
    attribute INIT_19 of inst : label is "3CC978BBA0F41F7C89C23BBB3331102076323A1C748F8685AB5D4955C8D1294A";
    attribute INIT_1A of inst : label is "4EC4A50DC3161719C62E24A5216DB6C1527B3C06A1BA3C3C337DD7900C673C3C";
    attribute INIT_1B of inst : label is "1884B08618A1F864C4ED38E1F14F387C8F0E3CC30E3CC3020C0005218C8321A7";
    attribute INIT_1C of inst : label is "B1C4ECC6026CABE23310A1FFA6092C32476D9BA5B9E6DA47926533597585EB1D";
    attribute INIT_1D of inst : label is "98C84470229064BA635320A9CB03B45808608191560283022601000431FCD8F3";
    attribute INIT_1E of inst : label is "1371484F4200C95C993703079988D33040E318C6318C51182000000000173125";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000021104091000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "59108E9B849B6D71C6262000665B0F64C135FA8CA285C765084AC271211291FF";
    attribute INIT_23 of inst : label is "3396CEBA2E9B573C00C90C161025869924CB25A0CE94D08C54490422334BF5A6";
    attribute INIT_24 of inst : label is "C08B02511C92F85BEF570BC19863628D34C932004800899988800135A5996814";
    attribute INIT_25 of inst : label is "000000001B73716E12CA869814500000000000000000000000002361B2749400";
    attribute INIT_26 of inst : label is "50C2C462111ECCCC500B0489FE6F505FC010E6E534237096E123299281090000";
    attribute INIT_27 of inst : label is "0A1044726120A0AAAB5008808036DB6D4ACBA444516A6A57216DECFF7B3160A4";
    attribute INIT_28 of inst : label is "75715369AB04AC60034C06A66AEE2A2DB704AC68834C0013BA035531087091CC";
    attribute INIT_29 of inst : label is "92016330B1406A66AEE2F2C13B6EC60034C064CDD5C54DA6AC13B1822D301933";
    attribute INIT_2A of inst : label is "015201179960D999844C9DE4EE2660040880C025C452FA5F96E7DB6D808A89CD";
    attribute INIT_2B of inst : label is "035424E022032C0F879413E618C321112A0493015090880CB03E0B941321152A";
    attribute INIT_2C of inst : label is "0684CA4DE4201810E7FFFFFBCC4CF36A5896A20DA2380420000000005024CA12";
    attribute INIT_2D of inst : label is "330001755228980F0A5792C96151000005DB9ED529196AA453910311602908C6";
    attribute INIT_2E of inst : label is "1145FFFFDCA6598CC8E5960880230148605214400E2F34846E12330C0A52676D";
    attribute INIT_2F of inst : label is "AE00C6EA2C44E018C2C448B1A98344E8440D448163A334D329124C5A440E91C7";
    attribute INIT_30 of inst : label is "651CAD6523498C49552C1C8180118E84450A0031AEA2C44E031B0B112AC6B112";
    attribute INIT_31 of inst : label is "4991A3180471D481A06461D0AB21C819A074D23B6D831C3E3213A68E9A4D0CE4";
    attribute INIT_32 of inst : label is "D2D1239D481A0643A100D1D101CA67948C4323107401444E4489100F7E937801";
    attribute INIT_33 of inst : label is "0C18A811409288319093122A4449893522A0C40A810400A2748CDEC15A466DA8";
    attribute INIT_34 of inst : label is "2C6EAC1D29AA5302280802C70228074C303868E0156064163805581ED86070D0";
    attribute INIT_35 of inst : label is "94829E1096014887604560C5604560556045008B021002022A903AC224230580";
    attribute INIT_36 of inst : label is "0001FF012CA3C5A6C81674C3A9B0B606C0D840540000C0050400EC3402862924";
    attribute INIT_37 of inst : label is "D2A074A807100400701A5480394A00118804622201811440B162000000000660";
    attribute INIT_38 of inst : label is "0000000000000008880011000020000800112040002080008A0A030A443A5E45";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "68E9A887D82A8DB515ABB655515A529DFF049161DE4EF9347130285071F94781";
    attribute INIT_3B of inst : label is "4F646812249A0124D00EE258649A71D9B339A2C462113333B3B31100083D28ED";
    attribute INIT_3C of inst : label is "6567D38AD0E33349497193D38807A20B708078407D18AC892CCCB0C9D8912C84";
    attribute INIT_3D of inst : label is "1F57DFCDC59BE2E5F1629BE2F2E5E5F16AECFAFAB62E72F2F8EFBA7EE272B1C4";
    attribute INIT_3E of inst : label is "000000040000001000000040000000800000020000810AAABA94A5294A480248";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFF96ECC2754B0503820D8D1E9119606201F000000080000009";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "D0DC82F1755759E85681976EA6637B6065AE84FFFFA0BD0842FC8B13FD00D7AB";
    attribute INIT_01 of inst : label is "952651D51015CCA7D61A78A834BE60A2A170141381AD346FC28907F72DA628BF";
    attribute INIT_02 of inst : label is "D6C14D1E54E118763CB4440442C498004E36314AC510A2BE600BC6EADCB93BAE";
    attribute INIT_03 of inst : label is "B07C051252941325A40480120913404240573236BA623150FFFFD1F4164FAB14";
    attribute INIT_04 of inst : label is "03000580027010FE31AD662820AA90A2059C911249210066178137204D6485E4";
    attribute INIT_05 of inst : label is "A1551B10553345C02E02829870900C0000000000001314C40100028AB8214053";
    attribute INIT_06 of inst : label is "00002AAAAA80002AA02A82A08288A208A02A80882A828208A0028C5300002935";
    attribute INIT_07 of inst : label is "A5294A5294A5294A5294A5294A50294A5294A5294A5294A5294A52AAA954F800";
    attribute INIT_08 of inst : label is "680000978012F0025F06D0025E004BC009785A004BC2E0A0828A0A0AA5555294";
    attribute INIT_09 of inst : label is "00085B0025D0364009720E0DA06D0025F005B40097C1B4009780000978012F83";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFEAAA0022A288A00A22A8A82A2288800000000001000000";
    attribute INIT_0B of inst : label is "FFFFFCA91249248828459694F236D32A7494F236D3A7752EBB63999F4554C60B";
    attribute INIT_0C of inst : label is "2A1A22AB60780193200B02B4FE902665940881932029CB02B5FCE91C9ACCCB2B";
    attribute INIT_0D of inst : label is "55703980B11A00000E640040130AE3A6A001E62012130CCA1A674CD3FFFF8002";
    attribute INIT_0E of inst : label is "B0000000000005503C3450060026810DE9AC005BFF000355974101088490B300";
    attribute INIT_0F of inst : label is "00000000000080080000000000000000000000000050FFFFFE00000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000002002000000000000000000000000041000000000000";
    attribute INIT_11 of inst : label is "4104104104104104104104104020800000000000000000000000000010400400";
    attribute INIT_12 of inst : label is "8200020820828820A20A20828A28828828A20A20A28820100000410410410010";
    attribute INIT_13 of inst : label is "1002004008010004001101101101101101100440111501105411054110444420";
    attribute INIT_14 of inst : label is "B65BFFFFE44220A804415000882A001105400220220044044008801100004202";
    attribute INIT_15 of inst : label is "0082001040401000196B0051054EA204B820A4334200820A0CC14C3001D0AE1E";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000208208000200";
    attribute INIT_17 of inst : label is "743392739245B30B548180A49F61815EF8862000FD36064AE802A0208188FFFE";
    attribute INIT_18 of inst : label is "73B670664D26B04182DBB58BE00000000E104A0004074044C0000D4001A800B0";
    attribute INIT_19 of inst : label is "A4CB5AA056524A4A9952133A222274F001780E184179292939DB597D99037BCE";
    attribute INIT_1A of inst : label is "58091AA12A55B630846915AA00AD3682A6412516E5A130A0A35076880464B4A4";
    attribute INIT_1B of inst : label is "3985BA2B0403687DCCAA21A53389695A9D0F3CC30B2C82030C000A5B7DD64B75";
    attribute INIT_1C of inst : label is "20EC88820C482AE61220836C10036C527C149565B9A6DA659665F3887D8D8B71";
    attribute INIT_1D of inst : label is "B0413CC004C003F66BD0015994620FDC0CC04FA9560820200810830833B5FCD2";
    attribute INIT_1E of inst : label is "027558681821155387181A34196AE324CAC2108421085689B6000000001E3B75";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD000000010000100000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "51204C9B491B6D61004A604866D8044943BD89D96DF3ABC37496D6DD216493FF";
    attribute INIT_23 of inst : label is "3396CF9ECF1DCE9D54522915A645C71964DBE599CD98A11CF4C9842C328A91F4";
    attribute INIT_24 of inst : label is "1988A1B31026AF466DE87B0280C276C0AD5B72069B819911938208358CAB9019";
    attribute INIT_25 of inst : label is "82082082125A484924B5D09D5EE8000000000000000000000005D26592BDBDD0";
    attribute INIT_26 of inst : label is "727249E6DBBE8888A2790D8BFEC1BD4F8010A58F34224924924859CBA5930820";
    attribute INIT_27 of inst : label is "42C7477ED2593937D1EB3466DE269A6A48DB65CAFB3672711B6D04DB413D63EC";
    attribute INIT_28 of inst : label is "754A6D553A4CE855D9EF46864EE94DAAA74CA85559AF0219B8CB55BC6B692CB9";
    attribute INIT_29 of inst : label is "A5D662252A746864EE94DA93394E85771EE670C9D529B554E933A17DC6B99C32";
    attribute INIT_2A of inst : label is "03A6A1648563D9998589916C8B64488649D11C2E1572DAE08680DA6D0395CD89";
    attribute INIT_2B of inst : label is "0E1248AC2C436D9A0422A420309721632EC932864920B10DB6680822A521672E";
    attribute INIT_2C of inst : label is "0995D84FC420100B0A01008FCEC88257DF4FA6097E63843440000000FF4D16B7";
    attribute INIT_2D of inst : label is "F3FFCE8557D5401452CD2F978D55557FF5DB98557F0A8AAEBC81035560FB5988";
    attribute INIT_2E of inst : label is "01C4FFFFCDEED18C9DAD350BB77B76D9CA14CC400B683A84492483AC3256656D";
    attribute INIT_2F of inst : label is "AF2076F98CC7640EF8CC56B159828508088A969B6723A41E3B324863CE05D0A7";
    attribute INIT_30 of inst : label is "AB18E9C34D61345955CE95D0A0B198808D1A281D8F98CC7481DBE3315AC55314";
    attribute INIT_31 of inst : label is "5B9BE7348EF1FD91CC78211CD66298EBCC7F7623A90330127137249AD2498A30";
    attribute INIT_32 of inst : label is "607723BFD91CC782390093D342EADF0D34D78140BE024C56E49F105778B25C0B";
    attribute INIT_33 of inst : label is "10011C05804A900303C2784F09E13C0784749E83D22668E644DC84D3C26E4963";
    attribute INIT_34 of inst : label is "394CEE18290AE8004C14424C004D03AFA01C29802660821260099A071F403858";
    attribute INIT_35 of inst : label is "B0430208E002624F0019800880098009800991088800400A72E6340C10504400";
    attribute INIT_36 of inst : label is "03490000ECE2C0E2C4292E95E0104208410808088010A40944004C38CC922B6C";
    attribute INIT_37 of inst : label is "810860420000101000A039880206231088C42200100000001122000000000562";
    attribute INIT_38 of inst : label is "0000000000000000000800000000004880000000800000000002000000403F01";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "484010C0FA59ABB9313B45D572DE77BFFF4DC802C4C1530D6272D55C8D6C4CC3";
    attribute INIT_3B of inst : label is "2164A12071371189B818525C6C984141B2253AC9E6488332A222274C1010C9D4";
    attribute INIT_3C of inst : label is "656657351CC333CEC961B313488CCA21AA88C9446530BE89ACC4B8D90019AC92";
    attribute INIT_3D of inst : label is "1FFD5FE9C1D3E0C5F872D3E2E0C1C1E870EEE2F4B70F62E0F444A292866D4186";
    attribute INIT_3E of inst : label is "000000040000001000000040000000800000020000800EEEEA10842108400200";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFB6CDD4EFDB0F0E042EC099119B60E60BF000000080000001";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "83FF90FC6AA08CE813821D0376E0086087BFD2FFFFD17E9141FCE1E8F9C5F29E";
    attribute INIT_01 of inst : label is "C091BCD5401341D2404FFE56466C20E1C5D04C98900FB408A48490A7E71669AA";
    attribute INIT_02 of inst : label is "9CD73981F3BC6CDDD41F0C139872086422059420702241170004F224165491C1";
    attribute INIT_03 of inst : label is "211F338B69C6D9B6B67259C96DCE28E7D82FCBFEFFF87C11FFFFD8AA00655373";
    attribute INIT_04 of inst : label is "26080D040C82362AD6B5B2FB26BEDB43B4E4488B6DB77672DDEDB19B6CC6DCC6";
    attribute INIT_05 of inst : label is "D0AAC6392A987CB24E8888BC3DBCC324449932650A311C472699116785144517";
    attribute INIT_06 of inst : label is "00000000002AAAAAA0002AA02A82A08288A208A02A808AA0A81B40AFCCC2970D";
    attribute INIT_07 of inst : label is "000000000000000000000000000000000000000000000000000000000000F800";
    attribute INIT_08 of inst : label is "1800009080121002460230024200484009084600484200AA02A00AA000000000";
    attribute INIT_09 of inst : label is "00084700243011C0090AA4046023002420048C0090808C009080000908012101";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFE82202008000028A8002200082A8000000000000000000";
    attribute INIT_0B of inst : label is "FFFFF8448B65B458983042582310C91116582318C91193C2C3D980C02223B324";
    attribute INIT_0C of inst : label is "0E09E40C5F319C4892004BEC3048D21341E10C48962DC84BED133C9263742686";
    attribute INIT_0D of inst : label is "7F333860EC360000339648884E6184F821223832297CA2027320470CFFFF8000";
    attribute INIT_0E of inst : label is "400000000000055574121244409CC93048344226FF07440671C5B019CF461C21";
    attribute INIT_0F of inst : label is "1861871C71410410638E38E38C30E38E30C30E389005FFFFFE000000000000D0";
    attribute INIT_10 of inst : label is "C61861861C71C71C71C50410610C38E30E30E38C38E30E38E2830C20C71C71C6";
    attribute INIT_11 of inst : label is "61871C61861C71861871871850610418E38E38E38E38E38C30C30C30A0820831";
    attribute INIT_12 of inst : label is "8610638C30E38E38C30E38E38E30E38C30C38E38C38C2820820C71C71C71C318";
    attribute INIT_13 of inst : label is "1002004008010004001101101101101101100440111541105411054110544441";
    attribute INIT_14 of inst : label is "4524FFFFE4422002844005508800A81100140220088044011008801100004202";
    attribute INIT_15 of inst : label is "1F663F31BC9FEF325454651E51C27146DE246D9C7980C921240AC0A902723241";
    attribute INIT_16 of inst : label is "00000000000000000000000000000000000000000000000000002A02A3F27DF3";
    attribute INIT_17 of inst : label is "DF70987098640D237604A4320E054AE328C39106376E0000F908F27210E4FFFE";
    attribute INIT_18 of inst : label is "D6BAF989E0F94224598640E6EF9BE6F981EFB5F20941D8A408080FC805F9027C";
    attribute INIT_19 of inst : label is "B26130E80B8B633180D0C999111DD99108888A08087D0503EB58EB858EAD6B5A";
    attribute INIT_1A of inst : label is "632DF55342844CF6BDECC67EA24180CDEF77B2C2308CB6B6B1745666022232B2";
    attribute INIT_1B of inst : label is "C8330859034D2327404613109085C421840F3CD30B2C920F3CD308131AAC0310";
    attribute INIT_1C of inst : label is "16404459242C81A0C1D64D200B036D14E445B12DB5B2C998B0EC0BA821C4B3D7";
    attribute INIT_1D of inst : label is "42430C08131903F221C080F885E2471E1A48B48C4623DE6455E1487590936941";
    attribute INIT_1E of inst : label is "29E06324D38116100B18DBB708CAE11B62C4310C4310FD8F0C000000001A5081";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001E21CDEF2000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "9ED985DB2D8B6D64016E1F36321D8CEDD13DD09F274F83CDD2DEDD836C09B9FF";
    attribute INIT_23 of inst : label is "11B6C4309A7E7662AB1BACB65991A24B2E432C8C2CB85ECC0C3631811123A1A7";
    attribute INIT_24 of inst : label is "0CE4B90994A3FD87CEF48362C2797E12FB5B6603653C8088EEC93690C1B9CEC2";
    attribute INIT_25 of inst : label is "000020005B7B676CB6EAA9581410000000000000000000000000ACF5863DB299";
    attribute INIT_26 of inst : label is "1B1B3761966244475CC5B0E6FFA8BBA000067294B42B65B6CB74A583A1010020";
    attribute INIT_27 of inst : label is "3871F1B94B6C8C8A0905EC3C3316DB6D98432F74512966F90F01FAC07FB164F7";
    attribute INIT_28 of inst : label is "336129709BB66E20A90CB242262C252E91B66E20094DC930BF62ABB7BDE5B6AE";
    attribute INIT_29 of inst : label is "360B7110810B242262C252ED9826E28094CB2844CD84A5D22ED8B8A2A432CA11";
    attribute INIT_2A of inst : label is "07D90C0C816488C8B03808C046023330987C219F844AC1FA8022030184EFC545";
    attribute INIT_2B of inst : label is "98B96C5181B90E70C679B7B09E5D6C0D7B6DE14CE5B606E439C30079B76C097A";
    attribute INIT_2C of inst : label is "304623DE818052459F31388D040461709806E105A204319F0000000000B320EC";
    attribute INIT_2D of inst : label is "0BFFFB4818956C6CAB397C3E501110400CCBBA018B65903004819111613C4E10";
    attribute INIT_2E of inst : label is "DE38FFFFEF3988C47319E67E6CC5CC3571C267002E0CB4856CB74B4584C2EC64";
    attribute INIT_2F of inst : label is "2DB2226EF408B6446F4088B2AD644898271530487278DB288B8CB3053A225452";
    attribute INIT_30 of inst : label is "91C3BB1DD8A363A2AAA22044121C818277CF8C89AEEF4088C889BD0222CAD02A";
    attribute INIT_31 of inst : label is "0430B9033420F5C2A7158C2B5E0781F0A712E38516D906C30C88DBC36DB28591";
    attribute INIT_32 of inst : label is "6908790F5C2A71585600307864030677631888190300E08C0BC1C907210DC724";
    attribute INIT_33 of inst : label is "4204E4419260C2486646C8D91B23646C8D91322446913E118B83214C25C19234";
    attribute INIT_34 of inst : label is "6C26245909230481324319408131901024819C109DD218CA042773202049032E";
    attribute INIT_35 of inst : label is "498664311909C071902710271026102710266620204108271B538A1981BCF200";
    attribute INIT_36 of inst : label is "00010002AE61C261C3BDFBA1F2C198330460310700685554F00325066A4B0C13";
    attribute INIT_37 of inst : label is "7EF79FBDEF31EF31F91FC610FDF84021100C463F31F27CD92246000000000450";
    attribute INIT_38 of inst : label is "000000000000000000000020200000000000040000000000AAA8AA9BCC3FC090";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "F9824781780C89BB0BEB4AAAFB5AD6B1FF3EA3C0D467D19C66CFAAE889B3C026";
    attribute INIT_3B of inst : label is "785234852073C1039C4A090302482420911082F76125E1119111DD9A46225856";
    attribute INIT_3C of inst : label is "1052612B2A388414241C08D92804C201A0804C40660269640A32060400440A49";
    attribute INIT_3D of inst : label is "60000FC9CD93E4CDF36493E6E6CDCDF364CCE4F9266E64E4F914E59393EACC71";
    attribute INIT_3E of inst : label is "0000001C00000070000001C00000038000000E000380305056739CE739C00E00";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFF6C775E54337CEC4AE12DD50C8736136F000000380000007";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "07FF90F0600180681101150322E0104047BFC87FFF807C1043FCC1A1F9C1F1BA";
    attribute INIT_01 of inst : label is "0040A8C000174542800FFE54244420C34D80D9DD384FB04D6E0DB0172234E380";
    attribute INIT_02 of inst : label is "08551098F1300415141A2C02082000E0201800002032E384000CE22E483008C7";
    attribute INIT_03 of inst : label is "733D138921CEC89213721DC864CE28EF982F89FE7F904810FFFFCCAA14255151";
    attribute INIT_04 of inst : label is "66181D0C0C1226004210B0FB249E4A433447588924937670DDECA3BB28E24CE2";
    attribute INIT_05 of inst : label is "00AA8220AA892C76059898946D2DA32CCC9B366C182308C3679B316D8F3C4F12";
    attribute INIT_06 of inst : label is "00000000000000000AAAAAA0002AA02A82A08288A208A2AA001A002FDD861709";
    attribute INIT_07 of inst : label is "AD2B4AD2B4AD2B4AD2B4AD2B4AD2AB4AD2B4AD2B4AD2B4AD2B4AD2AAA954F800";
    attribute INIT_08 of inst : label is "680000968012D0025A02D0025A004B4009685A004B42CA0002AAA00AA55552B4";
    attribute INIT_09 of inst : label is "00085B0025B016C0096AAC05A02D0025A004B4009680B4009680000968012D01";
    attribute INIT_0A of inst : label is "FFFFFFFFFFFFFFFFFFE820000080000002000020002808000000000000000000";
    attribute INIT_0B of inst : label is "FFFFF044893C9418482822CC7112491132C821124993B106491580AC23222B10";
    attribute INIT_0C of inst : label is "AE08B40A5A239A245A08EF302328EA082B418A245A35C8EF3111129521941050";
    attribute INIT_0D of inst : label is "E4733820B20400002B57C4A82A20F0D427121471296A91023220028AFFFFAAAA";
    attribute INIT_0E of inst : label is "200000000000055564121E254055C5A9483C2A12FF05000571C1D219CF220825";
    attribute INIT_0F of inst : label is "0000010410020A288082082082080000002002080444FFFFFE00000000000080";
    attribute INIT_10 of inst : label is "410000400400410400400A288280082080002080002082082045144100000001";
    attribute INIT_11 of inst : label is "41441451041041041451041040820A2800020800820000800820820811451050";
    attribute INIT_12 of inst : label is "8A20A28820A20828A28820820828A28820828A28A28A20510414514514514010";
    attribute INIT_13 of inst : label is "9012024048090104041141141141141141140450115541145411454114544522";
    attribute INIT_14 of inst : label is "448AFFFFE4522000244005048800A09100001220000244000048A09100005202";
    attribute INIT_15 of inst : label is "0000001000400003545A255E51C271464E346C997501C401042AC2AD007A2B61";
    attribute INIT_16 of inst : label is "00000000000000000000000000000000000000000000000000002AA800000000";
    attribute INIT_17 of inst : label is "5F70A870A86405237400A0200E146890B88100383D2E0020D908FE700040FFFE";
    attribute INIT_18 of inst : label is "529A7D40C0C12A344882A040E0080200800000010D41F80428080FE805FD007C";
    attribute INIT_19 of inst : label is "92C070802989416380C04999991158B028580A0C08350506C949A91488B5294A";
    attribute INIT_1A of inst : label is "53A4F00B02042ED7BDE4453EA2E49241CB259646318592929120026E06222292";
    attribute INIT_1B of inst : label is "8811580B084121AC40461711D084C463848F3CC30B2C82030C000A133B360330";
    attribute INIT_1C of inst : label is "12404449142583A0411341210D012516E445B10C9CB25820B2CC39A824C49952";
    attribute INIT_1D of inst : label is "26430C280AB883F223C280F886E1424E0068450CCC0000054680C4C4D0904841";
    attribute INIT_1E of inst : label is "39A05126D61F07108A1AD1A308CA6119624010800108348D0400000015521051";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000004001000000";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "081807C9E4C9273405261A36324E8EE4801C801725CF82A51E4E5407641B35FF";
    attribute INIT_23 of inst : label is "11B26492925427CAAA89A43249B0E2CB0E490C84E43848AC0C0090C311610082";
    attribute INIT_24 of inst : label is "0440F5188361DDCFC4E281A34E103E3BCC5136036C6880888AC506B0C4A08647";
    attribute INIT_25 of inst : label is "8000008049293F27926005C8145000000000000000000000000205B492289638";
    attribute INIT_26 of inst : label is "1A0A856092A266445C4E8840FFEC23D78006D65194293C9279228C8285810000";
    attribute INIT_27 of inst : label is "1420A1B9792585888154A41413124925D8490D4400232CF907249649259122E2";
    attribute INIT_28 of inst : label is "31232B3099966620A944B642262465669196262AA104C5109F22AB9294FC92A0";
    attribute INIT_29 of inst : label is "12293111830B642262465665982662AA90597864C48CACD22658988004165E11";
    attribute INIT_2A of inst : label is "07DB061C81208888907808C046023011B868E8DF845A49FA82224924808FA323";
    attribute INIT_2B of inst : label is "81FF2448C3B926C1437F9353841564186BA4A1C1FC930EE49B05017F9364186A";
    attribute INIT_2C of inst : label is "10C5139CA0C05E25FFC1E08944046132920661048A1D10DA0000000000B7A0A5";
    attribute INIT_2D of inst : label is "39FFEA2814803422AAAF6FB7C15100000CC9B0014320D0291C83D111203A4558";
    attribute INIT_2E of inst : label is "5A28FFFFEC6008C444008272244E445500A0223024269085279229048EC2CC2C";
    attribute INIT_2F of inst : label is "24F02266442A9E046442A89AAD3468D80451300922D059E8860D923D3E02D040";
    attribute INIT_30 of inst : label is "0086A93502E90A92AA9610C210088580468D1C08A66442A9C089910AA26AD0AA";
    attribute INIT_31 of inst : label is "0230910B0420630A220486E95E1785F42200C11D524D0E420E9459832D9384B4";
    attribute INIT_32 of inst : label is "60A4510630A2204DD2003870E24286D40A9584389100E28C39808887A70CC312";
    attribute INIT_33 of inst : label is "2A00AC01F0408E0072D25A0B48612C2584B09612C24334128983218424C19212";
    attribute INIT_34 of inst : label is "4000042909228E80AA2E8D4280AB89743C4898505451746A14151712E8789126";
    attribute INIT_35 of inst : label is "AD40A0051D054029D015500550155005500560A0014028061D510A0A90B8A000";
    attribute INIT_36 of inst : label is "91490002A4218021812FCFA15B60AC1582B0070400400552A0020006290D0A29";
    attribute INIT_37 of inst : label is "0000000000100000008000000000001008000000000000008100000000000540";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000004000000";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "B1012A00784C999B0EC96AAAE24A5291FF0D90C09423909846CB802089134020";
    attribute INIT_3B of inst : label is "28403000207181038C00000204482C249111C2456000A9919911158A0A01585B";
    attribute INIT_3C of inst : label is "0042A221A8100414400810512004C001A00054006A100B2088100C0800088800";
    attribute INIT_3D of inst : label is "80000C0002000102018300010306060183000100403003030095439501E86822";
    attribute INIT_3E of inst : label is "0400028408880A1044400241110000814420020504814055039CE739CE71B38D";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFF24585E54917CF47A63BCD5049316112F444440482000001";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
