library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity stargate_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of stargate_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7E",X"D0",X"0C",X"7E",X"D0",X"0C",X"7E",X"D2",X"C8",X"7E",X"D0",X"3A",X"8E",X"BF",X"10",X"10",
		X"8E",X"D0",X"04",X"5F",X"EB",X"A4",X"31",X"29",X"10",X"8C",X"F0",X"00",X"25",X"F6",X"E7",X"88",
		X"B2",X"12",X"BD",X"01",X"57",X"8E",X"D0",X"58",X"86",X"01",X"BD",X"01",X"30",X"96",X"F8",X"26",
		X"06",X"96",X"36",X"10",X"26",X"00",X"8C",X"7E",X"D2",X"C8",X"34",X"12",X"8E",X"9C",X"3B",X"AE",
		X"84",X"27",X"13",X"9C",X"3F",X"27",X"F8",X"A6",X"05",X"81",X"02",X"27",X"F2",X"81",X"01",X"27",
		X"EE",X"BD",X"00",X"EE",X"20",X"E9",X"35",X"92",X"96",X"36",X"A7",X"47",X"6F",X"48",X"6F",X"49",
		X"96",X"36",X"A1",X"47",X"27",X"19",X"A7",X"47",X"96",X"F8",X"81",X"50",X"26",X"05",X"BD",X"D2",
		X"2D",X"20",X"0C",X"BD",X"01",X"57",X"B6",X"00",X"00",X"8E",X"D0",X"C3",X"BD",X"01",X"19",X"96",
		X"57",X"84",X"08",X"A1",X"48",X"27",X"16",X"A7",X"48",X"27",X"12",X"96",X"F8",X"81",X"10",X"27",
		X"0C",X"BD",X"01",X"57",X"B6",X"00",X"00",X"8E",X"D2",X"C8",X"BD",X"01",X"19",X"96",X"57",X"84",
		X"40",X"A1",X"49",X"27",X"16",X"A7",X"49",X"27",X"12",X"96",X"F8",X"81",X"40",X"27",X"0C",X"BD",
		X"01",X"57",X"B6",X"00",X"00",X"8E",X"D2",X"37",X"BD",X"01",X"19",X"86",X"02",X"8E",X"D0",X"60",
		X"7E",X"00",X"A8",X"86",X"50",X"97",X"F8",X"86",X"FF",X"97",X"91",X"BD",X"D0",X"3A",X"BD",X"13",
		X"BD",X"BD",X"08",X"3A",X"BD",X"1F",X"69",X"BD",X"5F",X"DE",X"BD",X"19",X"43",X"D5",X"B9",X"BD",
		X"D2",X"2D",X"DE",X"3F",X"96",X"36",X"A7",X"4B",X"86",X"02",X"97",X"68",X"86",X"08",X"A7",X"4A",
		X"8E",X"14",X"AC",X"BD",X"D2",X"19",X"8E",X"3E",X"E0",X"86",X"17",X"BD",X"70",X"52",X"8E",X"35",
		X"E8",X"86",X"18",X"BD",X"70",X"52",X"86",X"7B",X"8E",X"2B",X"CC",X"BD",X"70",X"52",X"8E",X"33",
		X"C0",X"86",X"7C",X"BD",X"70",X"52",X"8E",X"CC",X"02",X"BD",X"14",X"1A",X"ED",X"48",X"F6",X"CC",
		X"15",X"C4",X"0F",X"27",X"02",X"6F",X"49",X"E6",X"49",X"26",X"05",X"8E",X"38",X"58",X"20",X"0F",
		X"8E",X"59",X"58",X"1F",X"98",X"C6",X"02",X"BD",X"D1",X"BD",X"A6",X"48",X"8E",X"19",X"58",X"C6",
		X"01",X"BD",X"D1",X"BD",X"96",X"36",X"81",X"01",X"27",X"0B",X"BD",X"D2",X"0B",X"86",X"0A",X"8E",
		X"D1",X"55",X"7E",X"00",X"A8",X"C6",X"01",X"8E",X"35",X"14",X"86",X"7F",X"BD",X"70",X"58",X"96",
		X"36",X"81",X"02",X"25",X"04",X"A6",X"49",X"26",X"02",X"A6",X"48",X"5F",X"8D",X"78",X"86",X"80",
		X"8E",X"D1",X"76",X"7E",X"00",X"A8",X"96",X"36",X"81",X"02",X"25",X"27",X"BD",X"D2",X"0B",X"86",
		X"0A",X"8E",X"D1",X"87",X"7E",X"00",X"A8",X"C6",X"02",X"8E",X"35",X"14",X"86",X"7F",X"BD",X"70",
		X"58",X"E6",X"48",X"96",X"36",X"81",X"04",X"25",X"06",X"6D",X"49",X"27",X"02",X"E6",X"49",X"1F",
		X"98",X"8D",X"43",X"6A",X"4A",X"10",X"27",X"01",X"1F",X"96",X"36",X"A1",X"4B",X"27",X"06",X"A7",
		X"4B",X"86",X"08",X"A7",X"4A",X"86",X"80",X"8E",X"D1",X"44",X"7E",X"00",X"A8",X"34",X"12",X"86",
		X"80",X"BD",X"70",X"58",X"E6",X"E4",X"AE",X"61",X"30",X"88",X"18",X"86",X"81",X"BD",X"70",X"58",
		X"AE",X"61",X"30",X"88",X"28",X"86",X"82",X"BD",X"70",X"58",X"AE",X"61",X"30",X"88",X"38",X"86",
		X"83",X"BD",X"70",X"58",X"35",X"92",X"B7",X"BD",X"DE",X"B7",X"BD",X"E0",X"34",X"04",X"C6",X"0A",
		X"3D",X"F7",X"BD",X"E1",X"35",X"04",X"F7",X"BE",X"1D",X"F7",X"BE",X"1F",X"86",X"0A",X"3D",X"F7",
		X"BE",X"20",X"BD",X"1E",X"35",X"BD",X"1E",X"CB",X"7E",X"1D",X"F7",X"CC",X"00",X"00",X"8D",X"D6",
		X"8E",X"2E",X"13",X"CC",X"3D",X"08",X"7E",X"13",X"B9",X"34",X"10",X"8E",X"CC",X"00",X"BD",X"14",
		X"1C",X"5D",X"27",X"07",X"AE",X"E4",X"86",X"84",X"BD",X"70",X"52",X"35",X"90",X"8E",X"3E",X"40",
		X"D6",X"36",X"86",X"7A",X"7E",X"70",X"58",X"86",X"40",X"97",X"F8",X"86",X"FF",X"97",X"91",X"BD",
		X"D0",X"3A",X"86",X"01",X"BD",X"5F",X"EA",X"BD",X"13",X"BD",X"8E",X"0E",X"10",X"CC",X"08",X"01",
		X"BD",X"D6",X"5D",X"DE",X"3F",X"86",X"85",X"8E",X"40",X"44",X"BD",X"70",X"58",X"8E",X"CC",X"24",
		X"BD",X"14",X"1C",X"4F",X"1F",X"02",X"BD",X"14",X"1C",X"86",X"86",X"BD",X"70",X"58",X"CC",X"11",
		X"11",X"DD",X"D3",X"CC",X"44",X"44",X"DD",X"D5",X"CC",X"77",X"77",X"DD",X"D7",X"CC",X"33",X"8F",
		X"BD",X"19",X"8F",X"8E",X"14",X"CA",X"BD",X"D2",X"19",X"8E",X"3E",X"E0",X"BD",X"D2",X"30",X"BD",
		X"19",X"43",X"D5",X"B9",X"BD",X"19",X"43",X"D5",X"D6",X"BD",X"19",X"43",X"1C",X"CF",X"DE",X"3F",
		X"CC",X"10",X"40",X"ED",X"47",X"6A",X"48",X"27",X"18",X"6A",X"47",X"27",X"08",X"86",X"3C",X"8E",
		X"D2",X"A5",X"7E",X"00",X"A8",X"96",X"57",X"84",X"40",X"27",X"06",X"86",X"01",X"A7",X"47",X"20",
		X"EC",X"96",X"36",X"27",X"03",X"7E",X"D0",X"C3",X"86",X"FF",X"97",X"91",X"86",X"66",X"97",X"DE",
		X"86",X"10",X"97",X"F8",X"BD",X"D0",X"3A",X"4F",X"8E",X"D2",X"E1",X"BD",X"01",X"19",X"7E",X"00",
		X"E4",X"8E",X"9C",X"26",X"6F",X"80",X"8C",X"9C",X"36",X"25",X"F9",X"BD",X"70",X"28",X"BD",X"13",
		X"BD",X"BD",X"19",X"72",X"BD",X"19",X"43",X"D5",X"B9",X"86",X"8A",X"BD",X"70",X"55",X"8E",X"D4",
		X"4A",X"4F",X"BD",X"01",X"19",X"86",X"AA",X"97",X"10",X"8E",X"CD",X"64",X"BD",X"14",X"0B",X"30",
		X"1C",X"81",X"3A",X"26",X"05",X"8C",X"CD",X"3E",X"24",X"F2",X"30",X"02",X"34",X"10",X"8E",X"0E",
		X"47",X"86",X"31",X"BD",X"70",X"31",X"86",X"5C",X"BD",X"70",X"31",X"30",X"89",X"03",X"00",X"10",
		X"8E",X"CD",X"3E",X"1E",X"12",X"BD",X"14",X"0B",X"1E",X"12",X"BD",X"70",X"31",X"10",X"AC",X"E4",
		X"23",X"F1",X"30",X"89",X"02",X"00",X"10",X"8E",X"CD",X"66",X"CE",X"70",X"55",X"BD",X"D4",X"56",
		X"30",X"89",X"05",X"00",X"86",X"5B",X"BD",X"70",X"31",X"10",X"8E",X"CD",X"38",X"C6",X"03",X"1E",
		X"12",X"BD",X"14",X"0B",X"1E",X"12",X"BD",X"70",X"31",X"5A",X"26",X"F3",X"86",X"5C",X"BD",X"70",
		X"31",X"DE",X"3F",X"86",X"02",X"A7",X"47",X"CC",X"0C",X"56",X"ED",X"4A",X"10",X"8E",X"CD",X"6E",
		X"10",X"AF",X"4C",X"86",X"0D",X"A7",X"4E",X"7E",X"D3",X"A3",X"DE",X"3F",X"86",X"01",X"A7",X"47",
		X"CC",X"0C",X"D0",X"ED",X"4A",X"10",X"8E",X"CF",X"9E",X"10",X"AF",X"4C",X"86",X"02",X"A7",X"4E",
		X"7E",X"D3",X"A3",X"86",X"03",X"A7",X"49",X"0F",X"11",X"A6",X"4E",X"A7",X"48",X"86",X"01",X"8E",
		X"D3",X"B5",X"7E",X"00",X"A8",X"96",X"10",X"8B",X"11",X"81",X"88",X"23",X"02",X"86",X"11",X"97",
		X"10",X"AE",X"4A",X"E6",X"47",X"86",X"8B",X"BD",X"70",X"4F",X"10",X"AE",X"4C",X"C6",X"03",X"1E",
		X"12",X"BD",X"14",X"0B",X"1E",X"12",X"BD",X"70",X"2B",X"5A",X"26",X"F3",X"AE",X"4A",X"30",X"89",
		X"0E",X"00",X"CE",X"70",X"4F",X"BD",X"D4",X"56",X"DE",X"3F",X"10",X"AE",X"4C",X"31",X"2E",X"10",
		X"AF",X"4C",X"AE",X"4A",X"30",X"07",X"AF",X"4A",X"A6",X"47",X"8B",X"01",X"19",X"A7",X"47",X"6A",
		X"48",X"26",X"AA",X"30",X"89",X"30",X"00",X"86",X"07",X"E6",X"4E",X"3D",X"50",X"30",X"85",X"AF",
		X"4A",X"6A",X"49",X"26",X"94",X"10",X"8C",X"CF",X"AC",X"10",X"23",X"FF",X"6D",X"BD",X"19",X"43",
		X"D5",X"D6",X"DE",X"3F",X"86",X"08",X"A7",X"47",X"6A",X"47",X"27",X"08",X"86",X"3C",X"8E",X"D4",
		X"28",X"7E",X"00",X"A8",X"86",X"78",X"A7",X"47",X"96",X"57",X"84",X"08",X"27",X"4F",X"6A",X"47",
		X"27",X"4B",X"86",X"1E",X"8E",X"D4",X"38",X"7E",X"00",X"A8",X"8E",X"0E",X"10",X"CC",X"0A",X"01",
		X"BD",X"D6",X"5D",X"7E",X"00",X"E4",X"34",X"20",X"1E",X"12",X"BD",X"14",X"0B",X"BD",X"14",X"1C",
		X"1E",X"12",X"84",X"0F",X"26",X"07",X"5D",X"26",X"04",X"86",X"8D",X"20",X"0C",X"34",X"20",X"1F",
		X"02",X"86",X"8C",X"AD",X"C4",X"35",X"20",X"86",X"3F",X"34",X"02",X"1E",X"12",X"BD",X"14",X"0B",
		X"BD",X"14",X"1C",X"1E",X"12",X"1F",X"02",X"35",X"02",X"AD",X"C4",X"35",X"A0",X"BD",X"D0",X"3A",
		X"86",X"20",X"97",X"F8",X"86",X"01",X"BD",X"5F",X"EA",X"BD",X"13",X"BD",X"BD",X"19",X"43",X"D5",
		X"B9",X"6F",X"4D",X"BD",X"E0",X"06",X"27",X"07",X"8E",X"D5",X"6F",X"6C",X"4D",X"20",X"03",X"8E",
		X"CC",X"36",X"AF",X"47",X"8E",X"CC",X"9A",X"C6",X"20",X"BD",X"D5",X"A1",X"AF",X"49",X"86",X"19",
		X"A7",X"4B",X"A7",X"4C",X"86",X"AA",X"97",X"10",X"0F",X"11",X"AE",X"47",X"A6",X"4D",X"27",X"04",
		X"A6",X"80",X"20",X"03",X"BD",X"14",X"0B",X"AF",X"47",X"AE",X"49",X"BD",X"70",X"31",X"AF",X"49",
		X"6A",X"4B",X"27",X"08",X"86",X"03",X"8E",X"D4",X"CA",X"7E",X"00",X"A8",X"A6",X"4C",X"27",X"14",
		X"6F",X"4C",X"86",X"19",X"A7",X"4B",X"8E",X"CC",X"9C",X"C6",X"30",X"BD",X"D5",X"A1",X"AF",X"49",
		X"0F",X"11",X"20",X"E0",X"BD",X"19",X"43",X"D6",X"2F",X"8E",X"0E",X"58",X"CC",X"01",X"02",X"BD",
		X"D6",X"5D",X"86",X"28",X"8E",X"D5",X"1A",X"7E",X"00",X"A8",X"BD",X"D0",X"3A",X"0F",X"26",X"BD",
		X"19",X"43",X"D5",X"B9",X"BD",X"19",X"43",X"D5",X"D6",X"86",X"17",X"8E",X"34",X"98",X"BD",X"70",
		X"58",X"86",X"18",X"8E",X"25",X"A8",X"BD",X"70",X"58",X"8E",X"3A",X"BC",X"BD",X"D2",X"30",X"86",
		X"7B",X"8E",X"28",X"CC",X"BD",X"70",X"52",X"86",X"7C",X"8E",X"30",X"D4",X"BD",X"70",X"52",X"86",
		X"28",X"8E",X"D5",X"57",X"7E",X"00",X"A8",X"AE",X"C8",X"11",X"31",X"89",X"88",X"24",X"86",X"07",
		X"97",X"2F",X"86",X"99",X"BD",X"D7",X"0F",X"86",X"FF",X"8E",X"DA",X"00",X"7E",X"00",X"A8",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",
		X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"3D",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"3F",X"20",X"20",X"20",X"20",
		X"20",X"86",X"25",X"6D",X"4D",X"26",X"0F",X"BD",X"14",X"0B",X"81",X"10",X"24",X"02",X"86",X"10",
		X"81",X"3C",X"23",X"02",X"86",X"3C",X"1F",X"01",X"39",X"6C",X"47",X"A6",X"47",X"84",X"07",X"8E",
		X"D5",X"CE",X"A6",X"86",X"97",X"30",X"86",X"05",X"8E",X"D5",X"B9",X"7E",X"00",X"A8",X"07",X"87",
		X"FF",X"FF",X"C7",X"C7",X"FF",X"FF",X"8E",X"D6",X"07",X"AF",X"47",X"AE",X"47",X"10",X"8E",X"9C",
		X"27",X"A6",X"80",X"26",X"05",X"8E",X"D6",X"07",X"20",X"F7",X"A7",X"A0",X"10",X"8C",X"9C",X"2F",
		X"26",X"EF",X"AE",X"47",X"30",X"01",X"A6",X"84",X"26",X"03",X"8E",X"D6",X"07",X"AF",X"47",X"86",
		X"03",X"8E",X"D5",X"DB",X"7E",X"00",X"A8",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",
		X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",X"CA",X"C0",X"D0",X"98",X"38",X"33",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",
		X"D6",X"4D",X"BD",X"07",X"EC",X"84",X"0F",X"A6",X"86",X"97",X"26",X"86",X"05",X"8E",X"D6",X"43",
		X"7E",X"00",X"A8",X"0F",X"26",X"86",X"03",X"8E",X"D6",X"2F",X"7E",X"00",X"A8",X"07",X"0F",X"17",
		X"1E",X"25",X"2C",X"2B",X"2A",X"28",X"60",X"D0",X"C0",X"C3",X"85",X"47",X"87",X"AF",X"C8",X"11",
		X"A7",X"48",X"E7",X"C8",X"14",X"35",X"10",X"AF",X"C8",X"15",X"8E",X"D8",X"2D",X"AF",X"4F",X"6F",
		X"C8",X"13",X"AE",X"4F",X"10",X"AE",X"81",X"27",X"14",X"A6",X"80",X"ED",X"49",X"A6",X"80",X"A7",
		X"47",X"EC",X"81",X"E3",X"C8",X"11",X"AF",X"4F",X"1F",X"01",X"7E",X"D6",X"90",X"6E",X"D8",X"15",
		X"6F",X"4A",X"AF",X"4B",X"A6",X"A4",X"27",X"43",X"2A",X"0C",X"85",X"40",X"26",X"08",X"84",X"3F",
		X"A7",X"4A",X"31",X"21",X"20",X"EE",X"34",X"20",X"BD",X"D6",X"DE",X"A6",X"4A",X"27",X"07",X"6A",
		X"4A",X"27",X"03",X"10",X"AE",X"E4",X"32",X"62",X"63",X"47",X"2A",X"02",X"6C",X"4B",X"10",X"AF",
		X"4D",X"6A",X"C8",X"13",X"2A",X"0E",X"A6",X"48",X"A7",X"C8",X"13",X"8E",X"D6",X"D4",X"A6",X"C8",
		X"14",X"7E",X"00",X"A8",X"AE",X"4B",X"10",X"AE",X"4D",X"20",X"B9",X"7E",X"D6",X"72",X"34",X"06",
		X"A6",X"A0",X"34",X"02",X"85",X"40",X"26",X"06",X"84",X"3F",X"30",X"86",X"20",X"1B",X"84",X"3F",
		X"27",X"17",X"E6",X"47",X"E4",X"49",X"1A",X"10",X"7F",X"C9",X"00",X"EA",X"84",X"E7",X"80",X"C6",
		X"01",X"F7",X"C9",X"00",X"1C",X"EF",X"4A",X"26",X"E9",X"A6",X"E0",X"2A",X"D3",X"35",X"86",X"10",
		X"9F",X"4F",X"35",X"20",X"DE",X"3F",X"AF",X"47",X"10",X"AF",X"4D",X"5F",X"8D",X"61",X"5D",X"27",
		X"18",X"DE",X"3F",X"ED",X"49",X"AF",X"4B",X"86",X"01",X"8E",X"D7",X"2F",X"7E",X"00",X"A8",X"EC",
		X"49",X"AE",X"4B",X"30",X"89",X"01",X"00",X"C6",X"FF",X"5C",X"1E",X"10",X"91",X"4F",X"1E",X"10",
		X"25",X"DA",X"DE",X"3F",X"AE",X"47",X"86",X"4B",X"97",X"4F",X"BD",X"D7",X"F3",X"AF",X"4B",X"86",
		X"01",X"8E",X"D7",X"57",X"7E",X"00",X"A8",X"86",X"8C",X"97",X"4F",X"E6",X"4C",X"86",X"4B",X"1F",
		X"01",X"BD",X"D7",X"F3",X"86",X"01",X"8E",X"D7",X"6C",X"7E",X"00",X"A8",X"AE",X"4B",X"30",X"01",
		X"1E",X"10",X"86",X"0E",X"D1",X"50",X"1E",X"10",X"25",X"CC",X"DE",X"3F",X"6E",X"D8",X"0D",X"34",
		X"16",X"8D",X"20",X"26",X"04",X"8D",X"39",X"20",X"F8",X"8D",X"43",X"8D",X"33",X"8D",X"3F",X"8D",
		X"12",X"27",X"04",X"8D",X"2B",X"20",X"F8",X"30",X"1E",X"8D",X"33",X"30",X"01",X"8D",X"2F",X"30",
		X"01",X"20",X"DE",X"34",X"06",X"1A",X"10",X"7F",X"C9",X"00",X"8D",X"0C",X"A4",X"84",X"C6",X"01",
		X"F7",X"C9",X"00",X"1C",X"EF",X"4D",X"35",X"86",X"86",X"F0",X"5D",X"27",X"02",X"86",X"0F",X"39",
		X"30",X"01",X"1E",X"10",X"D1",X"50",X"1E",X"10",X"25",X"F5",X"32",X"62",X"35",X"96",X"34",X"06",
		X"1A",X"10",X"7F",X"C9",X"00",X"8D",X"E1",X"A4",X"84",X"27",X"0F",X"8D",X"DB",X"84",X"99",X"34",
		X"02",X"8D",X"D5",X"43",X"A4",X"84",X"AA",X"E0",X"A7",X"84",X"86",X"01",X"B7",X"C9",X"00",X"1C",
		X"EF",X"35",X"86",X"34",X"16",X"5F",X"8D",X"AB",X"26",X"04",X"8D",X"1E",X"20",X"F8",X"8D",X"CE",
		X"8D",X"18",X"8D",X"CA",X"8D",X"9D",X"27",X"04",X"8D",X"10",X"20",X"F8",X"30",X"89",X"FF",X"00",
		X"8D",X"BC",X"8D",X"06",X"8D",X"B8",X"8D",X"02",X"20",X"DC",X"5D",X"27",X"0E",X"30",X"89",X"01",
		X"00",X"1E",X"10",X"91",X"4F",X"1E",X"10",X"24",X"A1",X"C6",X"FF",X"5C",X"39",X"D8",X"5F",X"11",
		X"F0",X"00",X"00",X"D8",X"89",X"22",X"F0",X"10",X"00",X"D8",X"92",X"33",X"F0",X"1F",X"00",X"D8",
		X"DF",X"44",X"F0",X"2F",X"00",X"D9",X"06",X"55",X"F0",X"3F",X"00",X"D8",X"92",X"66",X"F0",X"4F",
		X"00",X"D8",X"89",X"77",X"F0",X"5F",X"00",X"D9",X"30",X"88",X"F0",X"6F",X"00",X"00",X"00",X"06",
		X"44",X"09",X"D0",X"04",X"48",X"07",X"D0",X"03",X"4A",X"06",X"D0",X"02",X"4C",X"05",X"D0",X"82",
		X"01",X"4E",X"04",X"D0",X"8D",X"50",X"03",X"D0",X"82",X"50",X"04",X"CE",X"50",X"05",X"CC",X"50",
		X"06",X"CA",X"50",X"07",X"C8",X"50",X"09",X"C4",X"00",X"87",X"CA",X"8A",X"4A",X"02",X"D7",X"87",
		X"CA",X"00",X"0F",X"42",X"02",X"D0",X"0D",X"44",X"02",X"D0",X"0B",X"46",X"02",X"D0",X"09",X"48",
		X"02",X"D0",X"07",X"4A",X"02",X"D0",X"05",X"4C",X"02",X"D0",X"03",X"4E",X"02",X"D0",X"01",X"50",
		X"02",X"D0",X"82",X"51",X"02",X"D0",X"85",X"4C",X"07",X"C5",X"82",X"51",X"02",X"D0",X"01",X"50",
		X"02",X"D0",X"03",X"4E",X"02",X"D0",X"05",X"4C",X"02",X"D0",X"07",X"4A",X"02",X"D0",X"09",X"48",
		X"02",X"D0",X"0B",X"46",X"02",X"D0",X"0D",X"44",X"02",X"D0",X"0F",X"42",X"02",X"D0",X"00",X"8A",
		X"E3",X"C0",X"C0",X"84",X"56",X"02",X"CB",X"82",X"01",X"55",X"02",X"CB",X"82",X"02",X"54",X"02",
		X"CB",X"03",X"53",X"04",X"C9",X"04",X"51",X"07",X"C7",X"05",X"4F",X"0A",X"C5",X"07",X"4B",X"0E",
		X"C3",X"09",X"47",X"12",X"C1",X"00",X"0C",X"CB",X"0A",X"CF",X"08",X"D3",X"07",X"D5",X"05",X"D8",
		X"04",X"DA",X"03",X"DC",X"02",X"DE",X"02",X"DF",X"01",X"4F",X"03",X"CE",X"01",X"4D",X"07",X"CD",
		X"4C",X"0B",X"CC",X"82",X"4B",X"0D",X"CB",X"82",X"4A",X"0F",X"CA",X"89",X"4A",X"02",X"D7",X"00",
		X"89",X"4A",X"02",X"D7",X"8F",X"4A",X"02",X"4A",X"03",X"CA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"86",X"FF",X"97",X"91",X"86",X"30",X"97",X"F8",X"7F",X"BD",X"DE",X"7F",X"BE",X"1D",X"7F",X"BD",
		X"E0",X"7F",X"BE",X"1F",X"7F",X"BD",X"E1",X"7F",X"BE",X"20",X"BD",X"D0",X"09",X"BD",X"13",X"BD",
		X"BD",X"08",X"3A",X"86",X"01",X"DE",X"3F",X"BD",X"5F",X"EA",X"8E",X"00",X"00",X"BD",X"DC",X"CB",
		X"86",X"05",X"BD",X"70",X"4F",X"86",X"01",X"BD",X"5F",X"F0",X"CC",X"30",X"00",X"ED",X"0A",X"86",
		X"80",X"A7",X"0C",X"CC",X"19",X"35",X"ED",X"08",X"0F",X"F1",X"0F",X"F2",X"BD",X"45",X"60",X"86",
		X"80",X"97",X"91",X"86",X"02",X"DE",X"3F",X"BD",X"5F",X"ED",X"BD",X"5F",X"DE",X"CC",X"02",X"00",
		X"DD",X"F1",X"86",X"60",X"8E",X"DA",X"6A",X"7E",X"00",X"A8",X"86",X"FF",X"97",X"91",X"C6",X"1C",
		X"BD",X"45",X"52",X"86",X"02",X"DE",X"3F",X"BD",X"5F",X"EA",X"BD",X"13",X"DD",X"BD",X"5F",X"DB",
		X"8E",X"80",X"00",X"9F",X"20",X"9F",X"22",X"BD",X"2C",X"00",X"0F",X"F1",X"86",X"80",X"97",X"91",
		X"DE",X"3F",X"BD",X"10",X"CA",X"86",X"02",X"DE",X"3F",X"BD",X"5F",X"ED",X"0F",X"D2",X"86",X"14",
		X"B7",X"BE",X"7C",X"8E",X"DA",X"EF",X"AF",X"47",X"AE",X"47",X"EC",X"81",X"27",X"3F",X"81",X"FF",
		X"26",X"0E",X"B6",X"BE",X"7C",X"D6",X"D2",X"30",X"01",X"10",X"A3",X"1E",X"26",X"2F",X"20",X"EA",
		X"AF",X"47",X"34",X"06",X"C5",X"20",X"27",X"0A",X"8E",X"0D",X"CF",X"86",X"04",X"BD",X"01",X"30",
		X"EC",X"E4",X"C5",X"10",X"27",X"07",X"BD",X"19",X"43",X"17",X"E2",X"EC",X"E4",X"C4",X"01",X"D7",
		X"F2",X"35",X"06",X"C4",X"82",X"D7",X"F1",X"8E",X"DA",X"A8",X"7E",X"00",X"A8",X"20",X"52",X"30",
		X"02",X"0C",X"A2",X"FF",X"13",X"00",X"05",X"82",X"18",X"00",X"FF",X"13",X"01",X"20",X"01",X"0C",
		X"A2",X"FF",X"12",X"01",X"18",X"02",X"FF",X"12",X"02",X"1A",X"01",X"0D",X"A2",X"FF",X"11",X"02",
		X"1C",X"02",X"FF",X"11",X"03",X"1A",X"01",X"07",X"22",X"FF",X"10",X"03",X"19",X"02",X"2C",X"92",
		X"28",X"02",X"1C",X"12",X"FF",X"10",X"04",X"09",X"01",X"98",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"8E",X"DC",X"A9",X"AF",X"47",X"86",X"FF",X"97",X"91",X"BD",X"D0",X"09",X"86",X"03",X"BD",
		X"5F",X"EA",X"10",X"AE",X"47",X"AE",X"A1",X"8C",X"FF",X"FF",X"10",X"27",X"01",X"BE",X"34",X"60",
		X"BD",X"DC",X"CB",X"0F",X"F1",X"0F",X"F2",X"8E",X"BE",X"7C",X"6F",X"80",X"8C",X"BE",X"83",X"26",
		X"F9",X"86",X"01",X"97",X"67",X"BD",X"07",X"D9",X"9F",X"69",X"86",X"02",X"A7",X"09",X"BD",X"5F",
		X"E1",X"BD",X"5F",X"E4",X"BD",X"07",X"EC",X"84",X"3F",X"8B",X"E0",X"9B",X"9C",X"97",X"9C",X"97",
		X"97",X"97",X"99",X"96",X"B8",X"84",X"3F",X"8B",X"E0",X"8B",X"50",X"97",X"96",X"97",X"98",X"97",
		X"9A",X"96",X"B7",X"2B",X"0B",X"DC",X"92",X"43",X"53",X"C3",X"00",X"01",X"DD",X"92",X"DD",X"94",
		X"86",X"80",X"97",X"91",X"35",X"60",X"A6",X"A0",X"34",X"60",X"AD",X"B4",X"35",X"60",X"31",X"22",
		X"A6",X"A0",X"AE",X"A1",X"10",X"AF",X"47",X"BD",X"70",X"4F",X"86",X"03",X"BD",X"5F",X"ED",X"BD",
		X"5F",X"DE",X"DE",X"3F",X"CC",X"03",X"00",X"ED",X"49",X"86",X"01",X"A7",X"4B",X"A7",X"4C",X"96",
		X"B6",X"44",X"A7",X"4D",X"AE",X"49",X"86",X"10",X"97",X"88",X"30",X"1F",X"AF",X"49",X"10",X"27",
		X"00",X"85",X"96",X"91",X"81",X"DA",X"10",X"27",X"00",X"92",X"96",X"9C",X"81",X"48",X"23",X"1A",
		X"81",X"C0",X"24",X"11",X"6A",X"4B",X"27",X"17",X"BD",X"07",X"EC",X"81",X"FC",X"25",X"27",X"BD",
		X"07",X"EC",X"44",X"25",X"05",X"CC",X"00",X"01",X"20",X"08",X"CC",X"80",X"00",X"20",X"03",X"CC",
		X"00",X"00",X"D7",X"F2",X"D6",X"F1",X"C4",X"02",X"D7",X"F1",X"9A",X"F1",X"97",X"F1",X"BD",X"07",
		X"EC",X"44",X"44",X"12",X"A7",X"4B",X"6A",X"4C",X"26",X"17",X"BD",X"07",X"EC",X"D6",X"F1",X"81",
		X"80",X"22",X"04",X"CA",X"02",X"20",X"02",X"C4",X"FD",X"D7",X"F1",X"96",X"B6",X"44",X"44",X"A7",
		X"4C",X"BD",X"07",X"EC",X"81",X"0C",X"22",X"08",X"8E",X"0D",X"CF",X"86",X"04",X"BD",X"01",X"30",
		X"6A",X"4D",X"26",X"0B",X"BD",X"19",X"43",X"17",X"E2",X"96",X"B6",X"8A",X"10",X"A7",X"4D",X"86",
		X"01",X"8E",X"DB",X"E4",X"7E",X"00",X"A8",X"BD",X"D0",X"09",X"86",X"08",X"9A",X"91",X"97",X"91",
		X"86",X"02",X"BD",X"5F",X"EA",X"86",X"FF",X"97",X"91",X"7E",X"DB",X"52",X"BD",X"19",X"43",X"DC",
		X"A1",X"86",X"6C",X"8E",X"DC",X"77",X"7E",X"00",X"A8",X"8E",X"DC",X"A9",X"AF",X"47",X"7E",X"DB",
		X"52",X"9E",X"98",X"BD",X"2C",X"09",X"7E",X"00",X"E4",X"B0",X"00",X"08",X"4F",X"40",X"13",X"32",
		X"27",X"80",X"00",X"14",X"4F",X"43",X"14",X"36",X"27",X"80",X"00",X"0A",X"5A",X"D0",X"16",X"33",
		X"27",X"00",X"00",X"00",X"DD",X"06",X"15",X"2D",X"27",X"FF",X"FF",X"34",X"76",X"86",X"FF",X"97",
		X"91",X"BD",X"13",X"BD",X"86",X"66",X"97",X"DE",X"BD",X"1E",X"96",X"8E",X"2C",X"27",X"CC",X"40",
		X"05",X"BD",X"13",X"B9",X"BD",X"08",X"4A",X"EC",X"62",X"DD",X"20",X"DD",X"22",X"BD",X"2C",X"00",
		X"BD",X"08",X"FB",X"BD",X"0E",X"EC",X"BD",X"0A",X"9C",X"BD",X"5F",X"DB",X"BD",X"19",X"72",X"BD",
		X"19",X"43",X"10",X"21",X"35",X"F6",X"86",X"18",X"B7",X"BE",X"78",X"BD",X"19",X"43",X"DD",X"11",
		X"39",X"BD",X"38",X"4F",X"86",X"32",X"8E",X"DD",X"11",X"7E",X"00",X"A8",X"BD",X"13",X"BD",X"BD",
		X"08",X"3A",X"BD",X"19",X"72",X"BD",X"08",X"4A",X"BD",X"5F",X"DE",X"4F",X"5F",X"DD",X"20",X"DD",
		X"22",X"86",X"DB",X"97",X"91",X"DE",X"3F",X"8E",X"DE",X"4B",X"AF",X"47",X"10",X"AE",X"47",X"EC",
		X"A4",X"27",X"0E",X"BD",X"DD",X"E4",X"10",X"AF",X"47",X"86",X"08",X"8E",X"DD",X"3C",X"7E",X"00",
		X"A8",X"86",X"01",X"8E",X"DD",X"59",X"7E",X"00",X"A8",X"8E",X"DE",X"A9",X"AF",X"47",X"10",X"AE",
		X"47",X"A6",X"A0",X"27",X"10",X"AE",X"A1",X"10",X"AF",X"47",X"BD",X"70",X"52",X"86",X"04",X"8E",
		X"DD",X"5E",X"7E",X"00",X"A8",X"86",X"1E",X"A7",X"49",X"6F",X"4A",X"8E",X"2F",X"76",X"AF",X"4B",
		X"8E",X"DD",X"D2",X"AF",X"4D",X"8E",X"DE",X"A9",X"AF",X"47",X"6A",X"49",X"10",X"27",X"F2",X"76",
		X"10",X"AE",X"47",X"A6",X"A0",X"81",X"93",X"27",X"EC",X"AE",X"A1",X"10",X"AF",X"47",X"BD",X"70",
		X"52",X"86",X"04",X"8E",X"DD",X"A9",X"7E",X"00",X"A8",X"A6",X"4A",X"97",X"11",X"AE",X"4B",X"10",
		X"AE",X"4D",X"10",X"8C",X"DD",X"E4",X"27",X"C1",X"A6",X"A0",X"C6",X"AA",X"D7",X"10",X"BD",X"70",
		X"31",X"96",X"11",X"A7",X"4A",X"AF",X"4B",X"10",X"AF",X"4D",X"86",X"02",X"8E",X"DD",X"90",X"7E",
		X"00",X"A8",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"20",X"20",X"45",X"4E",X"45",
		X"4D",X"49",X"45",X"53",X"34",X"50",X"BD",X"19",X"43",X"DE",X"1C",X"1F",X"13",X"BD",X"01",X"88",
		X"EC",X"B1",X"ED",X"02",X"ED",X"49",X"AF",X"47",X"EC",X"A1",X"ED",X"4B",X"6F",X"4D",X"4F",X"5F",
		X"ED",X"0E",X"ED",X"88",X"10",X"EC",X"A1",X"E7",X"0C",X"6F",X"0D",X"5F",X"44",X"56",X"44",X"56",
		X"ED",X"0A",X"86",X"01",X"A7",X"88",X"14",X"BD",X"27",X"00",X"35",X"D0",X"A6",X"4B",X"81",X"01",
		X"10",X"27",X"22",X"C0",X"AE",X"47",X"EC",X"02",X"10",X"83",X"20",X"10",X"27",X"15",X"A6",X"4D",
		X"4C",X"A1",X"4B",X"25",X"01",X"4F",X"A7",X"4D",X"C6",X"0A",X"3D",X"10",X"AE",X"49",X"31",X"AB",
		X"10",X"AF",X"02",X"A6",X"4C",X"8E",X"DE",X"24",X"7E",X"00",X"A8",X"DE",X"A5",X"01",X"00",X"66",
		X"96",X"4F",X"4F",X"05",X"08",X"1D",X"4A",X"45",X"5E",X"04",X"03",X"68",X"48",X"DE",X"A7",X"04",
		X"08",X"13",X"72",X"38",X"56",X"03",X"08",X"47",X"BA",X"DE",X"A3",X"01",X"00",X"7D",X"70",X"4F",
		X"4B",X"04",X"01",X"3C",X"3C",X"5A",X"D3",X"04",X"02",X"12",X"94",X"38",X"52",X"07",X"02",X"7E",
		X"4A",X"4F",X"4D",X"08",X"02",X"56",X"3C",X"5A",X"D5",X"02",X"04",X"2C",X"98",X"DE",X"A1",X"01",
		X"00",X"7C",X"9A",X"38",X"54",X"03",X"08",X"36",X"BA",X"38",X"5C",X"03",X"08",X"5D",X"BC",X"00",
		X"00",X"20",X"9F",X"1F",X"F2",X"20",X"1B",X"20",X"4D",X"14",X"0C",X"58",X"91",X"60",X"58",X"8E",
		X"0C",X"7E",X"15",X"2D",X"C8",X"92",X"76",X"7E",X"13",X"30",X"30",X"90",X"60",X"A2",X"16",X"0C",
		X"A2",X"8F",X"78",X"58",X"93",X"2F",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"E2",X"AC",X"7E",X"E6",X"82",X"7E",X"E6",X"F6",X"7E",X"E7",X"04",X"7E",X"E0",X"0F",X"34",
		X"02",X"A6",X"80",X"1E",X"12",X"BD",X"14",X"24",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",X"8E",
		X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",X"36",X"8E",X"E0",X"51",X"10",
		X"8E",X"CC",X"00",X"C6",X"1B",X"8D",X"D8",X"35",X"B6",X"34",X"36",X"8E",X"E0",X"6C",X"10",X"8E",
		X"CC",X"36",X"C6",X"34",X"8D",X"C9",X"BD",X"E6",X"5B",X"8E",X"CC",X"A0",X"BD",X"14",X"24",X"35",
		X"B6",X"10",X"03",X"07",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"00",X"03",X"05",X"30",X"00",
		X"00",X"00",X"10",X"04",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"49",X"4C",X"4C",
		X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",
		X"20",X"49",X"4E",X"43",X"3D",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"3F",X"20",X"20",X"20",X"20",X"20",X"25",X"25",
		X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",
		X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",
		X"01",X"02",X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",
		X"01",X"00",X"02",X"02",X"00",X"00",X"05",X"30",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"03",X"13",X"00",X"00",X"00",X"05",X"30",X"00",X"00",X"00",X"05",X"50",X"02",X"06",X"01",X"05",
		X"99",X"02",X"07",X"02",X"00",X"50",X"E1",X"96",X"00",X"2C",X"01",X"20",X"E1",X"9F",X"00",X"38",
		X"00",X"50",X"E1",X"AD",X"00",X"44",X"00",X"08",X"E1",X"BE",X"00",X"57",X"00",X"99",X"E1",X"AA",
		X"01",X"62",X"00",X"99",X"E1",X"AA",X"01",X"6C",X"00",X"99",X"E1",X"AA",X"01",X"76",X"00",X"99",
		X"E1",X"AA",X"01",X"80",X"00",X"99",X"E1",X"AA",X"01",X"8A",X"00",X"99",X"E1",X"AA",X"01",X"94",
		X"00",X"01",X"E1",X"D1",X"00",X"A7",X"00",X"05",X"E1",X"DB",X"00",X"17",X"00",X"30",X"E1",X"E8",
		X"02",X"23",X"00",X"99",X"E1",X"F3",X"02",X"2E",X"00",X"20",X"E1",X"AA",X"02",X"3C",X"00",X"99",
		X"E1",X"AA",X"02",X"46",X"00",X"10",X"E1",X"FE",X"02",X"50",X"05",X"20",X"E2",X"05",X"00",X"63",
		X"02",X"09",X"E2",X"10",X"00",X"6F",X"01",X"99",X"E2",X"1B",X"00",X"7B",X"03",X"20",X"E2",X"22",
		X"00",X"87",X"00",X"01",X"E1",X"D6",X"00",X"9A",X"00",X"01",X"E1",X"D6",X"00",X"A6",X"00",X"01",
		X"E1",X"D6",X"00",X"B2",X"00",X"01",X"E1",X"D6",X"00",X"BE",X"00",X"01",X"E1",X"D6",X"00",X"CA",
		X"00",X"01",X"E1",X"D6",X"00",X"D6",X"00",X"78",X"01",X"5E",X"10",X"5F",X"11",X"5E",X"FF",X"00",
		X"60",X"02",X"61",X"03",X"62",X"04",X"63",X"05",X"60",X"FF",X"00",X"60",X"FF",X"00",X"6C",X"01",
		X"60",X"05",X"61",X"06",X"60",X"07",X"62",X"08",X"60",X"09",X"63",X"10",X"60",X"FF",X"00",X"64",
		X"01",X"70",X"02",X"71",X"03",X"72",X"04",X"73",X"05",X"74",X"06",X"75",X"07",X"76",X"08",X"77",
		X"FF",X"00",X"66",X"01",X"65",X"FF",X"00",X"66",X"01",X"6F",X"FF",X"00",X"64",X"01",X"67",X"02",
		X"68",X"03",X"62",X"04",X"6A",X"05",X"6B",X"FF",X"00",X"67",X"03",X"68",X"05",X"69",X"07",X"6A",
		X"10",X"6B",X"FF",X"00",X"67",X"13",X"68",X"26",X"69",X"39",X"6A",X"60",X"6B",X"FF",X"00",X"69",
		X"01",X"6A",X"02",X"6B",X"FF",X"00",X"6B",X"07",X"6A",X"10",X"62",X"11",X"68",X"15",X"67",X"FF",
		X"00",X"67",X"03",X"68",X"04",X"62",X"05",X"6A",X"06",X"6B",X"FF",X"00",X"60",X"10",X"62",X"11",
		X"60",X"FF",X"00",X"60",X"20",X"62",X"FF",X"34",X"22",X"86",X"11",X"6D",X"44",X"27",X"02",X"86",
		X"16",X"E6",X"45",X"1F",X"01",X"A6",X"E4",X"BD",X"70",X"52",X"8D",X"02",X"35",X"A2",X"34",X"36",
		X"1E",X"12",X"BD",X"14",X"1C",X"1E",X"12",X"1E",X"10",X"86",X"59",X"E6",X"45",X"1E",X"10",X"34",
		X"06",X"CC",X"3C",X"05",X"BD",X"13",X"B9",X"35",X"06",X"8D",X"05",X"BD",X"70",X"52",X"35",X"B6",
		X"34",X"20",X"10",X"AE",X"42",X"E1",X"A1",X"24",X"FC",X"A6",X"3D",X"35",X"A0",X"BD",X"13",X"BD",
		X"CE",X"E0",X"F4",X"10",X"8E",X"CC",X"00",X"86",X"43",X"8E",X"CC",X"16",X"8D",X"1E",X"86",X"42",
		X"BD",X"70",X"4F",X"CE",X"E1",X"30",X"10",X"8E",X"CC",X"14",X"86",X"4D",X"39",X"BD",X"13",X"BD",
		X"CE",X"E1",X"36",X"10",X"8E",X"CC",X"16",X"86",X"4E",X"8E",X"CC",X"36",X"34",X"76",X"8D",X"87",
		X"33",X"46",X"31",X"22",X"4C",X"10",X"AC",X"62",X"26",X"F4",X"35",X"F6",X"8E",X"CC",X"2A",X"6F",
		X"80",X"8C",X"CC",X"36",X"25",X"F9",X"BD",X"E6",X"42",X"8D",X"B2",X"CE",X"E0",X"F4",X"10",X"8E",
		X"CC",X"00",X"86",X"43",X"BD",X"E5",X"CD",X"BD",X"E3",X"7A",X"BD",X"19",X"43",X"E4",X"31",X"BD",
		X"E3",X"99",X"8D",X"08",X"86",X"01",X"8E",X"E2",X"CF",X"7E",X"00",X"A8",X"35",X"06",X"DE",X"3F",
		X"ED",X"4D",X"86",X"20",X"A7",X"47",X"B6",X"C8",X"04",X"46",X"25",X"06",X"46",X"25",X"1E",X"6E",
		X"D8",X"0D",X"BD",X"E3",X"29",X"86",X"01",X"8E",X"E2",X"FD",X"7E",X"00",X"A8",X"B6",X"C8",X"04",
		X"46",X"24",X"EC",X"6A",X"47",X"26",X"EE",X"86",X"05",X"A7",X"47",X"20",X"E5",X"BD",X"E3",X"49",
		X"86",X"01",X"8E",X"E3",X"18",X"7E",X"00",X"A8",X"B6",X"C8",X"04",X"85",X"02",X"27",X"D0",X"6A",
		X"47",X"26",X"ED",X"86",X"05",X"A7",X"47",X"20",X"E4",X"BD",X"E5",X"D8",X"1F",X"21",X"BD",X"14",
		X"0B",X"8B",X"01",X"19",X"25",X"12",X"A1",X"41",X"22",X"0E",X"1F",X"21",X"BD",X"14",X"24",X"BD",
		X"E6",X"42",X"BD",X"E2",X"3E",X"BD",X"E5",X"E3",X"39",X"BD",X"E5",X"D8",X"1F",X"21",X"BD",X"14",
		X"0B",X"4D",X"27",X"F4",X"8B",X"99",X"19",X"A1",X"C4",X"25",X"ED",X"20",X"DD",X"34",X"12",X"A6",
		X"44",X"27",X"13",X"8E",X"CC",X"06",X"4A",X"27",X"03",X"8E",X"CC",X"16",X"BD",X"14",X"0B",X"4D",
		X"27",X"04",X"1A",X"01",X"35",X"92",X"1C",X"FE",X"35",X"92",X"34",X"16",X"E6",X"45",X"86",X"0C",
		X"1F",X"01",X"86",X"41",X"BD",X"70",X"52",X"35",X"96",X"34",X"16",X"E6",X"45",X"86",X"0C",X"1F",
		X"01",X"CC",X"03",X"05",X"BD",X"13",X"B9",X"35",X"96",X"35",X"06",X"DE",X"3F",X"ED",X"4D",X"86",
		X"30",X"A7",X"47",X"B6",X"C8",X"04",X"2B",X"09",X"B6",X"C8",X"06",X"46",X"25",X"1D",X"6E",X"D8",
		X"0D",X"BD",X"E3",X"E6",X"86",X"01",X"8E",X"E3",X"BC",X"7E",X"00",X"A8",X"B6",X"C8",X"04",X"2A",
		X"ED",X"6A",X"47",X"26",X"EF",X"86",X"08",X"A7",X"47",X"20",X"E6",X"BD",X"E4",X"0C",X"86",X"01",
		X"8E",X"E3",X"D6",X"7E",X"00",X"A8",X"B6",X"C8",X"06",X"46",X"24",X"D2",X"6A",X"47",X"26",X"EE",
		X"86",X"08",X"A7",X"47",X"20",X"E5",X"BD",X"E5",X"D8",X"BD",X"E3",X"89",X"10",X"8C",X"CC",X"34",
		X"27",X"16",X"31",X"22",X"4C",X"33",X"46",X"10",X"8C",X"CC",X"16",X"26",X"03",X"BD",X"E2",X"8D",
		X"BD",X"E3",X"5D",X"25",X"E7",X"BD",X"E5",X"CD",X"BD",X"E3",X"7A",X"39",X"BD",X"E5",X"D8",X"BD",
		X"E3",X"89",X"10",X"8C",X"CC",X"00",X"27",X"F0",X"31",X"3E",X"4A",X"33",X"5A",X"10",X"8C",X"CC",
		X"14",X"26",X"03",X"BD",X"E2",X"6D",X"BD",X"E3",X"5D",X"25",X"E7",X"BD",X"E5",X"CD",X"7E",X"E3",
		X"7A",X"86",X"01",X"8E",X"E4",X"39",X"7E",X"00",X"A8",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F1",
		X"BD",X"01",X"57",X"BD",X"13",X"BD",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"2D",
		X"84",X"0F",X"27",X"14",X"7F",X"CC",X"2D",X"BD",X"E6",X"42",X"BD",X"13",X"BD",X"BD",X"E6",X"DF",
		X"86",X"40",X"8E",X"E4",X"68",X"7E",X"00",X"A8",X"B6",X"CC",X"2F",X"84",X"0F",X"27",X"11",X"7F",
		X"CC",X"2F",X"BD",X"E6",X"42",X"BD",X"E9",X"49",X"86",X"40",X"8E",X"E4",X"80",X"7E",X"00",X"A8",
		X"B6",X"CC",X"33",X"84",X"0F",X"27",X"5E",X"7F",X"CC",X"33",X"BD",X"E6",X"42",X"86",X"3A",X"8E",
		X"CC",X"36",X"C6",X"32",X"BD",X"14",X"24",X"5A",X"26",X"FA",X"BD",X"13",X"BD",X"86",X"7D",X"BD",
		X"70",X"55",X"10",X"8E",X"CC",X"36",X"8E",X"25",X"30",X"CC",X"19",X"80",X"BD",X"E7",X"04",X"C6",
		X"30",X"8E",X"CC",X"9A",X"10",X"8E",X"CC",X"36",X"BD",X"E5",X"24",X"86",X"7D",X"BD",X"70",X"55",
		X"BD",X"E5",X"A7",X"10",X"8E",X"CC",X"68",X"8E",X"25",X"40",X"CC",X"19",X"80",X"BD",X"E7",X"04",
		X"C6",X"40",X"8E",X"CC",X"9C",X"10",X"8E",X"CC",X"68",X"BD",X"E5",X"24",X"BD",X"E6",X"5B",X"8E",
		X"CC",X"A0",X"BD",X"14",X"24",X"B6",X"CC",X"35",X"84",X"0F",X"27",X"09",X"7F",X"CC",X"35",X"BD",
		X"E6",X"42",X"BD",X"E9",X"46",X"B6",X"CC",X"31",X"84",X"0F",X"27",X"0B",X"7F",X"CC",X"31",X"BD",
		X"E6",X"42",X"8D",X"0F",X"7E",X"F4",X"8C",X"8D",X"0A",X"CC",X"00",X"00",X"DD",X"5E",X"DD",X"62",
		X"7E",X"5F",X"D6",X"B6",X"CC",X"2B",X"84",X"0F",X"27",X"09",X"7C",X"CC",X"9E",X"7C",X"CC",X"9E",
		X"7F",X"CC",X"2B",X"39",X"DE",X"3F",X"86",X"25",X"ED",X"47",X"35",X"06",X"ED",X"4D",X"AF",X"4B",
		X"10",X"AF",X"49",X"86",X"25",X"BD",X"14",X"24",X"86",X"95",X"BD",X"70",X"55",X"86",X"04",X"8E",
		X"E5",X"45",X"7E",X"00",X"A8",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F1",X"B6",X"C8",X"04",X"46",
		X"24",X"10",X"AE",X"4B",X"BD",X"14",X"0B",X"AE",X"4B",X"4C",X"81",X"3C",X"23",X"15",X"86",X"3C",
		X"20",X"11",X"46",X"24",X"1E",X"AE",X"4B",X"BD",X"14",X"0B",X"AE",X"4B",X"4A",X"81",X"10",X"24",
		X"02",X"86",X"10",X"BD",X"14",X"24",X"A7",X"47",X"BD",X"E5",X"A7",X"86",X"10",X"8E",X"E5",X"4C",
		X"7E",X"00",X"A8",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"08",X"86",X"04",X"8E",X"E5",X"4C",X"7E",
		X"00",X"A8",X"BD",X"13",X"BD",X"86",X"04",X"8E",X"E5",X"9D",X"7E",X"00",X"A8",X"B6",X"C8",X"0C",
		X"85",X"02",X"26",X"F1",X"6E",X"D8",X"0D",X"0F",X"11",X"AE",X"47",X"30",X"89",X"FF",X"00",X"86",
		X"5A",X"C6",X"09",X"BD",X"13",X"B9",X"AE",X"47",X"0F",X"11",X"10",X"AE",X"49",X"C6",X"19",X"1E",
		X"12",X"BD",X"14",X"0B",X"1E",X"12",X"BD",X"70",X"31",X"5A",X"26",X"F3",X"39",X"10",X"BF",X"9D",
		X"02",X"FF",X"9D",X"05",X"B7",X"9D",X"04",X"39",X"10",X"BE",X"9D",X"02",X"FE",X"9D",X"05",X"B6",
		X"9D",X"04",X"39",X"10",X"8C",X"CC",X"16",X"27",X"07",X"10",X"8C",X"CC",X"06",X"27",X"2B",X"39",
		X"1F",X"21",X"BD",X"14",X"0B",X"34",X"02",X"48",X"48",X"AB",X"E0",X"8E",X"E0",X"D6",X"30",X"86",
		X"33",X"46",X"31",X"22",X"A6",X"80",X"34",X"10",X"1F",X"21",X"BD",X"14",X"24",X"35",X"10",X"BD",
		X"E2",X"3E",X"10",X"8C",X"CC",X"20",X"25",X"E8",X"20",X"28",X"1F",X"21",X"BD",X"14",X"0B",X"48",
		X"34",X"02",X"48",X"AB",X"E0",X"8E",X"E0",X"A0",X"30",X"86",X"33",X"46",X"31",X"22",X"A6",X"80",
		X"34",X"10",X"1F",X"21",X"BD",X"14",X"24",X"35",X"10",X"BD",X"E2",X"3E",X"10",X"8C",X"CC",X"12",
		X"25",X"E8",X"34",X"12",X"8D",X"08",X"8E",X"CC",X"9E",X"BD",X"14",X"24",X"35",X"92",X"34",X"34",
		X"8E",X"CC",X"00",X"10",X"8E",X"CC",X"36",X"8D",X"09",X"35",X"B4",X"8E",X"CC",X"36",X"10",X"8E",
		X"CC",X"9E",X"10",X"9F",X"4F",X"4F",X"E6",X"80",X"C4",X"0F",X"34",X"04",X"AB",X"E0",X"9C",X"4F",
		X"26",X"F4",X"8B",X"37",X"39",X"8D",X"D7",X"34",X"02",X"8E",X"CC",X"9E",X"BD",X"14",X"0B",X"A1",
		X"E0",X"39",X"8D",X"6B",X"8D",X"EF",X"27",X"3A",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"E0",X"2A",
		X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"AB",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"13",X"BD",X"86",
		X"39",X"B7",X"CB",X"FF",X"8D",X"23",X"BD",X"E9",X"4C",X"BD",X"E9",X"40",X"8D",X"C7",X"27",X"15",
		X"86",X"6D",X"BD",X"70",X"55",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"27",
		X"F4",X"39",X"7E",X"E9",X"40",X"86",X"6E",X"20",X"E9",X"8E",X"CD",X"02",X"C6",X"04",X"A6",X"80",
		X"84",X"0F",X"81",X"09",X"23",X"03",X"5A",X"27",X"06",X"8C",X"CD",X"38",X"26",X"F0",X"39",X"86",
		X"79",X"BD",X"70",X"55",X"8E",X"CD",X"02",X"6F",X"80",X"8C",X"CD",X"38",X"26",X"F9",X"39",X"8D",
		X"05",X"27",X"FB",X"7E",X"E0",X"39",X"BD",X"E6",X"5B",X"34",X"02",X"8E",X"CC",X"A0",X"BD",X"14",
		X"0B",X"A1",X"E0",X"39",X"DE",X"3F",X"ED",X"47",X"AF",X"49",X"10",X"AF",X"4B",X"35",X"06",X"ED",
		X"4D",X"86",X"04",X"8E",X"E7",X"19",X"7E",X"00",X"A8",X"B6",X"C8",X"04",X"46",X"25",X"F2",X"BD",
		X"19",X"43",X"E8",X"ED",X"EC",X"4D",X"ED",X"0D",X"EC",X"47",X"ED",X"07",X"EF",X"09",X"9F",X"F9",
		X"86",X"99",X"97",X"10",X"0F",X"11",X"7F",X"BE",X"BF",X"7F",X"BE",X"C0",X"7F",X"BE",X"C1",X"BD",
		X"E7",X"CF",X"BD",X"E7",X"DB",X"86",X"3A",X"BD",X"E8",X"06",X"86",X"02",X"8E",X"E7",X"52",X"7E",
		X"00",X"A8",X"BD",X"E8",X"2C",X"B6",X"C8",X"04",X"46",X"24",X"EF",X"A6",X"48",X"8B",X"0A",X"A7",
		X"48",X"86",X"02",X"8E",X"E7",X"69",X"7E",X"00",X"A8",X"B6",X"C8",X"04",X"46",X"24",X"0A",X"6A",
		X"48",X"27",X"06",X"A6",X"48",X"81",X"80",X"26",X"E8",X"A6",X"48",X"84",X"80",X"A7",X"48",X"8D",
		X"70",X"81",X"5E",X"27",X"22",X"96",X"11",X"B7",X"BE",X"C1",X"8D",X"62",X"8D",X"63",X"AE",X"49",
		X"BF",X"BE",X"BF",X"BD",X"70",X"31",X"AF",X"49",X"BD",X"E8",X"1B",X"6A",X"47",X"26",X"A0",X"9E",
		X"F9",X"BD",X"00",X"EE",X"6E",X"D8",X"0D",X"8D",X"45",X"8D",X"24",X"86",X"3A",X"BD",X"E8",X"06",
		X"BE",X"BE",X"BF",X"AF",X"49",X"F6",X"BE",X"C1",X"D7",X"11",X"6C",X"47",X"10",X"AE",X"4B",X"31",
		X"3F",X"10",X"8C",X"C0",X"00",X"25",X"02",X"31",X"3F",X"10",X"AF",X"4B",X"7E",X"E7",X"36",X"34",
		X"06",X"AE",X"49",X"CC",X"04",X"07",X"BD",X"13",X"B9",X"35",X"86",X"86",X"99",X"AE",X"49",X"A7",
		X"08",X"A7",X"89",X"01",X"08",X"A7",X"89",X"02",X"08",X"A7",X"89",X"03",X"08",X"39",X"4F",X"20",
		X"EC",X"10",X"AE",X"4B",X"10",X"8C",X"C0",X"00",X"24",X"03",X"A6",X"A4",X"39",X"34",X"10",X"AE",
		X"4B",X"BD",X"14",X"0B",X"35",X"90",X"10",X"AE",X"4B",X"10",X"8C",X"C0",X"00",X"24",X"03",X"A7",
		X"A4",X"39",X"34",X"10",X"AE",X"4B",X"BD",X"14",X"24",X"35",X"90",X"10",X"AE",X"4B",X"31",X"21",
		X"10",X"8C",X"C0",X"00",X"25",X"02",X"31",X"21",X"10",X"AF",X"4B",X"39",X"B6",X"C8",X"04",X"2B",
		X"07",X"B6",X"C8",X"06",X"46",X"25",X"14",X"39",X"86",X"0A",X"8D",X"6C",X"BD",X"E8",X"E5",X"F6",
		X"C8",X"04",X"2A",X"F3",X"4A",X"26",X"F5",X"86",X"01",X"20",X"EF",X"86",X"0A",X"8D",X"10",X"BD",
		X"E8",X"E5",X"F6",X"C8",X"06",X"56",X"24",X"DF",X"4A",X"26",X"F4",X"86",X"01",X"20",X"EE",X"34",
		X"02",X"8D",X"8E",X"4C",X"6D",X"48",X"27",X"16",X"7D",X"BE",X"BF",X"27",X"04",X"81",X"5E",X"23",
		X"06",X"81",X"5D",X"23",X"02",X"86",X"30",X"81",X"3E",X"26",X"1C",X"4C",X"20",X"19",X"81",X"5A",
		X"23",X"0F",X"7D",X"BE",X"BF",X"27",X"08",X"81",X"5E",X"22",X"04",X"86",X"5E",X"20",X"02",X"86",
		X"3A",X"81",X"3B",X"26",X"02",X"86",X"41",X"BD",X"E8",X"06",X"BD",X"E7",X"CF",X"D6",X"11",X"AE",
		X"49",X"BD",X"70",X"31",X"D7",X"11",X"35",X"82",X"34",X"02",X"BD",X"E7",X"F1",X"4A",X"6D",X"48",
		X"27",X"16",X"81",X"30",X"24",X"0B",X"7D",X"BE",X"BF",X"27",X"04",X"86",X"5E",X"20",X"02",X"86",
		X"5D",X"81",X"3E",X"26",X"1E",X"4A",X"20",X"1B",X"81",X"39",X"26",X"0B",X"7D",X"BE",X"BF",X"27",
		X"04",X"86",X"5E",X"20",X"02",X"86",X"5A",X"81",X"40",X"26",X"02",X"86",X"3A",X"81",X"5D",X"26",
		X"02",X"86",X"5A",X"20",X"B2",X"8E",X"20",X"00",X"30",X"1F",X"26",X"FC",X"39",X"6D",X"48",X"26",
		X"34",X"86",X"FF",X"8E",X"E8",X"F9",X"7E",X"00",X"A8",X"86",X"FF",X"8E",X"E9",X"01",X"7E",X"00",
		X"A8",X"86",X"82",X"8E",X"E9",X"09",X"7E",X"00",X"A8",X"6A",X"47",X"26",X"E4",X"AE",X"49",X"33",
		X"84",X"BD",X"E7",X"F1",X"81",X"5E",X"26",X"05",X"86",X"3A",X"BD",X"E8",X"06",X"DE",X"3F",X"BD",
		X"00",X"EE",X"6E",X"D8",X"0D",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"E1",X"86",X"01",X"8E",X"E9",
		X"25",X"7E",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"EB",X"6B",X"7E",X"EC",X"6D",X"7E",X"EE",X"0C",X"7E",X"E9",X"A3",X"7E",X"E9",X"83",X"7E",
		X"E9",X"52",X"86",X"18",X"A7",X"47",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"08",X"8E",X"E9",X"63",
		X"7E",X"00",X"A8",X"B6",X"C8",X"0C",X"85",X"08",X"27",X"16",X"6A",X"47",X"26",X"ED",X"10",X"8E",
		X"CD",X"38",X"8E",X"E9",X"DC",X"C6",X"17",X"BD",X"E0",X"0C",X"BD",X"EB",X"32",X"7F",X"C8",X"0E",
		X"7E",X"00",X"E4",X"10",X"8E",X"CD",X"6E",X"C6",X"08",X"BD",X"EB",X"59",X"A8",X"26",X"84",X"0F",
		X"27",X"03",X"5A",X"27",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"9E",
		X"25",X"E7",X"39",X"86",X"39",X"B7",X"CB",X"FF",X"8E",X"E9",X"DC",X"10",X"8E",X"CD",X"38",X"C6",
		X"7D",X"BD",X"E0",X"0C",X"8E",X"EA",X"59",X"10",X"8E",X"CE",X"32",X"C6",X"B6",X"BD",X"E0",X"0C",
		X"BD",X"EB",X"32",X"10",X"8E",X"CD",X"6E",X"BD",X"EB",X"51",X"86",X"39",X"B7",X"CB",X"FF",X"31",
		X"2E",X"10",X"8C",X"CF",X"9E",X"25",X"F0",X"86",X"7E",X"7E",X"70",X"55",X"50",X"48",X"52",X"50",
		X"48",X"52",X"45",X"44",X"3A",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"00",X"10",X"21",X"81",X"56",X"49",X"44",X"00",X"04",X"16",X"45",X"4B",X"49",
		X"44",X"00",X"04",X"16",X"35",X"4C",X"54",X"44",X"00",X"04",X"16",X"30",X"44",X"52",X"4A",X"00",
		X"03",X"64",X"40",X"4C",X"45",X"44",X"00",X"02",X"18",X"57",X"53",X"41",X"4D",X"00",X"01",X"95",
		X"55",X"53",X"53",X"52",X"00",X"01",X"45",X"65",X"45",X"50",X"4A",X"00",X"01",X"27",X"55",X"4A",
		X"45",X"52",X"00",X"01",X"27",X"50",X"43",X"52",X"42",X"00",X"01",X"21",X"50",X"50",X"47",X"44",
		X"00",X"01",X"11",X"10",X"4B",X"4A",X"46",X"00",X"01",X"04",X"20",X"4D",X"52",X"53",X"00",X"00",
		X"92",X"35",X"4D",X"4C",X"47",X"00",X"00",X"91",X"90",X"43",X"48",X"4F",X"00",X"00",X"84",X"05",
		X"54",X"4D",X"48",X"00",X"00",X"76",X"55",X"57",X"49",X"5A",X"00",X"00",X"75",X"35",X"4D",X"48",
		X"53",X"00",X"00",X"67",X"85",X"4D",X"44",X"52",X"00",X"00",X"66",X"65",X"4D",X"50",X"54",X"00",
		X"00",X"59",X"60",X"57",X"3A",X"52",X"00",X"00",X"56",X"70",X"44",X"47",X"59",X"00",X"00",X"55",
		X"60",X"47",X"48",X"48",X"00",X"00",X"54",X"30",X"45",X"4A",X"53",X"00",X"00",X"53",X"20",X"42",
		X"41",X"43",X"00",X"00",X"52",X"40",X"47",X"3A",X"57",X"00",X"00",X"52",X"20",X"4A",X"4A",X"4B",
		X"00",X"00",X"52",X"10",X"53",X"3A",X"4D",X"00",X"00",X"51",X"80",X"52",X"3A",X"47",X"00",X"00",
		X"51",X"55",X"4C",X"3A",X"52",X"00",X"00",X"51",X"30",X"53",X"46",X"44",X"00",X"00",X"51",X"15",
		X"41",X"4B",X"44",X"00",X"00",X"51",X"05",X"43",X"57",X"4B",X"00",X"00",X"50",X"70",X"4C",X"49",
		X"55",X"00",X"00",X"50",X"45",X"54",X"49",X"4D",X"00",X"00",X"50",X"20",X"4B",X"52",X"44",X"00",
		X"00",X"48",X"65",X"4E",X"48",X"44",X"00",X"00",X"47",X"85",X"52",X"41",X"59",X"00",X"00",X"47",
		X"65",X"47",X"41",X"59",X"00",X"00",X"47",X"65",X"52",X"4B",X"4D",X"00",X"00",X"45",X"55",X"3A",
		X"3A",X"3A",X"00",X"00",X"40",X"00",X"FF",X"01",X"01",X"1B",X"01",X"01",X"02",X"00",X"FF",X"01",
		X"01",X"1B",X"01",X"01",X"01",X"00",X"34",X"34",X"8E",X"EB",X"0F",X"C6",X"07",X"BD",X"E0",X"0C",
		X"35",X"B4",X"34",X"02",X"8D",X"05",X"B7",X"CD",X"66",X"35",X"82",X"34",X"10",X"8E",X"CD",X"38",
		X"4F",X"AB",X"84",X"30",X"01",X"8C",X"CD",X"66",X"27",X"F9",X"8C",X"CD",X"6E",X"26",X"F2",X"35",
		X"90",X"34",X"02",X"8D",X"04",X"A7",X"26",X"35",X"82",X"34",X"24",X"C6",X"0E",X"4F",X"C1",X"08",
		X"27",X"02",X"AB",X"A4",X"31",X"21",X"5A",X"26",X"F5",X"35",X"A4",X"86",X"32",X"34",X"02",X"10",
		X"8E",X"CD",X"6E",X"8D",X"E4",X"A8",X"26",X"84",X"0F",X"27",X"0F",X"BD",X"EC",X"42",X"7F",X"CD",
		X"00",X"7F",X"CD",X"01",X"6A",X"E4",X"27",X"12",X"20",X"E9",X"86",X"03",X"C6",X"04",X"8D",X"68",
		X"25",X"E9",X"31",X"2E",X"10",X"8C",X"CF",X"9E",X"25",X"D9",X"35",X"02",X"8E",X"EA",X"0C",X"10",
		X"8E",X"CF",X"9E",X"C6",X"2A",X"BD",X"E0",X"0C",X"8D",X"91",X"B8",X"CD",X"66",X"84",X"0F",X"27",
		X"02",X"8D",X"0F",X"10",X"8E",X"CD",X"38",X"86",X"17",X"C6",X"04",X"8D",X"3B",X"24",X"02",X"8D",
		X"01",X"39",X"8E",X"CD",X"3E",X"86",X"3A",X"BD",X"14",X"24",X"8C",X"CD",X"66",X"25",X"F8",X"8E",
		X"CD",X"6E",X"10",X"8E",X"CD",X"3E",X"86",X"06",X"BD",X"EC",X"62",X"10",X"8E",X"CD",X"38",X"BD",
		X"EC",X"62",X"8E",X"CD",X"74",X"10",X"8E",X"CD",X"66",X"86",X"08",X"BD",X"EC",X"62",X"BD",X"EB",
		X"32",X"10",X"8E",X"CD",X"6E",X"7E",X"EC",X"42",X"34",X"16",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",
		X"21",X"BD",X"14",X"1C",X"C1",X"41",X"24",X"04",X"C1",X"3A",X"26",X"32",X"C1",X"5A",X"22",X"2E",
		X"4A",X"26",X"EE",X"A6",X"61",X"BD",X"14",X"1C",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",
		X"14",X"1C",X"34",X"04",X"C4",X"0F",X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",
		X"22",X"0C",X"4A",X"26",X"EA",X"1C",X"FE",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"96",X"1A",X"01",
		X"20",X"F5",X"34",X"36",X"30",X"2E",X"8C",X"CF",X"9E",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",
		X"2E",X"30",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"EC",X"BD",X"EB",X"26",X"BD",X"EB",X"51",
		X"35",X"B6",X"34",X"36",X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"0F",X"F8",X"BD",
		X"13",X"BD",X"BD",X"15",X"15",X"8E",X"BD",X"D6",X"C6",X"01",X"8D",X"20",X"D6",X"68",X"5A",X"27",
		X"18",X"BD",X"13",X"BD",X"B6",X"C8",X"06",X"2A",X"03",X"BD",X"15",X"1F",X"8E",X"BE",X"15",X"C6",
		X"02",X"8D",X"09",X"BD",X"13",X"BD",X"BD",X"15",X"15",X"7E",X"D0",X"03",X"35",X"20",X"10",X"BF",
		X"BE",X"BB",X"9F",X"69",X"D7",X"67",X"BD",X"EE",X"63",X"24",X"50",X"BD",X"EE",X"1C",X"10",X"8E",
		X"CD",X"6E",X"8E",X"CF",X"90",X"BD",X"ED",X"F6",X"8E",X"CD",X"66",X"10",X"8E",X"CD",X"74",X"86",
		X"08",X"BD",X"EC",X"62",X"8E",X"CD",X"38",X"10",X"8E",X"CD",X"6E",X"86",X"06",X"BD",X"EC",X"62",
		X"10",X"8E",X"CD",X"6E",X"BD",X"EB",X"51",X"9E",X"69",X"10",X"8E",X"CD",X"66",X"C6",X"04",X"BD",
		X"E0",X"0C",X"BD",X"EB",X"32",X"8E",X"EB",X"0F",X"10",X"8E",X"CD",X"38",X"C6",X"03",X"BD",X"E0",
		X"0C",X"BD",X"13",X"BD",X"86",X"89",X"B7",X"BE",X"BD",X"20",X"22",X"BD",X"EE",X"6F",X"25",X"09",
		X"BD",X"EE",X"8B",X"25",X"04",X"6E",X"9F",X"BE",X"BB",X"7F",X"BE",X"BD",X"CC",X"EB",X"1E",X"10",
		X"8C",X"CF",X"9E",X"26",X"03",X"CC",X"EB",X"16",X"BD",X"06",X"FD",X"86",X"88",X"D6",X"67",X"0C",
		X"F8",X"BD",X"13",X"BD",X"BD",X"70",X"55",X"CC",X"3A",X"3A",X"FD",X"A1",X"00",X"B7",X"A1",X"02",
		X"CC",X"03",X"00",X"8E",X"46",X"80",X"10",X"8E",X"A1",X"00",X"BD",X"E0",X"09",X"BD",X"EE",X"6F",
		X"24",X"06",X"8E",X"CF",X"E4",X"BD",X"ED",X"DD",X"BD",X"EE",X"8B",X"24",X"43",X"7D",X"BE",X"BD",
		X"27",X"1C",X"8E",X"A1",X"00",X"10",X"8E",X"CD",X"38",X"C6",X"03",X"BD",X"E0",X"0C",X"BD",X"EB",
		X"32",X"86",X"05",X"8D",X"2F",X"24",X"29",X"1F",X"12",X"BD",X"EC",X"42",X"20",X"12",X"BD",X"ED",
		X"98",X"34",X"01",X"34",X"10",X"10",X"AC",X"E1",X"22",X"02",X"8D",X"61",X"35",X"01",X"24",X"10",
		X"BD",X"13",X"BD",X"86",X"94",X"BD",X"70",X"55",X"86",X"60",X"8E",X"ED",X"90",X"7E",X"00",X"A8",
		X"6E",X"9F",X"BE",X"BB",X"34",X"26",X"20",X"0C",X"34",X"26",X"8E",X"CD",X"38",X"8D",X"24",X"86",
		X"04",X"25",X"01",X"4C",X"97",X"4F",X"8E",X"CD",X"6E",X"8D",X"18",X"24",X"04",X"0A",X"4F",X"27",
		X"0E",X"30",X"0E",X"8C",X"CF",X"9E",X"25",X"F1",X"8E",X"CF",X"90",X"1C",X"FE",X"35",X"A6",X"1A",
		X"01",X"35",X"A6",X"34",X"10",X"10",X"8E",X"A1",X"00",X"C6",X"03",X"BD",X"14",X"0B",X"A1",X"A0",
		X"26",X"07",X"5A",X"26",X"F6",X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",X"34",X"20",X"BD",
		X"ED",X"F6",X"8E",X"A1",X"00",X"C6",X"03",X"BD",X"E0",X"0C",X"9E",X"69",X"C6",X"04",X"BD",X"E0",
		X"0C",X"35",X"20",X"7E",X"EB",X"51",X"34",X"30",X"1F",X"12",X"10",X"AC",X"62",X"27",X"0B",X"30",
		X"32",X"86",X"0E",X"BD",X"EC",X"62",X"31",X"32",X"20",X"F0",X"35",X"B0",X"35",X"06",X"FD",X"BE",
		X"BB",X"C6",X"01",X"8D",X"07",X"BD",X"EB",X"32",X"6E",X"9F",X"BE",X"BB",X"35",X"20",X"10",X"BF",
		X"BE",X"BD",X"4F",X"1F",X"02",X"CC",X"EB",X"16",X"BD",X"06",X"FD",X"8E",X"CC",X"28",X"BD",X"14",
		X"1C",X"86",X"87",X"BD",X"13",X"BD",X"BD",X"70",X"55",X"1F",X"98",X"BD",X"08",X"D1",X"8E",X"2D",
		X"80",X"10",X"8E",X"A1",X"14",X"C6",X"3A",X"E7",X"A2",X"10",X"8C",X"A1",X"00",X"22",X"F8",X"5F",
		X"BD",X"E0",X"09",X"8E",X"A1",X"00",X"10",X"8E",X"CD",X"3E",X"C6",X"14",X"BD",X"E0",X"0C",X"6E",
		X"9F",X"BE",X"BD",X"34",X"30",X"10",X"8E",X"CD",X"66",X"9E",X"69",X"8D",X"36",X"35",X"B0",X"34",
		X"10",X"10",X"8E",X"CF",X"A4",X"9E",X"69",X"8D",X"2A",X"25",X"0C",X"31",X"2E",X"10",X"8C",X"CF",
		X"F2",X"25",X"F4",X"1C",X"FE",X"35",X"90",X"31",X"3A",X"35",X"90",X"34",X"10",X"10",X"8E",X"CD",
		X"66",X"9E",X"69",X"8D",X"0E",X"25",X"F0",X"31",X"2E",X"10",X"8C",X"CF",X"90",X"25",X"F4",X"1C",
		X"FE",X"35",X"90",X"34",X"36",X"1E",X"12",X"C6",X"04",X"BD",X"14",X"0B",X"C1",X"04",X"26",X"02",
		X"84",X"0F",X"A1",X"A0",X"22",X"05",X"25",X"07",X"5A",X"26",X"EE",X"1C",X"FE",X"35",X"B6",X"1A",
		X"01",X"35",X"B6",X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"2D",X"20",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"28",X"43",X"29",X"20",X"31",X"39",
		X"38",X"31",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",
		X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",
		X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",
		X"44",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",
		X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"31",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",
		X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"F4",X"95",X"7E",X"F4",X"8F",X"7E",X"F4",X"D3",X"7E",X"F5",X"42",X"7E",X"F6",X"9E",X"34",
		X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"0F",X"58",X"34",X"04",X"58",X"EB",X"E0",X"8E",
		X"CC",X"FC",X"3A",X"BD",X"14",X"1C",X"34",X"04",X"BD",X"14",X"1C",X"34",X"04",X"BD",X"14",X"1C",
		X"34",X"04",X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",
		X"89",X"00",X"19",X"30",X"1A",X"BD",X"14",X"24",X"35",X"04",X"35",X"02",X"BD",X"14",X"30",X"35",
		X"02",X"35",X"96",X"1A",X"FF",X"10",X"CE",X"BF",X"FF",X"7F",X"C8",X"0D",X"7F",X"C8",X"0C",X"86",
		X"3C",X"B7",X"C8",X"0D",X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",X"B7",X"C8",
		X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"1F",X"D2",X"10",X"8E",
		X"C0",X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"1F",X"E2",X"25",X"F7",X"86",X"02",X"10",X"8E",X"F5",
		X"17",X"8E",X"00",X"00",X"7E",X"FC",X"6D",X"10",X"8E",X"F5",X"1E",X"7E",X"FE",X"4C",X"86",X"34",
		X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"7F",X"C8",X"0E",X"86",X"9C",X"1F",X"8B",X"10",X"CE",X"BF",
		X"FF",X"BD",X"13",X"BD",X"86",X"10",X"BD",X"70",X"55",X"10",X"8E",X"5F",X"D6",X"86",X"07",X"7E",
		X"FD",X"88",X"96",X"F3",X"26",X"0F",X"86",X"02",X"8E",X"F5",X"4E",X"7E",X"00",X"A8",X"B6",X"C8",
		X"0C",X"85",X"02",X"26",X"03",X"7E",X"00",X"E4",X"BD",X"01",X"57",X"BD",X"15",X"15",X"86",X"FF",
		X"97",X"F3",X"97",X"91",X"BD",X"F6",X"8D",X"B6",X"C8",X"0C",X"46",X"10",X"25",X"05",X"D8",X"BD",
		X"13",X"BD",X"1A",X"BF",X"10",X"8E",X"F5",X"7B",X"7E",X"FE",X"1A",X"86",X"39",X"B7",X"CB",X"FF",
		X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"10",X"8E",X"F5",X"8E",X"7E",X"FE",X"4C",X"86",X"9C",
		X"1F",X"8B",X"BD",X"13",X"BD",X"86",X"19",X"BD",X"70",X"55",X"C6",X"03",X"8E",X"70",X"00",X"86",
		X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"16",X"30",X"1F",X"8C",X"00",X"00",
		X"26",X"ED",X"5A",X"26",X"E7",X"10",X"8E",X"F5",X"C1",X"8E",X"00",X"00",X"86",X"FF",X"7E",X"FC",
		X"6D",X"86",X"01",X"B7",X"C9",X"00",X"86",X"9C",X"1F",X"8B",X"BD",X"13",X"BD",X"86",X"1A",X"BD",
		X"70",X"55",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"8E",X"9C",
		X"00",X"6F",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"C0",X"00",X"26",X"F4",X"CC",X"A5",X"5A",
		X"DD",X"B7",X"97",X"F3",X"BD",X"08",X"0B",X"BD",X"5F",X"E7",X"BD",X"15",X"15",X"03",X"91",X"BD",
		X"19",X"43",X"F6",X"0B",X"8D",X"7A",X"1C",X"00",X"7E",X"00",X"0C",X"BD",X"FB",X"0C",X"BD",X"FC",
		X"08",X"1C",X"01",X"86",X"1B",X"24",X"28",X"C6",X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",
		X"1A",X"10",X"10",X"CE",X"F6",X"2B",X"86",X"03",X"7E",X"FD",X"9C",X"10",X"CE",X"BF",X"FF",X"8D",
		X"4F",X"86",X"9C",X"1F",X"8B",X"1C",X"EF",X"86",X"1C",X"C1",X"1F",X"22",X"02",X"86",X"1D",X"BD",
		X"13",X"BD",X"BD",X"70",X"55",X"DE",X"3F",X"BD",X"FB",X"0C",X"6F",X"49",X"BD",X"FB",X"98",X"BD",
		X"FB",X"A1",X"BD",X"FB",X"3A",X"24",X"F8",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"F6",
		X"64",X"7E",X"00",X"A8",X"86",X"0C",X"B7",X"C8",X"0E",X"BD",X"FB",X"0C",X"BD",X"F9",X"85",X"BD",
		X"FB",X"0C",X"BD",X"F8",X"E2",X"BD",X"FB",X"3A",X"24",X"03",X"BD",X"FB",X"0C",X"7E",X"F6",X"E8",
		X"7F",X"C8",X"0E",X"86",X"34",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"39",X"8E",X"1F",X"D2",
		X"10",X"8E",X"9C",X"26",X"EC",X"81",X"ED",X"A1",X"8C",X"1F",X"E2",X"25",X"F7",X"39",X"86",X"3F",
		X"1F",X"8A",X"86",X"8F",X"BE",X"A3",X"00",X"30",X"89",X"12",X"34",X"10",X"8E",X"F6",X"B2",X"7E",
		X"FC",X"6D",X"10",X"8E",X"F6",X"B9",X"7E",X"FE",X"4C",X"86",X"9C",X"1F",X"8B",X"10",X"CE",X"BF",
		X"FF",X"BD",X"FC",X"08",X"24",X"16",X"86",X"1D",X"8C",X"CD",X"00",X"23",X"02",X"86",X"1C",X"BD",
		X"13",X"BD",X"BD",X"70",X"55",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"F9",X"BD",X"F7",X"0F",X"10",
		X"8E",X"F6",X"9E",X"86",X"04",X"7E",X"FD",X"88",X"BD",X"F7",X"64",X"BD",X"FB",X"0C",X"BD",X"13",
		X"BD",X"86",X"07",X"97",X"26",X"BD",X"FB",X"0C",X"86",X"38",X"97",X"26",X"BD",X"FB",X"0C",X"86",
		X"C0",X"97",X"26",X"BD",X"FB",X"0C",X"BD",X"F7",X"0F",X"BD",X"FB",X"0C",X"7E",X"FB",X"47",X"8E",
		X"9C",X"26",X"10",X"8E",X"F7",X"54",X"CE",X"C0",X"00",X"EC",X"A1",X"ED",X"81",X"ED",X"C1",X"86",
		X"39",X"B7",X"CB",X"FF",X"8C",X"9C",X"36",X"25",X"F0",X"CC",X"00",X"00",X"8E",X"00",X"00",X"9F",
		X"4F",X"30",X"89",X"0F",X"00",X"ED",X"83",X"34",X"02",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"02",
		X"9C",X"4F",X"26",X"F1",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",
		X"11",X"24",X"DC",X"39",X"05",X"05",X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",
		X"A8",X"A8",X"85",X"85",X"BD",X"13",X"BD",X"4F",X"BD",X"F9",X"7A",X"86",X"FF",X"97",X"27",X"86",
		X"C0",X"97",X"28",X"86",X"38",X"97",X"29",X"86",X"07",X"97",X"2A",X"10",X"8E",X"F8",X"6A",X"CC",
		X"01",X"01",X"AE",X"A4",X"ED",X"81",X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"F8",X"92",
		X"26",X"F0",X"86",X"11",X"10",X"8E",X"F8",X"4A",X"AE",X"A4",X"9F",X"4F",X"A7",X"84",X"0C",X"4F",
		X"9E",X"4F",X"AC",X"22",X"26",X"F6",X"31",X"24",X"10",X"8C",X"F8",X"6A",X"26",X"EA",X"10",X"8E",
		X"F8",X"92",X"AE",X"A4",X"9F",X"4F",X"A6",X"24",X"A7",X"84",X"0C",X"4F",X"9E",X"4F",X"AC",X"22",
		X"26",X"F6",X"31",X"25",X"10",X"8C",X"F8",X"CE",X"26",X"E8",X"10",X"8E",X"F8",X"CE",X"AE",X"A4",
		X"A6",X"24",X"A7",X"80",X"AC",X"22",X"26",X"FA",X"31",X"25",X"10",X"8C",X"F8",X"E2",X"26",X"EE",
		X"86",X"21",X"B7",X"43",X"7E",X"86",X"20",X"B7",X"93",X"7E",X"8E",X"4B",X"0A",X"1A",X"10",X"7F",
		X"C9",X"00",X"A6",X"84",X"C6",X"01",X"F7",X"C9",X"00",X"1C",X"EF",X"84",X"F0",X"8A",X"02",X"A7",
		X"80",X"8C",X"4B",X"6D",X"26",X"E7",X"8E",X"4B",X"90",X"1A",X"10",X"7F",X"C9",X"00",X"A6",X"84",
		X"C6",X"01",X"F7",X"C9",X"00",X"1C",X"EF",X"84",X"F0",X"8A",X"02",X"A7",X"80",X"8C",X"4B",X"F3",
		X"26",X"E7",X"8E",X"0B",X"18",X"9F",X"4F",X"9E",X"4F",X"A6",X"84",X"84",X"F0",X"8A",X"01",X"A7",
		X"84",X"D6",X"50",X"CB",X"22",X"25",X"04",X"D7",X"50",X"20",X"EC",X"C6",X"18",X"D7",X"50",X"D6",
		X"4F",X"CB",X"10",X"D7",X"4F",X"C1",X"9B",X"26",X"DE",X"39",X"04",X"07",X"94",X"07",X"04",X"29",
		X"94",X"29",X"04",X"4B",X"94",X"4B",X"04",X"6D",X"94",X"6D",X"04",X"8F",X"94",X"8F",X"04",X"B1",
		X"94",X"B1",X"04",X"D3",X"94",X"D3",X"04",X"F5",X"94",X"F5",X"03",X"07",X"03",X"F5",X"13",X"07",
		X"13",X"F5",X"23",X"07",X"23",X"F5",X"33",X"07",X"33",X"F5",X"43",X"07",X"43",X"F5",X"53",X"07",
		X"53",X"F5",X"63",X"07",X"63",X"F5",X"73",X"07",X"73",X"F5",X"83",X"07",X"83",X"F5",X"93",X"07",
		X"93",X"F5",X"45",X"05",X"52",X"05",X"44",X"45",X"06",X"52",X"06",X"44",X"45",X"07",X"52",X"07",
		X"00",X"45",X"08",X"52",X"08",X"33",X"45",X"09",X"52",X"09",X"33",X"45",X"F3",X"52",X"F3",X"33",
		X"45",X"F4",X"52",X"F4",X"33",X"45",X"F5",X"52",X"F5",X"00",X"45",X"F6",X"52",X"F6",X"44",X"45",
		X"F7",X"52",X"F7",X"44",X"04",X"7E",X"43",X"7E",X"22",X"54",X"7E",X"93",X"7E",X"22",X"02",X"6F",
		X"02",X"8E",X"04",X"03",X"6F",X"03",X"8E",X"30",X"93",X"6F",X"93",X"8E",X"00",X"94",X"6F",X"94",
		X"8E",X"34",X"35",X"06",X"DE",X"3F",X"ED",X"4D",X"BD",X"13",X"BD",X"86",X"33",X"BD",X"70",X"55",
		X"86",X"80",X"A7",X"47",X"86",X"01",X"8E",X"F8",X"FC",X"7E",X"00",X"A8",X"BD",X"FB",X"3A",X"25",
		X"34",X"6A",X"47",X"26",X"EF",X"B6",X"F9",X"62",X"8D",X"70",X"8D",X"2E",X"8E",X"F9",X"62",X"A6",
		X"80",X"DE",X"3F",X"AF",X"49",X"8D",X"63",X"86",X"80",X"A7",X"47",X"86",X"01",X"8E",X"F9",X"23",
		X"7E",X"00",X"A8",X"BD",X"FB",X"3A",X"25",X"0D",X"6A",X"47",X"26",X"EF",X"AE",X"49",X"8C",X"F9",
		X"6A",X"25",X"DC",X"20",X"D7",X"DE",X"3F",X"6E",X"D8",X"0D",X"8E",X"00",X"00",X"10",X"8E",X"F9",
		X"6A",X"9F",X"4F",X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"9C",X"4F",X"26",
		X"FA",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"10",X"8C",X"F9",X"7A",X"26",
		X"E0",X"39",X"02",X"03",X"04",X"10",X"18",X"20",X"40",X"80",X"00",X"FF",X"11",X"EE",X"22",X"DD",
		X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",X"8E",X"9C",X"26",X"A7",X"80",X"8C",
		X"9C",X"36",X"25",X"F9",X"39",X"35",X"06",X"DE",X"3F",X"ED",X"4D",X"86",X"0A",X"A7",X"4B",X"BD",
		X"13",X"BD",X"86",X"21",X"BD",X"70",X"55",X"CE",X"9D",X"00",X"6F",X"C0",X"11",X"83",X"9D",X"0A",
		X"23",X"F8",X"CE",X"FA",X"3E",X"8D",X"26",X"86",X"34",X"B7",X"C8",X"07",X"8D",X"1F",X"86",X"3C",
		X"B7",X"C8",X"07",X"8D",X"28",X"BD",X"FB",X"3A",X"24",X"06",X"DE",X"3F",X"6A",X"4B",X"27",X"08",
		X"86",X"01",X"8E",X"F9",X"A2",X"7E",X"00",X"A8",X"DE",X"3F",X"6E",X"D8",X"0D",X"AE",X"C1",X"27",
		X"0B",X"10",X"AE",X"C1",X"A6",X"84",X"A8",X"A4",X"A7",X"21",X"20",X"F1",X"39",X"CE",X"FA",X"56",
		X"10",X"8E",X"9D",X"00",X"C6",X"01",X"E5",X"21",X"27",X"02",X"8D",X"19",X"33",X"43",X"58",X"24",
		X"F5",X"31",X"22",X"10",X"8C",X"9D",X"09",X"22",X"0B",X"B6",X"C8",X"06",X"2B",X"E6",X"10",X"8C",
		X"9D",X"05",X"23",X"E0",X"39",X"34",X"14",X"86",X"3F",X"B7",X"C8",X"0E",X"E8",X"A4",X"E7",X"A4",
		X"E6",X"E4",X"E5",X"A4",X"26",X"10",X"E6",X"42",X"27",X"22",X"86",X"40",X"1F",X"01",X"CC",X"30",
		X"06",X"BD",X"13",X"B9",X"35",X"94",X"E6",X"42",X"27",X"12",X"86",X"40",X"1F",X"01",X"C6",X"BB",
		X"D7",X"10",X"EC",X"C4",X"BD",X"70",X"52",X"86",X"17",X"B7",X"C8",X"0E",X"35",X"94",X"C8",X"0C",
		X"9D",X"00",X"C8",X"04",X"9D",X"02",X"C8",X"06",X"9D",X"04",X"00",X"00",X"C8",X"04",X"9D",X"06",
		X"C8",X"06",X"9D",X"08",X"00",X"00",X"22",X"00",X"2C",X"23",X"00",X"33",X"24",X"00",X"3A",X"25",
		X"00",X"41",X"26",X"00",X"48",X"27",X"00",X"4F",X"28",X"00",X"56",X"00",X"00",X"00",X"29",X"01",
		X"5D",X"2A",X"01",X"64",X"2B",X"01",X"6B",X"2C",X"01",X"72",X"2D",X"00",X"79",X"2E",X"00",X"80",
		X"2F",X"01",X"87",X"30",X"01",X"8E",X"31",X"01",X"95",X"32",X"01",X"9C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"29",X"02",
		X"A3",X"2A",X"02",X"AA",X"2B",X"02",X"B1",X"2C",X"02",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2F",X"02",X"BF",X"30",X"02",X"C6",X"31",X"02",X"CD",X"32",X"02",X"D4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F5",
		X"DE",X"20",X"03",X"CE",X"F5",X"B5",X"10",X"CE",X"BF",X"FF",X"10",X"8E",X"FA",X"E3",X"86",X"01",
		X"7E",X"FD",X"88",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"10",X"8E",X"FA",X"F3",X"86",X"01",
		X"7E",X"FD",X"88",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F0",X"10",X"8E",X"FB",X"03",X"86",X"01",
		X"7E",X"FD",X"88",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"6E",X"C4",X"35",X"06",X"DE",X"3F",
		X"ED",X"4D",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"08",X"86",X"01",X"8E",X"FB",X"12",X"7E",X"00",
		X"A8",X"0F",X"26",X"BD",X"13",X"BD",X"20",X"07",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"08",X"86",
		X"02",X"8E",X"FB",X"28",X"7E",X"00",X"A8",X"6E",X"D8",X"0D",X"B6",X"C8",X"0C",X"85",X"02",X"27",
		X"03",X"1A",X"01",X"39",X"1C",X"FE",X"39",X"86",X"FF",X"97",X"91",X"BD",X"F6",X"8D",X"BD",X"FB",
		X"3A",X"24",X"03",X"BD",X"FB",X"0C",X"86",X"34",X"BD",X"70",X"55",X"CE",X"CD",X"02",X"86",X"35",
		X"34",X"02",X"BD",X"70",X"55",X"1E",X"31",X"BD",X"14",X"1C",X"34",X"04",X"BD",X"14",X"1A",X"1F",
		X"02",X"35",X"04",X"1E",X"31",X"5D",X"27",X"0C",X"86",X"3E",X"BD",X"70",X"55",X"86",X"3F",X"BD",
		X"70",X"55",X"20",X"05",X"86",X"40",X"BD",X"70",X"55",X"35",X"02",X"4C",X"11",X"83",X"CD",X"32",
		X"23",X"CE",X"BD",X"FB",X"0C",X"7E",X"E0",X"00",X"BD",X"13",X"BD",X"CC",X"FE",X"01",X"ED",X"47",
		X"39",X"35",X"06",X"ED",X"4D",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"FB",X"B2",X"7E",
		X"00",X"A8",X"86",X"0C",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"FB",X"BF",X"7E",X"00",X"A8",X"86",
		X"3F",X"B7",X"C8",X"0E",X"86",X"01",X"8E",X"FB",X"CC",X"7E",X"00",X"A8",X"EC",X"47",X"84",X"3F",
		X"B7",X"C8",X"0E",X"86",X"1E",X"BD",X"70",X"55",X"86",X"40",X"A7",X"4B",X"86",X"01",X"8E",X"FB",
		X"E4",X"7E",X"00",X"A8",X"BD",X"FB",X"3A",X"25",X"04",X"6A",X"4B",X"26",X"EF",X"A6",X"49",X"26",
		X"06",X"B6",X"C8",X"0C",X"46",X"24",X"0E",X"EC",X"47",X"1A",X"01",X"49",X"5C",X"C1",X"06",X"25",
		X"02",X"8D",X"98",X"ED",X"47",X"6E",X"D8",X"0D",X"8E",X"CC",X"00",X"10",X"8E",X"9D",X"00",X"A6",
		X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",X"C6",X"06",X"1A",X"3F",X"DE",X"B7",X"10",X"9E",
		X"B6",X"8E",X"CC",X"00",X"BD",X"07",X"EC",X"A7",X"80",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",
		X"00",X"26",X"F1",X"10",X"9F",X"B6",X"DF",X"B7",X"8E",X"CC",X"00",X"BD",X"07",X"EC",X"A8",X"80",
		X"84",X"0F",X"26",X"24",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"ED",X"5A",X"26",
		X"CB",X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"9D",X"00",X"10",X"8E",X"CC",X"00",X"A6",X"C0",X"A7",
		X"A0",X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",X"8D",X"EC",X"1A",X"01",X"39",X"1A",X"3F",X"7F",
		X"C9",X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",
		X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",
		X"ED",X"81",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",
		X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",
		X"00",X"26",X"C8",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",
		X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"10",X"A3",X"81",
		X"26",X"43",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",
		X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",X"8C",X"C0",
		X"00",X"26",X"C5",X"1F",X"03",X"1F",X"B8",X"81",X"FF",X"26",X"05",X"1F",X"30",X"7E",X"FC",X"78",
		X"4A",X"1F",X"8B",X"81",X"80",X"27",X"07",X"4D",X"1F",X"30",X"10",X"26",X"FF",X"6A",X"C6",X"01",
		X"F7",X"C9",X"00",X"6E",X"A4",X"30",X"1E",X"A8",X"84",X"E8",X"01",X"4D",X"26",X"07",X"5D",X"26",
		X"04",X"30",X"02",X"20",X"AD",X"CE",X"00",X"30",X"1E",X"10",X"5F",X"1E",X"10",X"8C",X"00",X"00",
		X"27",X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",X"10",X"11",X"83",X"00",X"30",X"23",X"EE",X"CE",
		X"00",X"10",X"20",X"E9",X"33",X"41",X"47",X"25",X"05",X"57",X"25",X"02",X"20",X"F6",X"1F",X"30",
		X"86",X"01",X"B7",X"C9",X"00",X"10",X"CE",X"FD",X"5C",X"7E",X"FD",X"9C",X"86",X"9C",X"1F",X"8B",
		X"1F",X"A8",X"43",X"85",X"C0",X"27",X"04",X"86",X"20",X"20",X"02",X"86",X"11",X"10",X"CE",X"BF",
		X"FF",X"BD",X"13",X"BD",X"BD",X"70",X"55",X"1F",X"A8",X"85",X"40",X"26",X"03",X"7E",X"FA",X"CE",
		X"10",X"8E",X"5F",X"D6",X"20",X"00",X"86",X"20",X"8E",X"58",X"00",X"30",X"1F",X"C6",X"39",X"F7",
		X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",X"EE",X"6E",X"A4",X"1F",X"03",X"86",X"02",
		X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"FD",X"AB",X"7E",X"FE",X"2A",X"86",X"02",X"10",X"8E",X"FD",
		X"B4",X"7E",X"FD",X"88",X"10",X"8E",X"FD",X"BB",X"7E",X"FE",X"1A",X"86",X"01",X"10",X"8E",X"FD",
		X"C4",X"7E",X"FD",X"88",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",X"8E",X"FD",X"D2",
		X"20",X"58",X"86",X"02",X"10",X"8E",X"FD",X"DA",X"20",X"AE",X"10",X"8E",X"FD",X"E0",X"20",X"3A",
		X"86",X"01",X"10",X"8E",X"FD",X"E8",X"20",X"A0",X"1F",X"30",X"1F",X"98",X"10",X"8E",X"FD",X"F2",
		X"20",X"38",X"86",X"02",X"10",X"8E",X"FD",X"FA",X"20",X"8E",X"10",X"8E",X"FE",X"00",X"20",X"1A",
		X"86",X"05",X"10",X"8E",X"FE",X"09",X"7E",X"FD",X"88",X"1F",X"B8",X"4A",X"1F",X"8B",X"26",X"92",
		X"10",X"8E",X"FE",X"16",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",X"B7",X"C8",X"0D",X"4C",
		X"B7",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",X"46",X"46",X"46",X"84",
		X"C0",X"B7",X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0F",X"86",
		X"34",X"C5",X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",X"1A",X"3F",X"8E",X"FE",
		X"C2",X"8C",X"FE",X"E2",X"27",X"6A",X"A6",X"01",X"27",X"18",X"A6",X"84",X"5F",X"1F",X"03",X"86",
		X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",X"1E",X"03",X"26",X"F3",X"E1",X"01",
		X"26",X"04",X"30",X"02",X"20",X"DB",X"A6",X"84",X"44",X"44",X"44",X"44",X"81",X"0D",X"25",X"02",
		X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",X"CE",X"FE",X"90",X"7E",X"FD",X"9C",
		X"86",X"9C",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"BF",X"FF",X"BD",X"13",X"BD",
		X"1F",X"A8",X"43",X"85",X"C0",X"27",X"04",X"86",X"1F",X"20",X"02",X"86",X"12",X"BD",X"70",X"55",
		X"1F",X"A9",X"C5",X"40",X"26",X"03",X"7E",X"FA",X"D3",X"10",X"8E",X"5F",X"D6",X"7E",X"FD",X"86",
		X"6E",X"A4",X"00",X"BC",X"10",X"0B",X"20",X"CA",X"30",X"21",X"40",X"FB",X"50",X"97",X"60",X"43",
		X"70",X"B3",X"80",X"15",X"90",X"00",X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",X"2F",X"E0",X"1F",
		X"F0",X"01",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F4",X"86",X"F4",X"86",X"F4",X"86",X"F4",X"86",X"9C",X"6B",X"F4",X"86",X"F4",X"86",X"F4",X"86",
		X"34",X"76",X"EC",X"04",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"35",X"F6",X"8E",X"9C",X"3B",X"9F",
		X"3F",X"96",X"39",X"27",X"FC",X"0F",X"39",X"D6",X"91",X"C5",X"69",X"27",X"04",X"0F",X"3A",X"20",
		X"46",X"48",X"9B",X"3A",X"80",X"04",X"2A",X"01",X"4F",X"97",X"3A",X"81",X"02",X"25",X"38",X"C6",
		X"03",X"D7",X"88",X"81",X"02",X"23",X"30",X"86",X"02",X"97",X"3A",X"10",X"8E",X"9C",X"41",X"AE",
		X"A4",X"27",X"24",X"A6",X"88",X"14",X"27",X"04",X"31",X"84",X"20",X"F3",X"EE",X"84",X"EF",X"A4",
		X"DC",X"B6",X"84",X"3F",X"8B",X"60",X"E3",X"0A",X"ED",X"0A",X"8D",X"A4",X"CC",X"00",X"00",X"ED",
		X"04",X"DE",X"47",X"9F",X"47",X"EF",X"84",X"8D",X"50",X"BD",X"27",X"06",X"BD",X"07",X"EC",X"BD",
		X"37",X"46",X"96",X"59",X"85",X"02",X"7E",X"2B",X"70",X"12",X"12",X"9E",X"5E",X"26",X"0C",X"9E",
		X"62",X"27",X"17",X"DC",X"64",X"0F",X"62",X"0F",X"63",X"20",X"06",X"DC",X"60",X"0F",X"5E",X"0F",
		X"5F",X"D4",X"91",X"26",X"E6",X"BD",X"01",X"30",X"20",X"E1",X"CE",X"9C",X"3B",X"20",X"0F",X"6A",
		X"44",X"26",X"0B",X"DF",X"3F",X"6E",X"D8",X"02",X"DE",X"3F",X"A7",X"44",X"AF",X"42",X"EE",X"C4",
		X"26",X"ED",X"10",X"CE",X"BF",X"FF",X"7E",X"00",X"0C",X"96",X"91",X"85",X"09",X"26",X"22",X"DC",
		X"96",X"CE",X"20",X"A9",X"0D",X"94",X"2A",X"03",X"CE",X"20",X"B3",X"34",X"46",X"0C",X"B5",X"BD",
		X"0F",X"07",X"35",X"46",X"26",X"08",X"8E",X"9C",X"49",X"BD",X"0F",X"0A",X"27",X"03",X"BD",X"5F",
		X"B8",X"0F",X"B5",X"39",X"9E",X"3F",X"8D",X"06",X"33",X"84",X"20",X"C2",X"AE",X"06",X"34",X"46",
		X"CE",X"9C",X"3B",X"AC",X"C4",X"26",X"18",X"EC",X"84",X"ED",X"C4",X"A6",X"06",X"27",X"06",X"DC",
		X"45",X"9F",X"45",X"20",X"04",X"DC",X"3D",X"9F",X"3D",X"ED",X"84",X"30",X"C4",X"35",X"C6",X"EE",
		X"C4",X"26",X"E0",X"8D",X"00",X"1A",X"10",X"20",X"FE",X"34",X"62",X"DE",X"45",X"26",X"01",X"BD",
		X"01",X"15",X"10",X"AE",X"C4",X"10",X"9F",X"45",X"86",X"01",X"A7",X"46",X"A6",X"E4",X"20",X"11",
		X"34",X"62",X"DE",X"3D",X"26",X"03",X"BD",X"01",X"15",X"10",X"AE",X"C4",X"10",X"9F",X"3D",X"6F",
		X"46",X"AF",X"42",X"A7",X"45",X"86",X"01",X"A7",X"44",X"AE",X"9F",X"9C",X"3F",X"EF",X"9F",X"9C",
		X"3F",X"AF",X"C4",X"30",X"C4",X"35",X"E2",X"34",X"12",X"8E",X"9C",X"3B",X"AE",X"84",X"27",X"0E",
		X"9C",X"3F",X"27",X"F8",X"A6",X"05",X"81",X"02",X"27",X"F2",X"8D",X"82",X"20",X"EE",X"35",X"92",
		X"8D",X"16",X"34",X"66",X"EF",X"06",X"EE",X"66",X"37",X"26",X"ED",X"02",X"10",X"AF",X"08",X"37",
		X"06",X"ED",X"88",X"12",X"EF",X"66",X"35",X"E6",X"34",X"46",X"9E",X"43",X"26",X"03",X"BD",X"01",
		X"15",X"EC",X"84",X"DD",X"43",X"DC",X"41",X"ED",X"84",X"4F",X"5F",X"ED",X"04",X"A7",X"88",X"14",
		X"35",X"C6",X"34",X"70",X"CE",X"9C",X"41",X"AC",X"C4",X"26",X"10",X"10",X"AE",X"D4",X"10",X"AF",
		X"C4",X"10",X"9E",X"43",X"9F",X"43",X"10",X"AF",X"84",X"35",X"F0",X"EE",X"C4",X"26",X"E8",X"CE",
		X"9C",X"47",X"AC",X"C4",X"27",X"E5",X"EE",X"C4",X"26",X"F8",X"BD",X"01",X"15",X"34",X"70",X"CE",
		X"9C",X"49",X"20",X"EE",X"34",X"18",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",
		X"CB",X"08",X"1F",X"03",X"20",X"4E",X"34",X"18",X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",
		X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"20",X"6A",X"34",X"18",X"CB",X"08",X"1F",X"03",
		X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"36",X"3F",X"33",X"C9",
		X"01",X"08",X"20",X"44",X"34",X"18",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",
		X"CB",X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"35",X"3F",X"36",X"3F",
		X"33",X"C9",X"01",X"08",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"35",X"3F",X"36",X"3F",
		X"10",X"FE",X"9C",X"53",X"35",X"98",X"34",X"18",X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",
		X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",X"3F",
		X"33",X"C9",X"01",X"08",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",X"3F",X"35",X"98",X"34",X"18",
		X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"08",X"1F",X"03",X"35",X"3F",
		X"36",X"3F",X"33",X"C9",X"01",X"08",X"20",X"9C",X"24",X"02",X"31",X"22",X"10",X"AE",X"22",X"1F",
		X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",X"ED",X"42",X"EC",X"24",X"ED",X"C9",X"01",X"00",X"EC",
		X"26",X"ED",X"C9",X"01",X"02",X"EC",X"28",X"ED",X"C9",X"02",X"00",X"EC",X"2A",X"ED",X"C9",X"02",
		X"02",X"39",X"1F",X"03",X"CC",X"00",X"00",X"ED",X"C4",X"ED",X"42",X"ED",X"C9",X"01",X"00",X"ED",
		X"C9",X"01",X"02",X"ED",X"C9",X"02",X"00",X"ED",X"C9",X"02",X"02",X"39",X"24",X"02",X"31",X"22",
		X"10",X"AE",X"22",X"1F",X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",X"A7",X"42",X"E7",X"C9",X"01",
		X"00",X"EC",X"24",X"ED",X"C9",X"01",X"01",X"39",X"1F",X"03",X"CC",X"00",X"00",X"ED",X"C4",X"A7",
		X"42",X"ED",X"C9",X"01",X"00",X"A7",X"C9",X"01",X"02",X"39",X"34",X"56",X"10",X"DF",X"53",X"24",
		X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"04",X"1F",X"03",X"35",X"16",X"36",X"16",X"33",X"C9",
		X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",
		X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",
		X"01",X"04",X"35",X"16",X"36",X"16",X"10",X"DE",X"53",X"35",X"D6",X"34",X"56",X"CB",X"04",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"33",
		X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",
		X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"35",X"D6",X"34",X"10",X"10",X"DF",X"53",X"24",X"02",
		X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"35",X"36",X"36",X"36",X"10",X"DE",X"53",X"35",X"90",X"34",X"10",X"CB",X"06",X"1F",X"03",
		X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",
		X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",
		X"01",X"06",X"36",X"36",X"35",X"90",X"34",X"10",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",
		X"EE",X"22",X"CB",X"06",X"1F",X"03",X"20",X"89",X"34",X"10",X"CB",X"06",X"1F",X"03",X"CC",X"00",
		X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"C2",X"34",X"10",X"10",X"DF",X"53",X"24",X"02",X"31",
		X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"7E",X"03",X"89",X"34",X"10",X"CB",X"06",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"99",X"34",X"10",X"10",X"DF",X"53",
		X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"07",X"1F",X"03",X"20",X"2A",X"34",X"10",X"CB",
		X"07",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1C",X"00",X"20",X"4F",X"34",
		X"10",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"07",X"1F",X"03",X"35",
		X"37",X"36",X"37",X"33",X"C9",X"01",X"07",X"35",X"37",X"36",X"37",X"33",X"C9",X"01",X"07",X"35",
		X"37",X"36",X"37",X"33",X"C9",X"01",X"07",X"35",X"37",X"36",X"37",X"33",X"C9",X"01",X"07",X"35",
		X"37",X"36",X"37",X"10",X"DE",X"53",X"35",X"90",X"34",X"10",X"CB",X"07",X"1F",X"03",X"CC",X"00",
		X"00",X"8E",X"00",X"00",X"31",X"84",X"1C",X"00",X"36",X"37",X"33",X"C9",X"01",X"07",X"36",X"37",
		X"33",X"C9",X"01",X"07",X"36",X"37",X"33",X"C9",X"01",X"07",X"36",X"37",X"33",X"C9",X"01",X"07",
		X"36",X"37",X"35",X"90",X"34",X"18",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",
		X"CB",X"09",X"1F",X"03",X"A6",X"E0",X"A7",X"57",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",
		X"A6",X"E0",X"A7",X"57",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"A6",X"E0",X"A7",X"57",
		X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"A6",X"E0",X"A7",X"57",X"35",X"3F",X"36",X"3F",
		X"33",X"C9",X"01",X"08",X"A6",X"E0",X"A7",X"57",X"35",X"3F",X"36",X"3F",X"10",X"FE",X"9C",X"53",
		X"35",X"98",X"34",X"10",X"CB",X"09",X"1F",X"03",X"8E",X"00",X"00",X"31",X"84",X"4F",X"36",X"32",
		X"36",X"30",X"33",X"C9",X"01",X"09",X"36",X"32",X"36",X"30",X"33",X"C9",X"01",X"09",X"36",X"32",
		X"36",X"30",X"33",X"C9",X"01",X"09",X"36",X"32",X"36",X"30",X"33",X"C9",X"01",X"09",X"36",X"32",
		X"36",X"30",X"35",X"90",X"34",X"10",X"10",X"DF",X"53",X"25",X"09",X"10",X"EE",X"22",X"CB",X"05",
		X"1F",X"03",X"20",X"0F",X"10",X"EE",X"24",X"CB",X"05",X"1F",X"03",X"35",X"32",X"36",X"32",X"33",
		X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"33",
		X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"10",X"DE",X"53",X"35",X"90",X"34",X"12",X"9B",X"36",
		X"19",X"24",X"02",X"86",X"99",X"97",X"36",X"8E",X"CD",X"00",X"BD",X"14",X"24",X"35",X"92",X"34",
		X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",X"C6",X"01",X"BD",
		X"F4",X"83",X"58",X"8E",X"CC",X"06",X"3A",X"BD",X"14",X"1C",X"8D",X"62",X"96",X"38",X"34",X"04",
		X"AB",X"E4",X"97",X"38",X"96",X"37",X"AB",X"E0",X"97",X"37",X"8E",X"CC",X"12",X"BD",X"14",X"1C",
		X"8D",X"4C",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",X"96",X"8E",X"CC",X"0E",X"BD",X"14",X"1C",
		X"8D",X"3C",X"8D",X"24",X"34",X"02",X"D7",X"37",X"8E",X"CC",X"10",X"BD",X"14",X"1C",X"96",X"38",
		X"8D",X"2C",X"8D",X"14",X"4D",X"27",X"04",X"0F",X"37",X"0F",X"38",X"AB",X"E0",X"19",X"C6",X"04",
		X"BD",X"F4",X"80",X"BD",X"05",X"7C",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",
		X"1E",X"89",X"86",X"99",X"8B",X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",
		X"1E",X"89",X"5F",X"4D",X"26",X"02",X"35",X"82",X"8B",X"99",X"19",X"5C",X"20",X"F5",X"8E",X"9C",
		X"5B",X"10",X"8E",X"05",X"9B",X"20",X"10",X"8E",X"9C",X"5C",X"10",X"8E",X"05",X"8F",X"20",X"07",
		X"8E",X"9C",X"5D",X"10",X"8E",X"05",X"95",X"96",X"5A",X"26",X"20",X"A6",X"84",X"26",X"1C",X"86",
		X"16",X"A7",X"84",X"10",X"AF",X"49",X"86",X"0A",X"8E",X"06",X"4E",X"7E",X"00",X"A8",X"96",X"5A",
		X"26",X"09",X"CC",X"06",X"5E",X"BD",X"06",X"FD",X"AD",X"D8",X"09",X"7E",X"00",X"E4",X"FF",X"01",
		X"18",X"19",X"00",X"EF",X"01",X"20",X"1E",X"00",X"EE",X"02",X"08",X"11",X"01",X"20",X"17",X"00",
		X"F0",X"01",X"40",X"0A",X"00",X"F0",X"01",X"10",X"0B",X"00",X"E8",X"01",X"04",X"14",X"02",X"06",
		X"11",X"02",X"0A",X"17",X"00",X"E8",X"06",X"04",X"11",X"01",X"10",X"17",X"00",X"E0",X"03",X"0A",
		X"08",X"00",X"E0",X"01",X"18",X"1F",X"00",X"E0",X"01",X"18",X"11",X"00",X"D8",X"01",X"10",X"1A",
		X"00",X"D0",X"01",X"30",X"15",X"00",X"D0",X"01",X"10",X"05",X"00",X"D0",X"01",X"08",X"17",X"00",
		X"D0",X"01",X"08",X"07",X"00",X"D0",X"01",X"0A",X"01",X"00",X"D0",X"01",X"0A",X"06",X"00",X"E1",
		X"01",X"10",X"0B",X"00",X"C8",X"0A",X"01",X"0E",X"00",X"C0",X"01",X"08",X"07",X"00",X"C0",X"01",
		X"30",X"14",X"00",X"C0",X"01",X"20",X"18",X"00",X"C0",X"01",X"08",X"03",X"00",X"C0",X"01",X"30",
		X"09",X"00",X"C0",X"01",X"08",X"03",X"00",X"C0",X"01",X"18",X"0C",X"00",X"34",X"07",X"1A",X"FF",
		X"86",X"3F",X"B7",X"C8",X"0E",X"53",X"C4",X"3F",X"F7",X"C8",X"0E",X"35",X"87",X"7E",X"26",X"46",
		X"12",X"1F",X"01",X"A6",X"84",X"91",X"8C",X"25",X"0D",X"97",X"8C",X"30",X"1E",X"1A",X"10",X"9F",
		X"8A",X"CC",X"01",X"01",X"DD",X"8D",X"35",X"97",X"96",X"8D",X"27",X"14",X"0A",X"8D",X"26",X"38",
		X"9E",X"8A",X"0A",X"8E",X"26",X"2C",X"30",X"03",X"9F",X"8A",X"A6",X"84",X"26",X"22",X"97",X"8C",
		X"96",X"57",X"85",X"02",X"26",X"0A",X"96",X"87",X"27",X"1E",X"0F",X"87",X"C6",X"0F",X"20",X"16",
		X"96",X"87",X"26",X"14",X"96",X"91",X"85",X"98",X"26",X"0E",X"C6",X"16",X"D7",X"87",X"20",X"06",
		X"97",X"8E",X"EC",X"01",X"97",X"8D",X"8D",X"94",X"B6",X"C8",X"0C",X"85",X"40",X"27",X"04",X"86",
		X"3C",X"97",X"5A",X"96",X"5A",X"27",X"02",X"0A",X"5A",X"96",X"5B",X"27",X"02",X"0A",X"5B",X"96",
		X"5D",X"27",X"02",X"0A",X"5D",X"96",X"5C",X"27",X"02",X"0A",X"5C",X"96",X"57",X"9A",X"58",X"43",
		X"D6",X"57",X"D7",X"58",X"7E",X"26",X"5C",X"D7",X"57",X"F6",X"C8",X"06",X"D7",X"59",X"94",X"57",
		X"27",X"1B",X"CE",X"5F",X"7C",X"5F",X"CB",X"04",X"44",X"24",X"FB",X"34",X"46",X"33",X"C5",X"37",
		X"16",X"DE",X"5E",X"7E",X"2B",X"B2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"55",X"9A",
		X"56",X"43",X"D6",X"55",X"D7",X"56",X"F6",X"C8",X"0C",X"C4",X"3F",X"D7",X"55",X"95",X"55",X"27",
		X"17",X"8E",X"00",X"78",X"30",X"1F",X"26",X"FC",X"F6",X"C8",X"0C",X"D4",X"55",X"D7",X"55",X"94",
		X"55",X"27",X"05",X"CE",X"5F",X"9C",X"8D",X"BD",X"39",X"34",X"02",X"96",X"67",X"8E",X"BD",X"D6",
		X"4A",X"27",X"03",X"8E",X"BE",X"15",X"35",X"82",X"34",X"02",X"20",X"F1",X"34",X"04",X"D6",X"B6",
		X"86",X"03",X"3D",X"CB",X"11",X"96",X"B8",X"44",X"44",X"44",X"98",X"B8",X"44",X"06",X"B7",X"06",
		X"B8",X"DB",X"B8",X"D9",X"B7",X"D7",X"B6",X"96",X"B6",X"35",X"84",X"34",X"16",X"4F",X"5F",X"8E",
		X"B5",X"F5",X"9F",X"3D",X"30",X"0F",X"AF",X"11",X"8C",X"BA",X"E1",X"26",X"F7",X"ED",X"84",X"DD",
		X"3B",X"8E",X"BA",X"F0",X"9F",X"45",X"30",X"88",X"17",X"AF",X"88",X"E9",X"8C",X"BB",X"4C",X"26",
		X"F5",X"ED",X"84",X"8E",X"9C",X"3B",X"9F",X"3F",X"35",X"96",X"8E",X"1F",X"D2",X"CE",X"9C",X"26",
		X"C6",X"10",X"A6",X"80",X"A7",X"C0",X"5A",X"26",X"F9",X"39",X"34",X"17",X"1A",X"FF",X"8E",X"AD",
		X"6C",X"9F",X"43",X"30",X"88",X"17",X"AF",X"88",X"E9",X"8C",X"B5",X"DE",X"26",X"F5",X"4F",X"5F",
		X"ED",X"84",X"DD",X"47",X"DD",X"41",X"DD",X"49",X"35",X"97",X"34",X"56",X"EC",X"A4",X"ED",X"C4",
		X"3D",X"30",X"4A",X"AF",X"42",X"30",X"8B",X"AF",X"44",X"34",X"10",X"30",X"8B",X"34",X"10",X"EC",
		X"26",X"ED",X"46",X"EC",X"28",X"ED",X"48",X"AE",X"22",X"33",X"4A",X"8D",X"0E",X"AE",X"24",X"EE",
		X"62",X"EC",X"E4",X"ED",X"62",X"8D",X"04",X"32",X"64",X"35",X"D6",X"EC",X"81",X"85",X"F0",X"27",
		X"02",X"8A",X"F0",X"85",X"0F",X"27",X"02",X"8A",X"0F",X"C5",X"F0",X"27",X"02",X"CA",X"F0",X"C5",
		X"0F",X"27",X"02",X"CA",X"0F",X"84",X"BB",X"C4",X"BB",X"ED",X"C1",X"11",X"A3",X"64",X"25",X"DB",
		X"39",X"34",X"02",X"BD",X"07",X"EC",X"A1",X"E4",X"23",X"03",X"44",X"20",X"F9",X"4C",X"32",X"61",
		X"39",X"34",X"04",X"5F",X"81",X"10",X"25",X"06",X"CB",X"0A",X"80",X"10",X"20",X"F6",X"34",X"04",
		X"AB",X"E0",X"35",X"84",X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",X"19",
		X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"8E",X"BB",X"C3",X"C6",X"10",
		X"D7",X"88",X"5F",X"BD",X"07",X"EC",X"81",X"9C",X"24",X"F9",X"A7",X"84",X"BD",X"07",X"EC",X"81",
		X"A0",X"22",X"F9",X"81",X"2C",X"23",X"F5",X"A7",X"01",X"E7",X"02",X"CB",X"11",X"C4",X"77",X"30",
		X"04",X"8C",X"BC",X"03",X"26",X"DD",X"39",X"96",X"91",X"85",X"20",X"26",X"F9",X"8E",X"BB",X"C3",
		X"DC",X"20",X"C4",X"80",X"DD",X"4B",X"DC",X"22",X"C4",X"80",X"93",X"4B",X"58",X"49",X"97",X"4B",
		X"C6",X"F0",X"96",X"21",X"85",X"40",X"26",X"01",X"53",X"D7",X"4D",X"4F",X"A7",X"94",X"A7",X"98",
		X"04",X"A7",X"98",X"08",X"A7",X"98",X"0C",X"A7",X"98",X"10",X"A7",X"98",X"14",X"A7",X"98",X"18",
		X"A7",X"98",X"1C",X"A7",X"98",X"20",X"A7",X"98",X"24",X"A7",X"98",X"28",X"A7",X"98",X"2C",X"A7",
		X"98",X"30",X"A7",X"98",X"34",X"A7",X"98",X"38",X"A7",X"98",X"3C",X"D6",X"88",X"A6",X"84",X"9B",
		X"4B",X"81",X"9C",X"25",X"0A",X"81",X"C0",X"23",X"04",X"86",X"9B",X"20",X"02",X"86",X"00",X"A7",
		X"84",X"A6",X"02",X"94",X"4D",X"A7",X"98",X"00",X"30",X"04",X"5A",X"26",X"E0",X"D6",X"B6",X"C4",
		X"3C",X"8E",X"BB",X"C3",X"3A",X"A6",X"02",X"8B",X"11",X"84",X"77",X"A7",X"02",X"96",X"B6",X"85",
		X"01",X"26",X"1C",X"81",X"98",X"25",X"02",X"80",X"84",X"6F",X"98",X"00",X"A7",X"84",X"96",X"91",
		X"85",X"02",X"27",X"0B",X"96",X"B8",X"84",X"3F",X"C6",X"03",X"3D",X"CB",X"2C",X"E7",X"01",X"86",
		X"87",X"90",X"20",X"81",X"26",X"23",X"25",X"96",X"EE",X"27",X"20",X"4F",X"5F",X"97",X"EE",X"8E",
		X"BE",X"97",X"ED",X"98",X"06",X"ED",X"98",X"12",X"ED",X"98",X"1E",X"ED",X"98",X"2A",X"A7",X"0B",
		X"A7",X"88",X"17",X"A7",X"88",X"23",X"A7",X"88",X"2F",X"97",X"EF",X"39",X"D6",X"3A",X"C1",X"02",
		X"24",X"D5",X"96",X"91",X"85",X"02",X"26",X"CF",X"CC",X"87",X"AA",X"97",X"EE",X"93",X"20",X"58",
		X"49",X"58",X"49",X"DD",X"4B",X"CC",X"00",X"00",X"8E",X"BE",X"97",X"ED",X"98",X"06",X"ED",X"98",
		X"12",X"ED",X"98",X"1E",X"ED",X"98",X"2A",X"A6",X"0B",X"27",X"2D",X"6A",X"0B",X"27",X"29",X"EC",
		X"84",X"E3",X"04",X"ED",X"04",X"D3",X"4B",X"81",X"9A",X"25",X"04",X"7E",X"2B",X"E4",X"12",X"A7",
		X"06",X"EC",X"02",X"C3",X"00",X"10",X"ED",X"02",X"E3",X"07",X"ED",X"07",X"8B",X"10",X"81",X"3C",
		X"23",X"E9",X"CC",X"44",X"44",X"ED",X"98",X"06",X"30",X"0C",X"8C",X"BE",X"BB",X"26",X"C8",X"0A",
		X"EF",X"2A",X"38",X"DC",X"B6",X"C4",X"3F",X"D7",X"EF",X"84",X"03",X"4C",X"97",X"4B",X"8E",X"BE",
		X"97",X"A6",X"0B",X"26",X"1B",X"6F",X"04",X"D6",X"B6",X"1D",X"ED",X"84",X"86",X"03",X"BD",X"08",
		X"C1",X"40",X"D6",X"B8",X"ED",X"02",X"C4",X"3F",X"CB",X"38",X"E7",X"0B",X"86",X"9C",X"A7",X"07",
		X"30",X"0C",X"8C",X"BE",X"BB",X"27",X"04",X"0A",X"4B",X"26",X"D6",X"39",X"8E",X"BB",X"83",X"9F",
		X"7B",X"BD",X"07",X"EC",X"A7",X"88",X"20",X"A7",X"80",X"8C",X"BB",X"A3",X"26",X"F3",X"39",X"9E",
		X"7B",X"DE",X"96",X"33",X"C9",X"FF",X"01",X"EC",X"84",X"ED",X"C4",X"A6",X"05",X"E6",X"09",X"ED",
		X"42",X"A6",X"0C",X"A7",X"44",X"96",X"57",X"85",X"02",X"27",X"22",X"A6",X"03",X"E6",X"06",X"ED",
		X"C9",X"FF",X"01",X"A6",X"0A",X"A7",X"C9",X"FF",X"03",X"A6",X"04",X"E6",X"07",X"ED",X"C9",X"FE",
		X"01",X"A6",X"0B",X"A7",X"C9",X"FE",X"03",X"A6",X"08",X"A7",X"C9",X"FD",X"02",X"39",X"DE",X"7B",
		X"9E",X"96",X"30",X"89",X"08",X"01",X"37",X"26",X"ED",X"84",X"10",X"AF",X"02",X"37",X"26",X"A7",
		X"04",X"96",X"57",X"85",X"02",X"27",X"18",X"E7",X"89",X"01",X"01",X"10",X"AF",X"89",X"01",X"02",
		X"37",X"26",X"10",X"AF",X"89",X"02",X"01",X"A7",X"89",X"02",X"03",X"E7",X"89",X"03",X"02",X"39",
		X"DE",X"96",X"5F",X"8E",X"00",X"00",X"31",X"84",X"33",X"C9",X"08",X"06",X"36",X"34",X"AF",X"C9",
		X"01",X"01",X"E7",X"C9",X"01",X"03",X"AF",X"C9",X"02",X"01",X"E7",X"C9",X"02",X"03",X"E7",X"C9",
		X"03",X"02",X"39",X"DE",X"96",X"5F",X"8E",X"00",X"00",X"31",X"84",X"33",X"C9",X"FF",X"06",X"36",
		X"34",X"AF",X"C9",X"FF",X"01",X"E7",X"C9",X"FF",X"03",X"AF",X"C9",X"FE",X"01",X"E7",X"C9",X"FE",
		X"03",X"E7",X"C9",X"FD",X"02",X"39",X"97",X"53",X"96",X"91",X"85",X"10",X"27",X"09",X"DC",X"92",
		X"DD",X"94",X"DC",X"98",X"DD",X"96",X"39",X"96",X"53",X"91",X"97",X"23",X"F9",X"D1",X"97",X"22",
		X"F5",X"96",X"94",X"2B",X"06",X"8D",X"2C",X"8D",X"BA",X"20",X"04",X"8D",X"26",X"8D",X"91",X"DC",
		X"92",X"DD",X"94",X"2B",X"05",X"8D",X"08",X"7E",X"0A",X"AF",X"8D",X"11",X"7E",X"0A",X"EE",X"10",
		X"8E",X"20",X"A9",X"96",X"9B",X"48",X"DC",X"98",X"DD",X"96",X"7E",X"03",X"69",X"10",X"8E",X"20",
		X"B3",X"20",X"F0",X"DC",X"96",X"7E",X"03",X"BA",X"96",X"91",X"85",X"40",X"10",X"26",X"01",X"0A",
		X"0F",X"4B",X"DC",X"9E",X"43",X"53",X"C3",X"00",X"01",X"2A",X"02",X"03",X"4B",X"58",X"49",X"58",
		X"49",X"D3",X"9F",X"DD",X"9F",X"96",X"4B",X"99",X"9E",X"97",X"9E",X"DC",X"9E",X"96",X"57",X"85",
		X"02",X"27",X"12",X"0F",X"4B",X"DC",X"94",X"2A",X"02",X"03",X"4B",X"D3",X"9F",X"DD",X"9F",X"96",
		X"4B",X"99",X"9E",X"97",X"9E",X"DC",X"9E",X"47",X"56",X"47",X"56",X"4F",X"57",X"46",X"97",X"70",
		X"D7",X"6F",X"96",X"94",X"2B",X"07",X"86",X"20",X"5D",X"2B",X"07",X"20",X"09",X"86",X"70",X"5D",
		X"2B",X"04",X"0F",X"70",X"0F",X"6F",X"D6",X"70",X"9B",X"6F",X"97",X"6F",X"93",X"9A",X"27",X"26",
		X"25",X"12",X"10",X"83",X"01",X"00",X"23",X"1E",X"CC",X"00",X"40",X"DD",X"71",X"CC",X"01",X"00",
		X"D3",X"9A",X"20",X"18",X"10",X"83",X"FF",X"00",X"2E",X"0C",X"CC",X"FF",X"C0",X"DD",X"71",X"CC",
		X"FF",X"00",X"D3",X"9A",X"20",X"06",X"4F",X"5F",X"DD",X"71",X"DC",X"6F",X"DD",X"9A",X"97",X"98",
		X"DC",X"20",X"DD",X"22",X"DC",X"9E",X"10",X"83",X"01",X"00",X"2D",X"03",X"CC",X"01",X"00",X"10",
		X"83",X"FF",X"00",X"2E",X"03",X"CC",X"FF",X"00",X"DD",X"9E",X"D3",X"20",X"93",X"71",X"DD",X"20",
		X"DC",X"9A",X"44",X"56",X"44",X"56",X"C4",X"E0",X"D3",X"20",X"DD",X"A3",X"D6",X"9C",X"96",X"59",
		X"44",X"25",X"09",X"96",X"57",X"2B",X"20",X"CC",X"00",X"00",X"20",X"36",X"C1",X"2D",X"23",X"3A",
		X"DC",X"A1",X"2A",X"0E",X"C3",X"FF",X"F8",X"10",X"83",X"FE",X"00",X"2C",X"25",X"CC",X"FE",X"00",
		X"20",X"20",X"CC",X"FF",X"00",X"20",X"1B",X"C1",X"EE",X"24",X"1F",X"DC",X"A1",X"2F",X"0E",X"C3",
		X"00",X"08",X"10",X"83",X"02",X"00",X"23",X"0A",X"CC",X"02",X"00",X"20",X"05",X"CC",X"01",X"00",
		X"20",X"00",X"DD",X"A1",X"D3",X"9C",X"DD",X"9C",X"97",X"99",X"39",X"96",X"91",X"85",X"20",X"26",
		X"22",X"8E",X"9C",X"41",X"20",X"19",X"EC",X"0A",X"E3",X"0E",X"ED",X"0A",X"EC",X"0C",X"E3",X"88",
		X"10",X"81",X"2C",X"24",X"02",X"86",X"F0",X"81",X"F0",X"23",X"02",X"86",X"2C",X"ED",X"0C",X"AE",
		X"84",X"26",X"E3",X"39",X"DD",X"4D",X"96",X"91",X"85",X"20",X"26",X"4B",X"8E",X"9C",X"41",X"20",
		X"42",X"EC",X"04",X"27",X"13",X"D1",X"4D",X"22",X"3A",X"D1",X"4E",X"23",X"36",X"10",X"AE",X"02",
		X"AD",X"B8",X"08",X"CC",X"00",X"00",X"ED",X"04",X"E6",X"0C",X"D1",X"4D",X"22",X"25",X"D1",X"4E",
		X"23",X"21",X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",X"80",X"24",X"17",X"10",X"AE",X"02",X"58",
		X"49",X"58",X"49",X"AB",X"A4",X"81",X"9C",X"22",X"0A",X"A0",X"A4",X"58",X"E6",X"0C",X"ED",X"04",
		X"AD",X"B8",X"06",X"AE",X"84",X"26",X"BA",X"39",X"34",X"66",X"96",X"75",X"81",X"14",X"24",X"4F",
		X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",X"80",X"24",X"45",X"58",X"49",X"58",X"49",X"E6",X"0C",
		X"C1",X"2C",X"23",X"3B",X"9E",X"43",X"27",X"37",X"ED",X"04",X"ED",X"0A",X"1E",X"89",X"ED",X"0C",
		X"EF",X"06",X"4F",X"5F",X"ED",X"0E",X"ED",X"88",X"10",X"EE",X"66",X"37",X"26",X"ED",X"88",X"12",
		X"10",X"AF",X"02",X"37",X"06",X"EF",X"66",X"ED",X"08",X"86",X"14",X"A7",X"88",X"15",X"A7",X"88",
		X"16",X"EC",X"84",X"DD",X"43",X"DC",X"49",X"ED",X"84",X"0C",X"75",X"9F",X"49",X"35",X"E6",X"EE",
		X"66",X"33",X"46",X"EF",X"66",X"4F",X"35",X"E6",X"8E",X"9C",X"49",X"20",X"1B",X"A6",X"88",X"16",
		X"27",X"05",X"6A",X"88",X"15",X"26",X"11",X"EE",X"84",X"EF",X"A4",X"DE",X"43",X"EF",X"84",X"9F",
		X"43",X"BD",X"00",X"00",X"0A",X"75",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"DF",X"39",X"BD",
		X"26",X"99",X"12",X"12",X"12",X"0C",X"8F",X"CC",X"06",X"CE",X"BD",X"06",X"FD",X"9E",X"98",X"96",
		X"92",X"2A",X"06",X"7E",X"0E",X"6B",X"7E",X"00",X"E4",X"30",X"89",X"07",X"04",X"AF",X"47",X"AF",
		X"49",X"AF",X"4B",X"96",X"91",X"85",X"40",X"26",X"63",X"AE",X"47",X"CC",X"99",X"11",X"8C",X"98",
		X"00",X"24",X"59",X"E7",X"84",X"E7",X"89",X"01",X"00",X"E7",X"89",X"02",X"00",X"E7",X"89",X"03",
		X"00",X"30",X"89",X"04",X"00",X"A7",X"84",X"AF",X"47",X"10",X"9E",X"80",X"10",X"8C",X"BB",X"80",
		X"25",X"04",X"10",X"8E",X"BB",X"63",X"AE",X"49",X"EC",X"A1",X"A7",X"84",X"E7",X"89",X"01",X"00",
		X"E6",X"A0",X"E7",X"89",X"02",X"00",X"30",X"89",X"03",X"00",X"10",X"9F",X"80",X"AF",X"49",X"6F",
		X"D8",X"0B",X"6C",X"4B",X"EC",X"47",X"80",X"06",X"34",X"40",X"CE",X"20",X"93",X"BD",X"0F",X"07",
		X"35",X"40",X"26",X"08",X"86",X"01",X"8E",X"0D",X"F3",X"7E",X"00",X"A8",X"AE",X"4B",X"4F",X"A7",
		X"84",X"30",X"89",X"01",X"00",X"AC",X"47",X"23",X"F6",X"20",X"7C",X"30",X"04",X"AF",X"47",X"AF",
		X"49",X"AF",X"4B",X"96",X"91",X"85",X"40",X"26",X"61",X"AE",X"47",X"CC",X"99",X"11",X"8C",X"05",
		X"00",X"23",X"57",X"E7",X"84",X"E7",X"89",X"FF",X"00",X"E7",X"89",X"FE",X"00",X"E7",X"89",X"FD",
		X"00",X"30",X"89",X"FC",X"00",X"A7",X"84",X"AF",X"47",X"10",X"9E",X"80",X"10",X"8C",X"BB",X"80",
		X"25",X"04",X"10",X"8E",X"BB",X"63",X"AE",X"49",X"EC",X"A0",X"A7",X"84",X"E7",X"89",X"FF",X"00",
		X"E6",X"A0",X"E7",X"89",X"FE",X"00",X"30",X"89",X"FD",X"00",X"10",X"9F",X"80",X"AF",X"49",X"6F",
		X"D8",X"0B",X"6A",X"4B",X"EC",X"47",X"34",X"40",X"CE",X"20",X"93",X"BD",X"0F",X"07",X"35",X"40",
		X"26",X"08",X"86",X"01",X"8E",X"0E",X"73",X"7E",X"00",X"A8",X"AE",X"4B",X"4F",X"A7",X"84",X"30",
		X"89",X"FF",X"00",X"AC",X"47",X"24",X"F6",X"0A",X"8F",X"7E",X"00",X"E4",X"8E",X"BB",X"63",X"9F",
		X"80",X"BD",X"07",X"EC",X"5F",X"44",X"24",X"02",X"CB",X"01",X"44",X"24",X"02",X"CB",X"10",X"E7",
		X"80",X"8C",X"BB",X"83",X"26",X"EB",X"39",X"8E",X"9C",X"41",X"DD",X"AD",X"E3",X"C4",X"DD",X"AF",
		X"20",X"17",X"EC",X"04",X"27",X"13",X"91",X"AF",X"24",X"0F",X"D1",X"B0",X"24",X"0B",X"E3",X"98",
		X"02",X"91",X"AD",X"23",X"04",X"D1",X"AE",X"22",X"05",X"AE",X"84",X"26",X"E5",X"39",X"DF",X"B3",
		X"10",X"AE",X"02",X"A3",X"A4",X"DD",X"4F",X"4F",X"5F",X"DD",X"A7",X"DD",X"A9",X"DC",X"4F",X"D0",
		X"AE",X"22",X"05",X"50",X"D7",X"A8",X"20",X"02",X"D7",X"AA",X"90",X"AD",X"22",X"05",X"40",X"97",
		X"A7",X"20",X"02",X"97",X"A9",X"DC",X"4F",X"E3",X"A4",X"D0",X"B0",X"22",X"01",X"5F",X"90",X"AF",
		X"22",X"01",X"4F",X"DD",X"B1",X"EC",X"A4",X"93",X"A7",X"93",X"B1",X"DD",X"A5",X"A6",X"41",X"97",
		X"AC",X"D6",X"A9",X"3D",X"EE",X"42",X"33",X"CB",X"A6",X"21",X"97",X"AB",X"10",X"AE",X"22",X"D6",
		X"A7",X"3D",X"31",X"AB",X"96",X"A8",X"31",X"A6",X"96",X"AA",X"33",X"C6",X"D6",X"A6",X"5A",X"A6",
		X"C5",X"27",X"2A",X"A6",X"A5",X"27",X"26",X"31",X"A5",X"1F",X"20",X"EE",X"02",X"A3",X"42",X"10",
		X"AE",X"04",X"E0",X"41",X"82",X"00",X"25",X"06",X"31",X"A9",X"01",X"00",X"20",X"F4",X"EB",X"41",
		X"89",X"00",X"31",X"A5",X"10",X"9F",X"D0",X"AD",X"98",X"08",X"86",X"01",X"39",X"5A",X"2A",X"CF",
		X"DC",X"AB",X"31",X"A6",X"33",X"C5",X"0A",X"A5",X"26",X"C2",X"DE",X"B3",X"7E",X"0F",X"29",X"0F",
		X"90",X"8E",X"0F",X"E6",X"96",X"90",X"E6",X"86",X"27",X"F5",X"0C",X"90",X"D7",X"27",X"86",X"02",
		X"8E",X"0F",X"D1",X"7E",X"00",X"A8",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",X"3F",X"37",X"2F",
		X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",X"CA",X"DA",X"E8",
		X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"3C",X"00",X"9E",X"7B",X"30",X"01",X"8C",
		X"BB",X"A3",X"23",X"03",X"8E",X"BB",X"83",X"9F",X"7B",X"86",X"04",X"8E",X"10",X"0B",X"7E",X"00",
		X"A8",X"BD",X"10",X"6E",X"86",X"02",X"8E",X"10",X"2C",X"7E",X"00",X"A8",X"BD",X"10",X"45",X"BD",
		X"0D",X"A8",X"86",X"02",X"8E",X"10",X"3A",X"7E",X"00",X"A8",X"BD",X"10",X"CA",X"86",X"04",X"8E",
		X"10",X"21",X"7E",X"00",X"A8",X"DC",X"20",X"83",X"0C",X"80",X"DD",X"4F",X"8E",X"9C",X"41",X"20",
		X"16",X"EC",X"0A",X"93",X"4F",X"10",X"83",X"3E",X"80",X"25",X"0C",X"EE",X"84",X"EF",X"A4",X"DE",
		X"47",X"EF",X"84",X"9F",X"47",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"E4",X"39",X"DC",X"20",
		X"83",X"0C",X"80",X"DD",X"4F",X"8E",X"9C",X"47",X"20",X"49",X"96",X"91",X"85",X"20",X"26",X"29",
		X"EC",X"88",X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"E3",X"0C",X"81",X"2C",X"24",X"06",X"81",
		X"0E",X"23",X"06",X"86",X"F0",X"81",X"F0",X"23",X"02",X"86",X"2C",X"ED",X"0C",X"EC",X"0E",X"58",
		X"49",X"58",X"49",X"58",X"49",X"E3",X"0A",X"ED",X"0A",X"EC",X"0A",X"93",X"4F",X"10",X"83",X"3E",
		X"80",X"24",X"10",X"EE",X"84",X"EF",X"A4",X"DE",X"41",X"EF",X"84",X"9F",X"41",X"4F",X"5F",X"ED",
		X"04",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"B1",X"39",X"CE",X"00",X"00",X"C6",X"08",X"8E",
		X"BC",X"83",X"EF",X"94",X"EF",X"98",X"02",X"EF",X"98",X"04",X"EF",X"98",X"06",X"3A",X"9C",X"73",
		X"25",X"F0",X"AE",X"9F",X"9C",X"73",X"27",X"08",X"EF",X"84",X"6F",X"02",X"EF",X"89",X"FF",X"00",
		X"DC",X"20",X"83",X"6D",X"40",X"DD",X"4F",X"44",X"44",X"CE",X"11",X"B6",X"C6",X"03",X"3D",X"33",
		X"CB",X"96",X"91",X"85",X"02",X"26",X"22",X"86",X"2C",X"10",X"8E",X"BD",X"4B",X"8E",X"00",X"00",
		X"AF",X"B4",X"37",X"14",X"ED",X"A4",X"AF",X"B1",X"4C",X"8E",X"00",X"00",X"AF",X"B4",X"37",X"14",
		X"ED",X"A4",X"AF",X"B1",X"4C",X"81",X"6C",X"26",X"E4",X"8E",X"48",X"08",X"CC",X"90",X"90",X"ED",
		X"84",X"ED",X"88",X"1A",X"8E",X"4F",X"08",X"CC",X"09",X"09",X"ED",X"84",X"ED",X"88",X"1A",X"7E",
		X"25",X"B0",X"CE",X"BC",X"83",X"8D",X"6A",X"8E",X"9C",X"47",X"8D",X"65",X"DF",X"73",X"DC",X"96",
		X"44",X"44",X"44",X"44",X"54",X"54",X"54",X"C3",X"47",X"03",X"ED",X"C4",X"AE",X"C4",X"CC",X"90",
		X"99",X"ED",X"84",X"A7",X"02",X"86",X"09",X"A7",X"89",X"FF",X"01",X"39",X"EC",X"0A",X"93",X"4F",
		X"44",X"44",X"E6",X"0C",X"54",X"54",X"54",X"C3",X"2C",X"03",X"ED",X"C4",X"EC",X"88",X"12",X"81",
		X"1F",X"26",X"2C",X"EC",X"C4",X"81",X"6B",X"26",X"03",X"4A",X"A7",X"C4",X"10",X"8E",X"FF",X"F0",
		X"10",X"AF",X"D1",X"5C",X"ED",X"C4",X"10",X"8E",X"F0",X"FF",X"10",X"AF",X"D1",X"4C",X"ED",X"C4",
		X"10",X"8E",X"F0",X"F0",X"10",X"AF",X"D1",X"5A",X"ED",X"C4",X"10",X"AF",X"D1",X"20",X"02",X"ED",
		X"D1",X"AE",X"84",X"26",X"B7",X"39",X"1B",X"08",X"80",X"1A",X"80",X"08",X"1C",X"80",X"08",X"1E",
		X"80",X"08",X"1F",X"88",X"00",X"1F",X"88",X"00",X"1E",X"88",X"00",X"1C",X"88",X"00",X"1A",X"88",
		X"00",X"1C",X"88",X"00",X"1E",X"88",X"00",X"1F",X"80",X"08",X"20",X"88",X"00",X"20",X"88",X"00",
		X"1F",X"88",X"00",X"1E",X"88",X"00",X"1C",X"08",X"80",X"1C",X"88",X"00",X"1D",X"80",X"08",X"1F",
		X"88",X"00",X"1F",X"88",X"00",X"1F",X"02",X"20",X"1F",X"22",X"00",X"1F",X"02",X"20",X"1E",X"22",
		X"00",X"1F",X"22",X"00",X"1E",X"02",X"20",X"1C",X"02",X"20",X"1A",X"02",X"20",X"1C",X"20",X"02",
		X"1D",X"02",X"20",X"1C",X"02",X"20",X"19",X"02",X"20",X"16",X"02",X"20",X"18",X"20",X"02",X"1B",
		X"20",X"02",X"1D",X"20",X"02",X"1F",X"20",X"02",X"1F",X"22",X"00",X"1F",X"22",X"00",X"1F",X"20",
		X"02",X"20",X"22",X"00",X"1F",X"0B",X"B0",X"1D",X"0B",X"B0",X"1C",X"BB",X"00",X"1E",X"BB",X"00",
		X"1E",X"0B",X"B0",X"1B",X"0B",X"B0",X"1D",X"B0",X"0B",X"1F",X"0B",X"B0",X"20",X"BB",X"00",X"1F",
		X"0B",X"B0",X"1F",X"B0",X"0B",X"1F",X"BB",X"00",X"1F",X"B0",X"0B",X"20",X"BB",X"00",X"1F",X"0B",
		X"B0",X"1F",X"B0",X"0B",X"1F",X"BB",X"00",X"1F",X"0B",X"B0",X"1F",X"BB",X"00",X"1F",X"BB",X"00",
		X"1E",X"0B",X"B0",X"1D",X"0B",X"B0",X"1B",X"08",X"80",X"1A",X"80",X"08",X"1C",X"80",X"08",X"1E",
		X"80",X"08",X"1F",X"88",X"00",X"1F",X"88",X"00",X"1E",X"88",X"00",X"1C",X"88",X"00",X"1A",X"88",
		X"00",X"1C",X"88",X"00",X"1E",X"88",X"00",X"1F",X"80",X"08",X"20",X"88",X"00",X"20",X"88",X"00",
		X"1F",X"88",X"00",X"1E",X"88",X"00",X"1C",X"08",X"80",X"1C",X"88",X"00",X"1D",X"80",X"08",X"1F",
		X"88",X"00",X"1F",X"88",X"00",X"1F",X"02",X"20",X"1F",X"22",X"00",X"1F",X"02",X"20",X"1E",X"22",
		X"00",X"1F",X"22",X"00",X"1E",X"02",X"20",X"1C",X"02",X"20",X"1A",X"02",X"20",X"1C",X"20",X"02",
		X"1D",X"02",X"20",X"1C",X"02",X"20",X"19",X"02",X"20",X"16",X"02",X"20",X"18",X"20",X"02",X"1B",
		X"20",X"02",X"1D",X"20",X"02",X"1F",X"20",X"02",X"1F",X"22",X"00",X"1F",X"22",X"00",X"1F",X"20",
		X"02",X"20",X"22",X"00",X"1F",X"0B",X"B0",X"1D",X"0B",X"B0",X"1C",X"BB",X"00",X"1E",X"BB",X"00",
		X"1E",X"0B",X"B0",X"1B",X"0B",X"B0",X"1D",X"B0",X"0B",X"1F",X"0B",X"B0",X"20",X"BB",X"00",X"1F",
		X"0B",X"B0",X"1F",X"B0",X"0B",X"1F",X"BB",X"00",X"1F",X"B0",X"0B",X"20",X"BB",X"00",X"1F",X"0B",
		X"B0",X"1F",X"B0",X"0B",X"1F",X"BB",X"00",X"1F",X"0B",X"B0",X"1F",X"BB",X"00",X"1F",X"BB",X"00",
		X"1E",X"0B",X"B0",X"1D",X"0B",X"B0",X"34",X"76",X"1F",X"01",X"EC",X"A4",X"10",X"AE",X"22",X"34",
		X"06",X"C5",X"01",X"26",X"17",X"C0",X"02",X"EE",X"A5",X"EF",X"85",X"C0",X"02",X"2A",X"F8",X"E6",
		X"61",X"30",X"89",X"01",X"00",X"31",X"A5",X"4A",X"26",X"EB",X"20",X"1D",X"5A",X"A6",X"A5",X"A7",
		X"85",X"C0",X"02",X"2B",X"08",X"EE",X"A5",X"EF",X"85",X"C0",X"02",X"2A",X"F8",X"E6",X"61",X"30",
		X"89",X"01",X"00",X"31",X"A5",X"6A",X"E4",X"26",X"E3",X"32",X"62",X"35",X"F6",X"34",X"56",X"1F",
		X"01",X"EC",X"A4",X"CE",X"00",X"00",X"34",X"04",X"C5",X"01",X"26",X"13",X"C0",X"02",X"EF",X"85",
		X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",X"89",X"01",X"00",X"4A",X"26",X"EF",X"20",X"16",X"5A",
		X"6F",X"85",X"C0",X"02",X"2B",X"06",X"EF",X"85",X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",X"89",
		X"01",X"00",X"4A",X"26",X"EA",X"32",X"61",X"35",X"D6",X"34",X"56",X"20",X"C6",X"34",X"76",X"CE",
		X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"36",X"36",X"36",X"36",X"36",X"36",X"36",
		X"36",X"36",X"36",X"36",X"10",X"11",X"83",X"00",X"00",X"26",X"EE",X"35",X"F6",X"34",X"7E",X"CE",
		X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"1F",X"8B",X"C6",X"08",X"36",X"3A",X"36",
		X"3A",X"36",X"3A",X"36",X"3A",X"5A",X"26",X"F5",X"36",X"3A",X"36",X"3A",X"36",X"3A",X"36",X"10",
		X"33",X"C8",X"D4",X"11",X"83",X"00",X"00",X"26",X"E2",X"35",X"FE",X"A6",X"01",X"84",X"0F",X"34",
		X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",X"8D",X"EF",X"34",X"02",X"8D",X"EB",
		X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",X"A7",X"81",X"35",X"82",
		X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",X"7E",X"26",X"7C",X"12",X"09",X"66",
		X"44",X"34",X"02",X"86",X"00",X"24",X"08",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"BD",
		X"07",X"D9",X"DD",X"4F",X"C6",X"03",X"E0",X"E0",X"A6",X"85",X"9B",X"50",X"19",X"A7",X"85",X"5A",
		X"2B",X"0E",X"A6",X"85",X"99",X"4F",X"19",X"A7",X"85",X"86",X"00",X"97",X"4F",X"5A",X"2A",X"F2",
		X"DC",X"85",X"27",X"2F",X"31",X"04",X"8D",X"30",X"25",X"29",X"A6",X"22",X"9B",X"86",X"19",X"A7",
		X"22",X"A6",X"21",X"99",X"85",X"19",X"A7",X"21",X"A6",X"A4",X"89",X"00",X"19",X"A7",X"A4",X"BD",
		X"5F",X"C7",X"BD",X"5F",X"BB",X"BD",X"5F",X"BE",X"CC",X"06",X"63",X"BD",X"06",X"FD",X"C6",X"05",
		X"BD",X"F4",X"83",X"8D",X"13",X"35",X"76",X"39",X"34",X"06",X"EC",X"84",X"10",X"A3",X"A4",X"26",
		X"05",X"EC",X"02",X"10",X"A3",X"22",X"35",X"86",X"96",X"DB",X"27",X"01",X"39",X"96",X"67",X"8E",
		X"70",X"00",X"D6",X"91",X"2B",X"07",X"91",X"67",X"26",X"03",X"8E",X"70",X"5B",X"34",X"12",X"4A",
		X"26",X"08",X"8E",X"07",X"23",X"CE",X"BD",X"D6",X"20",X"06",X"8E",X"6D",X"23",X"CE",X"BE",X"15",
		X"0F",X"4F",X"C6",X"07",X"A6",X"C0",X"10",X"AE",X"61",X"C5",X"01",X"26",X"06",X"33",X"5F",X"44",
		X"44",X"44",X"44",X"84",X"0F",X"26",X"08",X"C1",X"02",X"23",X"04",X"0D",X"4F",X"27",X"0D",X"0C",
		X"4F",X"48",X"48",X"31",X"A6",X"1E",X"10",X"BD",X"13",X"36",X"1E",X"10",X"30",X"89",X"04",X"00",
		X"5A",X"26",X"D1",X"35",X"A2",X"34",X"16",X"8E",X"15",X"BA",X"CC",X"01",X"3C",X"20",X"0D",X"34",
		X"16",X"B6",X"C8",X"06",X"2A",X"F1",X"8E",X"16",X"4C",X"CC",X"03",X"34",X"9F",X"6C",X"F7",X"C8",
		X"07",X"B7",X"C9",X"00",X"86",X"7E",X"97",X"6B",X"35",X"96",X"34",X"10",X"9E",X"3B",X"27",X"09",
		X"10",X"AC",X"02",X"27",X"06",X"AE",X"84",X"26",X"F7",X"1C",X"FB",X"35",X"90",X"BD",X"13",X"DD",
		X"9E",X"69",X"A6",X"09",X"BD",X"08",X"E4",X"1F",X"89",X"81",X"05",X"23",X"02",X"86",X"05",X"34",
		X"02",X"86",X"03",X"BD",X"70",X"58",X"35",X"82",X"0F",X"26",X"DE",X"3F",X"35",X"10",X"AF",X"4D",
		X"5F",X"1F",X"02",X"1F",X"89",X"86",X"02",X"ED",X"4B",X"86",X"02",X"BD",X"70",X"58",X"8E",X"38",
		X"A0",X"B6",X"BE",X"54",X"A7",X"49",X"27",X"22",X"1F",X"10",X"10",X"8E",X"20",X"39",X"BD",X"13",
		X"36",X"30",X"89",X"04",X"00",X"EC",X"4B",X"BD",X"14",X"3A",X"AF",X"47",X"86",X"04",X"8E",X"15",
		X"A4",X"7E",X"00",X"A8",X"AE",X"47",X"6A",X"49",X"26",X"DE",X"9E",X"69",X"BD",X"5F",X"C1",X"86",
		X"80",X"8E",X"15",X"B7",X"7E",X"00",X"A8",X"6E",X"D8",X"0D",X"86",X"9C",X"1F",X"8B",X"86",X"34",
		X"B7",X"C8",X"0F",X"B6",X"C8",X"0E",X"B6",X"CB",X"00",X"81",X"80",X"25",X"2B",X"96",X"6E",X"26",
		X"6C",X"0C",X"6E",X"BD",X"07",X"18",X"BD",X"0B",X"B8",X"BD",X"09",X"27",X"B6",X"CB",X"00",X"80",
		X"08",X"81",X"A8",X"23",X"02",X"86",X"A8",X"97",X"7E",X"DC",X"7E",X"BD",X"0C",X"F4",X"DC",X"7E",
		X"BD",X"0B",X"66",X"BD",X"16",X"C8",X"20",X"45",X"D6",X"6E",X"27",X"41",X"0F",X"6E",X"0C",X"39",
		X"C6",X"39",X"F7",X"CB",X"FF",X"81",X"04",X"22",X"1B",X"CE",X"C0",X"10",X"DC",X"30",X"9E",X"32",
		X"10",X"9E",X"34",X"36",X"36",X"DC",X"2A",X"9E",X"2C",X"10",X"9E",X"2E",X"36",X"36",X"DC",X"26",
		X"9E",X"28",X"36",X"16",X"BD",X"07",X"AD",X"96",X"91",X"85",X"02",X"26",X"03",X"BD",X"2C",X"03",
		X"DC",X"7D",X"BD",X"0B",X"66",X"DC",X"7D",X"BD",X"0C",X"F4",X"BD",X"0C",X"CB",X"1A",X"FF",X"86",
		X"35",X"B7",X"C8",X"0F",X"A6",X"E4",X"84",X"6F",X"A7",X"E4",X"35",X"FF",X"86",X"9C",X"1F",X"8B",
		X"86",X"34",X"B7",X"C8",X"0F",X"B6",X"C8",X"0E",X"B6",X"CB",X"00",X"81",X"60",X"25",X"21",X"D6",
		X"6E",X"26",X"DA",X"0C",X"6E",X"43",X"97",X"7E",X"BD",X"07",X"AD",X"96",X"91",X"85",X"02",X"26",
		X"03",X"BD",X"2C",X"03",X"DC",X"7D",X"BD",X"0B",X"66",X"DC",X"7D",X"BD",X"0C",X"F4",X"20",X"BD",
		X"D6",X"6E",X"27",X"B9",X"0F",X"6E",X"0C",X"39",X"C6",X"39",X"F7",X"CB",X"FF",X"81",X"04",X"22",
		X"1B",X"CE",X"C0",X"10",X"DC",X"30",X"9E",X"32",X"10",X"9E",X"34",X"36",X"36",X"DC",X"2A",X"9E",
		X"2C",X"10",X"9E",X"2E",X"36",X"36",X"DC",X"26",X"9E",X"28",X"36",X"16",X"BD",X"07",X"18",X"BD",
		X"0B",X"B8",X"BD",X"09",X"27",X"DC",X"7E",X"BD",X"0B",X"66",X"DC",X"7E",X"BD",X"0C",X"F4",X"BD",
		X"16",X"C8",X"BD",X"0C",X"CB",X"7E",X"16",X"3D",X"96",X"91",X"85",X"20",X"26",X"3D",X"DC",X"20",
		X"C4",X"E0",X"DD",X"79",X"DC",X"22",X"C4",X"E0",X"93",X"79",X"58",X"49",X"58",X"49",X"DD",X"79",
		X"8E",X"9C",X"49",X"20",X"22",X"10",X"AE",X"04",X"EC",X"88",X"10",X"E3",X"0C",X"81",X"2C",X"23",
		X"47",X"ED",X"0C",X"EC",X"0E",X"D3",X"79",X"E3",X"0A",X"81",X"97",X"24",X"3B",X"ED",X"0A",X"58",
		X"E6",X"0C",X"ED",X"04",X"6E",X"98",X"12",X"AE",X"84",X"26",X"DA",X"39",X"DE",X"82",X"24",X"02",
		X"33",X"46",X"CC",X"00",X"00",X"ED",X"A4",X"A7",X"22",X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",
		X"02",X"10",X"AE",X"04",X"EC",X"C4",X"ED",X"A4",X"EC",X"42",X"A7",X"22",X"E7",X"A9",X"01",X"00",
		X"EC",X"44",X"ED",X"A9",X"01",X"01",X"20",X"CF",X"4F",X"5F",X"A7",X"88",X"16",X"ED",X"A4",X"A7",
		X"22",X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"20",X"BC",X"CC",X"00",X"00",X"ED",X"A4",
		X"A7",X"22",X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"EE",X"04",X"CC",X"99",X"99",X"25",
		X"0E",X"84",X"0F",X"ED",X"C4",X"A7",X"42",X"C4",X"F0",X"E7",X"C9",X"01",X"01",X"20",X"98",X"84",
		X"F0",X"ED",X"C9",X"01",X"00",X"A7",X"C9",X"01",X"02",X"C4",X"0F",X"E7",X"41",X"20",X"88",X"EE",
		X"04",X"CC",X"00",X"99",X"A7",X"A4",X"A7",X"A9",X"01",X"00",X"A7",X"A9",X"02",X"00",X"25",X"09",
		X"E7",X"C4",X"E7",X"C9",X"01",X"00",X"7E",X"17",X"07",X"86",X"09",X"A7",X"C4",X"E7",X"C9",X"01",
		X"00",X"86",X"90",X"A7",X"C9",X"02",X"00",X"7E",X"17",X"07",X"02",X"01",X"17",X"B4",X"17",X"B4",
		X"02",X"88",X"02",X"B2",X"FF",X"FF",X"CC",X"00",X"25",X"BD",X"14",X"3A",X"0A",X"75",X"BD",X"01",
		X"CD",X"BD",X"00",X"00",X"EC",X"0A",X"44",X"56",X"44",X"56",X"D3",X"20",X"ED",X"0A",X"A6",X"0C",
		X"80",X"02",X"A7",X"0C",X"CC",X"20",X"75",X"ED",X"02",X"BD",X"27",X"03",X"CC",X"06",X"97",X"7E",
		X"06",X"FD",X"96",X"89",X"26",X"23",X"0C",X"89",X"DC",X"94",X"53",X"43",X"C3",X"00",X"01",X"DD",
		X"92",X"86",X"02",X"8E",X"17",X"F9",X"7E",X"00",X"A8",X"96",X"57",X"85",X"40",X"26",X"F2",X"86",
		X"05",X"8E",X"18",X"07",X"7E",X"00",X"A8",X"0F",X"89",X"7E",X"00",X"E4",X"96",X"76",X"26",X"5F",
		X"9E",X"69",X"A6",X"0A",X"27",X"59",X"0C",X"76",X"6A",X"0A",X"BD",X"5F",X"BE",X"CC",X"06",X"85",
		X"BD",X"06",X"FD",X"9E",X"41",X"27",X"1A",X"EC",X"0A",X"93",X"20",X"10",X"83",X"27",X"00",X"24",
		X"0C",X"A6",X"88",X"14",X"81",X"02",X"24",X"05",X"7E",X"26",X"89",X"20",X"E6",X"AE",X"84",X"20",
		X"E4",X"DE",X"3F",X"86",X"04",X"A7",X"47",X"03",X"26",X"86",X"02",X"8E",X"18",X"51",X"7E",X"00",
		X"A8",X"6A",X"47",X"26",X"F2",X"0F",X"26",X"86",X"0A",X"8E",X"18",X"5F",X"7E",X"00",X"A8",X"96",
		X"57",X"85",X"04",X"26",X"F2",X"86",X"0A",X"8E",X"18",X"6D",X"7E",X"00",X"A8",X"0F",X"76",X"7E",
		X"00",X"E4",X"96",X"91",X"85",X"FD",X"10",X"26",X"00",X"9D",X"84",X"02",X"A7",X"4B",X"86",X"77",
		X"97",X"91",X"BD",X"13",X"DD",X"86",X"0F",X"8E",X"18",X"8D",X"7E",X"00",X"A8",X"9E",X"49",X"27",
		X"05",X"BD",X"01",X"CD",X"20",X"F7",X"0F",X"75",X"DC",X"B6",X"DD",X"20",X"DD",X"22",X"54",X"24",
		X"08",X"CC",X"20",X"00",X"8E",X"03",X"00",X"20",X"06",X"8E",X"FD",X"00",X"CC",X"70",X"00",X"DD",
		X"9A",X"9F",X"92",X"D6",X"B7",X"54",X"CB",X"2C",X"D7",X"9C",X"DD",X"98",X"4F",X"5F",X"97",X"A0",
		X"DD",X"9E",X"DD",X"A1",X"BD",X"2C",X"00",X"C6",X"50",X"8D",X"6E",X"BD",X"01",X"70",X"20",X"A9",
		X"19",X"35",X"00",X"00",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",X"10",X"DC",X"9C",X"ED",X"0C",
		X"DC",X"9A",X"44",X"56",X"44",X"56",X"D3",X"20",X"ED",X"0A",X"96",X"92",X"2A",X"05",X"CE",X"20",
		X"B3",X"EF",X"02",X"DE",X"3F",X"AF",X"47",X"BD",X"27",X"00",X"86",X"28",X"8E",X"19",X"02",X"7E",
		X"00",X"A8",X"BD",X"19",X"43",X"19",X"1A",X"EC",X"47",X"ED",X"07",X"A6",X"4B",X"97",X"91",X"96",
		X"B8",X"81",X"C0",X"10",X"22",X"12",X"C3",X"7E",X"00",X"E4",X"AE",X"47",X"BD",X"1C",X"71",X"BD",
		X"01",X"88",X"86",X"0A",X"8E",X"19",X"2A",X"7E",X"00",X"A8",X"AE",X"47",X"DC",X"43",X"ED",X"84",
		X"9F",X"43",X"7E",X"00",X"E4",X"4F",X"35",X"86",X"5F",X"B6",X"BE",X"54",X"26",X"02",X"CA",X"02",
		X"D7",X"91",X"39",X"34",X"42",X"EE",X"63",X"37",X"10",X"EF",X"63",X"86",X"00",X"BD",X"01",X"30",
		X"35",X"C2",X"08",X"05",X"08",X"05",X"07",X"05",X"06",X"04",X"05",X"03",X"04",X"03",X"03",X"02",
		X"02",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"00",X"01",X"8E",X"9D",X"00",X"9F",X"DF",X"30",X"88",X"40",X"AF",X"88",X"C0",X"8C",X"A0",X"C0",
		X"26",X"F5",X"4F",X"5F",X"ED",X"84",X"DD",X"E1",X"DD",X"E3",X"DD",X"E5",X"97",X"DB",X"39",X"34",
		X"11",X"CB",X"08",X"1F",X"03",X"44",X"44",X"44",X"84",X"FE",X"8E",X"19",X"52",X"EC",X"86",X"DD",
		X"D9",X"35",X"01",X"DC",X"D3",X"25",X"06",X"84",X"F0",X"C4",X"F0",X"20",X"04",X"84",X"0F",X"C4",
		X"0F",X"1F",X"01",X"31",X"84",X"36",X"36",X"36",X"36",X"33",X"C9",X"07",X"0C",X"36",X"36",X"36",
		X"36",X"25",X"04",X"33",X"C9",X"FF",X"00",X"96",X"D3",X"A7",X"C4",X"A7",X"C9",X"FF",X"00",X"A7",
		X"C9",X"FE",X"00",X"A7",X"C9",X"FD",X"00",X"A7",X"C9",X"FC",X"00",X"A7",X"C9",X"FB",X"00",X"A7",
		X"C9",X"FA",X"00",X"A7",X"4B",X"A7",X"C9",X"FF",X"0B",X"A7",X"C9",X"FE",X"0B",X"A7",X"C9",X"FD",
		X"0B",X"A7",X"C9",X"FC",X"0B",X"A7",X"C9",X"FB",X"0B",X"A7",X"C9",X"FA",X"0B",X"96",X"D9",X"24",
		X"07",X"4C",X"44",X"56",X"8B",X"F9",X"20",X"04",X"44",X"56",X"8B",X"FA",X"59",X"C6",X"03",X"33",
		X"CB",X"DC",X"D5",X"25",X"2A",X"A7",X"C4",X"A7",X"45",X"A7",X"C9",X"01",X"00",X"A7",X"C9",X"01",
		X"05",X"A7",X"C9",X"02",X"00",X"A7",X"C9",X"02",X"05",X"84",X"F0",X"C4",X"F0",X"ED",X"41",X"ED",
		X"43",X"ED",X"C9",X"03",X"00",X"ED",X"C9",X"03",X"02",X"ED",X"C9",X"03",X"04",X"20",X"2A",X"A7",
		X"C9",X"01",X"00",X"A7",X"C9",X"01",X"05",X"A7",X"C9",X"02",X"00",X"A7",X"C9",X"02",X"05",X"A7",
		X"C9",X"03",X"00",X"A7",X"C9",X"03",X"05",X"84",X"0F",X"C4",X"0F",X"ED",X"C9",X"03",X"01",X"ED",
		X"C9",X"03",X"03",X"ED",X"C4",X"ED",X"42",X"ED",X"44",X"96",X"DA",X"C6",X"02",X"89",X"00",X"44",
		X"33",X"CB",X"DC",X"D7",X"25",X"08",X"84",X"F0",X"C4",X"F0",X"ED",X"C4",X"35",X"90",X"84",X"0F",
		X"C4",X"0F",X"ED",X"C4",X"35",X"90",X"34",X"10",X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",
		X"00",X"00",X"31",X"84",X"36",X"36",X"36",X"36",X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",
		X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",
		X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",
		X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",X"33",X"C9",X"01",X"0C",X"36",X"36",X"36",X"36",
		X"35",X"90",X"08",X"04",X"1A",X"DC",X"1A",X"DC",X"19",X"8F",X"1A",X"86",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"14",X"EC",X"0A",
		X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"8E",X"A1",X"00",X"A6",
		X"8B",X"35",X"94",X"97",X"4F",X"F6",X"BE",X"64",X"03",X"84",X"2B",X"01",X"50",X"D7",X"50",X"8E",
		X"1B",X"6D",X"86",X"00",X"BD",X"01",X"19",X"33",X"84",X"96",X"4F",X"A7",X"4F",X"4F",X"5F",X"ED",
		X"47",X"ED",X"49",X"ED",X"4B",X"ED",X"4D",X"BD",X"01",X"70",X"20",X"4D",X"1C",X"32",X"88",X"88",
		X"D6",X"50",X"1D",X"ED",X"0E",X"4F",X"5F",X"ED",X"88",X"10",X"96",X"4F",X"44",X"56",X"9B",X"4F",
		X"D3",X"A3",X"8B",X"80",X"ED",X"0A",X"86",X"50",X"A7",X"0C",X"A7",X"C8",X"10",X"EF",X"06",X"9F",
		X"41",X"96",X"4F",X"48",X"8B",X"05",X"AF",X"C6",X"0A",X"4F",X"26",X"CB",X"39",X"96",X"B6",X"84",
		X"06",X"8B",X"07",X"AE",X"C6",X"10",X"27",X"00",X"B1",X"D6",X"B6",X"86",X"0A",X"C4",X"3F",X"CB",
		X"E0",X"2B",X"01",X"40",X"10",X"AE",X"02",X"31",X"A6",X"10",X"8C",X"20",X"4D",X"24",X"04",X"10",
		X"8E",X"20",X"4D",X"10",X"8C",X"20",X"6B",X"23",X"04",X"10",X"8E",X"20",X"6B",X"10",X"AF",X"02",
		X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"1F",X"89",X"50",
		X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"A6",X"05",X"26",X"3B",X"96",X"B6",X"81",X"40",X"22",
		X"16",X"84",X"03",X"8B",X"FE",X"AB",X"C8",X"10",X"81",X"40",X"24",X"02",X"86",X"40",X"81",X"68",
		X"25",X"02",X"86",X"68",X"A7",X"C8",X"10",X"A6",X"C8",X"10",X"A0",X"0C",X"8B",X"10",X"81",X"20",
		X"23",X"48",X"80",X"10",X"2B",X"05",X"CC",X"FF",X"F0",X"20",X"03",X"CC",X"00",X"10",X"E3",X"88",
		X"10",X"ED",X"88",X"10",X"20",X"34",X"90",X"97",X"2B",X"12",X"81",X"20",X"25",X"05",X"CC",X"FF",
		X"F0",X"20",X"19",X"81",X"10",X"22",X"1B",X"CC",X"00",X"10",X"20",X"10",X"81",X"E0",X"2E",X"05",
		X"CC",X"00",X"10",X"20",X"07",X"81",X"F0",X"2D",X"09",X"CC",X"FF",X"F0",X"E3",X"88",X"10",X"ED",
		X"88",X"10",X"96",X"B8",X"84",X"07",X"26",X"02",X"8D",X"28",X"86",X"01",X"8E",X"1B",X"6D",X"7E",
		X"00",X"A8",X"BD",X"1C",X"87",X"01",X"25",X"06",X"B5",X"7A",X"BE",X"56",X"EE",X"06",X"31",X"47",
		X"AC",X"A1",X"26",X"FC",X"4F",X"5F",X"ED",X"3E",X"6A",X"4F",X"26",X"05",X"30",X"C4",X"BD",X"00",
		X"EE",X"39",X"96",X"75",X"81",X"0A",X"24",X"18",X"BD",X"0D",X"48",X"17",X"0C",X"20",X"7F",X"17",
		X"B6",X"27",X"0D",X"D6",X"B7",X"1D",X"58",X"49",X"96",X"B6",X"84",X"1F",X"4C",X"A7",X"88",X"15",
		X"39",X"BD",X"01",X"A2",X"7E",X"00",X"00",X"34",X"10",X"BD",X"00",X"EC",X"35",X"10",X"20",X"0A",
		X"34",X"10",X"BD",X"00",X"EC",X"35",X"10",X"BD",X"01",X"A2",X"34",X"46",X"EE",X"64",X"37",X"06",
		X"BD",X"14",X"3A",X"8D",X"09",X"37",X"06",X"EF",X"64",X"BD",X"06",X"FD",X"35",X"C6",X"34",X"76",
		X"BD",X"00",X"00",X"BD",X"27",X"03",X"35",X"F6",X"8E",X"1C",X"C6",X"AF",X"47",X"86",X"06",X"8E",
		X"1C",X"B5",X"7E",X"00",X"A8",X"AE",X"47",X"EC",X"81",X"DD",X"33",X"A6",X"80",X"97",X"35",X"8C",
		X"1C",X"CF",X"25",X"E7",X"20",X"E2",X"81",X"81",X"2F",X"81",X"2F",X"07",X"2F",X"81",X"07",X"86",
		X"FF",X"97",X"30",X"0F",X"32",X"86",X"03",X"8E",X"1C",X"DD",X"7E",X"00",X"A8",X"96",X"B6",X"84",
		X"1F",X"8E",X"0F",X"E6",X"A6",X"86",X"97",X"30",X"97",X"32",X"8E",X"24",X"B7",X"9C",X"82",X"26",
		X"03",X"8E",X"24",X"C3",X"9F",X"82",X"86",X"06",X"8E",X"1C",X"CF",X"7E",X"00",X"A8",X"34",X"10",
		X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"05",X"1F",X"03",X"20",X"2A",
		X"34",X"10",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"05",X"1F",X"03",
		X"20",X"20",X"34",X"10",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"05",
		X"1F",X"03",X"35",X"32",X"36",X"32",X"33",X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",
		X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",
		X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",
		X"01",X"05",X"35",X"32",X"36",X"32",X"33",X"C9",X"01",X"05",X"35",X"32",X"36",X"32",X"10",X"DE",
		X"53",X"35",X"90",X"34",X"10",X"10",X"DF",X"53",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",
		X"05",X"1F",X"03",X"20",X"D5",X"34",X"10",X"CB",X"05",X"1F",X"03",X"4F",X"8E",X"00",X"00",X"31",
		X"84",X"20",X"46",X"34",X"10",X"CB",X"05",X"1F",X"03",X"4F",X"8E",X"00",X"00",X"31",X"84",X"20",
		X"20",X"34",X"10",X"CB",X"05",X"1F",X"03",X"4F",X"8E",X"00",X"00",X"31",X"84",X"20",X"18",X"34",
		X"10",X"CB",X"05",X"1F",X"03",X"4F",X"8E",X"00",X"00",X"31",X"84",X"36",X"32",X"33",X"C9",X"01",
		X"05",X"36",X"32",X"33",X"C9",X"01",X"05",X"36",X"32",X"33",X"C9",X"01",X"05",X"36",X"32",X"33",
		X"C9",X"01",X"05",X"36",X"32",X"33",X"C9",X"01",X"05",X"36",X"32",X"33",X"C9",X"01",X"05",X"36",
		X"32",X"33",X"C9",X"01",X"05",X"36",X"32",X"35",X"90",X"34",X"10",X"CB",X"05",X"1F",X"03",X"8E",
		X"00",X"00",X"31",X"84",X"4F",X"20",X"DC",X"34",X"76",X"96",X"DB",X"26",X"15",X"8E",X"07",X"20",
		X"B6",X"BD",X"E1",X"8D",X"0F",X"96",X"68",X"4A",X"27",X"08",X"8E",X"6D",X"20",X"B6",X"BE",X"20",
		X"8D",X"02",X"35",X"F6",X"34",X"02",X"CC",X"24",X"02",X"BD",X"13",X"B9",X"A6",X"E0",X"27",X"14",
		X"81",X"B4",X"23",X"02",X"86",X"B4",X"C6",X"FF",X"E7",X"84",X"E7",X"01",X"30",X"89",X"01",X"00",
		X"80",X"05",X"22",X"F2",X"39",X"34",X"76",X"96",X"DB",X"26",X"15",X"8E",X"07",X"13",X"B6",X"BD",
		X"DE",X"8D",X"0F",X"96",X"68",X"4A",X"27",X"08",X"8E",X"6D",X"13",X"B6",X"BE",X"1D",X"8D",X"02",
		X"35",X"F6",X"34",X"02",X"CC",X"24",X"06",X"BD",X"13",X"B9",X"A6",X"E4",X"81",X"11",X"23",X"02",
		X"86",X"11",X"81",X"0A",X"25",X"1B",X"80",X"0A",X"A7",X"E4",X"10",X"8E",X"20",X"A9",X"1F",X"10",
		X"BD",X"13",X"36",X"10",X"8E",X"1F",X"22",X"C3",X"00",X"02",X"BD",X"13",X"36",X"30",X"89",X"08",
		X"03",X"A6",X"E4",X"27",X"0F",X"1F",X"10",X"10",X"8E",X"1F",X"32",X"BD",X"13",X"36",X"8B",X"04",
		X"6A",X"E4",X"26",X"F7",X"35",X"82",X"34",X"76",X"CC",X"40",X"20",X"8E",X"2C",X"08",X"BD",X"13",
		X"B9",X"8E",X"00",X"08",X"CC",X"2F",X"28",X"BD",X"13",X"B9",X"8E",X"71",X"08",X"CC",X"2B",X"28",
		X"BD",X"13",X"B9",X"BD",X"1F",X"69",X"BD",X"1E",X"35",X"8D",X"10",X"BD",X"1D",X"F7",X"96",X"68",
		X"BD",X"14",X"BF",X"4A",X"26",X"FA",X"BD",X"37",X"43",X"35",X"F6",X"34",X"76",X"96",X"DB",X"26",
		X"15",X"8E",X"07",X"1A",X"B6",X"BD",X"E0",X"8D",X"0F",X"96",X"68",X"4A",X"27",X"08",X"8E",X"6D",
		X"1A",X"B6",X"BE",X"1F",X"8D",X"02",X"35",X"F6",X"34",X"02",X"CC",X"24",X"05",X"BD",X"13",X"B9",
		X"A6",X"E4",X"81",X"11",X"23",X"02",X"86",X"11",X"81",X"0A",X"25",X"11",X"80",X"0A",X"A7",X"E4",
		X"10",X"8E",X"1F",X"42",X"1F",X"10",X"BD",X"13",X"36",X"30",X"89",X"08",X"02",X"A6",X"E4",X"27",
		X"0F",X"10",X"8E",X"20",X"BD",X"1F",X"10",X"BD",X"13",X"36",X"8B",X"04",X"6A",X"E4",X"26",X"F7",
		X"35",X"82",X"04",X"03",X"1F",X"26",X"BB",X"0B",X"BB",X"9B",X"9B",X"96",X"99",X"90",X"99",X"9B",
		X"96",X"96",X"04",X"03",X"1F",X"36",X"BB",X"BB",X"B6",X"00",X"BE",X"66",X"00",X"F0",X"6F",X"00",
		X"00",X"F0",X"07",X"05",X"1F",X"46",X"99",X"00",X"00",X"00",X"99",X"00",X"90",X"99",X"90",X"00",
		X"09",X"92",X"92",X"92",X"09",X"99",X"92",X"92",X"92",X"99",X"99",X"22",X"92",X"22",X"99",X"90",
		X"9C",X"9C",X"9C",X"90",X"00",X"00",X"C0",X"00",X"00",X"96",X"DE",X"D6",X"DE",X"8E",X"00",X"2B",
		X"A7",X"84",X"30",X"89",X"01",X"00",X"8C",X"2C",X"08",X"25",X"F5",X"8E",X"6C",X"2B",X"A7",X"84",
		X"30",X"89",X"01",X"00",X"8C",X"9C",X"00",X"25",X"F5",X"B7",X"2C",X"07",X"B7",X"2D",X"07",X"B7",
		X"2C",X"24",X"B7",X"2D",X"24",X"84",X"0F",X"8E",X"2B",X"07",X"A7",X"80",X"8C",X"2B",X"2B",X"26",
		X"F9",X"96",X"DE",X"D6",X"DE",X"B7",X"6B",X"07",X"B7",X"6A",X"07",X"B7",X"6A",X"24",X"B7",X"6B",
		X"24",X"84",X"F0",X"8E",X"6C",X"07",X"A7",X"80",X"8C",X"6C",X"2B",X"26",X"F9",X"CC",X"99",X"99",
		X"8E",X"48",X"06",X"ED",X"84",X"ED",X"88",X"1E",X"30",X"89",X"01",X"00",X"8C",X"50",X"06",X"26",
		X"F2",X"39",X"00",X"F9",X"07",X"28",X"2F",X"00",X"A4",X"15",X"C7",X"FF",X"38",X"17",X"CC",X"81",
		X"81",X"2F",X"02",X"05",X"20",X"CB",X"02",X"10",X"20",X"D5",X"02",X"15",X"20",X"DF",X"02",X"20",
		X"20",X"E9",X"05",X"08",X"22",X"47",X"22",X"6F",X"02",X"6E",X"01",X"FA",X"04",X"08",X"22",X"97",
		X"22",X"97",X"02",X"14",X"02",X"46",X"04",X"08",X"22",X"B7",X"22",X"B7",X"02",X"14",X"02",X"46",
		X"01",X"01",X"20",X"1A",X"20",X"1A",X"14",X"19",X"14",X"19",X"00",X"04",X"08",X"22",X"D7",X"22",
		X"F7",X"02",X"14",X"02",X"46",X"02",X"08",X"23",X"17",X"23",X"27",X"01",X"D4",X"01",X"E6",X"02",
		X"08",X"23",X"37",X"23",X"47",X"01",X"D4",X"01",X"E6",X"02",X"08",X"23",X"57",X"23",X"67",X"01",
		X"D4",X"01",X"E6",X"02",X"08",X"23",X"77",X"23",X"87",X"01",X"D4",X"01",X"E6",X"04",X"08",X"23",
		X"97",X"23",X"B7",X"02",X"14",X"02",X"46",X"04",X"08",X"23",X"D7",X"23",X"F7",X"02",X"14",X"02",
		X"46",X"04",X"08",X"24",X"17",X"24",X"37",X"02",X"14",X"02",X"46",X"04",X"08",X"24",X"57",X"24",
		X"77",X"02",X"14",X"02",X"46",X"04",X"08",X"24",X"97",X"24",X"97",X"02",X"14",X"02",X"46",X"02",
		X"03",X"24",X"B7",X"24",X"BD",X"02",X"CC",X"02",X"E8",X"02",X"03",X"24",X"C3",X"24",X"C9",X"02",
		X"CC",X"02",X"E8",X"08",X"01",X"20",X"97",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",
		X"04",X"24",X"CF",X"24",X"DB",X"02",X"88",X"02",X"B2",X"08",X"06",X"24",X"E7",X"25",X"17",X"03",
		X"69",X"03",X"BA",X"08",X"06",X"25",X"47",X"25",X"77",X"03",X"69",X"03",X"BA",X"03",X"03",X"25",
		X"A7",X"06",X"05",X"20",X"F3",X"21",X"11",X"1D",X"10",X"1D",X"A1",X"06",X"05",X"21",X"2F",X"21",
		X"4D",X"1D",X"10",X"1D",X"A1",X"07",X"05",X"21",X"6B",X"21",X"8E",X"1C",X"FE",X"1D",X"93",X"07",
		X"05",X"21",X"B1",X"21",X"D4",X"1C",X"FE",X"1D",X"93",X"08",X"05",X"21",X"F7",X"22",X"1F",X"1D",
		X"22",X"1D",X"AF",X"11",X"00",X"11",X"10",X"11",X"10",X"10",X"10",X"00",X"10",X"11",X"10",X"11",
		X"00",X"11",X"10",X"00",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"10",
		X"10",X"01",X"00",X"01",X"01",X"01",X"11",X"01",X"11",X"00",X"11",X"01",X"01",X"01",X"00",X"01",
		X"11",X"00",X"11",X"01",X"11",X"01",X"01",X"01",X"01",X"01",X"11",X"01",X"01",X"01",X"11",X"FF",
		X"F0",X"FF",X"00",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",X"EE",X"E0",X"E0",X"E0",X"EE",X"E0",X"E0",
		X"E0",X"E0",X"E0",X"DD",X"D0",X"D0",X"D0",X"DD",X"D0",X"D0",X"D0",X"D0",X"D0",X"0F",X"0F",X"0F",
		X"00",X"0F",X"FF",X"00",X"FF",X"0F",X"FF",X"0E",X"0E",X"0E",X"0E",X"0E",X"EE",X"0E",X"0E",X"0E",
		X"EE",X"0D",X"0D",X"0D",X"0D",X"0D",X"DD",X"0D",X"0D",X"0D",X"DD",X"10",X"10",X"10",X"10",X"10",
		X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",
		X"10",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"10",X"10",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"01",X"01",X"01",X"11",X"01",X"01",X"01",
		X"01",X"01",X"11",X"01",X"01",X"01",X"11",X"01",X"01",X"01",X"01",X"01",X"11",X"01",X"01",X"01",
		X"11",X"C0",X"C0",X"C0",X"C0",X"C0",X"CC",X"C0",X"CC",X"00",X"CC",X"C0",X"00",X"C0",X"C0",X"C0",
		X"CC",X"C0",X"C0",X"C0",X"CC",X"C0",X"C0",X"C0",X"C0",X"C0",X"CC",X"C0",X"C0",X"C0",X"CC",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"0C",X"CC",X"00",
		X"CC",X"0C",X"CC",X"0C",X"0C",X"0C",X"0C",X"0C",X"CC",X"0C",X"0C",X"0C",X"CC",X"0C",X"0C",X"0C",
		X"0C",X"0C",X"CC",X"0C",X"0C",X"0C",X"CC",X"FF",X"00",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"00",
		X"F0",X"FF",X"F1",X"F1",X"F1",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"F1",X"F1",X"F1",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",
		X"00",X"0F",X"0F",X"0F",X"FF",X"0F",X"FF",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"1F",
		X"1F",X"1F",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"1F",X"1F",X"1F",X"FF",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"FF",X"1F",X"1F",X"1F",X"FF",X"00",X"03",X"F0",X"F0",X"F3",X"00",X"01",X"10",X"0C",
		X"0C",X"04",X"08",X"38",X"10",X"00",X"00",X"C0",X"C0",X"38",X"78",X"78",X"A0",X"A0",X"A0",X"00",
		X"33",X"03",X"03",X"33",X"10",X"01",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"10",X"00",
		X"00",X"0F",X"0F",X"0F",X"00",X"00",X"01",X"00",X"30",X"00",X"00",X"33",X"01",X"10",X"00",X"CC",
		X"CC",X"43",X"87",X"87",X"0A",X"0A",X"0A",X"00",X"03",X"80",X"80",X"83",X"01",X"00",X"00",X"00",
		X"30",X"3F",X"3F",X"3F",X"00",X"10",X"01",X"00",X"00",X"0D",X"6C",X"6C",X"0D",X"00",X"00",X"06",
		X"E6",X"C8",X"83",X"82",X"C8",X"EC",X"06",X"60",X"6D",X"8C",X"28",X"28",X"8C",X"6D",X"60",X"00",
		X"00",X"E0",X"C6",X"C6",X"E0",X"00",X"00",X"00",X"00",X"02",X"22",X"24",X"02",X"00",X"00",X"02",
		X"22",X"44",X"44",X"24",X"42",X"22",X"00",X"20",X"22",X"44",X"44",X"24",X"42",X"22",X"00",X"00",
		X"00",X"20",X"22",X"22",X"20",X"00",X"00",X"00",X"0E",X"00",X"D8",X"00",X"0E",X"00",X"00",X"0F",
		X"08",X"8C",X"C8",X"8C",X"08",X"0F",X"00",X"00",X"0E",X"80",X"C8",X"80",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"08",X"8C",X"08",X"E0",X"00",X"00",X"F0",X"80",X"C8",X"8C",X"C8",X"80",X"F0",X"00",X"00",
		X"E0",X"00",X"8D",X"00",X"E0",X"00",X"00",X"33",X"43",X"43",X"87",X"87",X"07",X"07",X"07",X"00",
		X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"03",X"04",X"04",X"08",X"08",X"00",X"00",X"00",X"30",
		X"30",X"38",X"78",X"78",X"70",X"70",X"70",X"33",X"43",X"43",X"87",X"87",X"77",X"77",X"77",X"00",
		X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"03",X"04",X"04",X"08",X"08",X"07",X"07",X"07",X"30",
		X"30",X"38",X"78",X"78",X"70",X"70",X"70",X"03",X"03",X"83",X"87",X"87",X"07",X"07",X"07",X"30",
		X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"33",
		X"34",X"34",X"78",X"78",X"70",X"70",X"70",X"03",X"03",X"83",X"87",X"87",X"07",X"07",X"07",X"30",
		X"40",X"40",X"80",X"80",X"70",X"70",X"70",X"00",X"00",X"08",X"08",X"08",X"00",X"00",X"00",X"33",
		X"34",X"34",X"78",X"78",X"77",X"77",X"77",X"08",X"08",X"DD",X"DE",X"DE",X"DE",X"DD",X"00",X"88",
		X"88",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"88",X"88",X"D8",X"D8",X"D8",X"D0",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"88",
		X"88",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"88",X"88",X"DD",X"ED",X"ED",X"ED",X"DD",X"00",X"80",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"DD",X"DE",X"DE",X"DE",X"DD",X"00",X"00",
		X"88",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"00",X"88",X"D8",X"D8",X"D8",X"D8",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"00",
		X"88",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"00",X"88",X"DD",X"ED",X"ED",X"ED",X"DD",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"DD",X"DE",X"DE",X"DE",X"DD",X"00",X"00",
		X"00",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"00",X"00",X"D8",X"D8",X"D8",X"D8",X"D8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"00",
		X"00",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"ED",X"ED",X"ED",X"DD",X"00",X"00",
		X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"DD",X"DE",X"DE",X"DE",X"DD",X"00",X"00",
		X"00",X"DD",X"EE",X"FE",X"EE",X"DD",X"88",X"00",X"00",X"D0",X"D8",X"D8",X"D8",X"D8",X"88",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"00",
		X"00",X"DD",X"EE",X"EF",X"EE",X"DD",X"88",X"00",X"00",X"DD",X"ED",X"ED",X"ED",X"DD",X"88",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"0C",X"CC",X"CC",X"CC",X"CC",X"0C",X"00",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",
		X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"00",X"A0",X"0A",X"A0",X"A0",X"00",X"A0",X"0A",X"00",X"0A",
		X"0A",X"A0",X"0A",X"0A",X"AA",X"0A",X"00",X"A0",X"00",X"00",X"0A",X"00",X"A0",X"AA",X"A0",X"00",
		X"02",X"23",X"02",X"20",X"22",X"23",X"22",X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"02",
		X"22",X"32",X"22",X"00",X"20",X"32",X"20",X"FB",X"0B",X"BB",X"0B",X"BB",X"06",X"00",X"B0",X"BB",
		X"B6",X"66",X"66",X"00",X"00",X"BB",X"66",X"66",X"FF",X"00",X"00",X"BB",X"66",X"66",X"F0",X"00",
		X"00",X"B0",X"6D",X"66",X"00",X"00",X"00",X"00",X"EF",X"66",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"0B",X"00",X"0B",X"00",X"B0",X"BB",X"BB",
		X"BB",X"B6",X"66",X"00",X"00",X"BB",X"66",X"66",X"6F",X"00",X"00",X"BB",X"66",X"66",X"FF",X"00",
		X"00",X"BB",X"66",X"66",X"00",X"00",X"00",X"00",X"DE",X"66",X"00",X"00",X"00",X"00",X"F0",X"6F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"0F",X"F6",X"00",X"00",X"00",X"00",X"ED",X"66",X"00",X"00",X"00",X"BB",X"66",X"66",X"00",X"00",
		X"00",X"BB",X"66",X"66",X"FF",X"00",X"00",X"BB",X"66",X"66",X"F6",X"0B",X"BB",X"BB",X"BB",X"6B",
		X"66",X"F0",X"00",X"B0",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"FE",X"66",X"00",X"00",X"00",X"0B",X"D6",X"66",X"00",X"00",
		X"00",X"BB",X"66",X"66",X"0F",X"00",X"00",X"BB",X"66",X"66",X"FF",X"00",X"0B",X"BB",X"6B",X"66",
		X"66",X"BF",X"B0",X"BB",X"B0",X"BB",X"60",X"90",X"09",X"90",X"99",X"99",X"99",X"90",X"CC",X"90",
		X"DE",X"3F",X"A6",X"47",X"4C",X"81",X"04",X"23",X"01",X"4F",X"A7",X"47",X"26",X"17",X"BD",X"5F",
		X"D0",X"81",X"05",X"22",X"10",X"8E",X"9C",X"41",X"CE",X"BC",X"83",X"8D",X"74",X"8E",X"9C",X"47",
		X"8D",X"6F",X"7E",X"11",X"4C",X"8E",X"9C",X"41",X"7E",X"11",X"42",X"EC",X"0A",X"93",X"4F",X"44",
		X"44",X"E6",X"0C",X"54",X"54",X"54",X"C3",X"2C",X"03",X"ED",X"C4",X"EC",X"88",X"12",X"27",X"4F",
		X"10",X"83",X"90",X"00",X"27",X"49",X"10",X"83",X"40",X"00",X"27",X"43",X"81",X"33",X"27",X"3F",
		X"10",X"83",X"66",X"66",X"27",X"39",X"10",X"83",X"44",X"33",X"27",X"33",X"81",X"1F",X"26",X"2C",
		X"EC",X"C4",X"81",X"6B",X"26",X"03",X"4A",X"A7",X"C4",X"10",X"8E",X"FF",X"F0",X"10",X"AF",X"D1",
		X"5C",X"ED",X"C4",X"10",X"8E",X"F0",X"FF",X"10",X"AF",X"D1",X"4C",X"ED",X"C4",X"10",X"8E",X"F0",
		X"F0",X"10",X"AF",X"D1",X"5A",X"ED",X"C4",X"10",X"AF",X"D1",X"20",X"05",X"CC",X"99",X"99",X"ED",
		X"D1",X"AE",X"84",X"26",X"96",X"39",X"34",X"17",X"0F",X"87",X"1F",X"01",X"A6",X"84",X"0D",X"91",
		X"10",X"2A",X"E0",X"B1",X"81",X"F0",X"10",X"24",X"E0",X"AB",X"35",X"97",X"D6",X"91",X"2A",X"16",
		X"54",X"25",X"13",X"F6",X"C8",X"04",X"C4",X"7D",X"DA",X"F1",X"D7",X"57",X"F6",X"C8",X"06",X"C4",
		X"FE",X"DA",X"F2",X"7E",X"07",X"8C",X"F6",X"C8",X"04",X"7E",X"07",X"87",X"34",X"76",X"0D",X"91",
		X"2B",X"05",X"1A",X"01",X"7E",X"14",X"3E",X"35",X"F6",X"EC",X"02",X"10",X"83",X"20",X"10",X"10",
		X"27",X"F1",X"AA",X"AD",X"98",X"08",X"7E",X"18",X"23",X"96",X"DB",X"26",X"07",X"96",X"8F",X"81",
		X"04",X"24",X"01",X"39",X"7E",X"00",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"27",X"09",X"7E",X"27",X"87",X"7E",X"28",X"45",X"34",X"66",X"10",X"8E",X"BE",X"6E",X"C6",
		X"56",X"0D",X"91",X"2B",X"13",X"E1",X"A8",X"54",X"27",X"0E",X"96",X"B7",X"81",X"0D",X"22",X"08",
		X"D6",X"B8",X"86",X"9C",X"1F",X"02",X"6A",X"A4",X"96",X"DB",X"26",X"1E",X"8D",X"4A",X"22",X"1A",
		X"96",X"91",X"85",X"04",X"26",X"14",X"EC",X"0A",X"93",X"20",X"10",X"83",X"26",X"00",X"22",X"0A",
		X"BD",X"27",X"DE",X"24",X"09",X"BD",X"28",X"22",X"24",X"F6",X"9F",X"41",X"35",X"E6",X"96",X"91",
		X"2B",X"06",X"CC",X"06",X"A1",X"BD",X"06",X"FD",X"A6",X"88",X"14",X"8A",X"02",X"A7",X"88",X"14",
		X"CC",X"2F",X"00",X"ED",X"22",X"6F",X"27",X"EC",X"02",X"ED",X"24",X"CC",X"20",X"10",X"ED",X"02",
		X"9F",X"41",X"6F",X"26",X"AF",X"2C",X"35",X"E6",X"EC",X"98",X"02",X"C1",X"0F",X"22",X"07",X"5C",
		X"54",X"3D",X"10",X"83",X"00",X"19",X"39",X"34",X"66",X"96",X"DB",X"26",X"4F",X"8D",X"E9",X"22",
		X"4B",X"96",X"91",X"85",X"04",X"26",X"45",X"EC",X"0A",X"93",X"20",X"81",X"26",X"22",X"3D",X"DD",
		X"BD",X"BD",X"27",X"F8",X"24",X"08",X"BD",X"28",X"22",X"25",X"31",X"BD",X"27",X"F8",X"CC",X"01",
		X"00",X"ED",X"22",X"6F",X"27",X"EE",X"02",X"EF",X"24",X"6F",X"26",X"DC",X"BD",X"58",X"49",X"58",
		X"49",X"E6",X"0C",X"ED",X"28",X"DC",X"D0",X"A3",X"28",X"A1",X"C4",X"24",X"04",X"E1",X"41",X"25",
		X"04",X"EC",X"C4",X"44",X"54",X"54",X"ED",X"2A",X"E3",X"28",X"ED",X"28",X"35",X"E6",X"34",X"10",
		X"10",X"9E",X"DF",X"27",X"0F",X"AE",X"A4",X"9F",X"DF",X"9E",X"E1",X"AF",X"A4",X"10",X"9F",X"E1",
		X"1C",X"FE",X"35",X"90",X"1A",X"01",X"35",X"90",X"34",X"10",X"10",X"9E",X"DF",X"27",X"F5",X"AE",
		X"A4",X"9F",X"DF",X"9E",X"E3",X"AF",X"A4",X"10",X"9F",X"E3",X"1C",X"FE",X"35",X"90",X"34",X"10",
		X"AE",X"A4",X"AF",X"9F",X"9C",X"B9",X"9E",X"DF",X"AF",X"A4",X"10",X"9F",X"DF",X"10",X"9E",X"B9",
		X"35",X"90",X"34",X"10",X"10",X"8E",X"9C",X"E3",X"10",X"9F",X"B9",X"10",X"9E",X"E3",X"27",X"C4",
		X"AE",X"A4",X"27",X"08",X"10",X"9F",X"B9",X"10",X"AE",X"A4",X"20",X"F4",X"BD",X"29",X"45",X"8D",
		X"CD",X"1C",X"FE",X"35",X"90",X"96",X"DB",X"27",X"01",X"39",X"96",X"91",X"85",X"04",X"27",X"33",
		X"10",X"8E",X"9C",X"E1",X"10",X"9F",X"B9",X"10",X"AE",X"A4",X"27",X"16",X"EC",X"24",X"AE",X"2C",
		X"ED",X"02",X"A6",X"88",X"14",X"84",X"FD",X"A7",X"88",X"14",X"BD",X"29",X"45",X"BD",X"28",X"0E",
		X"20",X"E2",X"10",X"8E",X"9C",X"E3",X"10",X"9F",X"B9",X"10",X"AE",X"A4",X"27",X"CB",X"BD",X"28",
		X"0E",X"20",X"F3",X"96",X"3A",X"81",X"02",X"C6",X"08",X"24",X"01",X"50",X"1D",X"D3",X"C5",X"10",
		X"83",X"01",X"40",X"23",X"03",X"CC",X"01",X"40",X"10",X"83",X"00",X"AA",X"24",X"03",X"CC",X"00",
		X"AA",X"DD",X"C5",X"10",X"9E",X"E3",X"27",X"3F",X"DC",X"20",X"C4",X"C0",X"DD",X"BD",X"DC",X"22",
		X"C4",X"C0",X"93",X"BD",X"58",X"49",X"58",X"49",X"97",X"C4",X"10",X"8E",X"9C",X"E3",X"10",X"9F",
		X"B9",X"10",X"AE",X"A4",X"27",X"21",X"EC",X"22",X"D3",X"C5",X"ED",X"22",X"81",X"30",X"23",X"08",
		X"BD",X"29",X"45",X"BD",X"28",X"0E",X"20",X"E6",X"D6",X"C4",X"1D",X"E3",X"27",X"ED",X"27",X"BD",
		X"29",X"45",X"BD",X"29",X"A5",X"20",X"D7",X"10",X"8E",X"9C",X"E1",X"10",X"9F",X"B9",X"10",X"AE",
		X"A4",X"27",X"51",X"EC",X"22",X"83",X"01",X"00",X"ED",X"22",X"2B",X"0C",X"AE",X"2C",X"EC",X"0A",
		X"93",X"20",X"8B",X"0C",X"85",X"C0",X"27",X"16",X"EC",X"24",X"AE",X"2C",X"ED",X"02",X"A6",X"88",
		X"14",X"84",X"FD",X"A7",X"88",X"14",X"BD",X"29",X"45",X"BD",X"28",X"0E",X"20",X"CD",X"80",X"0C",
		X"58",X"49",X"58",X"49",X"E6",X"0C",X"DD",X"4F",X"C6",X"DA",X"3D",X"48",X"EE",X"24",X"E6",X"C4",
		X"3D",X"E6",X"41",X"54",X"54",X"ED",X"2A",X"59",X"D3",X"4F",X"ED",X"28",X"BD",X"29",X"45",X"BD",
		X"29",X"A5",X"20",X"A7",X"39",X"E6",X"26",X"27",X"5B",X"C0",X"32",X"22",X"57",X"50",X"8E",X"29",
		X"59",X"3A",X"54",X"3A",X"CC",X"00",X"00",X"6E",X"84",X"ED",X"B8",X"3E",X"ED",X"B8",X"3C",X"ED",
		X"B8",X"3A",X"ED",X"B8",X"38",X"ED",X"B8",X"36",X"ED",X"B8",X"34",X"ED",X"B8",X"32",X"ED",X"B8",
		X"30",X"ED",X"B8",X"2E",X"ED",X"B8",X"2C",X"ED",X"B8",X"2A",X"ED",X"B8",X"28",X"ED",X"B8",X"26",
		X"ED",X"B8",X"24",X"ED",X"B8",X"22",X"ED",X"B8",X"20",X"ED",X"B8",X"1E",X"ED",X"B8",X"1C",X"ED",
		X"B8",X"1A",X"ED",X"B8",X"18",X"ED",X"B8",X"16",X"ED",X"B8",X"14",X"ED",X"B8",X"12",X"ED",X"B8",
		X"10",X"ED",X"B8",X"0E",X"39",X"EE",X"24",X"37",X"16",X"DD",X"C1",X"A6",X"22",X"97",X"BB",X"E6",
		X"2A",X"3D",X"DD",X"BD",X"EC",X"27",X"93",X"BD",X"4D",X"27",X"14",X"D7",X"BE",X"D6",X"C2",X"3A",
		X"0A",X"C1",X"26",X"03",X"7E",X"2B",X"1D",X"D6",X"BE",X"DB",X"BB",X"89",X"00",X"26",X"EC",X"DD",
		X"BD",X"C1",X"98",X"10",X"22",X"01",X"46",X"96",X"BB",X"48",X"97",X"BC",X"E6",X"2B",X"3D",X"DD",
		X"BF",X"E6",X"29",X"4F",X"97",X"C3",X"93",X"BF",X"4D",X"27",X"11",X"0C",X"C3",X"0A",X"C2",X"0A",
		X"C2",X"2E",X"03",X"7E",X"2B",X"1D",X"DB",X"BC",X"89",X"00",X"26",X"EF",X"C1",X"2C",X"25",X"EB",
		X"D7",X"C0",X"08",X"C3",X"CE",X"2B",X"20",X"96",X"C2",X"48",X"EE",X"C6",X"34",X"60",X"31",X"2E",
		X"96",X"C3",X"30",X"86",X"96",X"BE",X"6E",X"C4",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",
		X"25",X"4C",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"25",X"46",X"ED",X"A4",X"EE",X"81",
		X"EF",X"B1",X"DB",X"BC",X"25",X"40",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"25",X"3A",
		X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"25",X"34",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",
		X"DB",X"BC",X"25",X"2E",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"0A",X"C1",X"27",X"28",X"9B",X"BB",
		X"25",X"24",X"81",X"98",X"22",X"20",X"D6",X"C3",X"3A",X"D6",X"C0",X"6E",X"F8",X"02",X"C6",X"0C",
		X"20",X"7F",X"C6",X"0A",X"20",X"7B",X"C6",X"08",X"20",X"77",X"C6",X"06",X"20",X"73",X"C6",X"04",
		X"20",X"6F",X"C6",X"02",X"20",X"6B",X"20",X"7D",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",
		X"24",X"04",X"C6",X"0D",X"20",X"5B",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"24",X"04",
		X"C6",X"0B",X"20",X"4D",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"24",X"04",X"C6",X"09",
		X"20",X"3F",X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"24",X"04",X"C6",X"07",X"20",X"31",
		X"ED",X"A4",X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"24",X"04",X"C6",X"05",X"20",X"23",X"ED",X"A4",
		X"EE",X"81",X"EF",X"B1",X"DB",X"BC",X"24",X"04",X"C6",X"03",X"20",X"15",X"ED",X"A4",X"EE",X"81",
		X"EF",X"B1",X"DB",X"BC",X"24",X"04",X"C6",X"01",X"20",X"07",X"ED",X"A4",X"EE",X"80",X"EF",X"B1",
		X"5F",X"0A",X"C1",X"27",X"10",X"9B",X"BB",X"25",X"0C",X"81",X"98",X"22",X"08",X"DB",X"C3",X"3A",
		X"D6",X"C0",X"6E",X"F8",X"02",X"AE",X"E4",X"1F",X"20",X"A3",X"E4",X"C0",X"0E",X"E7",X"06",X"AE",
		X"08",X"8C",X"98",X"00",X"22",X"05",X"CC",X"00",X"00",X"ED",X"84",X"35",X"E0",X"6F",X"26",X"39",
		X"2A",X"5A",X"2A",X"EA",X"2A",X"54",X"2A",X"DC",X"2A",X"4A",X"2A",X"CE",X"2A",X"40",X"2A",X"C0",
		X"2A",X"36",X"2A",X"B2",X"2A",X"2C",X"2A",X"A4",X"2A",X"22",X"2A",X"96",X"2A",X"18",X"2A",X"88",
		X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"2E",X"20",X"31",X"39",X"38",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"27",X"03",X"BD",X"5F",X"CA",X"96",X"F3",X"26",X"36",X"9E",X"5E",X"26",X"0D",X"9E",X"62",X"27",
		X"12",X"DC",X"64",X"0F",X"62",X"0F",X"63",X"7E",X"00",X"91",X"DC",X"60",X"0F",X"5E",X"0F",X"5F",
		X"7E",X"00",X"91",X"9E",X"F4",X"27",X"09",X"DC",X"F6",X"0F",X"F4",X"0F",X"F5",X"7E",X"00",X"91",
		X"9E",X"FB",X"10",X"27",X"D4",X"F4",X"DC",X"FD",X"0F",X"FB",X"0F",X"FC",X"7E",X"00",X"91",X"7E",
		X"00",X"9A",X"26",X"06",X"DD",X"5E",X"9F",X"60",X"20",X"18",X"DE",X"62",X"26",X"06",X"DD",X"62",
		X"9F",X"64",X"20",X"0E",X"DE",X"F4",X"26",X"06",X"DD",X"F4",X"9F",X"F6",X"20",X"04",X"DD",X"FB",
		X"9F",X"FD",X"35",X"46",X"4D",X"10",X"26",X"DB",X"BD",X"39",X"96",X"66",X"26",X"03",X"7E",X"00",
		X"E4",X"7E",X"5F",X"CD",X"6F",X"0B",X"6F",X"06",X"7E",X"0A",X"58",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"2C",X"0C",X"7E",X"2C",X"C6",X"7E",X"2C",X"B9",X"7E",X"31",X"4A",X"8E",X"D0",X"04",X"96",
		X"91",X"2B",X"1C",X"4F",X"AB",X"84",X"30",X"09",X"8C",X"F0",X"00",X"25",X"F7",X"81",X"56",X"27",
		X"0E",X"D6",X"B7",X"C1",X"16",X"22",X"08",X"D6",X"B6",X"86",X"9C",X"1F",X"02",X"63",X"A4",X"BD",
		X"2C",X"7F",X"BD",X"2C",X"AC",X"8E",X"A6",X"34",X"9F",X"04",X"86",X"E0",X"97",X"08",X"C6",X"01",
		X"B6",X"30",X"49",X"48",X"25",X"01",X"50",X"CB",X"E0",X"D7",X"09",X"86",X"FF",X"97",X"07",X"86",
		X"80",X"97",X"06",X"0F",X"0A",X"86",X"4D",X"97",X"02",X"BD",X"2E",X"C4",X"0A",X"02",X"26",X"F9",
		X"8E",X"00",X"00",X"9F",X"02",X"9E",X"02",X"30",X"89",X"00",X"80",X"27",X"0B",X"9F",X"02",X"9C",
		X"20",X"24",X"05",X"BD",X"2E",X"C4",X"20",X"ED",X"DC",X"20",X"C4",X"80",X"DD",X"00",X"39",X"8E",
		X"30",X"49",X"CE",X"A1",X"00",X"C6",X"E0",X"E7",X"C0",X"10",X"8E",X"00",X"04",X"A6",X"80",X"48",
		X"24",X"03",X"5C",X"20",X"01",X"5A",X"48",X"24",X"03",X"5C",X"20",X"01",X"5A",X"11",X"83",X"A5",
		X"00",X"27",X"08",X"E7",X"C0",X"31",X"3F",X"26",X"E6",X"20",X"DE",X"39",X"8E",X"A5",X"00",X"4F",
		X"5F",X"ED",X"81",X"4C",X"81",X"99",X"23",X"F9",X"39",X"4F",X"5F",X"8E",X"A5",X"00",X"ED",X"91",
		X"8C",X"A6",X"34",X"26",X"F9",X"39",X"DC",X"20",X"C4",X"80",X"93",X"00",X"58",X"49",X"27",X"28",
		X"97",X"02",X"2B",X"10",X"96",X"0A",X"2A",X"03",X"BD",X"2D",X"F1",X"BD",X"2E",X"C4",X"0A",X"02",
		X"26",X"F9",X"20",X"0E",X"96",X"0A",X"2B",X"03",X"BD",X"2E",X"1A",X"BD",X"2E",X"3F",X"0C",X"02",
		X"26",X"F9",X"DC",X"20",X"C4",X"80",X"DD",X"00",X"10",X"DF",X"02",X"DC",X"20",X"10",X"DE",X"04",
		X"C5",X"20",X"27",X"04",X"32",X"E9",X"03",X"9C",X"C5",X"40",X"27",X"02",X"32",X"63",X"8E",X"00",
		X"00",X"86",X"09",X"10",X"8E",X"A5",X"04",X"32",X"66",X"AF",X"B4",X"35",X"44",X"E7",X"21",X"EF",
		X"B4",X"AF",X"B8",X"02",X"35",X"44",X"E7",X"23",X"EF",X"B8",X"02",X"AF",X"B8",X"04",X"35",X"44",
		X"E7",X"25",X"EF",X"B8",X"04",X"AF",X"B8",X"06",X"35",X"44",X"E7",X"27",X"EF",X"B8",X"06",X"AF",
		X"B8",X"08",X"35",X"44",X"E7",X"29",X"EF",X"B8",X"08",X"AF",X"B8",X"0A",X"35",X"44",X"E7",X"2B",
		X"EF",X"B8",X"0A",X"AF",X"B8",X"0C",X"35",X"44",X"E7",X"2D",X"EF",X"B8",X"0C",X"AF",X"B8",X"0E",
		X"35",X"44",X"E7",X"2F",X"EF",X"B8",X"0E",X"AF",X"B8",X"10",X"35",X"44",X"E7",X"A8",X"11",X"EF",
		X"B8",X"10",X"AF",X"B8",X"12",X"35",X"44",X"E7",X"A8",X"13",X"EF",X"B8",X"12",X"AF",X"B8",X"14",
		X"35",X"44",X"E7",X"A8",X"15",X"EF",X"B8",X"14",X"AF",X"B8",X"16",X"35",X"44",X"E7",X"A8",X"17",
		X"EF",X"B8",X"16",X"AF",X"B8",X"18",X"35",X"44",X"E7",X"A8",X"19",X"EF",X"B8",X"18",X"AF",X"B8",
		X"1A",X"35",X"44",X"E7",X"A8",X"1B",X"EF",X"B8",X"1A",X"AF",X"B8",X"1C",X"35",X"44",X"E7",X"A8",
		X"1D",X"EF",X"B8",X"1C",X"AF",X"B8",X"1E",X"35",X"44",X"E7",X"A8",X"1F",X"EF",X"B8",X"1E",X"31",
		X"A8",X"20",X"4A",X"10",X"26",X"FF",X"52",X"AF",X"B4",X"35",X"44",X"E7",X"21",X"EF",X"B4",X"AF",
		X"B8",X"02",X"35",X"44",X"E7",X"23",X"EF",X"B8",X"02",X"AF",X"B8",X"04",X"35",X"44",X"E7",X"25",
		X"EF",X"B8",X"04",X"AF",X"B8",X"06",X"35",X"44",X"E7",X"27",X"EF",X"B8",X"06",X"10",X"DE",X"02",
		X"39",X"03",X"0A",X"96",X"06",X"8B",X"27",X"97",X"06",X"9E",X"04",X"30",X"89",X"01",X"CB",X"A6",
		X"01",X"E6",X"84",X"84",X"0F",X"26",X"01",X"5C",X"D7",X"08",X"A6",X"89",X"03",X"9D",X"E6",X"89",
		X"03",X"9C",X"84",X"0F",X"26",X"01",X"5C",X"D7",X"09",X"39",X"03",X"0A",X"96",X"06",X"80",X"27",
		X"97",X"06",X"9E",X"04",X"A6",X"01",X"E6",X"84",X"84",X"0F",X"27",X"01",X"5C",X"D7",X"08",X"A6",
		X"89",X"03",X"9D",X"E6",X"89",X"03",X"9C",X"84",X"0F",X"27",X"01",X"5C",X"D7",X"09",X"39",X"8E",
		X"30",X"C9",X"D6",X"06",X"EC",X"85",X"58",X"49",X"58",X"49",X"1F",X"89",X"46",X"03",X"07",X"2B",
		X"0A",X"44",X"44",X"44",X"44",X"54",X"54",X"54",X"54",X"0A",X"06",X"84",X"0F",X"C4",X"0F",X"8E",
		X"2F",X"C9",X"48",X"48",X"48",X"58",X"58",X"58",X"31",X"85",X"30",X"86",X"DE",X"04",X"33",X"5A",
		X"11",X"83",X"A6",X"34",X"24",X"03",X"CE",X"A7",X"FC",X"DF",X"04",X"EC",X"02",X"DB",X"08",X"ED",
		X"42",X"ED",X"C9",X"01",X"D0",X"EC",X"84",X"AB",X"43",X"AB",X"07",X"ED",X"C4",X"ED",X"C9",X"01",
		X"CE",X"AB",X"06",X"97",X"08",X"EC",X"04",X"ED",X"44",X"ED",X"C9",X"01",X"D2",X"30",X"C9",X"03",
		X"9C",X"EC",X"22",X"DB",X"09",X"ED",X"02",X"ED",X"89",X"01",X"D0",X"EC",X"A4",X"AB",X"03",X"AB",
		X"27",X"ED",X"84",X"ED",X"89",X"01",X"CE",X"AB",X"26",X"97",X"09",X"EC",X"24",X"ED",X"04",X"ED",
		X"89",X"01",X"D2",X"39",X"8E",X"30",X"C9",X"D6",X"06",X"EC",X"85",X"58",X"49",X"1F",X"89",X"46",
		X"03",X"07",X"2B",X"0A",X"44",X"44",X"44",X"44",X"54",X"54",X"54",X"54",X"20",X"06",X"84",X"0F",
		X"C4",X"0F",X"0C",X"06",X"8E",X"2F",X"49",X"48",X"48",X"48",X"58",X"58",X"58",X"31",X"85",X"30",
		X"86",X"DE",X"04",X"EC",X"84",X"9B",X"08",X"ED",X"C4",X"ED",X"C9",X"01",X"CE",X"EC",X"02",X"EB",
		X"C4",X"EB",X"06",X"ED",X"42",X"ED",X"C9",X"01",X"D0",X"EB",X"07",X"D7",X"08",X"EC",X"04",X"ED",
		X"44",X"ED",X"C9",X"01",X"D2",X"30",X"C9",X"03",X"9C",X"EC",X"A4",X"9B",X"09",X"ED",X"84",X"ED",
		X"89",X"01",X"CE",X"EC",X"22",X"EB",X"84",X"EB",X"26",X"ED",X"02",X"ED",X"89",X"01",X"D0",X"EB",
		X"27",X"D7",X"09",X"EC",X"24",X"ED",X"04",X"ED",X"89",X"01",X"D2",X"33",X"46",X"11",X"83",X"A8",
		X"02",X"25",X"03",X"CE",X"A6",X"34",X"DF",X"04",X"39",X"FE",X"07",X"70",X"FE",X"07",X"70",X"00",
		X"00",X"FE",X"07",X"70",X"FF",X"70",X"07",X"00",X"01",X"FE",X"07",X"70",X"00",X"07",X"70",X"00",
		X"00",X"FE",X"07",X"70",X"01",X"70",X"07",X"00",X"01",X"FF",X"70",X"07",X"FE",X"07",X"70",X"01",
		X"00",X"FF",X"70",X"07",X"FF",X"70",X"07",X"01",X"01",X"FF",X"70",X"07",X"00",X"07",X"70",X"01",
		X"00",X"FF",X"70",X"07",X"01",X"70",X"07",X"01",X"01",X"00",X"07",X"70",X"FE",X"07",X"70",X"00",
		X"00",X"00",X"07",X"70",X"FF",X"70",X"07",X"00",X"01",X"00",X"07",X"70",X"00",X"07",X"70",X"00",
		X"00",X"00",X"07",X"70",X"01",X"70",X"07",X"00",X"01",X"01",X"70",X"07",X"FE",X"07",X"70",X"01",
		X"00",X"01",X"70",X"07",X"FF",X"70",X"07",X"01",X"01",X"01",X"70",X"07",X"00",X"07",X"70",X"01",
		X"00",X"01",X"70",X"07",X"01",X"70",X"07",X"01",X"01",X"01",X"07",X"70",X"01",X"07",X"70",X"01",
		X"01",X"01",X"07",X"70",X"FF",X"07",X"70",X"01",X"01",X"01",X"07",X"70",X"00",X"70",X"07",X"01",
		X"00",X"01",X"07",X"70",X"FE",X"70",X"07",X"01",X"00",X"FF",X"07",X"70",X"01",X"07",X"70",X"01",
		X"01",X"FF",X"07",X"70",X"FF",X"07",X"70",X"01",X"01",X"FF",X"07",X"70",X"00",X"70",X"07",X"01",
		X"00",X"FF",X"07",X"70",X"FE",X"70",X"07",X"01",X"00",X"00",X"70",X"07",X"01",X"07",X"70",X"00",
		X"01",X"00",X"70",X"07",X"FF",X"07",X"70",X"00",X"01",X"00",X"70",X"07",X"00",X"70",X"07",X"00",
		X"00",X"00",X"70",X"07",X"FE",X"70",X"07",X"00",X"00",X"FE",X"70",X"07",X"01",X"07",X"70",X"00",
		X"01",X"FE",X"70",X"07",X"FF",X"07",X"70",X"00",X"01",X"FE",X"70",X"07",X"00",X"70",X"07",X"00",
		X"00",X"FE",X"70",X"07",X"FE",X"70",X"07",X"00",X"00",X"55",X"40",X"00",X"00",X"00",X"00",X"3F",
		X"FF",X"FF",X"FF",X"FC",X"00",X"07",X"FF",X"FF",X"D3",X"D5",X"54",X"79",X"C7",X"55",X"4D",X"55",
		X"4A",X"AB",X"24",X"00",X"0A",X"A8",X"00",X"0A",X"A8",X"00",X"0A",X"AB",X"FF",X"F5",X"57",X"FF",
		X"F5",X"57",X"FF",X"F6",X"CD",X"55",X"AD",X"69",X"AA",X"AA",X"AA",X"AA",X"AE",X"21",X"BA",X"AA",
		X"AA",X"00",X"0F",X"FE",X"A8",X"08",X"81",X"01",X"FF",X"80",X"2A",X"00",X"05",X"12",X"51",X"DB",
		X"77",X"BF",X"BF",X"EF",X"FF",X"F5",X"55",X"55",X"55",X"54",X"15",X"55",X"55",X"F5",X"55",X"50",
		X"3A",X"AA",X"8E",X"6A",X"AA",X"7D",X"55",X"02",X"EA",X"A8",X"80",X"3A",X"AA",X"8F",X"FB",X"7C",
		X"A4",X"76",X"40",X"10",X"00",X"03",X"E2",X"08",X"BB",X"14",X"00",X"80",X"D3",X"FF",X"FD",X"E2",
		X"FE",X"D5",X"5F",X"A1",X"A5",X"6C",X"07",X"00",X"04",X"00",X"D0",X"00",X"0A",X"08",X"00",X"01",
		X"D4",X"3F",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"7F",X"FC",X"FF",X"FE",X"AA",X"87",X"EA",X"AA",
		X"81",X"F0",X"AA",X"AA",X"AA",X"8F",X"AA",X"AA",X"83",X"C0",X"7F",X"F5",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"40",X"AC",X"10",X"8C",X"04",X"02",X"20",X"03",X"F7",X"FF",X"FE",X"F9",
		X"AA",X"C2",X"77",X"8E",X"00",X"00",X"00",X"02",X"7B",X"DF",X"FF",X"DF",X"FE",X"FF",X"AA",X"AA",
		X"07",X"D5",X"55",X"50",X"7E",X"AA",X"AA",X"AA",X"A8",X"1A",X"AA",X"AB",X"7A",X"AA",X"80",X"0E",
		X"AA",X"AA",X"FC",X"8F",X"E3",X"A5",X"35",X"55",X"55",X"55",X"55",X"55",X"43",X"AA",X"AA",X"3E",
		X"AA",X"A8",X"1D",X"55",X"55",X"54",X"7E",X"AA",X"86",X"A5",X"55",X"69",X"55",X"55",X"55",X"2A",
		X"AB",X"26",X"A3",X"8C",X"00",X"00",X"0F",X"FF",X"FF",X"55",X"35",X"06",X"ED",X"4D",X"AF",X"4A",
		X"1F",X"10",X"BD",X"01",X"88",X"AF",X"47",X"E7",X"0C",X"44",X"56",X"44",X"56",X"D3",X"20",X"ED",
		X"0A",X"CC",X"31",X"A9",X"0D",X"92",X"2A",X"03",X"CC",X"31",X"B3",X"ED",X"02",X"86",X"0D",X"A7",
		X"49",X"BD",X"19",X"43",X"0F",X"CF",X"BD",X"19",X"43",X"1C",X"CF",X"BD",X"19",X"43",X"1C",X"A8",
		X"AE",X"47",X"96",X"B8",X"84",X"07",X"D6",X"B7",X"C4",X"03",X"5C",X"E3",X"4A",X"DD",X"D0",X"BD",
		X"27",X"03",X"6A",X"49",X"27",X"08",X"86",X"01",X"8E",X"31",X"80",X"7E",X"00",X"A8",X"86",X"60",
		X"8E",X"31",X"A6",X"7E",X"00",X"A8",X"6E",X"D8",X"0D",X"08",X"06",X"31",X"BD",X"31",X"BD",X"03",
		X"69",X"03",X"BA",X"08",X"06",X"31",X"ED",X"31",X"ED",X"03",X"69",X"03",X"BA",X"00",X"09",X"11",
		X"01",X"11",X"F1",X"11",X"19",X"AD",X"DD",X"A9",X"1F",X"19",X"10",X"9A",X"AF",X"A9",X"11",X"01",
		X"19",X"A9",X"11",X"A9",X"F1",X"00",X"11",X"91",X"1A",X"A9",X"1A",X"00",X"01",X"9F",X"1A",X"91",
		X"F1",X"00",X"00",X"19",X"F1",X"11",X"1A",X"00",X"00",X"01",X"F9",X"1A",X"19",X"00",X"00",X"00",
		X"1A",X"11",X"A9",X"00",X"00",X"11",X"A1",X"A1",X"A9",X"00",X"00",X"11",X"1F",X"F1",X"A9",X"00",
		X"01",X"19",X"19",X"A1",X"01",X"01",X"A1",X"91",X"19",X"A9",X"F1",X"11",X"11",X"9A",X"FD",X"AA",
		X"11",X"10",X"11",X"9A",X"DF",X"A9",X"F1",X"10",X"19",X"1F",X"A0",X"19",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"32",X"CD",X"11",X"22",X"33",X"44",X"55",X"66",X"77",X"88",X"FF",X"3F",X"F8",X"07",X"FF",
		X"38",X"C7",X"C0",X"5F",X"4F",X"FD",X"9D",X"06",X"ED",X"81",X"8D",X"43",X"ED",X"81",X"8D",X"54",
		X"FC",X"9D",X"06",X"ED",X"81",X"8D",X"38",X"43",X"53",X"C3",X"00",X"01",X"ED",X"81",X"8D",X"44",
		X"FC",X"9D",X"06",X"43",X"53",X"C3",X"00",X"01",X"ED",X"0E",X"ED",X"81",X"8D",X"21",X"ED",X"81",
		X"8D",X"32",X"30",X"02",X"8D",X"19",X"43",X"53",X"C3",X"00",X"01",X"ED",X"81",X"8D",X"25",X"FC",
		X"9D",X"06",X"C3",X"00",X"14",X"10",X"83",X"01",X"40",X"25",X"BA",X"BF",X"9D",X"0A",X"39",X"BD",
		X"33",X"FA",X"2A",X"04",X"CA",X"C0",X"20",X"02",X"C4",X"3F",X"1D",X"B3",X"9D",X"06",X"C3",X"01",
		X"40",X"47",X"56",X"39",X"4F",X"5F",X"ED",X"81",X"ED",X"81",X"CC",X"50",X"00",X"ED",X"81",X"CC",
		X"50",X"80",X"ED",X"81",X"6F",X"80",X"A6",X"9F",X"9D",X"08",X"A7",X"80",X"39",X"DE",X"3F",X"35",
		X"10",X"AF",X"4D",X"8E",X"9C",X"27",X"10",X"8E",X"9D",X"0E",X"CE",X"32",X"4B",X"EC",X"84",X"ED",
		X"A1",X"EC",X"C1",X"ED",X"81",X"8C",X"9C",X"2F",X"26",X"F3",X"CC",X"33",X"F2",X"BD",X"06",X"FD",
		X"FC",X"9D",X"0C",X"C3",X"34",X"56",X"FD",X"9D",X"0C",X"CC",X"32",X"43",X"FD",X"9D",X"08",X"86",
		X"07",X"B7",X"9D",X"03",X"86",X"09",X"B7",X"9D",X"02",X"86",X"07",X"B7",X"9D",X"01",X"86",X"01",
		X"B7",X"9D",X"00",X"8E",X"9D",X"16",X"BD",X"32",X"53",X"4F",X"7A",X"9D",X"00",X"26",X"0B",X"B6",
		X"9D",X"01",X"B7",X"9D",X"00",X"CE",X"32",X"49",X"A6",X"C6",X"97",X"26",X"B6",X"9D",X"02",X"4A",
		X"B7",X"9D",X"02",X"26",X"05",X"BD",X"33",X"C2",X"20",X"08",X"86",X"02",X"8E",X"33",X"42",X"7E",
		X"00",X"A8",X"10",X"8E",X"00",X"00",X"8E",X"9D",X"16",X"BC",X"9D",X"0A",X"26",X"18",X"0F",X"26",
		X"10",X"8E",X"9C",X"27",X"8E",X"9D",X"0E",X"EC",X"81",X"ED",X"A1",X"10",X"8C",X"9C",X"2F",X"26",
		X"F6",X"DE",X"3F",X"6E",X"D8",X"0D",X"BC",X"9D",X"0A",X"27",X"AE",X"10",X"AF",X"98",X"0A",X"EC",
		X"84",X"E3",X"06",X"ED",X"06",X"E3",X"0B",X"81",X"F6",X"24",X"21",X"81",X"0A",X"25",X"1D",X"ED",
		X"0B",X"EC",X"02",X"E3",X"04",X"ED",X"04",X"E3",X"08",X"81",X"9C",X"24",X"0F",X"ED",X"08",X"A7",
		X"0A",X"A6",X"0D",X"E6",X"0D",X"ED",X"98",X"0A",X"30",X"0E",X"20",X"CA",X"FE",X"9D",X"0A",X"33",
		X"52",X"FF",X"9D",X"0A",X"EC",X"C4",X"ED",X"84",X"EC",X"42",X"ED",X"02",X"EC",X"44",X"ED",X"04",
		X"EC",X"46",X"ED",X"06",X"EC",X"48",X"ED",X"08",X"EC",X"4A",X"ED",X"0A",X"EC",X"4C",X"ED",X"0C",
		X"20",X"A4",X"B6",X"9D",X"01",X"4A",X"81",X"05",X"25",X"03",X"B7",X"9D",X"01",X"86",X"09",X"B7",
		X"9D",X"02",X"7D",X"9D",X"03",X"27",X"3E",X"7A",X"9D",X"03",X"FC",X"9D",X"08",X"C3",X"00",X"01",
		X"10",X"83",X"32",X"4B",X"26",X"03",X"CC",X"32",X"43",X"FD",X"9D",X"08",X"BE",X"9D",X"0A",X"7E",
		X"32",X"53",X"FF",X"20",X"02",X"F2",X"60",X"01",X"F2",X"00",X"FC",X"9D",X"0C",X"46",X"56",X"B6",
		X"9D",X"0C",X"48",X"B8",X"9D",X"0C",X"F7",X"9D",X"0C",X"48",X"F6",X"9D",X"0D",X"56",X"46",X"B7",
		X"9D",X"0D",X"F6",X"9D",X"0D",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"35",X"50",X"11",X"22",X"33",X"44",X"55",X"66",X"77",X"88",X"07",X"F8",X"01",X"FE",X"03",
		X"FC",X"00",X"FF",X"03",X"FC",X"03",X"FC",X"01",X"FE",X"07",X"F8",X"34",X"67",X"34",X"6C",X"34",
		X"71",X"34",X"76",X"34",X"7B",X"34",X"6C",X"E8",X"01",X"08",X"17",X"00",X"E8",X"01",X"18",X"11",
		X"00",X"E8",X"01",X"0A",X"06",X"00",X"E8",X"01",X"08",X"14",X"00",X"E8",X"01",X"08",X"01",X"01",
		X"01",X"13",X"00",X"8C",X"AC",X"AD",X"24",X"75",X"BD",X"36",X"D9",X"C4",X"07",X"58",X"10",X"8E",
		X"34",X"4B",X"10",X"AE",X"A5",X"10",X"BF",X"9D",X"00",X"BD",X"36",X"D9",X"FC",X"9D",X"15",X"81",
		X"9C",X"24",X"F6",X"C1",X"0A",X"23",X"F2",X"C1",X"F6",X"24",X"EE",X"FD",X"9D",X"0E",X"4F",X"5F",
		X"FD",X"9D",X"06",X"ED",X"81",X"8D",X"4A",X"ED",X"81",X"8D",X"61",X"FC",X"9D",X"06",X"ED",X"81",
		X"8D",X"3F",X"43",X"53",X"C3",X"00",X"01",X"ED",X"81",X"8D",X"51",X"FC",X"9D",X"06",X"43",X"53",
		X"C3",X"00",X"01",X"34",X"06",X"ED",X"81",X"8D",X"28",X"ED",X"81",X"8D",X"3F",X"35",X"06",X"ED",
		X"81",X"8D",X"1E",X"43",X"53",X"C3",X"00",X"01",X"ED",X"81",X"8D",X"30",X"8C",X"AC",X"AD",X"24",
		X"0C",X"FC",X"9D",X"06",X"C3",X"00",X"60",X"10",X"83",X"08",X"00",X"25",X"B3",X"BF",X"9D",X"12",
		X"39",X"BD",X"36",X"D9",X"5F",X"B6",X"9D",X"16",X"2A",X"06",X"BA",X"9D",X"01",X"53",X"20",X"03",
		X"B4",X"9D",X"00",X"B3",X"9D",X"06",X"C3",X"08",X"00",X"47",X"56",X"39",X"FC",X"9D",X"0E",X"ED",
		X"81",X"A7",X"80",X"B6",X"9D",X"0F",X"ED",X"81",X"A6",X"9F",X"9D",X"10",X"A7",X"80",X"39",X"B6",
		X"9D",X"15",X"84",X"07",X"8B",X"02",X"B7",X"9D",X"09",X"BD",X"36",X"D9",X"CA",X"80",X"57",X"1D",
		X"83",X"00",X"80",X"FD",X"9D",X"0C",X"BD",X"36",X"D9",X"1D",X"58",X"49",X"FD",X"9D",X"0A",X"39",
		X"DE",X"3F",X"35",X"10",X"AF",X"4D",X"9E",X"6C",X"9F",X"DC",X"8E",X"36",X"F5",X"9F",X"6C",X"DC",
		X"B7",X"FD",X"9D",X"15",X"CC",X"34",X"43",X"FD",X"9D",X"10",X"86",X"10",X"B7",X"9D",X"03",X"86",
		X"30",X"B7",X"9D",X"02",X"86",X"01",X"B7",X"9D",X"08",X"86",X"FF",X"97",X"2D",X"8E",X"9D",X"17",
		X"10",X"8E",X"A5",X"00",X"8D",X"A9",X"FC",X"9D",X"0A",X"ED",X"02",X"FC",X"9D",X"0C",X"ED",X"84",
		X"EC",X"A1",X"ED",X"04",X"ED",X"06",X"86",X"77",X"A7",X"09",X"30",X"0A",X"10",X"8C",X"A6",X"34",
		X"24",X"07",X"7A",X"9D",X"09",X"26",X"DF",X"20",X"DB",X"BF",X"9D",X"12",X"B6",X"9D",X"03",X"81",
		X"10",X"26",X"2F",X"B6",X"9D",X"02",X"81",X"20",X"27",X"08",X"81",X"10",X"27",X"04",X"81",X"01",
		X"26",X"03",X"BD",X"36",X"AF",X"7A",X"9D",X"08",X"26",X"18",X"86",X"03",X"B7",X"9D",X"08",X"CC",
		X"34",X"7B",X"BD",X"06",X"FD",X"8E",X"0F",X"E6",X"BD",X"36",X"D9",X"C4",X"1F",X"A6",X"85",X"B7",
		X"9D",X"14",X"B6",X"9D",X"02",X"4A",X"B7",X"9D",X"02",X"26",X"05",X"BD",X"36",X"62",X"20",X"08",
		X"86",X"01",X"8E",X"35",X"F8",X"7E",X"00",X"A8",X"86",X"08",X"97",X"3A",X"BE",X"9D",X"12",X"8C",
		X"9D",X"7B",X"24",X"0B",X"9E",X"DC",X"9F",X"6C",X"0F",X"26",X"DE",X"3F",X"6E",X"D8",X"0D",X"8E",
		X"9D",X"17",X"10",X"8E",X"00",X"00",X"BC",X"9D",X"12",X"27",X"91",X"10",X"AF",X"98",X"06",X"EC",
		X"84",X"E3",X"07",X"81",X"F6",X"24",X"1D",X"81",X"0A",X"25",X"19",X"ED",X"07",X"EC",X"02",X"E3",
		X"04",X"81",X"9C",X"24",X"0F",X"ED",X"04",X"A7",X"06",X"A6",X"09",X"E6",X"09",X"ED",X"98",X"06",
		X"30",X"0A",X"20",X"D2",X"FE",X"9D",X"12",X"33",X"56",X"FF",X"9D",X"12",X"EC",X"42",X"ED",X"02",
		X"EC",X"C4",X"ED",X"84",X"EC",X"44",X"ED",X"04",X"EC",X"46",X"ED",X"06",X"EC",X"48",X"ED",X"08",
		X"20",X"B4",X"B6",X"9D",X"15",X"84",X"07",X"8B",X"02",X"B7",X"9D",X"02",X"7D",X"9D",X"03",X"27",
		X"3D",X"86",X"10",X"B0",X"9D",X"03",X"81",X"0A",X"23",X"09",X"81",X"14",X"22",X"05",X"86",X"04",
		X"B7",X"9D",X"02",X"7A",X"9D",X"03",X"FC",X"9D",X"10",X"C3",X"00",X"01",X"10",X"83",X"34",X"4B",
		X"26",X"03",X"CC",X"34",X"43",X"FD",X"9D",X"10",X"8D",X"2D",X"F6",X"9D",X"15",X"C4",X"1F",X"10",
		X"8E",X"0F",X"E6",X"E6",X"A5",X"F7",X"9D",X"14",X"BE",X"9D",X"12",X"7E",X"34",X"83",X"39",X"8E",
		X"9D",X"17",X"BC",X"9D",X"12",X"27",X"3D",X"EC",X"02",X"58",X"49",X"ED",X"02",X"EC",X"84",X"58",
		X"49",X"ED",X"84",X"30",X"0A",X"20",X"EB",X"BD",X"36",X"D9",X"C4",X"0E",X"C1",X"0C",X"24",X"F7",
		X"10",X"8E",X"34",X"5B",X"EC",X"A5",X"7E",X"06",X"FD",X"FC",X"9D",X"15",X"46",X"56",X"B6",X"9D",
		X"15",X"48",X"B8",X"9D",X"15",X"F7",X"9D",X"15",X"48",X"F6",X"9D",X"16",X"56",X"46",X"B7",X"9D",
		X"16",X"F6",X"9D",X"16",X"39",X"B6",X"CB",X"00",X"81",X"10",X"24",X"1F",X"B6",X"9D",X"14",X"26",
		X"15",X"96",X"26",X"85",X"C0",X"27",X"02",X"80",X"40",X"85",X"38",X"27",X"02",X"80",X"08",X"85",
		X"07",X"27",X"06",X"4A",X"20",X"03",X"7F",X"9D",X"14",X"97",X"26",X"6E",X"9F",X"9C",X"DC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"37",X"A3",X"7E",X"37",X"91",X"96",X"91",X"85",X"2C",X"26",X"2B",X"B6",X"BD",X"D0",X"27",
		X"26",X"7A",X"BD",X"D0",X"26",X"21",X"B6",X"BD",X"CF",X"85",X"10",X"27",X"0D",X"F6",X"BD",X"D3",
		X"10",X"BE",X"BD",X"D4",X"BE",X"BD",X"CD",X"7E",X"37",X"9C",X"8E",X"00",X"00",X"BF",X"BD",X"CD",
		X"8D",X"06",X"86",X"05",X"7E",X"38",X"34",X"39",X"34",X"72",X"8E",X"00",X"00",X"31",X"84",X"4F",
		X"CE",X"2C",X"2C",X"36",X"32",X"33",X"C9",X"01",X"05",X"11",X"83",X"6C",X"2C",X"25",X"F4",X"35",
		X"F2",X"CC",X"00",X"00",X"FD",X"BD",X"CD",X"B7",X"BD",X"D0",X"20",X"D4",X"34",X"16",X"BE",X"BD",
		X"CB",X"20",X"11",X"34",X"16",X"B6",X"BD",X"D0",X"27",X"08",X"A6",X"84",X"A1",X"9F",X"BD",X"CD",
		X"25",X"57",X"30",X"01",X"A6",X"80",X"B7",X"BD",X"CF",X"85",X"20",X"27",X"08",X"EC",X"81",X"10",
		X"B3",X"BD",X"CD",X"26",X"44",X"A6",X"80",X"B7",X"BD",X"D0",X"B6",X"BD",X"CF",X"85",X"04",X"27",
		X"02",X"8D",X"A5",X"A6",X"80",X"97",X"EC",X"BF",X"BD",X"CB",X"E6",X"61",X"AE",X"62",X"F7",X"BD",
		X"D3",X"10",X"BF",X"BD",X"D4",X"BF",X"BD",X"CD",X"BD",X"38",X"34",X"B6",X"BD",X"CF",X"85",X"08",
		X"27",X"0B",X"BE",X"BD",X"CB",X"AE",X"84",X"BF",X"BD",X"CD",X"BD",X"37",X"A3",X"B6",X"BD",X"CF",
		X"85",X"40",X"27",X"05",X"BD",X"19",X"43",X"38",X"0B",X"35",X"96",X"FC",X"BD",X"CD",X"ED",X"47",
		X"B6",X"BD",X"D2",X"97",X"2B",X"B6",X"BD",X"D1",X"8E",X"38",X"1E",X"7E",X"00",X"A8",X"FC",X"BD",
		X"CD",X"10",X"A3",X"47",X"26",X"0B",X"0F",X"2B",X"B6",X"BD",X"D1",X"8E",X"38",X"10",X"7E",X"00",
		X"A8",X"7E",X"00",X"E4",X"BD",X"70",X"52",X"86",X"01",X"97",X"39",X"39",X"00",X"00",X"00",X"00",
		X"7E",X"38",X"5E",X"7E",X"40",X"8F",X"7E",X"42",X"54",X"7E",X"41",X"DE",X"7E",X"39",X"39",X"7E",
		X"39",X"79",X"43",X"9F",X"3D",X"FB",X"3F",X"45",X"3B",X"A3",X"3C",X"6B",X"3D",X"33",X"96",X"B6",
		X"81",X"C0",X"10",X"23",X"01",X"13",X"BD",X"38",X"4C",X"38",X"91",X"43",X"9F",X"39",X"2E",X"33",
		X"33",X"27",X"1D",X"7C",X"BE",X"7F",X"86",X"03",X"A7",X"4C",X"DC",X"B6",X"84",X"1F",X"D3",X"20",
		X"ED",X"0A",X"54",X"CB",X"2C",X"E7",X"0C",X"86",X"08",X"A7",X"49",X"8D",X"6B",X"7E",X"27",X"00",
		X"39",X"AE",X"47",X"EC",X"02",X"10",X"83",X"20",X"10",X"27",X"3B",X"6A",X"49",X"26",X"13",X"B6",
		X"BE",X"6E",X"BD",X"08",X"C1",X"A7",X"49",X"BD",X"45",X"4C",X"27",X"06",X"CC",X"06",X"E2",X"BD",
		X"06",X"FD",X"6A",X"4C",X"26",X"06",X"86",X"03",X"A7",X"4C",X"8D",X"35",X"EC",X"04",X"27",X"16",
		X"86",X"06",X"A7",X"4B",X"86",X"01",X"8E",X"38",X"CC",X"7E",X"00",X"A8",X"AE",X"47",X"8D",X"0E",
		X"6A",X"4B",X"26",X"F0",X"20",X"BB",X"86",X"06",X"8E",X"38",X"91",X"7E",X"00",X"A8",X"10",X"AE",
		X"02",X"31",X"2A",X"10",X"8C",X"43",X"DB",X"23",X"04",X"10",X"8E",X"43",X"9F",X"10",X"AF",X"02",
		X"39",X"96",X"B6",X"B1",X"BE",X"6F",X"23",X"35",X"CC",X"40",X"01",X"DD",X"4F",X"EC",X"0A",X"93",
		X"A3",X"2B",X"02",X"00",X"4F",X"C3",X"02",X"80",X"10",X"83",X"05",X"00",X"23",X"07",X"D6",X"4F",
		X"1D",X"D3",X"9E",X"ED",X"0E",X"A6",X"0C",X"90",X"97",X"2B",X"02",X"00",X"50",X"8B",X"0A",X"81",
		X"14",X"23",X"0A",X"5F",X"96",X"50",X"D3",X"A1",X"47",X"56",X"ED",X"88",X"10",X"39",X"7A",X"BE",
		X"7F",X"BD",X"1C",X"80",X"01",X"20",X"06",X"B0",X"39",X"34",X"26",X"9E",X"43",X"27",X"31",X"9E",
		X"3D",X"27",X"2D",X"4F",X"EE",X"64",X"37",X"10",X"BD",X"01",X"30",X"31",X"84",X"BD",X"01",X"88",
		X"37",X"06",X"ED",X"02",X"37",X"06",X"ED",X"08",X"37",X"06",X"ED",X"88",X"12",X"EF",X"64",X"33",
		X"A4",X"EF",X"06",X"AF",X"47",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"0E",X"86",X"01",X"35",X"A6",
		X"EE",X"64",X"33",X"48",X"EF",X"64",X"4F",X"35",X"A6",X"BD",X"38",X"4C",X"39",X"BA",X"3D",X"FB",
		X"3A",X"AF",X"33",X"33",X"27",X"33",X"7C",X"BE",X"81",X"6F",X"49",X"DC",X"B6",X"84",X"1F",X"D3",
		X"20",X"ED",X"0A",X"54",X"CB",X"2C",X"E7",X"0C",X"B6",X"BE",X"78",X"BD",X"08",X"C1",X"A7",X"4D",
		X"10",X"8E",X"3B",X"67",X"96",X"B6",X"84",X"03",X"26",X"04",X"31",X"A9",X"00",X"0C",X"10",X"AF",
		X"4B",X"8D",X"4E",X"BD",X"3B",X"41",X"7E",X"27",X"00",X"39",X"AE",X"47",X"EC",X"02",X"10",X"83",
		X"20",X"10",X"27",X"2E",X"86",X"FF",X"D6",X"97",X"E0",X"0C",X"CB",X"14",X"C1",X"0A",X"24",X"02",
		X"86",X"FC",X"AB",X"4D",X"81",X"FC",X"25",X"13",X"BD",X"3A",X"38",X"B6",X"BE",X"78",X"10",X"AE",
		X"4B",X"10",X"8C",X"3B",X"73",X"26",X"01",X"44",X"BD",X"08",X"C1",X"A7",X"4D",X"8D",X"0B",X"BD",
		X"3B",X"41",X"86",X"06",X"8E",X"39",X"BA",X"7E",X"00",X"A8",X"96",X"B6",X"B1",X"BE",X"77",X"23",
		X"36",X"CC",X"20",X"01",X"DD",X"4F",X"EC",X"0A",X"93",X"A3",X"2B",X"02",X"00",X"4F",X"C3",X"02",
		X"80",X"10",X"83",X"05",X"00",X"23",X"07",X"D6",X"4F",X"1D",X"D3",X"9E",X"ED",X"0E",X"A6",X"0C",
		X"90",X"97",X"80",X"04",X"2B",X"02",X"00",X"50",X"8B",X"0A",X"81",X"14",X"23",X"09",X"96",X"50",
		X"D3",X"A1",X"47",X"56",X"ED",X"88",X"10",X"39",X"34",X"76",X"A6",X"0A",X"90",X"20",X"81",X"26",
		X"22",X"60",X"B6",X"BE",X"80",X"81",X"0C",X"24",X"59",X"31",X"84",X"BD",X"38",X"4C",X"3A",X"CF",
		X"3B",X"51",X"3A",X"A4",X"33",X"00",X"27",X"4A",X"7C",X"BE",X"80",X"CC",X"3A",X"BA",X"BD",X"06",
		X"FD",X"6F",X"49",X"96",X"B6",X"84",X"03",X"27",X"01",X"4A",X"C6",X"0C",X"3D",X"C3",X"3B",X"7F",
		X"ED",X"4B",X"C6",X"40",X"BD",X"08",X"C1",X"A6",X"2A",X"91",X"A3",X"2B",X"01",X"50",X"1D",X"D3",
		X"9E",X"ED",X"0E",X"B6",X"BE",X"79",X"44",X"BD",X"08",X"C1",X"A7",X"4A",X"BD",X"07",X"EC",X"D6",
		X"B7",X"1D",X"ED",X"88",X"10",X"EC",X"2A",X"ED",X"0A",X"EC",X"2C",X"ED",X"0C",X"BD",X"3B",X"41",
		X"9F",X"41",X"35",X"F6",X"7A",X"BE",X"80",X"BD",X"1C",X"80",X"00",X"50",X"3A",X"C7",X"39",X"7A",
		X"BE",X"81",X"BD",X"1C",X"80",X"01",X"20",X"3A",X"BF",X"39",X"D0",X"01",X"10",X"18",X"00",X"D0",
		X"01",X"0C",X"01",X"01",X"08",X"17",X"00",X"D0",X"01",X"0C",X"1A",X"01",X"08",X"17",X"00",X"AE",
		X"47",X"6A",X"4A",X"26",X"62",X"F6",X"BE",X"7A",X"4F",X"34",X"06",X"50",X"1D",X"34",X"06",X"B6",
		X"BE",X"7B",X"5F",X"34",X"06",X"40",X"34",X"06",X"DC",X"B7",X"84",X"01",X"D3",X"A3",X"A3",X"0A",
		X"DD",X"4F",X"DC",X"B6",X"84",X"07",X"D3",X"9C",X"A3",X"0C",X"DD",X"51",X"07",X"4F",X"06",X"50",
		X"07",X"51",X"06",X"52",X"DC",X"4F",X"2A",X"07",X"10",X"A3",X"64",X"2D",X"EF",X"20",X"05",X"10",
		X"A3",X"66",X"22",X"E8",X"DC",X"51",X"2A",X"07",X"10",X"A3",X"E4",X"2D",X"DF",X"20",X"05",X"10",
		X"A3",X"62",X"22",X"D8",X"32",X"68",X"ED",X"88",X"10",X"DC",X"4F",X"D3",X"9E",X"ED",X"0E",X"B6",
		X"BE",X"79",X"BD",X"08",X"C1",X"A7",X"4A",X"8D",X"08",X"86",X"06",X"8E",X"3A",X"CF",X"7E",X"00",
		X"A8",X"34",X"26",X"A6",X"49",X"4C",X"E6",X"0E",X"2B",X"07",X"81",X"02",X"23",X"0D",X"4F",X"20",
		X"0A",X"81",X"05",X"22",X"04",X"81",X"03",X"24",X"02",X"86",X"03",X"A7",X"49",X"10",X"AE",X"4B",
		X"48",X"EC",X"A6",X"ED",X"02",X"35",X"A6",X"3D",X"FB",X"3E",X"05",X"3E",X"0F",X"3D",X"FB",X"3E",
		X"19",X"3E",X"23",X"3F",X"45",X"3F",X"4F",X"3F",X"59",X"3F",X"45",X"3F",X"63",X"3F",X"6D",X"3D",
		X"33",X"3D",X"3D",X"3D",X"47",X"3D",X"33",X"3D",X"51",X"3D",X"5B",X"3C",X"6B",X"3C",X"75",X"3C",
		X"7F",X"3C",X"6B",X"3C",X"89",X"3C",X"93",X"3B",X"A3",X"3B",X"AD",X"3B",X"B7",X"3B",X"A3",X"3B",
		X"C1",X"3B",X"CB",X"03",X"05",X"3B",X"D5",X"3C",X"20",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3B",
		X"E4",X"3C",X"2F",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3B",X"F3",X"3C",X"3E",X"1D",X"73",X"1D",
		X"85",X"03",X"05",X"3C",X"02",X"3C",X"4D",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3C",X"11",X"3C",
		X"5C",X"1D",X"73",X"1D",X"85",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"40",
		X"40",X"40",X"40",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"44",X"40",X"00",
		X"00",X"00",X"40",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"00",X"44",X"44",X"40",X"40",X"00",
		X"40",X"40",X"44",X"00",X"00",X"00",X"44",X"44",X"04",X"04",X"04",X"44",X"40",X"40",X"40",X"40",
		X"40",X"44",X"44",X"00",X"44",X"44",X"44",X"44",X"04",X"44",X"44",X"40",X"40",X"40",X"40",X"40",
		X"04",X"04",X"04",X"04",X"04",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"04",
		X"04",X"04",X"04",X"04",X"44",X"40",X"40",X"40",X"44",X"44",X"00",X"00",X"00",X"44",X"04",X"04",
		X"04",X"04",X"04",X"44",X"44",X"40",X"44",X"44",X"44",X"44",X"00",X"44",X"44",X"04",X"00",X"00",
		X"00",X"04",X"44",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"04",X"04",X"00",X"04",
		X"04",X"44",X"44",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"03",X"05",X"3C",X"9D",X"3C",
		X"E8",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3C",X"AC",X"3C",X"F7",X"1D",X"73",X"1D",X"85",X"03",
		X"05",X"3C",X"BB",X"3D",X"06",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3C",X"CA",X"3D",X"15",X"1D",
		X"73",X"1D",X"85",X"03",X"05",X"3C",X"D9",X"3D",X"24",X"1D",X"73",X"1D",X"85",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"20",X"20",X"20",X"20",X"20",X"22",X"22",X"22",X"22",
		X"22",X"22",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"00",X"20",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"00",X"22",X"22",X"20",X"20",X"00",X"20",X"20",X"22",X"00",X"00",X"00",X"22",X"22",
		X"02",X"02",X"02",X"22",X"20",X"20",X"20",X"20",X"20",X"22",X"22",X"00",X"22",X"22",X"22",X"22",
		X"02",X"22",X"22",X"20",X"20",X"20",X"20",X"20",X"02",X"02",X"02",X"02",X"02",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"02",X"02",X"02",X"02",X"02",X"22",X"20",X"20",X"20",
		X"22",X"22",X"00",X"00",X"00",X"22",X"02",X"02",X"02",X"02",X"02",X"22",X"22",X"20",X"22",X"22",
		X"22",X"22",X"00",X"22",X"22",X"02",X"00",X"00",X"00",X"02",X"22",X"00",X"00",X"00",X"22",X"22",
		X"22",X"22",X"22",X"22",X"02",X"02",X"00",X"02",X"02",X"22",X"22",X"00",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"03",X"05",X"3D",X"65",X"3D",X"B0",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3D",
		X"74",X"3D",X"BF",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3D",X"83",X"3D",X"CE",X"1D",X"73",X"1D",
		X"85",X"03",X"05",X"3D",X"92",X"3D",X"DD",X"1D",X"73",X"1D",X"85",X"03",X"05",X"3D",X"A1",X"3D",
		X"EC",X"1D",X"73",X"1D",X"85",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"30",
		X"30",X"30",X"30",X"30",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"33",X"30",X"00",
		X"00",X"00",X"30",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"33",X"33",X"30",X"30",X"00",
		X"30",X"30",X"33",X"00",X"00",X"00",X"33",X"33",X"03",X"03",X"03",X"33",X"30",X"30",X"30",X"30",
		X"30",X"33",X"33",X"00",X"33",X"33",X"33",X"33",X"03",X"33",X"33",X"30",X"30",X"30",X"30",X"30",
		X"03",X"03",X"03",X"03",X"03",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"03",
		X"03",X"03",X"03",X"03",X"33",X"30",X"30",X"30",X"33",X"33",X"00",X"00",X"00",X"33",X"03",X"03",
		X"03",X"03",X"03",X"33",X"33",X"30",X"33",X"33",X"33",X"33",X"00",X"33",X"33",X"03",X"00",X"00",
		X"00",X"03",X"33",X"00",X"00",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"03",X"03",X"00",X"03",
		X"03",X"33",X"33",X"00",X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"03",X"07",X"3E",X"2D",X"3E",
		X"B9",X"04",X"3B",X"04",X"4D",X"04",X"07",X"3E",X"49",X"3E",X"D5",X"04",X"3B",X"04",X"4D",X"04",
		X"07",X"3E",X"65",X"3E",X"F1",X"04",X"3B",X"04",X"4D",X"04",X"07",X"3E",X"81",X"3F",X"0D",X"04",
		X"3B",X"04",X"4D",X"04",X"07",X"3E",X"9D",X"3F",X"29",X"04",X"3B",X"04",X"4D",X"99",X"98",X"98",
		X"98",X"98",X"98",X"99",X"99",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"88",
		X"88",X"99",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"99",X"98",X"98",X"98",X"98",X"98",X"99",
		X"99",X"90",X"90",X"90",X"90",X"90",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",
		X"00",X"00",X"00",X"00",X"90",X"99",X"98",X"98",X"98",X"98",X"98",X"99",X"99",X"88",X"99",X"90",
		X"99",X"88",X"99",X"99",X"88",X"99",X"00",X"99",X"88",X"99",X"90",X"90",X"90",X"00",X"90",X"90",
		X"90",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"99",
		X"98",X"98",X"98",X"98",X"98",X"99",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"99",X"98",X"99",
		X"00",X"99",X"98",X"99",X"99",X"88",X"99",X"00",X"99",X"88",X"99",X"99",X"88",X"98",X"98",X"98",
		X"88",X"99",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"09",X"09",X"09",X"09",X"09",X"09",X"09",
		X"99",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"88",X"88",X"88",X"88",X"88",X"99",X"99",X"89",
		X"89",X"89",X"89",X"89",X"99",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"99",X"89",X"89",X"89",
		X"89",X"89",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"99",X"09",X"09",X"09",X"09",X"09",X"09",X"09",X"99",X"88",X"89",X"89",X"89",X"88",X"99",X"99",
		X"88",X"99",X"00",X"99",X"88",X"99",X"99",X"89",X"99",X"00",X"99",X"89",X"99",X"09",X"00",X"00",
		X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"09",X"09",X"09",X"09",
		X"09",X"99",X"99",X"89",X"89",X"89",X"89",X"89",X"99",X"09",X"09",X"09",X"00",X"09",X"09",X"09",
		X"99",X"88",X"99",X"00",X"99",X"88",X"99",X"99",X"88",X"99",X"09",X"99",X"88",X"99",X"99",X"89",
		X"89",X"89",X"89",X"89",X"99",X"04",X"07",X"3F",X"77",X"40",X"03",X"04",X"3B",X"04",X"4D",X"04",
		X"07",X"3F",X"93",X"40",X"1F",X"04",X"3B",X"04",X"4D",X"04",X"07",X"3F",X"AF",X"40",X"3B",X"04",
		X"3B",X"04",X"4D",X"04",X"07",X"3F",X"CB",X"40",X"57",X"04",X"3B",X"04",X"4D",X"04",X"07",X"3F",
		X"E7",X"40",X"73",X"04",X"3B",X"04",X"4D",X"FF",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"FF",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",
		X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",X"FF",X"BB",X"FF",X"F0",X"FF",X"BB",X"FF",X"FF",X"BB",X"FF",
		X"00",X"FF",X"BB",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FB",X"FB",X"FB",X"FB",X"FB",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FB",X"FF",X"00",X"FF",X"FB",X"FF",X"FF",X"BB",
		X"FF",X"00",X"FF",X"BB",X"FF",X"FF",X"BB",X"FB",X"FB",X"FB",X"BB",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"FF",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"FF",X"BB",X"BF",X"BF",X"BF",X"BB",X"FF",X"FF",X"BB",X"FF",X"00",X"FF",X"BB",X"FF",
		X"FF",X"BF",X"FF",X"00",X"FF",X"BF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"BF",X"BF",X"BF",
		X"BF",X"BF",X"FF",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"FF",X"BB",X"FF",X"00",X"FF",X"BB",
		X"FF",X"FF",X"BB",X"FF",X"0F",X"FF",X"BB",X"FF",X"FF",X"BF",X"BF",X"BF",X"BF",X"BF",X"FF",X"97",
		X"4F",X"10",X"9E",X"B7",X"34",X"20",X"96",X"B6",X"84",X"01",X"D6",X"B7",X"C3",X"00",X"80",X"34",
		X"06",X"BD",X"19",X"43",X"41",X"23",X"EC",X"E4",X"ED",X"07",X"BD",X"01",X"70",X"20",X"1B",X"41",
		X"73",X"CC",X"CC",X"BD",X"07",X"EC",X"D6",X"B8",X"54",X"CB",X"2C",X"E7",X"0C",X"D6",X"B6",X"C4",
		X"3F",X"96",X"4F",X"46",X"24",X"01",X"50",X"1D",X"ED",X"0E",X"2A",X"05",X"50",X"8D",X"41",X"20",
		X"07",X"8D",X"3D",X"43",X"53",X"C3",X"00",X"01",X"34",X"06",X"D6",X"B7",X"1D",X"58",X"49",X"58",
		X"49",X"58",X"49",X"58",X"49",X"E3",X"64",X"E3",X"E4",X"E3",X"E4",X"ED",X"0A",X"32",X"62",X"D6",
		X"B8",X"C4",X"7F",X"C0",X"40",X"1D",X"2B",X"04",X"CA",X"20",X"20",X"02",X"C4",X"DF",X"ED",X"88",
		X"10",X"86",X"01",X"A7",X"88",X"14",X"BD",X"27",X"00",X"0A",X"4F",X"26",X"9D",X"32",X"64",X"39",
		X"34",X"04",X"A6",X"63",X"3D",X"34",X"04",X"A6",X"61",X"E6",X"65",X"3D",X"AB",X"E4",X"44",X"56",
		X"32",X"62",X"39",X"B6",X"BE",X"57",X"81",X"03",X"25",X"39",X"0F",X"4F",X"EC",X"47",X"83",X"00",
		X"40",X"25",X"04",X"0C",X"4F",X"20",X"F7",X"96",X"4F",X"BD",X"08",X"E4",X"A7",X"47",X"8E",X"41",
		X"67",X"E6",X"47",X"BD",X"37",X"40",X"86",X"40",X"8E",X"41",X"4E",X"7E",X"00",X"A8",X"B6",X"BE",
		X"57",X"81",X"03",X"25",X"0E",X"A6",X"47",X"8B",X"99",X"19",X"2B",X"07",X"A7",X"47",X"8E",X"41",
		X"6D",X"20",X"DE",X"7E",X"00",X"E4",X"76",X"A0",X"0C",X"50",X"0A",X"41",X"6D",X"A0",X"20",X"41",
		X"6D",X"50",X"0B",X"CC",X"43",X"75",X"ED",X"02",X"BD",X"1C",X"87",X"02",X"10",X"06",X"A6",X"7A",
		X"BE",X"57",X"86",X"06",X"BD",X"08",X"C1",X"10",X"AE",X"E4",X"10",X"8C",X"26",X"96",X"27",X"06",
		X"31",X"84",X"BD",X"38",X"46",X"39",X"C6",X"45",X"BD",X"07",X"EC",X"46",X"86",X"01",X"24",X"02",
		X"C6",X"60",X"BD",X"14",X"3A",X"BD",X"01",X"88",X"1F",X"12",X"BD",X"19",X"43",X"41",X"B3",X"10",
		X"AF",X"07",X"39",X"86",X"04",X"8E",X"41",X"BB",X"7E",X"00",X"A8",X"86",X"03",X"A7",X"49",X"AE",
		X"47",X"BD",X"27",X"03",X"FC",X"4F",X"49",X"ED",X"02",X"6A",X"49",X"27",X"08",X"86",X"03",X"8E",
		X"41",X"BF",X"7E",X"00",X"A8",X"DC",X"43",X"ED",X"84",X"9F",X"43",X"7E",X"00",X"E4",X"BD",X"01",
		X"57",X"86",X"FF",X"97",X"91",X"86",X"01",X"8E",X"41",X"ED",X"7E",X"00",X"A8",X"BD",X"13",X"BD",
		X"BD",X"70",X"28",X"C6",X"7F",X"D7",X"27",X"10",X"BE",X"5F",X"D9",X"31",X"A5",X"A6",X"A0",X"27",
		X"29",X"81",X"02",X"26",X"06",X"96",X"57",X"2A",X"2D",X"20",X"F2",X"81",X"01",X"26",X"06",X"AE",
		X"A1",X"0F",X"11",X"20",X"E8",X"8B",X"2E",X"CE",X"41",X"FD",X"34",X"40",X"FE",X"42",X"3D",X"F6",
		X"41",X"66",X"33",X"C5",X"33",X"C5",X"33",X"C5",X"6E",X"C4",X"86",X"01",X"8E",X"42",X"32",X"7E",
		X"00",X"A8",X"96",X"57",X"2B",X"F4",X"BD",X"13",X"BD",X"6E",X"9F",X"FF",X"FE",X"6E",X"CF",X"BD",
		X"07",X"EC",X"D6",X"B6",X"1D",X"58",X"49",X"ED",X"88",X"10",X"D6",X"B8",X"C4",X"3F",X"CB",X"E0",
		X"1D",X"ED",X"0E",X"39",X"34",X"76",X"97",X"4F",X"B6",X"BE",X"59",X"4C",X"81",X"14",X"22",X"33",
		X"BD",X"38",X"4C",X"42",X"C3",X"20",X"9F",X"42",X"95",X"24",X"24",X"27",X"26",X"B7",X"BE",X"59",
		X"EC",X"2A",X"ED",X"0A",X"EC",X"2C",X"ED",X"0C",X"8D",X"C5",X"DC",X"B7",X"F4",X"BE",X"6C",X"E7",
		X"49",X"84",X"1F",X"A7",X"44",X"B6",X"BE",X"6B",X"BD",X"08",X"C1",X"A7",X"4B",X"9F",X"41",X"0A",
		X"4F",X"26",X"C5",X"35",X"F6",X"7A",X"BE",X"59",X"BD",X"1C",X"71",X"34",X"10",X"BD",X"00",X"EC",
		X"35",X"10",X"EC",X"0A",X"83",X"00",X"40",X"ED",X"0A",X"A6",X"0C",X"80",X"02",X"A7",X"0C",X"CE",
		X"20",X"06",X"EF",X"02",X"CC",X"01",X"15",X"BD",X"14",X"3A",X"CC",X"06",X"C9",X"BD",X"06",X"FD",
		X"7E",X"27",X"03",X"AE",X"47",X"F6",X"BE",X"6A",X"10",X"9E",X"A3",X"10",X"AC",X"0A",X"24",X"01",
		X"50",X"1D",X"ED",X"0E",X"20",X"54",X"E6",X"49",X"AE",X"47",X"96",X"97",X"A1",X"0C",X"22",X"01",
		X"50",X"1D",X"E3",X"88",X"10",X"10",X"83",X"02",X"00",X"2D",X"03",X"CC",X"02",X"00",X"10",X"83",
		X"FE",X"00",X"2E",X"03",X"CC",X"FE",X"00",X"ED",X"88",X"10",X"43",X"53",X"58",X"49",X"58",X"49",
		X"1F",X"89",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"D6",X"B6",X"C4",X"1F",X"CB",X"F0",X"1D",
		X"E3",X"88",X"10",X"ED",X"88",X"10",X"DC",X"A3",X"A3",X"0A",X"C3",X"12",X"C0",X"10",X"83",X"25",
		X"80",X"22",X"A0",X"6A",X"4B",X"26",X"03",X"BD",X"43",X"32",X"86",X"03",X"8E",X"42",X"D6",X"7E",
		X"00",X"A8",X"34",X"10",X"DC",X"A3",X"A3",X"0A",X"A8",X"0E",X"2B",X"2F",X"31",X"84",X"BD",X"0D",
		X"48",X"17",X"4B",X"20",X"7F",X"17",X"B6",X"27",X"22",X"EC",X"2E",X"58",X"49",X"58",X"49",X"58",
		X"49",X"ED",X"0E",X"CC",X"06",X"E7",X"BD",X"06",X"FD",X"5F",X"96",X"97",X"A0",X"0C",X"47",X"56",
		X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",X"88",X"10",X"B6",X"BE",X"6B",X"BD",X"08",
		X"C1",X"A7",X"4B",X"35",X"90",X"04",X"08",X"43",X"7F",X"43",X"7F",X"02",X"14",X"02",X"46",X"00",
		X"0E",X"88",X"D8",X"F8",X"8E",X"08",X"00",X"D8",X"88",X"8C",X"C8",X"8C",X"88",X"EF",X"8F",X"F8",
		X"8E",X"88",X"C8",X"88",X"8E",X"8D",X"E8",X"00",X"80",X"E8",X"DD",X"D8",X"E8",X"80",X"00",X"06",
		X"04",X"43",X"E5",X"43",X"FD",X"02",X"FA",X"03",X"3B",X"06",X"04",X"44",X"15",X"44",X"2D",X"02",
		X"FA",X"03",X"3B",X"06",X"04",X"44",X"45",X"44",X"5D",X"02",X"FA",X"03",X"3B",X"06",X"04",X"44",
		X"75",X"44",X"8D",X"02",X"FA",X"03",X"3B",X"06",X"04",X"44",X"A5",X"44",X"BD",X"02",X"FA",X"03",
		X"3B",X"06",X"04",X"44",X"D5",X"44",X"ED",X"02",X"FA",X"03",X"3B",X"06",X"04",X"45",X"05",X"45",
		X"1D",X"02",X"FA",X"03",X"3B",X"00",X"03",X"31",X"03",X"33",X"11",X"11",X"33",X"33",X"00",X"00",
		X"33",X"33",X"01",X"01",X"33",X"30",X"13",X"11",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"31",X"11",X"33",X"33",X"10",X"10",X"33",X"33",X"00",X"00",X"33",X"33",X"11",X"11",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"11",X"11",X"33",X"33",X"10",X"10",
		X"33",X"33",X"00",X"00",X"33",X"30",X"13",X"11",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"31",X"11",X"33",X"33",X"11",X"11",X"33",X"33",X"00",X"00",X"33",X"33",X"01",X"01",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"11",X"11",X"33",X"33",X"11",X"11",
		X"33",X"33",X"00",X"00",X"33",X"30",X"03",X"01",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"31",X"11",X"33",X"33",X"11",X"11",X"33",X"33",X"10",X"10",X"33",X"33",X"00",X"00",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"01",X"01",X"33",X"33",X"11",X"11",
		X"33",X"33",X"10",X"10",X"33",X"30",X"03",X"01",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"30",X"10",X"33",X"33",X"11",X"11",X"33",X"33",X"11",X"11",X"33",X"33",X"00",X"00",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"00",X"00",X"33",X"33",X"11",X"11",
		X"33",X"33",X"11",X"11",X"33",X"30",X"03",X"01",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"30",X"10",X"33",X"33",X"01",X"01",X"33",X"33",X"11",X"11",X"33",X"33",X"10",X"10",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"00",X"00",X"33",X"33",X"01",X"01",
		X"33",X"33",X"11",X"11",X"33",X"30",X"13",X"11",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"30",X"10",X"33",X"33",X"00",X"00",X"33",X"33",X"11",X"11",X"33",X"33",X"11",X"11",
		X"33",X"00",X"30",X"13",X"30",X"00",X"03",X"31",X"03",X"33",X"10",X"10",X"33",X"33",X"00",X"00",
		X"33",X"33",X"11",X"11",X"33",X"30",X"13",X"11",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",
		X"00",X"03",X"31",X"11",X"33",X"33",X"00",X"00",X"33",X"33",X"01",X"01",X"33",X"33",X"11",X"11",
		X"33",X"00",X"30",X"13",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"49",X"8A",X"7E",X"49",X"1B",X"7E",X"45",X"63",X"7E",X"4D",X"12",X"7E",X"48",X"C0",X"7E",
		X"48",X"CB",X"7E",X"46",X"9F",X"7E",X"49",X"DB",X"46",X"EB",X"4C",X"89",X"45",X"9F",X"4D",X"2A",
		X"7E",X"4E",X"92",X"34",X"06",X"97",X"50",X"BD",X"01",X"70",X"20",X"25",X"45",X"9F",X"66",X"66",
		X"BD",X"07",X"EC",X"DC",X"B7",X"84",X"1F",X"AB",X"61",X"ED",X"0A",X"54",X"24",X"05",X"CC",X"20",
		X"39",X"ED",X"02",X"86",X"E0",X"A7",X"0C",X"86",X"10",X"A7",X"88",X"14",X"4F",X"5F",X"ED",X"88",
		X"10",X"ED",X"0E",X"ED",X"06",X"9F",X"41",X"AF",X"A1",X"0A",X"50",X"26",X"CA",X"35",X"86",X"96",
		X"B5",X"26",X"42",X"8D",X"48",X"BD",X"1C",X"71",X"CC",X"1F",X"FC",X"ED",X"02",X"EC",X"0A",X"83",
		X"00",X"40",X"ED",X"0A",X"BD",X"27",X"03",X"CC",X"06",X"97",X"7E",X"06",X"FD",X"EE",X"06",X"27",
		X"DE",X"EC",X"42",X"10",X"83",X"4C",X"BF",X"27",X"1C",X"96",X"B5",X"27",X"1B",X"CC",X"06",X"8D",
		X"BD",X"06",X"FD",X"34",X"10",X"BD",X"19",X"43",X"47",X"BA",X"31",X"84",X"35",X"10",X"AF",X"27",
		X"CC",X"4C",X"BF",X"ED",X"42",X"4F",X"35",X"86",X"8D",X"B9",X"7E",X"00",X"EC",X"31",X"84",X"34",
		X"52",X"0D",X"91",X"2B",X"2D",X"CE",X"BE",X"83",X"86",X"0A",X"10",X"AC",X"C1",X"27",X"06",X"4A",
		X"26",X"F8",X"BD",X"01",X"15",X"4F",X"5F",X"ED",X"5E",X"7A",X"BE",X"54",X"26",X"07",X"BD",X"19",
		X"43",X"46",X"3E",X"35",X"D2",X"F6",X"BE",X"54",X"C1",X"03",X"22",X"06",X"8E",X"46",X"24",X"BD",
		X"37",X"40",X"35",X"D2",X"E0",X"04",X"C0",X"09",X"D6",X"91",X"C5",X"74",X"27",X"08",X"86",X"04",
		X"8E",X"46",X"28",X"7E",X"00",X"A8",X"86",X"04",X"8E",X"46",X"3E",X"7E",X"00",X"A8",X"D6",X"91",
		X"C5",X"74",X"26",X"EA",X"CA",X"06",X"D7",X"91",X"9E",X"49",X"27",X"05",X"BD",X"01",X"CD",X"20",
		X"F7",X"C6",X"C0",X"8D",X"4A",X"86",X"01",X"8E",X"46",X"5D",X"7E",X"00",X"A8",X"8E",X"9C",X"47",
		X"10",X"AE",X"84",X"27",X"04",X"30",X"A4",X"20",X"F7",X"10",X"9E",X"41",X"10",X"AF",X"84",X"CC",
		X"00",X"00",X"DD",X"41",X"BD",X"13",X"BD",X"0C",X"DB",X"BD",X"34",X"40",X"BD",X"19",X"72",X"BD",
		X"13",X"BD",X"BD",X"5F",X"C4",X"6F",X"47",X"8E",X"9C",X"47",X"8D",X"2E",X"6C",X"47",X"8E",X"9C",
		X"41",X"8D",X"27",X"BD",X"10",X"45",X"96",X"91",X"84",X"FB",X"97",X"91",X"7E",X"00",X"E4",X"9E",
		X"3B",X"A6",X"05",X"81",X"02",X"27",X"0E",X"81",X"03",X"27",X"0A",X"81",X"04",X"27",X"06",X"81",
		X"05",X"27",X"02",X"E7",X"04",X"AE",X"84",X"26",X"E8",X"39",X"AE",X"84",X"27",X"2C",X"EC",X"0A",
		X"93",X"20",X"C3",X"0C",X"80",X"10",X"83",X"3E",X"80",X"24",X"EF",X"EC",X"02",X"10",X"83",X"1A",
		X"D2",X"27",X"E7",X"EC",X"0A",X"C3",X"80",X"00",X"ED",X"0A",X"6D",X"47",X"27",X"DC",X"EC",X"04",
		X"27",X"D8",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"20",X"D0",X"39",X"AE",X"47",X"30",X"02",X"8C",
		X"BE",X"97",X"25",X"03",X"8E",X"BE",X"83",X"AF",X"47",X"AE",X"84",X"27",X"77",X"EC",X"04",X"27",
		X"73",X"EC",X"08",X"10",X"83",X"45",X"9F",X"26",X"6B",X"EC",X"02",X"10",X"83",X"20",X"2F",X"22",
		X"2F",X"96",X"B6",X"81",X"08",X"23",X"51",X"BD",X"1A",X"FC",X"8B",X"04",X"81",X"E8",X"23",X"02",
		X"86",X"E8",X"C6",X"01",X"A1",X"0C",X"27",X"07",X"22",X"01",X"50",X"EB",X"0C",X"E7",X"0C",X"EE",
		X"02",X"33",X"4A",X"11",X"83",X"20",X"2F",X"23",X"03",X"CE",X"20",X"25",X"C6",X"E0",X"20",X"2D",
		X"96",X"B6",X"81",X"08",X"23",X"F3",X"BD",X"1A",X"FC",X"8B",X"0F",X"81",X"E8",X"23",X"02",X"86",
		X"E8",X"C6",X"01",X"A1",X"0C",X"27",X"07",X"22",X"01",X"50",X"EB",X"0C",X"E7",X"0C",X"EE",X"02",
		X"33",X"4A",X"11",X"83",X"20",X"43",X"23",X"03",X"CE",X"20",X"39",X"C6",X"20",X"EF",X"02",X"1D",
		X"E3",X"0A",X"ED",X"0A",X"86",X"02",X"8E",X"46",X"EB",X"7E",X"00",X"A8",X"CC",X"01",X"25",X"BD",
		X"14",X"3A",X"96",X"43",X"27",X"72",X"BD",X"01",X"70",X"20",X"C1",X"45",X"E5",X"00",X"00",X"10",
		X"AE",X"47",X"EC",X"24",X"10",X"26",X"00",X"74",X"EC",X"2A",X"93",X"A3",X"2B",X"0E",X"DC",X"20",
		X"C3",X"27",X"00",X"ED",X"0A",X"DC",X"9E",X"83",X"00",X"40",X"20",X"09",X"DC",X"20",X"ED",X"0A",
		X"DC",X"9E",X"C3",X"00",X"40",X"ED",X"0E",X"7E",X"48",X"1D",X"96",X"D2",X"48",X"48",X"81",X"0C",
		X"23",X"02",X"86",X"0C",X"10",X"8E",X"1F",X"E2",X"31",X"A6",X"0C",X"D2",X"0D",X"43",X"27",X"28",
		X"BD",X"01",X"88",X"EC",X"22",X"ED",X"02",X"EF",X"06",X"CC",X"45",X"E5",X"ED",X"08",X"CC",X"00",
		X"00",X"ED",X"88",X"12",X"EC",X"A4",X"20",X"1E",X"BD",X"5F",X"D0",X"26",X"09",X"10",X"BE",X"45",
		X"5A",X"BD",X"15",X"3A",X"26",X"55",X"96",X"43",X"27",X"4E",X"BD",X"01",X"70",X"20",X"CB",X"45",
		X"E5",X"00",X"00",X"CC",X"01",X"50",X"BD",X"14",X"3A",X"10",X"AE",X"47",X"BD",X"07",X"EC",X"D6",
		X"B6",X"57",X"57",X"57",X"1D",X"D3",X"9E",X"ED",X"0E",X"EC",X"2A",X"ED",X"0A",X"D6",X"B7",X"86",
		X"FF",X"ED",X"88",X"10",X"86",X"11",X"A7",X"88",X"14",X"EC",X"2C",X"2B",X"05",X"C3",X"18",X"00",
		X"20",X"03",X"83",X"20",X"00",X"ED",X"0C",X"9F",X"41",X"AF",X"47",X"86",X"64",X"8E",X"48",X"43",
		X"7E",X"00",X"A8",X"AE",X"47",X"BD",X"1C",X"71",X"7E",X"00",X"E4",X"BD",X"01",X"57",X"CC",X"02",
		X"20",X"BD",X"14",X"3A",X"0F",X"2B",X"86",X"76",X"97",X"91",X"86",X"01",X"8E",X"48",X"62",X"7E",
		X"00",X"A8",X"10",X"AE",X"47",X"EC",X"24",X"26",X"03",X"CC",X"50",X"B0",X"C0",X"15",X"80",X"08",
		X"1F",X"01",X"BD",X"70",X"28",X"86",X"0D",X"BD",X"70",X"55",X"CC",X"48",X"BB",X"BD",X"06",X"FD",
		X"86",X"18",X"A7",X"47",X"CC",X"08",X"00",X"ED",X"48",X"BD",X"07",X"EC",X"84",X"1F",X"8E",X"0F",
		X"E6",X"A6",X"86",X"97",X"26",X"86",X"02",X"8E",X"48",X"9D",X"7E",X"00",X"A8",X"0F",X"26",X"6A",
		X"47",X"10",X"27",X"17",X"2E",X"EC",X"48",X"10",X"83",X"01",X"60",X"22",X"03",X"CC",X"01",X"60",
		X"83",X"00",X"60",X"ED",X"48",X"8E",X"48",X"89",X"7E",X"00",X"A8",X"FF",X"01",X"30",X"0D",X"00",
		X"34",X"10",X"BD",X"0D",X"48",X"17",X"4B",X"20",X"7F",X"17",X"B6",X"27",X"35",X"D6",X"B6",X"C4",
		X"1F",X"CB",X"F0",X"DB",X"96",X"E0",X"04",X"1D",X"58",X"49",X"58",X"49",X"ED",X"0E",X"D6",X"B6",
		X"C1",X"78",X"23",X"0A",X"DC",X"9E",X"58",X"49",X"58",X"49",X"E3",X"0E",X"ED",X"0E",X"D6",X"B8",
		X"C4",X"1F",X"CB",X"F0",X"DB",X"97",X"E0",X"05",X"1D",X"58",X"49",X"58",X"49",X"ED",X"88",X"10",
		X"86",X"01",X"35",X"90",X"6A",X"4D",X"26",X"12",X"B6",X"BE",X"63",X"BD",X"08",X"C1",X"A7",X"4D",
		X"8D",X"AE",X"27",X"06",X"CC",X"06",X"D8",X"BD",X"06",X"FD",X"39",X"34",X"02",X"97",X"4F",X"BD",
		X"38",X"4C",X"4B",X"B7",X"1F",X"F2",X"49",X"5A",X"CC",X"33",X"27",X"2C",X"BD",X"07",X"EC",X"DC",
		X"20",X"83",X"25",X"80",X"DD",X"51",X"DC",X"B7",X"93",X"51",X"10",X"83",X"4B",X"00",X"24",X"03",
		X"C3",X"80",X"00",X"D3",X"51",X"ED",X"0A",X"96",X"B6",X"44",X"8B",X"2C",X"A7",X"0C",X"BD",X"27",
		X"00",X"7C",X"BE",X"58",X"0A",X"4F",X"26",X"C7",X"35",X"82",X"7A",X"BE",X"58",X"BD",X"1C",X"80",
		X"01",X"15",X"06",X"AB",X"39",X"34",X"10",X"B6",X"BE",X"54",X"27",X"1C",X"9E",X"77",X"30",X"02",
		X"8C",X"BE",X"97",X"25",X"03",X"8E",X"BE",X"83",X"EC",X"84",X"26",X"06",X"9C",X"77",X"26",X"EE",
		X"35",X"90",X"9F",X"77",X"ED",X"49",X"AF",X"4B",X"35",X"90",X"34",X"02",X"97",X"4F",X"7D",X"BE",
		X"54",X"26",X"03",X"7E",X"49",X"1F",X"BD",X"38",X"4C",X"4A",X"14",X"4D",X"2A",X"4C",X"5D",X"44",
		X"33",X"27",X"36",X"BD",X"07",X"EC",X"DC",X"B7",X"ED",X"0A",X"86",X"2E",X"A7",X"0C",X"FC",X"BE",
		X"61",X"ED",X"88",X"10",X"B6",X"BE",X"63",X"BD",X"08",X"C1",X"A7",X"4D",X"B6",X"BE",X"60",X"BD",
		X"08",X"C1",X"1F",X"89",X"4F",X"C5",X"01",X"27",X"02",X"53",X"43",X"ED",X"0E",X"BD",X"27",X"00",
		X"8D",X"93",X"7C",X"BE",X"7C",X"0A",X"4F",X"26",X"B5",X"35",X"82",X"34",X"76",X"CE",X"9C",X"3B",
		X"20",X"2C",X"10",X"AE",X"42",X"10",X"8C",X"4A",X"14",X"25",X"23",X"26",X"13",X"AE",X"47",X"B6",
		X"BE",X"60",X"BD",X"08",X"C1",X"1F",X"89",X"4F",X"6D",X"0E",X"2A",X"02",X"43",X"53",X"ED",X"0E",
		X"10",X"8C",X"4B",X"3A",X"22",X"08",X"B6",X"BE",X"63",X"BD",X"08",X"C1",X"A7",X"4D",X"EE",X"C4",
		X"26",X"D0",X"35",X"F6",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"27",X"16",X"A6",X"29",
		X"81",X"9F",X"26",X"10",X"A6",X"0A",X"84",X"FC",X"97",X"4F",X"A6",X"2A",X"84",X"FC",X"91",X"4F",
		X"27",X"6C",X"20",X"0F",X"A6",X"88",X"14",X"84",X"FE",X"A7",X"88",X"14",X"BD",X"49",X"65",X"10",
		X"27",X"01",X"3B",X"BD",X"1A",X"FC",X"80",X"32",X"A0",X"0C",X"22",X"0F",X"81",X"EC",X"2D",X"04",
		X"4F",X"5F",X"20",X"0A",X"FC",X"BE",X"61",X"43",X"53",X"20",X"03",X"FC",X"BE",X"61",X"ED",X"88",
		X"10",X"EC",X"02",X"10",X"83",X"20",X"10",X"27",X"1D",X"A6",X"05",X"27",X"19",X"BD",X"49",X"04",
		X"8D",X"1C",X"86",X"03",X"8E",X"4A",X"7A",X"7E",X"00",X"A8",X"AE",X"47",X"8D",X"10",X"86",X"03",
		X"8E",X"4A",X"14",X"7E",X"00",X"A8",X"86",X"06",X"8E",X"4A",X"14",X"7E",X"00",X"A8",X"EE",X"02",
		X"33",X"4A",X"11",X"83",X"4D",X"48",X"23",X"03",X"CE",X"4D",X"2A",X"EF",X"02",X"39",X"4F",X"5F",
		X"6C",X"88",X"14",X"ED",X"0E",X"ED",X"88",X"10",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",
		X"10",X"27",X"FF",X"80",X"A6",X"29",X"81",X"9F",X"10",X"26",X"FF",X"78",X"EC",X"2A",X"C4",X"E0",
		X"DD",X"51",X"EC",X"0A",X"C4",X"E0",X"10",X"93",X"51",X"27",X"0D",X"2D",X"04",X"C6",X"E0",X"20",
		X"02",X"C6",X"20",X"1D",X"E3",X"0A",X"ED",X"0A",X"A6",X"2C",X"80",X"0C",X"A1",X"0C",X"27",X"16",
		X"FC",X"BE",X"61",X"24",X"02",X"43",X"53",X"E3",X"0C",X"ED",X"0C",X"BD",X"49",X"04",X"86",X"01",
		X"8E",X"4A",X"A8",X"7E",X"00",X"A8",X"EC",X"0A",X"C3",X"00",X"40",X"A3",X"2A",X"10",X"83",X"00",
		X"80",X"22",X"E8",X"CC",X"4C",X"39",X"ED",X"08",X"FC",X"BE",X"61",X"53",X"43",X"ED",X"88",X"10",
		X"ED",X"A8",X"10",X"CC",X"06",X"BF",X"BD",X"06",X"FD",X"CC",X"45",X"BD",X"ED",X"28",X"DE",X"3F",
		X"AE",X"47",X"A6",X"0C",X"81",X"34",X"23",X"12",X"A6",X"05",X"27",X"06",X"BD",X"49",X"04",X"BD",
		X"4A",X"8E",X"86",X"03",X"8E",X"4B",X"1E",X"7E",X"00",X"A8",X"CC",X"06",X"C4",X"BD",X"06",X"FD",
		X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"26",X"0C",X"BD",X"1C",X"71",X"7A",X"BE",X"7C",
		X"7C",X"BE",X"55",X"7E",X"00",X"E4",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"A8",X"10",X"A6",X"2C",
		X"A1",X"0C",X"23",X"0F",X"6A",X"2C",X"86",X"12",X"BD",X"06",X"EC",X"86",X"01",X"8E",X"4B",X"40",
		X"7E",X"00",X"A8",X"30",X"A4",X"EC",X"24",X"8B",X"01",X"DD",X"D0",X"BD",X"45",X"A3",X"7A",X"BE",
		X"7C",X"26",X"17",X"B6",X"BE",X"55",X"26",X"12",X"96",X"91",X"85",X"02",X"26",X"0C",X"CC",X"08",
		X"FF",X"FD",X"BD",X"D1",X"8E",X"4C",X"85",X"BD",X"37",X"40",X"7C",X"BE",X"58",X"AE",X"47",X"6F",
		X"88",X"14",X"CC",X"1F",X"F2",X"ED",X"02",X"CC",X"CC",X"33",X"ED",X"88",X"12",X"CC",X"49",X"5A",
		X"ED",X"08",X"B6",X"BE",X"69",X"A7",X"49",X"AE",X"47",X"F6",X"BE",X"68",X"10",X"9E",X"A3",X"10",
		X"AC",X"0A",X"2C",X"01",X"50",X"1D",X"ED",X"0E",X"DC",X"A3",X"A3",X"0A",X"C3",X"01",X"7C",X"10",
		X"83",X"07",X"00",X"23",X"21",X"96",X"97",X"A0",X"0C",X"23",X"0B",X"81",X"08",X"22",X"0B",X"FC",
		X"BE",X"66",X"43",X"53",X"20",X"0B",X"81",X"F8",X"2E",X"04",X"4F",X"5F",X"20",X"03",X"FC",X"BE",
		X"66",X"ED",X"88",X"10",X"20",X"12",X"96",X"97",X"A1",X"0C",X"FC",X"BE",X"66",X"24",X"02",X"43",
		X"53",X"ED",X"88",X"10",X"EC",X"04",X"27",X"29",X"F6",X"BE",X"65",X"96",X"B6",X"2B",X"01",X"50",
		X"EB",X"0C",X"C1",X"2C",X"24",X"02",X"C6",X"F0",X"E7",X"0C",X"6A",X"49",X"26",X"13",X"B6",X"BE",
		X"69",X"BD",X"08",X"C1",X"A7",X"49",X"BD",X"48",X"C0",X"27",X"06",X"CC",X"06",X"DD",X"BD",X"06",
		X"FD",X"86",X"03",X"8E",X"4B",X"B7",X"7E",X"00",X"A8",X"EE",X"06",X"EC",X"D8",X"0B",X"27",X"1D",
		X"EE",X"06",X"34",X"10",X"BD",X"19",X"43",X"4C",X"89",X"EE",X"49",X"EF",X"07",X"CC",X"06",X"9C",
		X"BD",X"06",X"FD",X"CC",X"00",X"00",X"ED",X"C8",X"10",X"AF",X"46",X"35",X"10",X"7A",X"BE",X"7C",
		X"26",X"1B",X"B6",X"BE",X"55",X"26",X"16",X"96",X"91",X"85",X"02",X"26",X"10",X"CC",X"08",X"FF",
		X"FD",X"BD",X"D1",X"34",X"10",X"8E",X"4C",X"85",X"BD",X"37",X"40",X"35",X"10",X"BD",X"1C",X"80",
		X"01",X"15",X"06",X"BA",X"39",X"20",X"44",X"80",X"0C",X"AE",X"47",X"CC",X"00",X"08",X"E3",X"88",
		X"10",X"10",X"83",X"03",X"00",X"24",X"03",X"ED",X"88",X"10",X"BD",X"1A",X"FC",X"A1",X"0C",X"22",
		X"16",X"EC",X"88",X"10",X"10",X"83",X"00",X"E0",X"23",X"39",X"EC",X"04",X"C3",X"01",X"07",X"DD",
		X"D0",X"BD",X"45",X"A3",X"7E",X"00",X"E4",X"86",X"04",X"8E",X"4C",X"89",X"7E",X"00",X"A8",X"AE",
		X"47",X"CC",X"00",X"00",X"ED",X"88",X"10",X"96",X"9C",X"8B",X"0A",X"A7",X"0C",X"DC",X"A3",X"C3",
		X"00",X"80",X"ED",X"0A",X"BD",X"1A",X"FC",X"A1",X"0C",X"25",X"0F",X"86",X"01",X"8E",X"4C",X"BF",
		X"7E",X"00",X"A8",X"34",X"10",X"8E",X"47",X"7C",X"20",X"07",X"34",X"10",X"0A",X"D2",X"8E",X"47",
		X"E8",X"86",X"00",X"BD",X"01",X"30",X"31",X"84",X"35",X"10",X"AF",X"27",X"CC",X"00",X"00",X"ED",
		X"06",X"ED",X"88",X"10",X"CC",X"45",X"9F",X"ED",X"08",X"CC",X"06",X"92",X"BD",X"06",X"FD",X"7E",
		X"00",X"E4",X"8E",X"BE",X"83",X"10",X"AE",X"81",X"27",X"08",X"EC",X"28",X"10",X"83",X"45",X"9F",
		X"27",X"07",X"8C",X"BE",X"97",X"26",X"EE",X"86",X"01",X"39",X"05",X"08",X"4D",X"52",X"4D",X"7A",
		X"02",X"6E",X"01",X"FA",X"05",X"08",X"4D",X"A2",X"4D",X"CA",X"02",X"6E",X"01",X"FA",X"05",X"08",
		X"4D",X"F2",X"4E",X"1A",X"02",X"6E",X"01",X"FA",X"05",X"08",X"4E",X"42",X"4E",X"6A",X"02",X"6E",
		X"01",X"FA",X"00",X"03",X"30",X"30",X"23",X"00",X"03",X"30",X"23",X"44",X"03",X"03",X"33",X"30",
		X"00",X"00",X"33",X"44",X"30",X"30",X"23",X"30",X"30",X"30",X"20",X"43",X"03",X"03",X"33",X"30",
		X"03",X"00",X"00",X"00",X"30",X"30",X"20",X"00",X"00",X"30",X"00",X"00",X"03",X"03",X"02",X"00",
		X"00",X"03",X"02",X"34",X"00",X"00",X"33",X"03",X"30",X"00",X"33",X"44",X"33",X"33",X"32",X"03",
		X"03",X"03",X"32",X"44",X"00",X"00",X"33",X"03",X"00",X"00",X"00",X"30",X"33",X"33",X"32",X"00",
		X"30",X"03",X"00",X"03",X"30",X"20",X"33",X"00",X"03",X"30",X"32",X"44",X"33",X"33",X"32",X"30",
		X"00",X"00",X"33",X"44",X"00",X"00",X"33",X"30",X"30",X"30",X"30",X"42",X"33",X"33",X"32",X"30",
		X"03",X"00",X"00",X"00",X"30",X"30",X"30",X"00",X"00",X"30",X"00",X"00",X"03",X"02",X"03",X"00",
		X"00",X"03",X"03",X"34",X"03",X"03",X"33",X"03",X"30",X"00",X"23",X"44",X"30",X"30",X"23",X"03",
		X"03",X"03",X"33",X"44",X"03",X"03",X"33",X"03",X"00",X"00",X"00",X"20",X"33",X"33",X"23",X"00",
		X"30",X"03",X"00",X"03",X"23",X"33",X"33",X"00",X"03",X"30",X"33",X"33",X"30",X"30",X"23",X"30",
		X"00",X"00",X"23",X"33",X"03",X"03",X"33",X"30",X"30",X"30",X"30",X"33",X"30",X"30",X"23",X"30",
		X"03",X"00",X"00",X"00",X"20",X"30",X"30",X"00",X"00",X"30",X"00",X"00",X"02",X"03",X"03",X"00",
		X"00",X"03",X"03",X"33",X"33",X"33",X"32",X"03",X"30",X"00",X"32",X"33",X"00",X"00",X"33",X"03",
		X"03",X"03",X"33",X"33",X"33",X"33",X"32",X"03",X"00",X"00",X"00",X"30",X"02",X"03",X"33",X"00",
		X"30",X"03",X"00",X"02",X"33",X"33",X"32",X"00",X"03",X"30",X"33",X"33",X"00",X"00",X"33",X"30",
		X"00",X"00",X"32",X"33",X"33",X"33",X"32",X"30",X"30",X"30",X"30",X"33",X"00",X"00",X"33",X"30",
		X"03",X"00",X"00",X"00",X"30",X"20",X"30",X"00",X"00",X"30",X"00",X"00",X"03",X"03",X"03",X"00",
		X"00",X"03",X"03",X"23",X"30",X"30",X"23",X"03",X"30",X"00",X"33",X"33",X"03",X"03",X"33",X"03",
		X"03",X"03",X"23",X"33",X"30",X"30",X"23",X"03",X"00",X"00",X"00",X"30",X"03",X"02",X"33",X"00",
		X"30",X"03",X"CC",X"04",X"C0",X"8E",X"A0",X"00",X"34",X"16",X"BD",X"38",X"4C",X"4E",X"F2",X"4D",
		X"2A",X"4C",X"40",X"44",X"33",X"1F",X"12",X"9F",X"41",X"BD",X"01",X"70",X"20",X"25",X"45",X"BD",
		X"66",X"66",X"AF",X"49",X"9F",X"41",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"0E",X"ED",X"2E",X"EC",
		X"62",X"ED",X"0A",X"ED",X"2A",X"C3",X"18",X"00",X"ED",X"62",X"CC",X"E0",X"00",X"ED",X"0C",X"A6",
		X"61",X"ED",X"2C",X"80",X"28",X"A7",X"61",X"CC",X"02",X"00",X"ED",X"A8",X"10",X"ED",X"4B",X"86",
		X"01",X"A7",X"88",X"14",X"A7",X"A8",X"14",X"6A",X"E4",X"26",X"AF",X"86",X"0A",X"B7",X"BE",X"7C",
		X"35",X"96",X"AE",X"47",X"A6",X"0C",X"81",X"D0",X"24",X"08",X"86",X"01",X"8E",X"4E",X"F2",X"7E",
		X"00",X"A8",X"AE",X"47",X"CC",X"D4",X"00",X"ED",X"0C",X"CC",X"FF",X"80",X"ED",X"88",X"10",X"AE",
		X"49",X"ED",X"88",X"10",X"86",X"3C",X"8E",X"4F",X"14",X"7E",X"00",X"A8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"51",X"5D",X"7E",X"4F",X"51",X"7E",X"51",X"14",X"5A",X"78",X"57",X"21",X"58",X"E8",X"54",
		X"01",X"34",X"06",X"E6",X"E4",X"27",X"70",X"C1",X"02",X"23",X"0A",X"BD",X"07",X"EC",X"C6",X"02",
		X"44",X"24",X"02",X"CB",X"01",X"E7",X"61",X"DC",X"B7",X"47",X"47",X"D3",X"A3",X"8B",X"80",X"DD",
		X"51",X"B6",X"BE",X"72",X"34",X"02",X"44",X"44",X"40",X"AB",X"E0",X"BD",X"08",X"C1",X"85",X"01",
		X"27",X"01",X"40",X"97",X"50",X"96",X"B8",X"44",X"97",X"4F",X"BD",X"38",X"4C",X"50",X"64",X"54",
		X"01",X"50",X"59",X"22",X"22",X"27",X"30",X"BD",X"07",X"EC",X"DC",X"B7",X"84",X"03",X"D3",X"51",
		X"ED",X"0A",X"BD",X"1A",X"FC",X"90",X"4F",X"A7",X"0C",X"96",X"4F",X"8B",X"04",X"97",X"4F",X"A7",
		X"49",X"D6",X"50",X"1D",X"ED",X"0E",X"BD",X"4F",X"C9",X"BD",X"27",X"00",X"7C",X"BE",X"5A",X"6A",
		X"E4",X"6A",X"61",X"26",X"C5",X"20",X"8C",X"35",X"86",X"10",X"8E",X"54",X"01",X"A6",X"0E",X"2A",
		X"03",X"31",X"A8",X"32",X"EC",X"88",X"10",X"58",X"49",X"8B",X"02",X"2A",X"01",X"4F",X"81",X"04",
		X"23",X"02",X"86",X"04",X"C6",X"0A",X"3D",X"31",X"A5",X"10",X"AF",X"02",X"39",X"34",X"10",X"DC",
		X"A3",X"A3",X"0A",X"A8",X"0E",X"2B",X"5B",X"96",X"97",X"A0",X"0C",X"A8",X"88",X"10",X"2B",X"52",
		X"B6",X"BE",X"70",X"BD",X"08",X"C1",X"A7",X"4D",X"96",X"75",X"81",X"0F",X"22",X"44",X"31",X"84",
		X"BD",X"0D",X"48",X"17",X"7F",X"17",X"AA",X"17",X"B6",X"27",X"37",X"D6",X"B6",X"C4",X"1F",X"CB",
		X"F0",X"DB",X"96",X"E0",X"04",X"1D",X"58",X"49",X"58",X"49",X"ED",X"0E",X"EC",X"2E",X"58",X"49",
		X"58",X"49",X"E3",X"0E",X"ED",X"0E",X"D6",X"B8",X"C4",X"1F",X"CB",X"F0",X"DB",X"97",X"E0",X"05",
		X"1D",X"58",X"49",X"58",X"49",X"D3",X"A1",X"47",X"56",X"ED",X"88",X"10",X"CC",X"50",X"54",X"BD",
		X"06",X"FD",X"35",X"90",X"C0",X"03",X"08",X"02",X"00",X"7A",X"BE",X"5A",X"BD",X"1C",X"80",X"01",
		X"20",X"06",X"B0",X"39",X"AE",X"47",X"EC",X"02",X"10",X"83",X"20",X"10",X"26",X"08",X"86",X"06",
		X"8E",X"50",X"64",X"7E",X"00",X"A8",X"AE",X"47",X"A6",X"05",X"26",X"1F",X"BD",X"1A",X"FC",X"5F",
		X"A0",X"0C",X"A0",X"49",X"81",X"F6",X"2E",X"02",X"C6",X"FF",X"81",X"0A",X"2D",X"02",X"C6",X"01",
		X"E7",X"88",X"10",X"86",X"0A",X"8E",X"50",X"76",X"7E",X"00",X"A8",X"86",X"0F",X"BD",X"08",X"C1",
		X"8E",X"50",X"A6",X"7E",X"00",X"A8",X"AE",X"47",X"96",X"B6",X"84",X"1F",X"80",X"0F",X"A7",X"4A",
		X"96",X"B8",X"84",X"0F",X"8B",X"02",X"A7",X"4C",X"B6",X"BE",X"70",X"A7",X"4D",X"B6",X"BE",X"71",
		X"BD",X"08",X"C1",X"A7",X"4B",X"DC",X"A3",X"10",X"A3",X"0A",X"34",X"01",X"B6",X"BE",X"72",X"BD",
		X"08",X"C1",X"1F",X"89",X"35",X"01",X"24",X"01",X"50",X"1D",X"ED",X"0E",X"AE",X"47",X"E6",X"4B",
		X"96",X"97",X"AB",X"4A",X"A1",X"0C",X"22",X"01",X"50",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",
		X"43",X"53",X"47",X"56",X"47",X"56",X"47",X"56",X"E3",X"88",X"10",X"ED",X"88",X"10",X"6A",X"4D",
		X"26",X"03",X"BD",X"4F",X"ED",X"6A",X"4C",X"27",X"9D",X"BD",X"4F",X"C9",X"86",X"04",X"8E",X"50",
		X"DC",X"7E",X"00",X"A8",X"BD",X"19",X"43",X"51",X"1A",X"39",X"96",X"ED",X"26",X"3C",X"0C",X"ED",
		X"86",X"03",X"A7",X"47",X"86",X"08",X"8E",X"51",X"2C",X"7E",X"00",X"A8",X"96",X"57",X"81",X"51",
		X"27",X"0A",X"81",X"E2",X"27",X"EE",X"6A",X"47",X"26",X"EA",X"20",X"1C",X"86",X"03",X"A7",X"47",
		X"86",X"08",X"8E",X"51",X"48",X"7E",X"00",X"A8",X"96",X"57",X"81",X"A3",X"10",X"27",X"E6",X"F9",
		X"81",X"51",X"27",X"EC",X"6A",X"47",X"26",X"E8",X"0F",X"ED",X"7E",X"00",X"E4",X"34",X"02",X"8E",
		X"51",X"6D",X"86",X"00",X"BD",X"01",X"30",X"6A",X"E4",X"26",X"F4",X"35",X"82",X"BD",X"01",X"70",
		X"57",X"21",X"53",X"BB",X"AC",X"CA",X"BD",X"07",X"EC",X"C6",X"50",X"3D",X"8B",X"80",X"ED",X"0A",
		X"8B",X"AC",X"ED",X"0C",X"86",X"01",X"A7",X"88",X"14",X"AF",X"C9",X"00",X"07",X"9F",X"41",X"BD",
		X"53",X"39",X"D6",X"B6",X"C4",X"0F",X"CB",X"08",X"E7",X"49",X"BD",X"52",X"24",X"AE",X"47",X"96",
		X"91",X"85",X"20",X"26",X"11",X"BD",X"53",X"F5",X"23",X"0C",X"6A",X"49",X"2B",X"E1",X"86",X"0A",
		X"8E",X"51",X"9D",X"7E",X"00",X"A8",X"6F",X"4A",X"A6",X"4A",X"27",X"02",X"6A",X"4A",X"AE",X"47",
		X"A6",X"0C",X"90",X"97",X"97",X"4F",X"2B",X"23",X"81",X"09",X"22",X"06",X"10",X"8E",X"52",X"64",
		X"8D",X"61",X"81",X"0C",X"24",X"24",X"F6",X"BE",X"74",X"4F",X"0D",X"4F",X"2A",X"02",X"43",X"53",
		X"0D",X"E9",X"26",X"02",X"58",X"49",X"ED",X"88",X"10",X"20",X"1A",X"40",X"81",X"0C",X"22",X"06",
		X"10",X"8E",X"52",X"7F",X"8D",X"3D",X"81",X"0F",X"23",X"DC",X"6A",X"49",X"2B",X"02",X"20",X"0D",
		X"BD",X"53",X"39",X"8D",X"1F",X"96",X"B6",X"84",X"7F",X"8B",X"1E",X"A7",X"49",X"EC",X"04",X"26",
		X"08",X"86",X"01",X"8E",X"51",X"9D",X"7E",X"00",X"A8",X"BD",X"52",X"E5",X"86",X"01",X"8E",X"51",
		X"B8",X"7E",X"00",X"A8",X"D6",X"B8",X"1D",X"2A",X"03",X"83",X"00",X"A0",X"C3",X"00",X"50",X"ED",
		X"88",X"10",X"39",X"DE",X"69",X"A6",X"49",X"DE",X"3F",X"4A",X"27",X"20",X"81",X"02",X"22",X"12",
		X"4A",X"97",X"4F",X"BD",X"07",X"EC",X"81",X"E0",X"24",X"13",X"81",X"80",X"23",X"04",X"96",X"4F",
		X"27",X"0B",X"6D",X"4A",X"26",X"06",X"EC",X"04",X"27",X"02",X"6E",X"A4",X"39",X"B6",X"BE",X"73",
		X"43",X"A7",X"4A",X"39",X"BD",X"53",X"0C",X"EC",X"0A",X"93",X"A3",X"2B",X"09",X"BD",X"53",X"2D",
		X"10",X"8E",X"FF",X"A0",X"20",X"2E",X"BD",X"53",X"33",X"10",X"8E",X"00",X"60",X"20",X"25",X"BD",
		X"53",X"0C",X"EC",X"0A",X"93",X"A3",X"2B",X"09",X"BD",X"53",X"33",X"10",X"8E",X"FF",X"80",X"20",
		X"07",X"BD",X"53",X"2D",X"10",X"8E",X"00",X"80",X"96",X"B6",X"84",X"07",X"8B",X"12",X"97",X"51",
		X"EC",X"0C",X"20",X"0C",X"96",X"B6",X"8A",X"F8",X"80",X"EE",X"97",X"51",X"EC",X"0C",X"8B",X"04",
		X"DD",X"4F",X"EC",X"0A",X"C3",X"00",X"40",X"BD",X"38",X"4C",X"53",X"49",X"58",X"E8",X"53",X"AD",
		X"40",X"00",X"27",X"14",X"ED",X"0A",X"DC",X"4F",X"ED",X"0C",X"10",X"AF",X"0E",X"86",X"01",X"A7",
		X"88",X"14",X"9F",X"41",X"96",X"51",X"A7",X"49",X"B6",X"BE",X"73",X"43",X"DE",X"3F",X"A7",X"4A",
		X"AE",X"47",X"7E",X"52",X"0D",X"10",X"AE",X"02",X"A6",X"0E",X"2B",X"10",X"31",X"2A",X"10",X"8C",
		X"57",X"3F",X"23",X"04",X"10",X"8E",X"57",X"21",X"10",X"AF",X"02",X"39",X"31",X"36",X"10",X"8C",
		X"57",X"21",X"24",X"04",X"10",X"8E",X"57",X"3F",X"10",X"AF",X"02",X"39",X"A6",X"0C",X"91",X"97",
		X"22",X"0B",X"F6",X"BE",X"74",X"53",X"86",X"FF",X"83",X"00",X"10",X"20",X"06",X"F6",X"BE",X"74",
		X"CB",X"0A",X"4F",X"0D",X"E9",X"26",X"02",X"58",X"49",X"ED",X"88",X"10",X"39",X"CC",X"00",X"20",
		X"ED",X"0E",X"39",X"CC",X"FF",X"E0",X"ED",X"0E",X"39",X"D6",X"B8",X"57",X"57",X"57",X"57",X"2B",
		X"02",X"CB",X"14",X"C0",X"0A",X"1D",X"ED",X"0E",X"39",X"CC",X"06",X"DD",X"BD",X"06",X"FD",X"86",
		X"20",X"A7",X"4A",X"86",X"03",X"8E",X"53",X"5B",X"7E",X"00",X"A8",X"AE",X"47",X"BD",X"53",X"F5",
		X"22",X"23",X"6A",X"4A",X"27",X"1F",X"96",X"B6",X"84",X"07",X"C6",X"0A",X"3D",X"E3",X"02",X"10",
		X"83",X"59",X"2E",X"23",X"03",X"83",X"00",X"50",X"ED",X"02",X"E6",X"49",X"1D",X"E3",X"88",X"10",
		X"ED",X"88",X"10",X"20",X"CE",X"BD",X"01",X"A2",X"EC",X"04",X"27",X"06",X"10",X"AE",X"02",X"AD",
		X"B8",X"08",X"7E",X"00",X"E4",X"BD",X"14",X"3A",X"1F",X"20",X"BD",X"06",X"FD",X"34",X"10",X"BD",
		X"00",X"EC",X"35",X"10",X"BD",X"01",X"A2",X"BD",X"00",X"00",X"7E",X"01",X"88",X"CC",X"02",X"01",
		X"10",X"8E",X"06",X"97",X"8D",X"DF",X"CC",X"5A",X"78",X"20",X"0F",X"7A",X"BE",X"5C",X"CC",X"01",
		X"25",X"10",X"8E",X"06",X"97",X"8D",X"CE",X"CC",X"57",X"49",X"ED",X"02",X"1F",X"12",X"BD",X"19",
		X"43",X"53",X"D7",X"10",X"AF",X"07",X"39",X"86",X"03",X"A7",X"49",X"AE",X"47",X"BD",X"27",X"03",
		X"6A",X"49",X"27",X"08",X"86",X"05",X"8E",X"53",X"DB",X"7E",X"00",X"A8",X"DC",X"43",X"ED",X"84",
		X"9F",X"43",X"7E",X"00",X"E4",X"EC",X"0A",X"93",X"20",X"C3",X"09",X"60",X"10",X"83",X"38",X"40",
		X"39",X"05",X"07",X"54",X"65",X"54",X"88",X"04",X"5F",X"04",X"98",X"05",X"07",X"54",X"AB",X"54",
		X"CE",X"04",X"5F",X"04",X"98",X"05",X"07",X"54",X"F1",X"55",X"14",X"04",X"5F",X"04",X"98",X"05",
		X"07",X"55",X"37",X"55",X"5A",X"04",X"5F",X"04",X"98",X"05",X"07",X"55",X"7D",X"55",X"A0",X"04",
		X"5F",X"04",X"98",X"05",X"07",X"55",X"C3",X"55",X"E6",X"04",X"5F",X"04",X"98",X"05",X"07",X"56",
		X"09",X"56",X"2C",X"04",X"5F",X"04",X"98",X"05",X"07",X"56",X"4F",X"56",X"72",X"04",X"5F",X"04",
		X"98",X"05",X"07",X"56",X"95",X"56",X"B8",X"04",X"5F",X"04",X"98",X"05",X"07",X"56",X"DB",X"56",
		X"FE",X"04",X"5F",X"04",X"98",X"00",X"0A",X"06",X"66",X"00",X"0F",X"00",X"AA",X"A2",X"66",X"62",
		X"FF",X"88",X"FF",X"A0",X"AA",X"60",X"66",X"F0",X"8F",X"F0",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0A",
		X"AA",X"66",X"66",X"0F",X"F8",X"0F",X"AA",X"2A",X"66",X"26",X"FF",X"88",X"FF",X"00",X"A0",X"00",
		X"66",X"00",X"F0",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"0F",
		X"00",X"00",X"00",X"AA",X"66",X"FF",X"88",X"FF",X"00",X"00",X"A0",X"6A",X"F6",X"8F",X"F0",X"00",
		X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"0A",X"66",X"6F",X"F8",X"0F",X"00",X"00",X"AA",X"66",X"FF",
		X"88",X"FF",X"00",X"00",X"00",X"A0",X"66",X"F0",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"06",X"6F",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"00",X"00",
		X"00",X"F0",X"8F",X"F0",X"00",X"00",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"6F",X"F8",X"0F",
		X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"00",X"00",X"00",X"00",X"F6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"0F",X"66",X"0A",X"00",X"00",X"00",X"FF",
		X"88",X"FF",X"A2",X"AA",X"00",X"00",X"F0",X"8F",X"F6",X"AA",X"A0",X"00",X"00",X"00",X"00",X"61",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"0F",X"8F",X"6F",X"AA",X"0A",X"00",X"00",X"FF",X"88",X"FF",X"2A",X"AA",X"00",X"00",
		X"00",X"F0",X"66",X"A0",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"0F",X"06",
		X"66",X"00",X"0A",X"00",X"FF",X"88",X"FF",X"62",X"A2",X"A2",X"AA",X"F0",X"8F",X"F0",X"66",X"A0",
		X"AA",X"A0",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0F",X"F8",X"6F",X"66",X"0A",X"AA",X"0A",X"FF",X"88",
		X"FF",X"26",X"2A",X"2A",X"AA",X"00",X"F0",X"00",X"66",X"00",X"A0",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"0A",X"00",X"66",X"00",X"0F",
		X"00",X"AA",X"A2",X"66",X"62",X"FF",X"88",X"FF",X"A0",X"AA",X"66",X"66",X"F0",X"8F",X"F0",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"0A",X"AA",X"06",X"66",X"0F",X"F8",X"0F",X"AA",X"2A",X"66",X"26",X"FF",
		X"88",X"FF",X"00",X"A0",X"60",X"66",X"00",X"F0",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"66",X"0F",X"00",X"00",X"00",X"AA",X"66",X"FF",X"88",X"FF",X"00",X"00",X"A0",
		X"66",X"F6",X"8F",X"F0",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"0A",X"A6",X"6F",X"F8",X"0F",
		X"00",X"00",X"AA",X"66",X"FF",X"88",X"FF",X"00",X"00",X"00",X"60",X"66",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"88",X"FF",X"00",X"00",X"00",X"00",X"F6",X"8F",X"F0",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"F8",X"0F",X"00",X"00",X"00",X"00",X"FF",X"88",X"FF",X"00",X"00",X"00",X"00",
		X"60",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"0F",X"66",
		X"0A",X"00",X"00",X"00",X"FF",X"88",X"FF",X"A2",X"AA",X"00",X"00",X"F0",X"8F",X"F6",X"AA",X"A0",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"0F",X"F8",X"6F",X"AA",X"0A",X"00",X"00",X"FF",X"88",
		X"FF",X"2A",X"AA",X"00",X"00",X"00",X"F0",X"66",X"A0",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"66",X"00",X"0A",X"00",X"FF",X"88",X"FF",X"62",X"A2",X"A2",X"AA",
		X"F0",X"8F",X"F6",X"66",X"A0",X"AA",X"A0",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"0F",X"F8",X"0F",X"66",
		X"0A",X"AA",X"0A",X"FF",X"88",X"FF",X"26",X"2A",X"2A",X"AA",X"00",X"F0",X"60",X"66",X"00",X"A0",
		X"00",X"05",X"09",X"57",X"53",X"57",X"80",X"04",X"C4",X"05",X"12",X"05",X"09",X"57",X"AD",X"57",
		X"DA",X"04",X"C4",X"05",X"12",X"05",X"09",X"58",X"07",X"58",X"34",X"04",X"C4",X"05",X"12",X"05",
		X"09",X"58",X"61",X"58",X"8E",X"04",X"C4",X"05",X"12",X"05",X"09",X"58",X"BB",X"58",X"BB",X"04",
		X"C4",X"05",X"12",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"99",X"11",X"11",X"11",X"91",X"A9",X"AA",X"A0",X"A0",X"A0",X"90",X"10",X"10",X"11",
		X"91",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"19",
		X"11",X"01",X"01",X"09",X"0A",X"0A",X"0A",X"AA",X"9A",X"19",X"11",X"11",X"11",X"99",X"A9",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"11",X"11",X"11",X"11",X"01",X"00",X"00",X"00",X"00",X"90",X"9A",X"9A",X"90",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"01",X"91",X"91",X"91",X"91",X"01",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"01",X"00",X"00",X"00",X"00",X"10",X"19",X"19",X"19",X"19",X"10",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"09",X"A9",X"A9",X"09",X"00",X"00",X"00",X"00",X"10",
		X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"01",X"11",X"11",X"19",X"00",X"00",X"00",X"00",
		X"11",X"11",X"99",X"9A",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",X"09",
		X"01",X"01",X"00",X"00",X"00",X"00",X"A9",X"91",X"91",X"11",X"10",X"00",X"00",X"00",X"00",X"10",
		X"10",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"11",X"19",
		X"19",X"9A",X"00",X"00",X"00",X"00",X"10",X"10",X"90",X"A0",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"A9",X"99",X"11",X"11",X"00",X"00",X"00",X"00",X"91",X"11",X"11",X"10",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"99",X"0A",X"00",X"00",
		X"09",X"11",X"11",X"11",X"11",X"99",X"A0",X"A0",X"AA",X"99",X"11",X"11",X"10",X"10",X"00",X"00",
		X"00",X"00",X"90",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"09",X"00",X"00",X"00",X"00",X"01",X"01",
		X"11",X"11",X"99",X"AA",X"0A",X"0A",X"99",X"11",X"11",X"11",X"11",X"90",X"00",X"00",X"A0",X"99",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"11",X"11",X"19",
		X"11",X"11",X"01",X"00",X"11",X"11",X"99",X"9A",X"AA",X"9A",X"99",X"11",X"11",X"11",X"91",X"A9",
		X"AA",X"AA",X"AA",X"A9",X"91",X"11",X"10",X"11",X"91",X"91",X"A9",X"91",X"91",X"11",X"10",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"04",X"05",X"59",X"38",X"59",X"4C",X"05",X"44",
		X"1D",X"E9",X"04",X"05",X"59",X"60",X"59",X"74",X"05",X"44",X"1D",X"E9",X"04",X"05",X"59",X"88",
		X"59",X"9C",X"05",X"44",X"1D",X"E9",X"04",X"05",X"59",X"B0",X"59",X"C4",X"05",X"44",X"1D",X"E9",
		X"04",X"05",X"59",X"D8",X"59",X"EC",X"05",X"44",X"1D",X"E9",X"04",X"05",X"5A",X"00",X"5A",X"14",
		X"05",X"44",X"1D",X"E9",X"04",X"05",X"5A",X"28",X"5A",X"3C",X"05",X"44",X"1D",X"E9",X"04",X"05",
		X"5A",X"50",X"5A",X"64",X"05",X"44",X"1D",X"E9",X"00",X"02",X"02",X"20",X"02",X"00",X"40",X"44",
		X"04",X"02",X"20",X"20",X"40",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"24",X"24",X"00",X"20",X"02",X"02",X"44",X"42",X"20",X"00",X"00",X"00",X"20",X"00",
		X"02",X"20",X"04",X"02",X"00",X"02",X"20",X"40",X"24",X"00",X"00",X"02",X"40",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"02",X"44",X"22",X"00",X"20",X"00",
		X"04",X"40",X"02",X"00",X"20",X"00",X"00",X"00",X"00",X"02",X"24",X"02",X"00",X"20",X"02",X"04",
		X"40",X"20",X"00",X"20",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"02",X"20",X"40",X"24",X"02",X"00",X"22",X"40",X"02",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"02",X"00",X"20",X"02",X"00",X"40",X"44",X"02",X"00",X"20",X"22",X"20",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"24",X"04",X"00",X"20",X"02",X"02",
		X"42",X"20",X"00",X"00",X"20",X"00",X"20",X"00",X"00",X"20",X"02",X"00",X"00",X"20",X"44",X"00",
		X"44",X"00",X"00",X"00",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"02",X"04",X"20",X"04",X"00",X"00",X"40",X"04",X"40",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"20",X"02",X"02",X"02",X"24",X"44",X"40",X"02",X"00",X"20",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"04",X"24",X"20",X"20",X"42",
		X"40",X"02",X"20",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"04",X"20",X"00",X"00",X"00",X"04",
		X"24",X"00",X"20",X"20",X"42",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"20",X"20",X"40",X"02",X"00",X"02",X"02",X"44",X"42",X"00",X"00",X"00",X"20",X"20",X"00",
		X"00",X"20",X"04",X"02",X"00",X"20",X"44",X"40",X"42",X"20",X"00",X"02",X"20",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"02",X"04",X"44",X"24",X"02",X"00",X"40",
		X"02",X"20",X"02",X"00",X"20",X"00",X"00",X"00",X"05",X"08",X"5A",X"82",X"5A",X"82",X"02",X"6E",
		X"01",X"FA",X"00",X"02",X"22",X"22",X"22",X"22",X"02",X"00",X"22",X"22",X"22",X"24",X"24",X"22",
		X"22",X"22",X"22",X"22",X"44",X"44",X"44",X"44",X"22",X"22",X"22",X"22",X"22",X"42",X"42",X"22",
		X"22",X"22",X"00",X"20",X"22",X"22",X"22",X"22",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"5A",X"D7",X"5D",X"2E",X"5E",X"FF",X"34",X"02",X"BD",X"19",X"43",X"5A",X"E4",X"6A",X"E4",
		X"26",X"F7",X"35",X"82",X"BD",X"01",X"70",X"5D",X"2E",X"5C",X"3F",X"92",X"29",X"BD",X"07",X"EC",
		X"44",X"8B",X"40",X"ED",X"0A",X"8B",X"FC",X"ED",X"0C",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",
		X"10",X"AF",X"C9",X"00",X"07",X"9F",X"41",X"86",X"01",X"A7",X"C9",X"00",X"09",X"B6",X"BE",X"75",
		X"43",X"A7",X"C9",X"00",X"0A",X"BD",X"5B",X"E9",X"6D",X"49",X"26",X"57",X"96",X"B7",X"84",X"1F",
		X"8B",X"10",X"A7",X"49",X"EC",X"88",X"10",X"2A",X"0A",X"10",X"83",X"FF",X"80",X"22",X"0E",X"D6",
		X"B6",X"20",X"12",X"10",X"83",X"00",X"80",X"25",X"04",X"D6",X"B6",X"20",X"0C",X"D6",X"B6",X"A6",
		X"0C",X"81",X"6A",X"24",X"04",X"C4",X"3F",X"20",X"02",X"CA",X"C0",X"1D",X"E3",X"88",X"10",X"ED",
		X"88",X"10",X"EC",X"0E",X"2A",X"08",X"10",X"83",X"FF",X"D8",X"24",X"0C",X"20",X"06",X"10",X"83",
		X"00",X"28",X"23",X"04",X"47",X"56",X"ED",X"0E",X"D6",X"B8",X"57",X"57",X"57",X"57",X"1D",X"E3",
		X"0E",X"ED",X"0E",X"6D",X"4A",X"26",X"62",X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",X"80",X"24",
		X"58",X"DC",X"A3",X"A3",X"0A",X"2A",X"02",X"43",X"53",X"10",X"83",X"06",X"40",X"23",X"4A",X"86",
		X"18",X"BD",X"08",X"C1",X"97",X"4F",X"B6",X"BE",X"75",X"43",X"9B",X"4F",X"24",X"02",X"86",X"FF",
		X"A7",X"4A",X"B6",X"BE",X"82",X"81",X"06",X"24",X"30",X"31",X"84",X"BD",X"38",X"4C",X"5C",X"4F",
		X"5E",X"FF",X"5D",X"1E",X"90",X"00",X"27",X"21",X"10",X"AF",X"49",X"7C",X"BE",X"82",X"CC",X"5B",
		X"E1",X"BD",X"06",X"FD",X"EC",X"2A",X"10",X"93",X"A3",X"2A",X"06",X"EC",X"2E",X"2B",X"0A",X"20",
		X"04",X"EC",X"2E",X"2A",X"04",X"43",X"53",X"ED",X"2E",X"86",X"02",X"8E",X"5B",X"15",X"7E",X"00",
		X"A8",X"C0",X"01",X"40",X"19",X"01",X"01",X"16",X"00",X"AE",X"47",X"EC",X"0A",X"93",X"20",X"C3",
		X"06",X"40",X"10",X"83",X"32",X"00",X"24",X"36",X"FC",X"00",X"04",X"26",X"04",X"86",X"13",X"A7",
		X"4A",X"10",X"AE",X"02",X"EC",X"0E",X"2B",X"0E",X"31",X"36",X"10",X"8C",X"5D",X"2E",X"24",X"12",
		X"10",X"8E",X"5D",X"4C",X"20",X"0C",X"31",X"2A",X"10",X"8C",X"5D",X"4C",X"23",X"04",X"10",X"8E",
		X"5D",X"2E",X"10",X"AF",X"02",X"A6",X"4A",X"27",X"02",X"6A",X"4A",X"6A",X"49",X"39",X"86",X"13",
		X"A7",X"4A",X"86",X"10",X"8E",X"5C",X"3A",X"7E",X"00",X"A8",X"AE",X"47",X"7E",X"5B",X"1C",X"7A",
		X"BE",X"5D",X"CC",X"5D",X"56",X"ED",X"02",X"BD",X"1C",X"80",X"01",X"20",X"06",X"B5",X"39",X"10",
		X"AE",X"49",X"AE",X"47",X"EC",X"2A",X"93",X"A3",X"2A",X"07",X"EC",X"2A",X"C3",X"00",X"E0",X"20",
		X"05",X"EC",X"2A",X"83",X"00",X"60",X"ED",X"0A",X"EC",X"2C",X"8B",X"02",X"ED",X"0C",X"CC",X"00",
		X"00",X"ED",X"0E",X"ED",X"88",X"10",X"4C",X"A7",X"49",X"9F",X"41",X"AF",X"47",X"BD",X"5C",X"F7",
		X"6A",X"49",X"26",X"41",X"86",X"04",X"A7",X"49",X"8D",X"4A",X"23",X"0C",X"8D",X"59",X"22",X"08",
		X"CC",X"00",X"00",X"ED",X"88",X"10",X"20",X"16",X"DC",X"97",X"10",X"A3",X"0C",X"24",X"06",X"F6",
		X"BE",X"76",X"53",X"20",X"03",X"F6",X"BE",X"76",X"1D",X"58",X"49",X"ED",X"88",X"10",X"8D",X"24",
		X"23",X"1B",X"DC",X"A3",X"10",X"A3",X"0A",X"2A",X"06",X"F6",X"BE",X"76",X"53",X"20",X"03",X"F6",
		X"BE",X"76",X"1D",X"ED",X"0E",X"86",X"03",X"8E",X"5C",X"7D",X"7E",X"00",X"A8",X"CC",X"00",X"00",
		X"ED",X"0E",X"20",X"F1",X"DC",X"A3",X"C3",X"00",X"A0",X"A3",X"0A",X"2A",X"05",X"43",X"53",X"C3",
		X"00",X"01",X"10",X"83",X"01",X"20",X"39",X"DC",X"97",X"A3",X"0C",X"2A",X"05",X"43",X"53",X"C3",
		X"00",X"01",X"10",X"83",X"0A",X"00",X"39",X"AE",X"47",X"EC",X"0A",X"93",X"20",X"10",X"83",X"25",
		X"80",X"22",X"13",X"10",X"AE",X"02",X"31",X"2A",X"10",X"8C",X"5F",X"09",X"23",X"04",X"10",X"8E",
		X"5E",X"FF",X"10",X"AF",X"02",X"39",X"86",X"0C",X"8E",X"5C",X"7D",X"7E",X"00",X"A8",X"7A",X"BE",
		X"82",X"CC",X"5E",X"F5",X"ED",X"02",X"BD",X"1C",X"80",X"01",X"10",X"06",X"B5",X"39",X"05",X"09",
		X"5D",X"8D",X"5E",X"41",X"04",X"C4",X"05",X"12",X"05",X"09",X"5D",X"BA",X"5E",X"6E",X"04",X"C4",
		X"05",X"12",X"05",X"09",X"5D",X"E7",X"5E",X"9B",X"04",X"C4",X"05",X"12",X"05",X"09",X"5E",X"14",
		X"5E",X"C8",X"04",X"C4",X"05",X"12",X"05",X"09",X"5D",X"60",X"5D",X"60",X"04",X"C4",X"05",X"12",
		X"00",X"00",X"00",X"02",X"99",X"02",X"00",X"00",X"00",X"00",X"02",X"99",X"92",X"92",X"92",X"99",
		X"02",X"00",X"90",X"92",X"99",X"22",X"92",X"22",X"99",X"92",X"90",X"00",X"00",X"90",X"92",X"99",
		X"92",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",X"02",X"90",X"02",X"00",X"90",
		X"02",X"00",X"02",X"90",X"02",X"00",X"02",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"20",X"00",X"20",X"09",X"00",X"00",X"00",X"00",X"00",X"20",X"09",
		X"20",X"00",X"20",X"09",X"00",X"00",X"00",X"00",X"00",X"20",X"09",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",X"00",X"00",
		X"00",X"00",X"90",X"02",X"00",X"02",X"90",X"00",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",
		X"00",X"00",X"00",X"00",X"90",X"02",X"00",X"02",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"20",X"00",X"20",X"09",X"00",X"00",X"09",X"20",X"00",X"20",X"09",X"20",X"00",X"00",X"00",
		X"00",X"20",X"09",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"09",X"00",X"00",X"09",X"20",X"00",X"20",X"09",X"20",X"00",X"20",X"09",X"00",X"20",X"09",X"20",
		X"00",X"20",X"09",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",X"00",X"00",X"00",
		X"00",X"90",X"02",X"00",X"02",X"90",X"02",X"00",X"00",X"00",X"00",X"00",X"90",X"02",X"00",X"02",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"20",X"00",X"20",X"09",X"00",X"00",X"00",X"00",X"00",
		X"20",X"09",X"20",X"00",X"00",X"00",X"00",X"00",X"09",X"20",X"00",X"20",X"09",X"00",X"00",X"00",
		X"00",X"00",X"20",X"09",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",X"00",X"00",X"00",X"02",X"90",X"02",X"00",
		X"02",X"90",X"00",X"00",X"90",X"02",X"00",X"02",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"5F",X"4F",X"5F",X"4F",X"1D",X"73",X"1D",X"85",X"03",
		X"05",X"5F",X"13",X"5F",X"22",X"1D",X"73",X"1D",X"85",X"03",X"05",X"5F",X"31",X"5F",X"40",X"1D",
		X"73",X"1D",X"85",X"00",X"09",X"90",X"09",X"00",X"90",X"09",X"00",X"09",X"90",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"09",X"90",X"00",X"90",X"09",X"00",X"90",X"09",X"90",
		X"00",X"00",X"00",X"22",X"00",X"00",X"20",X"20",X"92",X"20",X"20",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"02",X"00",X"00",X"02",X"02",X"29",X"02",X"02",X"00",X"00",X"22",X"00",X"00",X"00",
		X"09",X"92",X"09",X"00",X"90",X"29",X"92",X"29",X"90",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"CF",X"04",X"E8",X"00",X"00",X"00",X"00",X"18",X"0C",X"05",X"E8",X"18",X"72",X"00",X"E8",
		X"61",X"0E",X"00",X"00",X"60",X"F4",X"00",X"00",X"17",X"E2",X"00",X"E8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F4",X"89",X"00",X"00",X"06",X"27",X"02",X"00",X"E9",X"4F",X"01",X"00",
		X"06",X"1E",X"02",X"00",X"06",X"30",X"02",X"00",X"7E",X"63",X"D5",X"7E",X"1E",X"35",X"7E",X"1E",
		X"CB",X"7E",X"68",X"E3",X"7E",X"1E",X"96",X"7E",X"60",X"35",X"7E",X"63",X"EA",X"7E",X"64",X"80",
		X"7E",X"68",X"8B",X"7E",X"67",X"1D",X"7E",X"60",X"5F",X"6B",X"C8",X"7E",X"63",X"96",X"7E",X"63",
		X"7C",X"7E",X"68",X"DF",X"7E",X"66",X"20",X"7E",X"60",X"E2",X"7E",X"6F",X"26",X"7E",X"8F",X"00",
		X"7E",X"6D",X"6D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"28",X"43",
		X"29",X"20",X"31",X"39",X"38",X"31",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",
		X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",
		X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",
		X"52",X"56",X"45",X"44",X"20",X"6C",X"08",X"6C",X"0A",X"34",X"10",X"8E",X"CC",X"22",X"BD",X"14",
		X"0B",X"BD",X"08",X"D1",X"35",X"10",X"AB",X"0B",X"25",X"02",X"A7",X"0B",X"7E",X"1D",X"F7",X"00",
		X"34",X"FF",X"35",X"00",X"34",X"00",X"3E",X"C8",X"0C",X"C8",X"0E",X"C8",X"04",X"C8",X"06",X"1A",
		X"FF",X"10",X"CE",X"BF",X"FF",X"86",X"9C",X"1F",X"8B",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"60",
		X"4F",X"4F",X"5F",X"ED",X"98",X"08",X"EC",X"81",X"ED",X"98",X"06",X"8C",X"60",X"57",X"26",X"F1",
		X"BD",X"13",X"BD",X"86",X"3F",X"B7",X"C8",X"0E",X"8E",X"9C",X"00",X"6F",X"80",X"C6",X"39",X"F7",
		X"CB",X"FF",X"8C",X"C0",X"00",X"26",X"F4",X"BD",X"E0",X"03",X"8E",X"CD",X"00",X"BD",X"14",X"1C",
		X"1F",X"98",X"81",X"20",X"22",X"06",X"84",X"0F",X"81",X"09",X"23",X"01",X"5F",X"D7",X"36",X"CC",
		X"A5",X"5A",X"DD",X"B7",X"CC",X"FF",X"70",X"DD",X"7D",X"0F",X"7F",X"C6",X"FF",X"DD",X"55",X"86",
		X"55",X"97",X"DE",X"BD",X"15",X"15",X"BD",X"08",X"0B",X"8D",X"17",X"BD",X"70",X"28",X"8E",X"D0",
		X"00",X"86",X"01",X"BD",X"01",X"30",X"86",X"0C",X"B7",X"C8",X"0E",X"03",X"91",X"1C",X"00",X"7E",
		X"00",X"0C",X"BD",X"08",X"3A",X"BD",X"0E",X"EC",X"BD",X"08",X"FB",X"BD",X"08",X"4A",X"BD",X"19",
		X"72",X"7E",X"0A",X"9C",X"96",X"91",X"2A",X"32",X"B6",X"CC",X"15",X"84",X"0F",X"27",X"04",X"86",
		X"01",X"97",X"36",X"96",X"36",X"27",X"23",X"8E",X"06",X"70",X"86",X"01",X"20",X"1A",X"96",X"91",
		X"2A",X"18",X"B6",X"CC",X"15",X"84",X"0F",X"27",X"04",X"86",X"02",X"97",X"36",X"96",X"36",X"81",
		X"02",X"25",X"07",X"8E",X"06",X"75",X"86",X"02",X"8D",X"03",X"7E",X"00",X"E4",X"CE",X"9C",X"B1",
		X"97",X"68",X"1F",X"10",X"BD",X"06",X"FD",X"0F",X"37",X"0F",X"38",X"BD",X"01",X"57",X"BD",X"13",
		X"BD",X"10",X"8E",X"00",X"00",X"4F",X"AB",X"A4",X"31",X"A8",X"10",X"10",X"8C",X"90",X"00",X"25",
		X"F5",X"A7",X"C8",X"4E",X"86",X"7F",X"97",X"91",X"86",X"01",X"97",X"67",X"97",X"25",X"8E",X"BD",
		X"D6",X"6F",X"80",X"8C",X"BE",X"54",X"26",X"F9",X"86",X"0A",X"B7",X"BD",X"E2",X"96",X"68",X"C6",
		X"08",X"BD",X"F4",X"80",X"34",X"10",X"8E",X"CC",X"04",X"BD",X"14",X"1C",X"35",X"10",X"5D",X"27",
		X"09",X"48",X"CE",X"CC",X"04",X"91",X"36",X"23",X"04",X"44",X"CE",X"CC",X"02",X"1F",X"89",X"96",
		X"36",X"8B",X"99",X"19",X"5A",X"26",X"FA",X"97",X"36",X"8E",X"CD",X"00",X"BD",X"14",X"24",X"1F",
		X"31",X"BD",X"14",X"0B",X"BD",X"08",X"D1",X"B7",X"BD",X"DE",X"B7",X"BD",X"E0",X"8E",X"CC",X"22",
		X"1F",X"89",X"BD",X"14",X"0B",X"BD",X"08",X"D1",X"3D",X"F7",X"BD",X"E1",X"8E",X"BD",X"D6",X"BD",
		X"68",X"E3",X"8E",X"CC",X"00",X"BD",X"14",X"1C",X"4F",X"58",X"49",X"58",X"49",X"58",X"49",X"58",
		X"49",X"DD",X"85",X"FD",X"BD",X"DB",X"8E",X"BD",X"D6",X"A6",X"80",X"A7",X"88",X"3E",X"8C",X"BE",
		X"15",X"26",X"F6",X"8E",X"61",X"EC",X"86",X"00",X"BD",X"01",X"30",X"39",X"C6",X"07",X"BD",X"F4",
		X"83",X"BD",X"13",X"DD",X"BD",X"60",X"E2",X"BD",X"01",X"57",X"86",X"7F",X"97",X"91",X"9E",X"3F",
		X"9C",X"3B",X"26",X"04",X"AE",X"84",X"27",X"10",X"86",X"0F",X"8E",X"62",X"10",X"7E",X"00",X"A8",
		X"96",X"5B",X"9A",X"5C",X"9A",X"5B",X"26",X"F0",X"BD",X"08",X"0B",X"8E",X"62",X"26",X"86",X"00",
		X"BD",X"01",X"30",X"7E",X"00",X"0C",X"B6",X"C8",X"06",X"2B",X"05",X"BD",X"15",X"15",X"20",X"16",
		X"BD",X"13",X"BD",X"96",X"67",X"4A",X"26",X"05",X"BD",X"15",X"15",X"20",X"03",X"BD",X"15",X"1F",
		X"86",X"FF",X"97",X"57",X"97",X"58",X"4F",X"5F",X"DD",X"20",X"DD",X"22",X"BD",X"2C",X"00",X"BD",
		X"63",X"96",X"8E",X"BE",X"83",X"9F",X"77",X"BD",X"07",X"D9",X"9F",X"69",X"A6",X"09",X"84",X"0F",
		X"CE",X"65",X"A1",X"A6",X"C6",X"97",X"DE",X"6A",X"08",X"BD",X"1E",X"96",X"FC",X"BD",X"D6",X"26",
		X"15",X"FC",X"BD",X"D8",X"26",X"10",X"7F",X"BD",X"CF",X"86",X"78",X"B7",X"BD",X"D0",X"8E",X"2E",
		X"27",X"86",X"96",X"BD",X"70",X"52",X"BD",X"19",X"43",X"10",X"21",X"BD",X"63",X"7C",X"96",X"25",
		X"27",X"22",X"D6",X"68",X"5A",X"27",X"1D",X"D6",X"67",X"86",X"00",X"8E",X"3F",X"80",X"8D",X"66",
		X"24",X"03",X"8E",X"3F",X"4A",X"BD",X"70",X"58",X"8D",X"5C",X"25",X"08",X"86",X"80",X"8E",X"62",
		X"B4",X"7E",X"00",X"A8",X"8D",X"50",X"24",X"0B",X"BD",X"63",X"40",X"86",X"80",X"8E",X"62",X"C3",
		X"7E",X"00",X"A8",X"BD",X"13",X"DD",X"C6",X"00",X"9E",X"69",X"A6",X"0C",X"BD",X"19",X"3C",X"BD",
		X"65",X"DD",X"8E",X"20",X"FB",X"10",X"8E",X"63",X"5F",X"A6",X"A0",X"88",X"5A",X"27",X"05",X"BD",
		X"70",X"2B",X"20",X"F5",X"0F",X"3A",X"0F",X"39",X"86",X"10",X"97",X"88",X"86",X"60",X"8E",X"62",
		X"F4",X"7E",X"00",X"A8",X"BD",X"66",X"34",X"0F",X"3A",X"0F",X"39",X"86",X"10",X"97",X"88",X"0F",
		X"25",X"0C",X"66",X"7E",X"66",X"E4",X"34",X"12",X"9E",X"69",X"A6",X"09",X"BD",X"08",X"E4",X"84",
		X"0F",X"27",X"08",X"81",X"05",X"27",X"0D",X"1C",X"FE",X"35",X"92",X"BD",X"63",X"2F",X"81",X"13",
		X"26",X"F5",X"20",X"07",X"BD",X"63",X"2F",X"81",X"24",X"26",X"EC",X"1A",X"01",X"35",X"92",X"9E",
		X"69",X"A6",X"0F",X"AB",X"88",X"11",X"AB",X"88",X"12",X"AB",X"88",X"15",X"AB",X"88",X"14",X"39",
		X"34",X"36",X"10",X"9E",X"69",X"A6",X"29",X"BD",X"08",X"E4",X"1F",X"89",X"84",X"0F",X"27",X"08",
		X"86",X"0E",X"9E",X"69",X"6F",X"0C",X"20",X"02",X"86",X"0F",X"BD",X"70",X"55",X"35",X"B6",X"01",
		X"19",X"06",X"7A",X"6B",X"63",X"62",X"6B",X"7A",X"0D",X"13",X"16",X"16",X"13",X"1B",X"17",X"09",
		X"7A",X"1F",X"16",X"1F",X"19",X"67",X"7A",X"13",X"14",X"19",X"67",X"5A",X"BD",X"19",X"43",X"0F",
		X"CF",X"BD",X"19",X"43",X"10",X"0B",X"BD",X"19",X"43",X"1C",X"CF",X"BD",X"19",X"43",X"1C",X"A8",
		X"BD",X"19",X"43",X"6D",X"05",X"39",X"CC",X"03",X"00",X"DD",X"94",X"DD",X"92",X"7F",X"BE",X"C3",
		X"0F",X"87",X"0F",X"8F",X"0F",X"66",X"0F",X"89",X"0F",X"76",X"0F",X"75",X"0F",X"D2",X"0F",X"EB",
		X"0F",X"ED",X"CC",X"20",X"80",X"DD",X"98",X"DD",X"96",X"CC",X"20",X"00",X"DD",X"9A",X"CC",X"08",
		X"00",X"D3",X"20",X"DD",X"A3",X"CC",X"80",X"00",X"DD",X"9C",X"4F",X"5F",X"DD",X"9E",X"97",X"A0",
		X"DD",X"A1",X"DD",X"E9",X"39",X"96",X"E9",X"26",X"0B",X"BD",X"19",X"43",X"64",X"80",X"96",X"91",
		X"8A",X"08",X"97",X"91",X"39",X"EC",X"01",X"10",X"08",X"00",X"96",X"91",X"85",X"E8",X"26",X"F4",
		X"96",X"E9",X"26",X"F0",X"4F",X"8E",X"63",X"FB",X"7E",X"01",X"30",X"9E",X"69",X"A6",X"0B",X"26",
		X"0F",X"96",X"F0",X"26",X"78",X"0C",X"F0",X"CC",X"63",X"E5",X"BD",X"06",X"FD",X"7E",X"00",X"E4",
		X"97",X"E9",X"96",X"91",X"8A",X"10",X"97",X"91",X"1A",X"10",X"BD",X"0B",X"43",X"BD",X"0B",X"20",
		X"BD",X"0B",X"B3",X"1C",X"EF",X"9E",X"43",X"27",X"1E",X"CC",X"20",X"A9",X"0D",X"94",X"2A",X"03",
		X"CC",X"20",X"B3",X"ED",X"02",X"DC",X"A3",X"ED",X"0A",X"DC",X"9C",X"ED",X"0C",X"DC",X"96",X"C3",
		X"04",X"03",X"DD",X"D0",X"BD",X"27",X"03",X"BD",X"1D",X"F7",X"9E",X"69",X"6A",X"0B",X"27",X"22",
		X"A6",X"0B",X"81",X"0A",X"22",X"04",X"86",X"07",X"97",X"26",X"86",X"03",X"8E",X"64",X"62",X"7E",
		X"00",X"A8",X"0F",X"26",X"96",X"59",X"85",X"02",X"27",X"08",X"86",X"03",X"8E",X"64",X"47",X"7E",
		X"00",X"A8",X"0F",X"E9",X"96",X"91",X"84",X"EF",X"97",X"91",X"BD",X"1D",X"F7",X"7E",X"00",X"E4",
		X"86",X"03",X"DE",X"3F",X"A7",X"45",X"96",X"91",X"2A",X"06",X"86",X"D8",X"97",X"91",X"20",X"05",
		X"C6",X"58",X"BD",X"19",X"39",X"DC",X"20",X"DD",X"22",X"9E",X"96",X"CC",X"08",X"06",X"BD",X"13",
		X"B9",X"BD",X"65",X"B1",X"CC",X"06",X"68",X"BD",X"06",X"FD",X"10",X"8E",X"20",X"A9",X"96",X"92",
		X"2A",X"04",X"10",X"8E",X"20",X"B3",X"8E",X"65",X"9A",X"AF",X"47",X"CE",X"BC",X"03",X"BD",X"08",
		X"6A",X"1F",X"31",X"DE",X"3F",X"AF",X"4B",X"DC",X"98",X"10",X"AE",X"4B",X"BD",X"13",X"7D",X"86",
		X"02",X"8E",X"64",X"D7",X"7E",X"00",X"A8",X"DC",X"98",X"10",X"AE",X"4B",X"BD",X"13",X"36",X"AE",
		X"47",X"A6",X"80",X"27",X"0E",X"97",X"31",X"0F",X"26",X"AF",X"47",X"86",X"02",X"8E",X"64",X"C7",
		X"7E",X"00",X"A8",X"0D",X"91",X"2A",X"07",X"86",X"DA",X"97",X"91",X"7E",X"00",X"E4",X"86",X"7B",
		X"97",X"91",X"86",X"FF",X"97",X"26",X"86",X"02",X"8E",X"65",X"0E",X"7E",X"00",X"A8",X"0F",X"26",
		X"BD",X"01",X"57",X"96",X"DB",X"27",X"03",X"BD",X"19",X"72",X"9E",X"98",X"0D",X"43",X"27",X"03",
		X"BD",X"2C",X"09",X"0F",X"8D",X"C6",X"13",X"BD",X"06",X"EC",X"BD",X"68",X"8B",X"26",X"06",X"BD",
		X"69",X"9E",X"BD",X"13",X"DD",X"96",X"67",X"9E",X"69",X"E6",X"08",X"26",X"28",X"D6",X"68",X"5A",
		X"27",X"3A",X"88",X"03",X"BD",X"07",X"E8",X"E6",X"08",X"27",X"31",X"D6",X"67",X"86",X"00",X"8E",
		X"3F",X"78",X"BD",X"70",X"58",X"86",X"01",X"8E",X"3D",X"88",X"BD",X"70",X"58",X"86",X"60",X"8E",
		X"65",X"65",X"7E",X"00",X"A8",X"96",X"67",X"4C",X"91",X"68",X"23",X"02",X"86",X"01",X"BD",X"07",
		X"E8",X"E6",X"08",X"27",X"F2",X"97",X"67",X"0C",X"25",X"7E",X"61",X"EC",X"86",X"FF",X"97",X"91",
		X"86",X"01",X"8E",X"3D",X"80",X"BD",X"70",X"58",X"0F",X"8D",X"C6",X"13",X"BD",X"06",X"EC",X"86",
		X"60",X"8E",X"65",X"97",X"7E",X"00",X"A8",X"7E",X"E9",X"43",X"07",X"0F",X"3F",X"7F",X"FF",X"17",
		X"00",X"00",X"BB",X"33",X"22",X"11",X"44",X"66",X"77",X"00",X"99",X"FF",X"88",X"11",X"77",X"99",
		X"44",X"34",X"56",X"DE",X"69",X"33",X"4C",X"86",X"33",X"6F",X"C0",X"4A",X"26",X"FB",X"DE",X"69",
		X"B6",X"BE",X"54",X"A7",X"4C",X"33",X"4D",X"8E",X"BE",X"55",X"A6",X"80",X"8C",X"BE",X"56",X"22",
		X"03",X"AB",X"88",X"26",X"A7",X"C0",X"8C",X"BE",X"7C",X"26",X"EF",X"35",X"D6",X"BE",X"45",X"58",
		X"86",X"00",X"BD",X"01",X"30",X"CE",X"BE",X"83",X"31",X"C4",X"EF",X"07",X"6F",X"C0",X"11",X"83",
		X"BE",X"97",X"26",X"F8",X"DE",X"69",X"A6",X"4C",X"B7",X"BE",X"54",X"27",X"22",X"81",X"07",X"23",
		X"11",X"44",X"44",X"5F",X"BD",X"45",X"46",X"CB",X"40",X"26",X"F9",X"48",X"48",X"40",X"AB",X"4C",
		X"27",X"0D",X"97",X"4F",X"D6",X"B7",X"86",X"01",X"BD",X"45",X"46",X"0A",X"4F",X"26",X"F5",X"39",
		X"34",X"50",X"CE",X"BE",X"5E",X"30",X"88",X"16",X"A6",X"80",X"A7",X"C0",X"11",X"83",X"BE",X"7C",
		X"26",X"F6",X"35",X"D0",X"DE",X"69",X"33",X"4D",X"8E",X"BE",X"55",X"A6",X"C0",X"A7",X"80",X"8C",
		X"BE",X"7C",X"26",X"F7",X"8E",X"BE",X"7C",X"6F",X"80",X"8C",X"BE",X"83",X"26",X"F9",X"9E",X"69",
		X"A6",X"09",X"4A",X"26",X"06",X"BD",X"68",X"DF",X"BD",X"66",X"20",X"B6",X"BE",X"59",X"7F",X"BE",
		X"59",X"20",X"2C",X"BD",X"01",X"88",X"96",X"B6",X"44",X"8B",X"2C",X"A7",X"0C",X"BD",X"07",X"EC",
		X"84",X"3F",X"8B",X"80",X"D3",X"20",X"ED",X"0A",X"96",X"51",X"81",X"06",X"23",X"02",X"86",X"06",
		X"31",X"84",X"BD",X"38",X"46",X"9E",X"43",X"AF",X"A4",X"10",X"9F",X"43",X"40",X"9B",X"51",X"97",
		X"51",X"26",X"D0",X"B6",X"BE",X"58",X"27",X"06",X"7F",X"BE",X"58",X"BD",X"45",X"43",X"B6",X"BE",
		X"57",X"27",X"03",X"BD",X"38",X"43",X"B6",X"BE",X"56",X"20",X"0F",X"81",X"03",X"23",X"02",X"86",
		X"03",X"34",X"02",X"BD",X"1B",X"13",X"96",X"51",X"A0",X"E0",X"97",X"51",X"26",X"ED",X"B6",X"BE",
		X"5B",X"27",X"03",X"BD",X"6D",X"6D",X"B6",X"BE",X"5A",X"27",X"06",X"7F",X"BE",X"5A",X"BD",X"4F",
		X"43",X"B6",X"BE",X"5C",X"27",X"03",X"BD",X"4F",X"40",X"B6",X"BE",X"5D",X"27",X"03",X"BD",X"5A",
		X"D0",X"0F",X"39",X"39",X"DE",X"3F",X"86",X"28",X"A7",X"47",X"B6",X"BE",X"6D",X"B7",X"BE",X"7E",
		X"86",X"01",X"B7",X"BE",X"7D",X"6F",X"49",X"96",X"59",X"85",X"02",X"26",X"02",X"0F",X"F0",X"96",
		X"91",X"85",X"08",X"10",X"26",X"00",X"BF",X"BD",X"68",X"8B",X"26",X"55",X"10",X"BE",X"45",X"5A",
		X"BD",X"15",X"3A",X"26",X"08",X"86",X"0F",X"8E",X"67",X"0C",X"7E",X"00",X"A8",X"86",X"77",X"97",
		X"91",X"BD",X"01",X"57",X"BD",X"65",X"B1",X"86",X"01",X"8E",X"67",X"2F",X"7E",X"00",X"A8",X"10",
		X"8E",X"9C",X"9D",X"BD",X"19",X"43",X"0F",X"CF",X"BD",X"19",X"43",X"1C",X"CF",X"BD",X"19",X"43",
		X"1C",X"A8",X"86",X"37",X"A1",X"A8",X"62",X"27",X"0E",X"96",X"B6",X"81",X"30",X"24",X"08",X"D6",
		X"B7",X"86",X"9C",X"1F",X"01",X"63",X"84",X"BD",X"69",X"9E",X"9E",X"69",X"6C",X"08",X"7E",X"61",
		X"F1",X"81",X"08",X"22",X"12",X"F6",X"BE",X"6D",X"54",X"81",X"03",X"22",X"01",X"54",X"5C",X"F1",
		X"BE",X"7E",X"24",X"03",X"F7",X"BE",X"7E",X"7A",X"BE",X"7E",X"26",X"19",X"81",X"04",X"B6",X"BE",
		X"6D",X"24",X"05",X"44",X"44",X"BD",X"08",X"C1",X"B7",X"BE",X"7E",X"B6",X"BE",X"7F",X"81",X"0C",
		X"24",X"03",X"BD",X"38",X"40",X"7A",X"BE",X"7D",X"27",X"05",X"B6",X"BE",X"7C",X"26",X"27",X"B6",
		X"BE",X"5E",X"B7",X"BE",X"7D",X"B6",X"BE",X"55",X"27",X"1C",X"B6",X"BE",X"7C",X"81",X"08",X"24",
		X"15",X"B6",X"BE",X"5F",X"B1",X"BE",X"55",X"23",X"03",X"B6",X"BE",X"55",X"BD",X"45",X"40",X"40",
		X"BB",X"BE",X"55",X"B7",X"BE",X"55",X"96",X"88",X"81",X"10",X"24",X"02",X"0C",X"88",X"96",X"24",
		X"4C",X"81",X"D2",X"23",X"06",X"C6",X"06",X"BD",X"F4",X"83",X"4F",X"97",X"24",X"DE",X"3F",X"6A",
		X"47",X"26",X"0D",X"C6",X"02",X"10",X"8E",X"BE",X"55",X"BD",X"69",X"75",X"86",X"28",X"A7",X"47",
		X"9E",X"69",X"A6",X"09",X"4A",X"26",X"31",X"A6",X"49",X"26",X"2D",X"96",X"D2",X"26",X"16",X"EC",
		X"01",X"10",X"83",X"00",X"20",X"24",X"0E",X"A6",X"08",X"81",X"01",X"23",X"1B",X"EC",X"01",X"10",
		X"83",X"00",X"10",X"25",X"13",X"96",X"91",X"85",X"08",X"26",X"0D",X"86",X"01",X"A7",X"49",X"BD",
		X"68",X"DF",X"BD",X"66",X"20",X"BD",X"45",X"55",X"B6",X"BE",X"54",X"27",X"3C",X"96",X"D2",X"26",
		X"38",X"BD",X"45",X"49",X"27",X"33",X"8E",X"68",X"87",X"BC",X"BD",X"CD",X"27",X"09",X"CC",X"18",
		X"FF",X"FD",X"BD",X"D1",X"BD",X"37",X"40",X"86",X"FF",X"97",X"2D",X"86",X"05",X"8E",X"68",X"53",
		X"7E",X"00",X"A8",X"86",X"FF",X"97",X"2D",X"86",X"04",X"8E",X"68",X"5F",X"7E",X"00",X"A8",X"0F",
		X"2D",X"86",X"06",X"8E",X"66",X"F7",X"7E",X"00",X"A8",X"8E",X"68",X"87",X"BC",X"BD",X"CD",X"26",
		X"05",X"86",X"01",X"B7",X"BD",X"D0",X"96",X"57",X"81",X"E2",X"26",X"03",X"BD",X"4F",X"46",X"86",
		X"0F",X"8E",X"66",X"F7",X"7E",X"00",X"A8",X"F0",X"44",X"FF",X"06",X"B6",X"BE",X"7C",X"BB",X"BE",
		X"55",X"BB",X"BE",X"56",X"BB",X"BE",X"57",X"BB",X"BE",X"59",X"BB",X"BE",X"58",X"BB",X"BE",X"5A",
		X"BB",X"BE",X"5C",X"BB",X"BE",X"5D",X"39",X"34",X"16",X"86",X"05",X"E6",X"09",X"5A",X"8D",X"08",
		X"26",X"04",X"86",X"0A",X"A7",X"0C",X"35",X"96",X"34",X"06",X"E0",X"E4",X"25",X"02",X"26",X"FA",
		X"35",X"86",X"34",X"76",X"CE",X"69",X"D7",X"BD",X"07",X"D9",X"30",X"0D",X"8B",X"04",X"10",X"8E",
		X"00",X"09",X"E6",X"C6",X"E7",X"80",X"33",X"C8",X"10",X"31",X"3F",X"26",X"F5",X"35",X"F6",X"34",
		X"56",X"20",X"08",X"34",X"56",X"6C",X"09",X"8D",X"BE",X"A6",X"09",X"34",X"02",X"81",X"0B",X"23",
		X"02",X"86",X"0B",X"CE",X"69",X"D7",X"8B",X"04",X"30",X"0D",X"E6",X"C6",X"E7",X"80",X"33",X"C8",
		X"10",X"11",X"83",X"6C",X"47",X"26",X"F3",X"E6",X"E4",X"86",X"05",X"8D",X"AB",X"26",X"0A",X"8D",
		X"B1",X"86",X"0A",X"8D",X"A3",X"26",X"02",X"8D",X"A9",X"A6",X"E4",X"80",X"0B",X"24",X"01",X"4F",
		X"97",X"4F",X"8E",X"CC",X"1C",X"BD",X"14",X"1A",X"BD",X"08",X"D1",X"A1",X"E4",X"22",X"1A",X"1E",
		X"89",X"BD",X"08",X"D1",X"A1",X"E4",X"23",X"02",X"A6",X"E4",X"34",X"04",X"A0",X"E0",X"4C",X"F6",
		X"CC",X"21",X"C4",X"0F",X"3D",X"DB",X"4F",X"D7",X"4F",X"32",X"61",X"8E",X"CC",X"18",X"BD",X"14",
		X"1A",X"BD",X"08",X"D1",X"9B",X"4F",X"97",X"4F",X"27",X"19",X"1F",X"98",X"BD",X"08",X"D1",X"91",
		X"4F",X"24",X"02",X"97",X"4F",X"96",X"4F",X"C6",X"03",X"BD",X"07",X"D9",X"31",X"0D",X"8D",X"05",
		X"4A",X"26",X"F4",X"35",X"D6",X"34",X"32",X"8E",X"69",X"D7",X"A6",X"85",X"2B",X"0A",X"AB",X"A4",
		X"25",X"10",X"A1",X"84",X"22",X"0C",X"20",X"08",X"AB",X"A4",X"24",X"06",X"A1",X"01",X"25",X"02",
		X"A7",X"A4",X"31",X"21",X"30",X"88",X"10",X"8C",X"6C",X"47",X"26",X"DE",X"35",X"B2",X"9E",X"69",
		X"A6",X"09",X"BD",X"08",X"E4",X"84",X"0F",X"81",X"05",X"26",X"26",X"CC",X"02",X"25",X"BD",X"14",
		X"3A",X"86",X"97",X"0F",X"26",X"BD",X"13",X"DD",X"BD",X"70",X"55",X"35",X"10",X"AF",X"47",X"86",
		X"C0",X"8E",X"69",X"C7",X"7E",X"00",X"A8",X"9E",X"69",X"BD",X"5F",X"C1",X"DE",X"3F",X"6E",X"D8",
		X"07",X"BD",X"15",X"4D",X"7E",X"15",X"68",X"14",X"00",X"00",X"00",X"0B",X"0B",X"0A",X"0A",X"12",
		X"00",X"11",X"11",X"11",X"11",X"00",X"12",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"02",X"03",X"03",X"03",X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"00",X"04",X"04",X"04",X"04",X"06",X"04",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"05",
		X"16",X"05",X"05",X"05",X"06",X"00",X"03",X"03",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",X"00",X"00",X"00",X"03",X"03",X"03",X"06",X"03",
		X"00",X"03",X"03",X"03",X"04",X"0D",X"04",X"03",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"03",
		X"06",X"03",X"03",X"03",X"03",X"00",X"04",X"1E",X"00",X"00",X"00",X"1E",X"1E",X"19",X"14",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"04",X"00",X"00",X"00",X"04",X"04",X"03",X"03",X"05",
		X"05",X"04",X"04",X"04",X"04",X"04",X"04",X"60",X"00",X"03",X"02",X"16",X"16",X"1E",X"24",X"2E",
		X"30",X"32",X"34",X"36",X"38",X"3A",X"3C",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"10",X"00",X"50",X"70",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"FC",X"FE",X"FF",X"4A",X"3A",X"2A",X"2A",
		X"28",X"26",X"24",X"22",X"20",X"1E",X"1C",X"30",X"00",X"00",X"00",X"20",X"20",X"28",X"2C",X"30",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"03",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",
		X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"08",X"06",X"40",X"62",X"E0",X"02",X"12",
		X"18",X"1E",X"24",X"2A",X"30",X"36",X"3C",X"60",X"00",X"08",X"04",X"08",X"0C",X"1C",X"24",X"28",
		X"2C",X"30",X"34",X"38",X"3C",X"40",X"44",X"FF",X"08",X"FE",X"FE",X"FF",X"2A",X"22",X"1E",X"1C",
		X"1A",X"18",X"16",X"14",X"12",X"10",X"0E",X"60",X"00",X"08",X"02",X"16",X"16",X"1E",X"20",X"22",
		X"24",X"26",X"28",X"2A",X"2C",X"2E",X"30",X"28",X"0A",X"FE",X"FF",X"19",X"19",X"19",X"19",X"18",
		X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"3F",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"3F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"FF",X"30",X"F8",X"FC",X"F0",X"D4",X"C4",X"A4",X"94",
		X"90",X"8C",X"8A",X"89",X"88",X"87",X"86",X"14",X"03",X"FF",X"FF",X"0F",X"0F",X"0D",X"0C",X"0A",
		X"09",X"08",X"07",X"06",X"05",X"04",X"03",X"C8",X"28",X"F4",X"F8",X"FA",X"F0",X"DC",X"C8",X"C8",
		X"C0",X"B8",X"B0",X"A8",X"A2",X"9A",X"92",X"FF",X"02",X"00",X"00",X"FF",X"60",X"0C",X"06",X"05",
		X"04",X"04",X"04",X"04",X"04",X"04",X"03",X"FF",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"68",X"18",X"01",X"01",X"20",X"20",X"38",X"48",X"58",
		X"58",X"58",X"58",X"58",X"58",X"58",X"58",X"F2",X"D0",X"01",X"02",X"80",X"80",X"C8",X"D3",X"D4",
		X"D7",X"DA",X"DD",X"E0",X"E3",X"E7",X"EA",X"FF",X"00",X"00",X"00",X"30",X"30",X"40",X"50",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"FF",X"00",X"04",X"08",X"28",X"28",X"38",X"50",X"50",
		X"F8",X"50",X"60",X"70",X"80",X"90",X"A0",X"50",X"00",X"02",X"02",X"01",X"08",X"20",X"24",X"28",
		X"2C",X"2C",X"30",X"30",X"30",X"30",X"3C",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"D0",X"C0",
		X"B0",X"A8",X"A0",X"98",X"90",X"88",X"80",X"FF",X"00",X"00",X"00",X"60",X"60",X"50",X"40",X"30",
		X"2C",X"28",X"24",X"20",X"1C",X"1C",X"1C",X"FF",X"00",X"00",X"00",X"10",X"10",X"10",X"0F",X"0E",
		X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"08",X"FF",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"FF",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0C",X"28",X"26",X"1A",X"1B",X"25",X"0C",X"1B",
		X"25",X"0C",X"25",X"26",X"13",X"24",X"19",X"13",X"26",X"17",X"02",X"01",X"0C",X"58",X"16",X"17",
		X"25",X"1B",X"19",X"20",X"17",X"16",X"0C",X"17",X"2A",X"15",X"1E",X"27",X"25",X"1B",X"28",X"17",
		X"1E",X"2B",X"0C",X"18",X"21",X"24",X"01",X"0C",X"68",X"29",X"1B",X"1E",X"1E",X"1B",X"13",X"1F",
		X"25",X"0C",X"17",X"1E",X"17",X"15",X"26",X"24",X"21",X"20",X"1B",X"15",X"25",X"0C",X"1B",X"20",
		X"15",X"0F",X"02",X"01",X"0C",X"78",X"14",X"2B",X"0C",X"17",X"27",X"19",X"17",X"20",X"17",X"0C",
		X"22",X"0F",X"0C",X"1C",X"13",X"24",X"28",X"1B",X"25",X"0C",X"13",X"20",X"16",X"0C",X"1E",X"13",
		X"29",X"24",X"17",X"20",X"15",X"17",X"0C",X"17",X"0F",X"0C",X"16",X"17",X"1F",X"13",X"24",X"02",
		X"01",X"0C",X"A8",X"15",X"21",X"22",X"2B",X"24",X"1B",X"19",X"1A",X"26",X"0C",X"03",X"0B",X"0A",
		X"03",X"0C",X"29",X"1B",X"1E",X"1E",X"1B",X"13",X"1F",X"25",X"0C",X"17",X"1E",X"17",X"15",X"26",
		X"24",X"21",X"20",X"1B",X"15",X"25",X"0C",X"1B",X"20",X"15",X"0F",X"01",X"0C",X"B8",X"13",X"1E",
		X"1E",X"0C",X"24",X"1B",X"19",X"1A",X"26",X"25",X"0C",X"24",X"17",X"25",X"17",X"24",X"28",X"17",
		X"16",X"00",X"17",X"22",X"30",X"96",X"20",X"8E",X"6D",X"4D",X"44",X"44",X"44",X"84",X"7F",X"E6",
		X"86",X"D7",X"2D",X"44",X"8E",X"6D",X"3D",X"E6",X"86",X"A6",X"86",X"DD",X"D3",X"DD",X"D5",X"DD",
		X"D7",X"E6",X"47",X"5C",X"C1",X"02",X"23",X"01",X"5F",X"E7",X"47",X"8E",X"9C",X"D3",X"58",X"3A",
		X"CC",X"AA",X"AA",X"ED",X"84",X"86",X"04",X"8E",X"6D",X"05",X"7E",X"00",X"A8",X"22",X"BB",X"BB",
		X"BB",X"BB",X"BB",X"88",X"88",X"88",X"88",X"88",X"88",X"22",X"22",X"22",X"22",X"C7",X"C7",X"C7",
		X"C7",X"C7",X"C7",X"87",X"47",X"47",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",
		X"1F",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"57",X"97",X"87",X"97",X"4F",X"86",
		X"55",X"D6",X"B6",X"C4",X"03",X"26",X"01",X"5C",X"3D",X"1F",X"98",X"1F",X"03",X"BD",X"01",X"70",
		X"1A",X"D2",X"6D",X"A8",X"1F",X"00",X"EF",X"0A",X"BD",X"07",X"EC",X"84",X"1F",X"8B",X"5C",X"A7",
		X"0C",X"86",X"11",X"A7",X"88",X"14",X"4F",X"5F",X"ED",X"0E",X"ED",X"88",X"10",X"9F",X"41",X"33",
		X"C9",X"50",X"00",X"0A",X"4F",X"26",X"D6",X"39",X"96",X"DB",X"26",X"14",X"B6",X"BE",X"C3",X"26",
		X"0F",X"96",X"91",X"85",X"08",X"26",X"09",X"96",X"B5",X"27",X"05",X"BD",X"19",X"43",X"6D",X"C3",
		X"4F",X"35",X"86",X"8E",X"BE",X"F4",X"96",X"91",X"84",X"02",X"A7",X"47",X"86",X"77",X"97",X"91",
		X"C6",X"56",X"E1",X"88",X"CE",X"27",X"0E",X"96",X"B7",X"81",X"19",X"24",X"08",X"D6",X"B8",X"86",
		X"9C",X"1F",X"01",X"6A",X"84",X"96",X"D2",X"10",X"27",X"00",X"84",X"8E",X"CC",X"26",X"BD",X"14",
		X"0B",X"BD",X"08",X"D1",X"9E",X"69",X"A1",X"09",X"25",X"75",X"F6",X"CC",X"25",X"C4",X"0F",X"D0",
		X"D2",X"22",X"0D",X"96",X"92",X"98",X"9E",X"2B",X"66",X"C6",X"09",X"BD",X"F4",X"83",X"20",X"0F",
		X"8E",X"6F",X"1E",X"C1",X"01",X"26",X"03",X"8E",X"6F",X"22",X"BD",X"37",X"40",X"20",X"50",X"BD",
		X"01",X"57",X"BD",X"13",X"BD",X"BD",X"65",X"B1",X"86",X"01",X"8E",X"6E",X"30",X"7E",X"00",X"A8",
		X"0C",X"DB",X"BD",X"32",X"40",X"BD",X"19",X"72",X"BD",X"19",X"43",X"0F",X"CF",X"BD",X"19",X"43",
		X"1C",X"CF",X"BD",X"19",X"43",X"1C",X"A8",X"BD",X"1E",X"96",X"9E",X"69",X"6C",X"09",X"BD",X"68",
		X"A7",X"6C",X"09",X"BD",X"68",X"A7",X"A6",X"09",X"4C",X"BD",X"08",X"E4",X"1F",X"89",X"86",X"04",
		X"BD",X"70",X"58",X"86",X"20",X"BD",X"15",X"68",X"9E",X"69",X"6C",X"08",X"7E",X"61",X"F1",X"C6",
		X"1D",X"BD",X"45",X"52",X"86",X"01",X"8E",X"6E",X"7C",X"7E",X"00",X"A8",X"9E",X"49",X"27",X"05",
		X"BD",X"01",X"CD",X"20",X"F7",X"86",X"02",X"BD",X"6F",X"26",X"BD",X"13",X"DD",X"CE",X"BE",X"83",
		X"86",X"FF",X"97",X"4F",X"8E",X"00",X"00",X"10",X"AE",X"C1",X"27",X"16",X"EC",X"28",X"10",X"B3",
		X"45",X"5C",X"27",X"0E",X"EC",X"26",X"26",X"0A",X"A6",X"2C",X"91",X"4F",X"22",X"04",X"97",X"4F",
		X"30",X"A4",X"11",X"83",X"BE",X"97",X"26",X"DF",X"30",X"84",X"27",X"33",X"4F",X"5F",X"DD",X"9E",
		X"DD",X"A1",X"96",X"B6",X"84",X"07",X"40",X"AB",X"0C",X"80",X"14",X"81",X"31",X"24",X"02",X"86",
		X"31",X"81",X"68",X"23",X"02",X"86",X"68",X"97",X"9C",X"CC",X"20",X"11",X"0D",X"94",X"2A",X"03",
		X"CC",X"70",X"15",X"97",X"9A",X"34",X"04",X"97",X"98",X"EC",X"0A",X"A0",X"E0",X"20",X"04",X"DC",
		X"20",X"8B",X"80",X"DD",X"20",X"BD",X"2C",X"00",X"86",X"01",X"8E",X"6F",X"83",X"7E",X"00",X"A8",
		X"5F",X"96",X"E9",X"27",X"02",X"C6",X"10",X"DE",X"3F",X"EA",X"47",X"D7",X"91",X"86",X"28",X"B7",
		X"BE",X"C3",X"8E",X"6F",X"18",X"7E",X"00",X"A8",X"7F",X"BE",X"C3",X"7E",X"00",X"E4",X"80",X"04",
		X"90",X"07",X"80",X"04",X"90",X"08",X"35",X"10",X"AF",X"4D",X"A7",X"4B",X"10",X"8E",X"BC",X"71",
		X"8E",X"9C",X"26",X"EC",X"81",X"ED",X"A1",X"8C",X"9C",X"36",X"26",X"F7",X"86",X"07",X"A7",X"4C",
		X"A6",X"4B",X"8E",X"6F",X"48",X"7E",X"00",X"A8",X"8E",X"9C",X"26",X"8D",X"0C",X"8C",X"9C",X"36",
		X"26",X"F9",X"6A",X"4C",X"2A",X"EA",X"6E",X"D8",X"0D",X"A6",X"84",X"E6",X"84",X"C4",X"07",X"E1",
		X"4C",X"23",X"01",X"4A",X"E6",X"84",X"54",X"54",X"54",X"C4",X"07",X"E1",X"4C",X"23",X"02",X"80",
		X"08",X"E6",X"84",X"54",X"54",X"54",X"54",X"54",X"C4",X"06",X"E1",X"4C",X"23",X"02",X"80",X"40",
		X"A7",X"80",X"39",X"A6",X"47",X"34",X"02",X"BD",X"10",X"6E",X"BD",X"10",X"45",X"BD",X"10",X"CA",
		X"DE",X"3F",X"35",X"02",X"A7",X"47",X"96",X"91",X"84",X"DD",X"AA",X"47",X"97",X"91",X"86",X"01",
		X"8E",X"6F",X"A6",X"7E",X"00",X"A8",X"96",X"91",X"8A",X"20",X"97",X"91",X"86",X"02",X"BD",X"8F",
		X"00",X"7E",X"6F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"08",X"70",X"83",X"03",X"08",X"70",X"9B",X"03",X"08",X"70",X"B3",X"03",X"08",X"70",X"CB",
		X"03",X"08",X"70",X"E3",X"03",X"08",X"70",X"FB",X"03",X"08",X"71",X"13",X"03",X"08",X"71",X"2B",
		X"03",X"08",X"71",X"43",X"03",X"08",X"71",X"5B",X"7E",X"72",X"98",X"7E",X"72",X"B4",X"7E",X"72",
		X"B2",X"7E",X"73",X"01",X"7E",X"72",X"FF",X"7E",X"73",X"D9",X"7E",X"73",X"E2",X"7E",X"73",X"F6",
		X"7E",X"73",X"EC",X"7E",X"73",X"9F",X"7E",X"73",X"A8",X"7E",X"73",X"BC",X"7E",X"73",X"B2",X"7E",
		X"74",X"53",X"7E",X"74",X"51",X"7E",X"74",X"5B",X"7E",X"74",X"59",X"03",X"08",X"71",X"73",X"03",
		X"08",X"71",X"8B",X"03",X"08",X"71",X"A3",X"03",X"08",X"71",X"BB",X"03",X"08",X"71",X"D3",X"03",
		X"08",X"71",X"EB",X"03",X"08",X"72",X"03",X"03",X"08",X"72",X"1B",X"03",X"08",X"72",X"33",X"03",
		X"08",X"72",X"4B",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"11",X"00",X"00",X"01",X"10",
		X"00",X"11",X"00",X"11",X"11",X"11",X"10",X"00",X"00",X"11",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"10",X"00",X"11",X"00",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"01",X"01",X"01",X"00",
		X"00",X"01",X"00",X"11",X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"01",
		X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"11",X"10",
		X"10",X"11",X"00",X"11",X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"01",X"00",X"00",X"00",X"00",
		X"01",X"01",X"00",X"11",X"00",X"00",X"01",X"11",X"10",X"10",X"00",X"11",X"11",X"11",X"10",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"11",X"10",
		X"10",X"11",X"00",X"11",X"01",X"01",X"10",X"01",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"00",
		X"00",X"01",X"00",X"11",X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"11",X"01",X"01",X"11",X"01",
		X"01",X"11",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"CC",X"C0",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"00",X"0C",X"0C",X"00",X"00",X"00",X"0C",X"0C",X"00",X"CC",X"00",X"00",X"0C",X"C0",
		X"00",X"CC",X"00",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"CC",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"CC",X"00",X"00",X"CC",X"00",X"00",X"CC",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"00",X"00",X"00",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"CC",X"00",
		X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"0C",X"0C",X"0C",X"0C",X"00",
		X"00",X"0C",X"00",X"CC",X"C0",X"C0",X"CC",X"00",X"00",X"CC",X"00",X"CC",X"00",X"00",X"CC",X"0C",
		X"0C",X"CC",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"CC",X"C0",X"C0",X"CC",X"C0",
		X"C0",X"CC",X"00",X"CC",X"00",X"00",X"CC",X"0C",X"0C",X"CC",X"00",X"0C",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"CC",X"00",X"00",X"0C",X"CC",X"C0",X"C0",X"00",X"CC",X"CC",X"CC",X"C0",X"00",
		X"00",X"00",X"00",X"0C",X"0C",X"0C",X"00",X"0C",X"0C",X"0C",X"00",X"CC",X"C0",X"C0",X"CC",X"C0",
		X"C0",X"CC",X"00",X"CC",X"0C",X"0C",X"C0",X"0C",X"0C",X"CC",X"00",X"0C",X"0C",X"0C",X"0C",X"00",
		X"00",X"0C",X"00",X"CC",X"C0",X"C0",X"CC",X"00",X"00",X"CC",X"00",X"CC",X"0C",X"0C",X"CC",X"0C",
		X"0C",X"CC",X"00",X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"2D",X"20",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"31",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"34",X"02",X"86",X"11",X"97",X"10",X"35",X"02",
		X"34",X"02",X"86",X"07",X"97",X"13",X"0F",X"11",X"0F",X"16",X"86",X"01",X"97",X"12",X"9F",X"14",
		X"35",X"82",X"0F",X"11",X"34",X"66",X"0D",X"11",X"27",X"06",X"0F",X"11",X"30",X"89",X"01",X"00",
		X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"05",X"D7",X"13",X"10",X"8E",X"75",X"A6",X"81",X"20",X"26",
		X"02",X"86",X"3A",X"81",X"5E",X"22",X"26",X"80",X"30",X"25",X"22",X"48",X"10",X"AE",X"A6",X"EC",
		X"A1",X"94",X"10",X"D4",X"10",X"ED",X"81",X"EC",X"A1",X"94",X"10",X"D4",X"10",X"ED",X"81",X"EC",
		X"A0",X"94",X"10",X"A7",X"84",X"30",X"89",X"00",X"FC",X"C1",X"33",X"26",X"E2",X"35",X"E6",X"0F",
		X"11",X"34",X"66",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"07",X"D7",X"13",X"10",X"8E",X"78",X"13",
		X"8D",X"07",X"44",X"31",X"A6",X"8D",X"18",X"35",X"E6",X"81",X"20",X"26",X"02",X"86",X"3A",X"81",
		X"5E",X"22",X"FA",X"80",X"30",X"25",X"F6",X"31",X"A6",X"48",X"31",X"A6",X"31",X"A6",X"39",X"D6",
		X"13",X"CE",X"9C",X"18",X"33",X"C5",X"DF",X"E7",X"6F",X"C2",X"5A",X"26",X"FB",X"CE",X"9C",X"18",
		X"A6",X"A4",X"48",X"D6",X"11",X"26",X"1B",X"48",X"24",X"06",X"D6",X"10",X"C4",X"F0",X"20",X"01",
		X"5F",X"E7",X"C0",X"11",X"93",X"E7",X"25",X"EF",X"8D",X"22",X"6D",X"A0",X"2B",X"DF",X"8D",X"2D",
		X"20",X"1A",X"48",X"24",X"08",X"D6",X"10",X"C4",X"0F",X"EA",X"C4",X"E7",X"C4",X"33",X"41",X"11",
		X"93",X"E7",X"26",X"EE",X"8D",X"17",X"8D",X"04",X"6D",X"A0",X"2B",X"C1",X"34",X"02",X"96",X"11",
		X"27",X"06",X"86",X"FF",X"30",X"89",X"01",X"00",X"4C",X"97",X"11",X"35",X"82",X"34",X"10",X"CE",
		X"9C",X"18",X"A6",X"C0",X"A7",X"84",X"30",X"01",X"11",X"93",X"E7",X"26",X"F5",X"35",X"90",X"0F",
		X"11",X"34",X"66",X"86",X"05",X"5F",X"20",X"1B",X"0F",X"11",X"34",X"66",X"86",X"05",X"C6",X"01",
		X"20",X"11",X"0F",X"11",X"34",X"66",X"86",X"07",X"C6",X"01",X"20",X"07",X"0F",X"11",X"34",X"66",
		X"86",X"07",X"5F",X"97",X"13",X"D7",X"12",X"A6",X"E4",X"20",X"02",X"34",X"66",X"0F",X"17",X"8D",
		X"4A",X"0C",X"17",X"A6",X"E4",X"8D",X"48",X"35",X"E6",X"0F",X"11",X"34",X"66",X"86",X"05",X"5F",
		X"20",X"1B",X"0F",X"11",X"34",X"66",X"86",X"05",X"C6",X"01",X"20",X"11",X"0F",X"11",X"34",X"66",
		X"86",X"07",X"C6",X"01",X"20",X"07",X"0F",X"11",X"34",X"66",X"86",X"07",X"5F",X"97",X"13",X"D7",
		X"12",X"A6",X"E4",X"20",X"02",X"34",X"66",X"0F",X"17",X"8D",X"10",X"A6",X"E4",X"8D",X"10",X"A6",
		X"61",X"8D",X"08",X"0C",X"17",X"A6",X"61",X"8D",X"06",X"35",X"E6",X"44",X"44",X"44",X"44",X"84",
		X"0F",X"26",X"08",X"D6",X"17",X"26",X"04",X"D6",X"12",X"26",X"0F",X"0C",X"17",X"8B",X"30",X"D6",
		X"13",X"C1",X"07",X"10",X"27",X"FE",X"CA",X"7E",X"72",X"B4",X"C1",X"02",X"26",X"0E",X"30",X"89",
		X"02",X"00",X"D6",X"13",X"C1",X"05",X"27",X"04",X"30",X"89",X"01",X"00",X"39",X"34",X"66",X"20",
		X"10",X"0F",X"11",X"34",X"66",X"C6",X"05",X"20",X"06",X"0F",X"11",X"34",X"66",X"C6",X"07",X"D7",
		X"13",X"34",X"42",X"CE",X"9D",X"57",X"C6",X"37",X"0D",X"91",X"2B",X"13",X"E1",X"C8",X"A8",X"27",
		X"0E",X"96",X"B7",X"81",X"12",X"22",X"08",X"D6",X"B6",X"86",X"9C",X"1F",X"03",X"63",X"C4",X"35",
		X"42",X"1F",X"89",X"4F",X"58",X"49",X"10",X"8E",X"79",X"2D",X"10",X"AE",X"AB",X"A6",X"A0",X"27",
		X"1F",X"81",X"16",X"24",X"0B",X"4A",X"48",X"CE",X"74",X"B2",X"EE",X"C6",X"AD",X"C4",X"20",X"ED",
		X"D6",X"13",X"C1",X"07",X"26",X"05",X"BD",X"73",X"01",X"20",X"E2",X"BD",X"72",X"B4",X"20",X"DD",
		X"35",X"E6",X"74",X"E6",X"74",X"E8",X"74",X"F3",X"74",X"FC",X"75",X"01",X"75",X"39",X"75",X"40",
		X"75",X"4D",X"75",X"5A",X"75",X"5F",X"75",X"67",X"75",X"6C",X"75",X"71",X"75",X"76",X"75",X"8A",
		X"75",X"7B",X"75",X"80",X"75",X"32",X"75",X"85",X"74",X"DC",X"75",X"62",X"B6",X"C8",X"06",X"10",
		X"2B",X"00",X"A7",X"EC",X"A1",X"39",X"8D",X"0B",X"1F",X"10",X"96",X"14",X"1F",X"01",X"96",X"16",
		X"97",X"11",X"39",X"1F",X"10",X"DB",X"13",X"CB",X"02",X"1F",X"01",X"39",X"A6",X"A0",X"97",X"10",
		X"39",X"1F",X"10",X"AB",X"A4",X"EB",X"21",X"1F",X"01",X"6D",X"22",X"27",X"22",X"6D",X"A4",X"2B",
		X"0F",X"96",X"11",X"27",X"06",X"30",X"89",X"01",X"00",X"86",X"FF",X"4C",X"97",X"11",X"20",X"0F",
		X"96",X"11",X"81",X"01",X"27",X"06",X"30",X"89",X"FF",X"00",X"86",X"02",X"4A",X"97",X"11",X"31",
		X"23",X"39",X"AE",X"A1",X"A6",X"A0",X"97",X"11",X"39",X"D6",X"11",X"D7",X"16",X"9F",X"14",X"39",
		X"96",X"13",X"81",X"07",X"27",X"06",X"86",X"07",X"97",X"13",X"30",X"1E",X"39",X"96",X"13",X"81",
		X"05",X"27",X"F9",X"86",X"05",X"97",X"13",X"30",X"02",X"39",X"86",X"01",X"97",X"12",X"39",X"0F",
		X"12",X"39",X"86",X"02",X"97",X"12",X"39",X"EC",X"A1",X"7E",X"74",X"05",X"EC",X"B1",X"7E",X"74",
		X"05",X"A6",X"A0",X"7E",X"73",X"CB",X"A6",X"B1",X"7E",X"73",X"CB",X"A6",X"63",X"7E",X"73",X"CB",
		X"EC",X"64",X"7E",X"74",X"05",X"A6",X"B1",X"97",X"10",X"39",X"32",X"78",X"E6",X"6B",X"E7",X"61",
		X"EC",X"6C",X"ED",X"62",X"CC",X"75",X"A3",X"ED",X"66",X"EC",X"A1",X"10",X"AF",X"64",X"1F",X"02",
		X"7E",X"74",X"8D",X"1F",X"32",X"39",X"76",X"04",X"76",X"0F",X"76",X"1A",X"76",X"25",X"76",X"30",
		X"76",X"3B",X"76",X"46",X"76",X"51",X"76",X"5C",X"76",X"67",X"76",X"72",X"76",X"78",X"76",X"83",
		X"76",X"8E",X"76",X"99",X"76",X"A9",X"76",X"B4",X"76",X"BF",X"76",X"CA",X"76",X"D5",X"76",X"E0",
		X"76",X"EB",X"76",X"F6",X"77",X"01",X"77",X"0C",X"77",X"17",X"77",X"1D",X"77",X"28",X"77",X"33",
		X"77",X"3E",X"77",X"4E",X"77",X"59",X"77",X"64",X"77",X"6F",X"77",X"7A",X"77",X"85",X"77",X"90",
		X"77",X"9B",X"77",X"A6",X"77",X"B1",X"77",X"C1",X"77",X"CC",X"77",X"D7",X"77",X"E2",X"77",X"ED",
		X"77",X"F3",X"78",X"03",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"00",X"FF",X"F0",X"FF",X"F0",
		X"F0",X"F0",X"00",X"F0",X"33",X"FF",X"00",X"0F",X"00",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",
		X"F0",X"F0",X"FF",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"00",X"FF",
		X"F0",X"00",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",
		X"33",X"FF",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",
		X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"00",X"00",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"33",X"00",X"00",X"00",X"00",X"00",X"33",X"0F",X"0F",X"0F",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"F0",X"33",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"0F",X"FF",X"00",X"00",X"F0",X"FF",
		X"FF",X"F0",X"F0",X"00",X"00",X"F0",X"00",X"00",X"33",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"33",X"FF",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",
		X"F0",X"00",X"F0",X"F0",X"33",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"00",X"00",X"00",X"F0",X"33",
		X"FF",X"F0",X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"00",X"33",X"FF",X"F0",X"FF",X"F0",X"FF",
		X"F0",X"00",X"F0",X"00",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"00",X"F0",X"00",X"00",
		X"33",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",X"33",X"F0",X"F0",X"FF",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"00",X"00",X"00",
		X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"00",
		X"F0",X"F0",X"33",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"00",X"00",X"F0",X"33",X"FF",X"F0",
		X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"33",X"FF",
		X"F0",X"F0",X"FF",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"F0",X"F0",X"F0",
		X"F0",X"00",X"F0",X"F0",X"33",X"FF",X"F0",X"FF",X"00",X"FF",X"F0",X"00",X"F0",X"F0",X"F0",X"33",
		X"FF",X"0F",X"0F",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"33",X"F0",X"F0",X"F0",X"F0",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"33",X"F0",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",X"00",
		X"33",X"F0",X"F0",X"F0",X"F0",X"FF",X"00",X"00",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"33",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"00",X"F0",X"F0",X"33",X"F0",X"F0",X"FF",X"0F",
		X"0F",X"F0",X"F0",X"F0",X"00",X"00",X"33",X"FF",X"00",X"0F",X"F0",X"FF",X"F0",X"F0",X"00",X"00",
		X"F0",X"33",X"00",X"0F",X"0F",X"0F",X"00",X"F0",X"00",X"00",X"00",X"F0",X"33",X"F0",X"0F",X"0F",
		X"0F",X"F0",X"33",X"00",X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"F0",X"FF",
		X"F0",X"00",X"33",X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"33",X"FF",X"C1",X"C1",X"FF",X"7F",X"00",X"90",X"B0",X"E0",X"FF",X"7F",X"00",X"C3",
		X"C7",X"C9",X"F9",X"71",X"00",X"C1",X"C9",X"C9",X"FF",X"7F",X"00",X"98",X"A8",X"C8",X"FF",X"7F",
		X"00",X"F9",X"F9",X"C9",X"C9",X"4F",X"00",X"FF",X"FF",X"C9",X"C9",X"4F",X"00",X"C3",X"C7",X"CC",
		X"F8",X"70",X"00",X"F7",X"FF",X"C9",X"C9",X"77",X"00",X"F9",X"F9",X"C9",X"C9",X"7F",X"00",X"80",
		X"80",X"00",X"00",X"00",X"00",X"FD",X"FD",X"80",X"00",X"00",X"00",X"86",X"87",X"80",X"00",X"00",
		X"00",X"83",X"83",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"B6",X"B6",
		X"00",X"00",X"00",X"98",X"98",X"98",X"18",X"00",X"00",X"FF",X"E8",X"E8",X"E8",X"FF",X"7F",X"FF",
		X"FF",X"EB",X"EB",X"FF",X"3E",X"FF",X"FF",X"C3",X"C3",X"C3",X"43",X"FF",X"C3",X"C3",X"C3",X"FF",
		X"3E",X"FF",X"FF",X"D3",X"D3",X"D3",X"43",X"FF",X"FF",X"D0",X"D0",X"D0",X"40",X"FF",X"FF",X"C3",
		X"CB",X"EB",X"6F",X"FF",X"FF",X"8C",X"8C",X"8C",X"7F",X"FF",X"7F",X"00",X"00",X"00",X"00",X"83",
		X"81",X"81",X"81",X"FF",X"7F",X"FF",X"FF",X"90",X"AC",X"E6",X"43",X"FF",X"83",X"83",X"83",X"83",
		X"03",X"FF",X"FF",X"E0",X"F8",X"E0",X"7F",X"FF",X"FF",X"E0",X"E0",X"E0",X"7F",X"FF",X"FF",X"C3",
		X"C3",X"C3",X"7F",X"FF",X"FF",X"D8",X"D8",X"D8",X"78",X"FF",X"FF",X"C3",X"C7",X"FF",X"01",X"FF",
		X"FF",X"D0",X"DC",X"D6",X"73",X"83",X"F3",X"D3",X"D3",X"DF",X"40",X"C0",X"C0",X"FF",X"FF",X"C0",
		X"40",X"FF",X"FF",X"83",X"83",X"83",X"7F",X"FC",X"FE",X"83",X"81",X"82",X"7C",X"FF",X"FF",X"83",
		X"8F",X"83",X"7F",X"E3",X"F7",X"9C",X"94",X"63",X"00",X"E0",X"F0",X"9F",X"8F",X"90",X"60",X"C3",
		X"C7",X"CB",X"D3",X"E3",X"43",X"9C",X"A2",X"41",X"00",X"00",X"00",X"C1",X"A2",X"1C",X"00",X"00",
		X"00",X"82",X"84",X"88",X"90",X"20",X"00",X"88",X"9C",X"BE",X"88",X"08",X"00",X"8B",X"0F",X"8B",
		X"1B",X"8B",X"62",X"8B",X"40",X"8B",X"27",X"8A",X"80",X"8A",X"95",X"8A",X"D1",X"8A",X"FF",X"8A",
		X"3C",X"8A",X"5B",X"8A",X"77",X"8A",X"B4",X"8A",X"34",X"89",X"FC",X"8A",X"17",X"89",X"8E",X"89",
		X"D8",X"89",X"CD",X"84",X"FC",X"85",X"1C",X"85",X"37",X"85",X"5F",X"85",X"DF",X"85",X"F0",X"83",
		X"E1",X"84",X"37",X"84",X"43",X"84",X"60",X"84",X"6A",X"84",X"E8",X"89",X"B7",X"89",X"C2",X"83",
		X"CF",X"83",X"0A",X"83",X"12",X"83",X"1A",X"83",X"25",X"83",X"36",X"83",X"40",X"83",X"4C",X"83",
		X"58",X"83",X"60",X"83",X"6A",X"83",X"78",X"83",X"86",X"83",X"8B",X"83",X"9E",X"83",X"A9",X"83",
		X"B1",X"83",X"B7",X"82",X"D5",X"81",X"CA",X"82",X"96",X"82",X"A6",X"82",X"B8",X"82",X"19",X"82",
		X"2E",X"82",X"42",X"82",X"5F",X"82",X"74",X"82",X"88",X"81",X"BD",X"81",X"C0",X"81",X"C3",X"7F",
		X"14",X"7F",X"1A",X"7F",X"BE",X"7F",X"CF",X"7F",X"EF",X"7F",X"F7",X"80",X"09",X"80",X"11",X"80",
		X"1B",X"80",X"30",X"80",X"3A",X"80",X"4A",X"80",X"7B",X"80",X"85",X"80",X"A3",X"80",X"AE",X"80",
		X"B9",X"80",X"C0",X"80",X"E8",X"81",X"05",X"81",X"1A",X"81",X"2D",X"81",X"44",X"81",X"67",X"81",
		X"72",X"81",X"7B",X"81",X"92",X"81",X"9D",X"81",X"B6",X"7C",X"D2",X"7C",X"D8",X"7C",X"FB",X"7C",
		X"FE",X"7D",X"15",X"7D",X"1B",X"7D",X"31",X"7D",X"70",X"7D",X"74",X"7D",X"77",X"7D",X"90",X"7D",
		X"97",X"7D",X"A3",X"7D",X"B7",X"7E",X"5D",X"7E",X"68",X"7E",X"CD",X"7D",X"4C",X"7D",X"D0",X"7D",
		X"E5",X"7D",X"F7",X"7E",X"0E",X"7E",X"1E",X"7E",X"33",X"7E",X"42",X"7E",X"53",X"7D",X"BE",X"81",
		X"D6",X"86",X"0A",X"86",X"18",X"86",X"3E",X"7B",X"30",X"81",X"E7",X"86",X"59",X"86",X"6B",X"86",
		X"7C",X"86",X"87",X"86",X"95",X"86",X"A4",X"86",X"E5",X"86",X"FB",X"7B",X"C6",X"7C",X"36",X"7C",
		X"94",X"7C",X"A7",X"7C",X"C2",X"7C",X"C8",X"7C",X"CB",X"85",X"7C",X"85",X"89",X"85",X"96",X"85",
		X"AF",X"85",X"BC",X"85",X"C9",X"7B",X"4E",X"7A",X"DD",X"89",X"4F",X"7A",X"5F",X"7A",X"A1",X"04",
		X"EE",X"12",X"1C",X"70",X"00",X"59",X"4C",X"4C",X"41",X"42",X"49",X"41",X"4E",X"20",X"53",X"54",
		X"41",X"52",X"46",X"4C",X"45",X"45",X"54",X"20",X"54",X"45",X"52",X"4D",X"49",X"4E",X"41",X"54",
		X"45",X"44",X"3D",X"3D",X"3D",X"04",X"FF",X"12",X"3C",X"90",X"00",X"32",X"35",X"30",X"30",X"3A",
		X"3A",X"04",X"DD",X"42",X"04",X"EE",X"4F",X"04",X"FF",X"4E",X"04",X"DD",X"55",X"04",X"EE",X"53",
		X"00",X"04",X"FF",X"12",X"28",X"70",X"00",X"46",X"49",X"52",X"45",X"42",X"4F",X"4D",X"42",X"45",
		X"52",X"20",X"53",X"54",X"52",X"49",X"4B",X"45",X"46",X"4F",X"52",X"43",X"45",X"20",X"41",X"4E",
		X"4E",X"49",X"48",X"49",X"4C",X"41",X"54",X"45",X"44",X"3A",X"3B",X"04",X"AA",X"12",X"38",X"90",
		X"00",X"35",X"30",X"30",X"30",X"20",X"20",X"42",X"4F",X"4E",X"55",X"53",X"00",X"04",X"99",X"12",
		X"13",X"70",X"00",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"54",X"48",X"45",X"20",X"4C",X"49",
		X"4E",X"45",X"20",X"55",X"53",X"49",X"4E",X"47",X"20",X"54",X"48",X"52",X"55",X"53",X"54",X"20",
		X"41",X"4E",X"44",X"20",X"46",X"49",X"52",X"45",X"12",X"1E",X"7E",X"00",X"50",X"52",X"45",X"53",
		X"53",X"20",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"57",X"48",X"45",X"4E",X"20",X"43",
		X"45",X"4E",X"54",X"45",X"52",X"45",X"44",X"04",X"BB",X"08",X"12",X"4B",X"50",X"00",X"3E",X"00",
		X"04",X"BB",X"12",X"2C",X"16",X"00",X"41",X"54",X"54",X"52",X"41",X"43",X"54",X"20",X"4D",X"4F",
		X"44",X"45",X"20",X"4D",X"45",X"53",X"53",X"41",X"47",X"45",X"0F",X"7B",X"8A",X"00",X"04",X"BB",
		X"12",X"20",X"70",X"00",X"35",X"20",X"45",X"4E",X"54",X"52",X"49",X"45",X"53",X"20",X"4D",X"41",
		X"58",X"49",X"4D",X"55",X"4D",X"20",X"50",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"12",X"28",X"90",X"01",X"4C",X"4F",X"57",X"45",X"53",X"54",X"20",X"45",X"4E",X"54",X"52",X"59",
		X"20",X"52",X"45",X"50",X"4C",X"41",X"43",X"45",X"44",X"00",X"08",X"04",X"33",X"12",X"2C",X"C0",
		X"00",X"0F",X"7F",X"A1",X"4C",X"45",X"54",X"54",X"45",X"52",X"12",X"37",X"CC",X"00",X"55",X"53",
		X"45",X"20",X"46",X"49",X"52",X"45",X"20",X"54",X"4F",X"20",X"45",X"4E",X"54",X"45",X"52",X"20",
		X"4C",X"45",X"54",X"54",X"45",X"52",X"04",X"44",X"00",X"00",X"12",X"40",X"10",X"00",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"00",X"04",X"BB",X"0F",X"7B",X"BA",X"09",X"11",X"12",X"20",X"28",
		X"00",X"59",X"4F",X"55",X"20",X"48",X"41",X"56",X"45",X"20",X"4A",X"55",X"53",X"54",X"20",X"43",
		X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"44",X"20",X"54",X"48",X"45",X"12",X"25",X"38",X"00",
		X"47",X"52",X"45",X"41",X"54",X"45",X"53",X"54",X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",
		X"45",X"20",X"4D",X"49",X"53",X"53",X"49",X"4F",X"4E",X"12",X"36",X"58",X"00",X"45",X"4E",X"54",
		X"45",X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"4E",X"41",X"4D",X"45",X"12",X"34",X"68",X"00",
		X"5B",X"55",X"50",X"20",X"54",X"4F",X"20",X"09",X"10",X"20",X"4C",X"45",X"54",X"54",X"45",X"52",
		X"53",X"5C",X"0F",X"7B",X"8A",X"00",X"04",X"44",X"0F",X"7B",X"BA",X"09",X"10",X"12",X"21",X"2C",
		X"00",X"59",X"4F",X"55",X"20",X"48",X"41",X"56",X"45",X"20",X"45",X"4E",X"54",X"45",X"52",X"45",
		X"44",X"20",X"54",X"48",X"45",X"20",X"52",X"45",X"41",X"4C",X"4D",X"12",X"23",X"38",X"01",X"4F",
		X"46",X"20",X"54",X"48",X"45",X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"49",
		X"4D",X"4D",X"4F",X"52",X"54",X"41",X"4C",X"53",X"12",X"2D",X"58",X"00",X"45",X"4E",X"54",X"45",
		X"52",X"20",X"59",X"4F",X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"3F",
		X"0F",X"7B",X"8A",X"00",X"04",X"99",X"0F",X"7B",X"BA",X"09",X"10",X"12",X"45",X"64",X"00",X"41",
		X"4C",X"53",X"4F",X"0F",X"7C",X"78",X"00",X"04",X"11",X"12",X"3D",X"3A",X"00",X"49",X"4D",X"4D",
		X"4F",X"52",X"54",X"41",X"4C",X"53",X"12",X"40",X"C0",X"00",X"4D",X"4F",X"52",X"54",X"41",X"4C",
		X"53",X"00",X"15",X"10",X"5C",X"3A",X"3A",X"00",X"15",X"11",X"00",X"05",X"08",X"00",X"00",X"15",
		X"11",X"00",X"15",X"10",X"30",X"30",X"30",X"00",X"15",X"10",X"30",X"30",X"30",X"20",X"20",X"0F",
		X"7C",X"E8",X"00",X"05",X"08",X"00",X"00",X"00",X"52",X"45",X"43",X"4F",X"4D",X"4D",X"45",X"4E",
		X"44",X"45",X"44",X"00",X"0F",X"7C",X"E3",X"0F",X"7C",X"E8",X"00",X"15",X"10",X"00",X"0F",X"7D",
		X"6A",X"48",X"49",X"47",X"48",X"20",X"56",X"4F",X"4C",X"55",X"4D",X"45",X"20",X"41",X"52",X"43",
		X"41",X"44",X"45",X"53",X"00",X"15",X"10",X"0F",X"7C",X"F4",X"00",X"0F",X"7D",X"6A",X"46",X"4F",
		X"52",X"20",X"57",X"45",X"41",X"4B",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",
		X"00",X"0F",X"7D",X"6A",X"43",X"55",X"53",X"54",X"4F",X"4D",X"20",X"40",X"3A",X"5B",X"41",X"44",
		X"4A",X"55",X"53",X"54",X"20",X"42",X"45",X"4C",X"4F",X"57",X"5C",X"00",X"59",X"45",X"53",X"0F",
		X"7C",X"E3",X"05",X"FE",X"00",X"00",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",
		X"20",X"41",X"43",X"54",X"49",X"56",X"41",X"54",X"45",X"00",X"15",X"10",X"0F",X"7C",X"E3",X"00",
		X"59",X"45",X"53",X"00",X"4E",X"4F",X"00",X"0F",X"7D",X"7E",X"0F",X"7D",X"88",X"00",X"0F",X"7D",
		X"6A",X"45",X"58",X"54",X"52",X"41",X"20",X"00",X"4C",X"49",X"42",X"45",X"52",X"41",X"4C",X"00",
		X"0F",X"7D",X"6A",X"0F",X"7D",X"88",X"00",X"0F",X"7D",X"6A",X"4D",X"4F",X"44",X"45",X"52",X"41",
		X"54",X"45",X"00",X"0F",X"7D",X"6A",X"0F",X"7D",X"AA",X"00",X"43",X"4F",X"4E",X"53",X"45",X"52",
		X"56",X"41",X"54",X"49",X"56",X"45",X"00",X"0F",X"7D",X"7E",X"0F",X"7D",X"AA",X"00",X"0F",X"7D",
		X"6A",X"4E",X"4F",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"53",X"48",X"49",X"50",X"53",X"00",
		X"0F",X"7D",X"6A",X"31",X"5E",X"46",X"49",X"46",X"54",X"59",X"20",X"20",X"33",X"5E",X"44",X"4F",
		X"4C",X"4C",X"41",X"52",X"00",X"0F",X"7D",X"6A",X"31",X"5E",X"31",X"20",X"44",X"4D",X"20",X"20",
		X"36",X"5E",X"35",X"20",X"44",X"4D",X"00",X"0F",X"7D",X"6A",X"31",X"5E",X"51",X"55",X"41",X"52",
		X"54",X"45",X"52",X"20",X"20",X"34",X"5E",X"44",X"4F",X"4C",X"4C",X"41",X"52",X"00",X"0F",X"7D",
		X"6A",X"31",X"5E",X"32",X"20",X"46",X"20",X"20",X"33",X"5E",X"35",X"20",X"46",X"00",X"0F",X"7D",
		X"6A",X"31",X"5E",X"46",X"49",X"46",X"54",X"59",X"20",X"20",X"32",X"5E",X"44",X"4F",X"4C",X"4C",
		X"41",X"52",X"00",X"0F",X"7D",X"6A",X"31",X"5E",X"32",X"35",X"20",X"20",X"34",X"5E",X"31",X"20",
		X"47",X"00",X"0F",X"7D",X"6A",X"31",X"5E",X"35",X"20",X"46",X"20",X"20",X"32",X"5E",X"31",X"30",
		X"20",X"46",X"00",X"0F",X"7D",X"6A",X"31",X"5E",X"31",X"30",X"20",X"46",X"00",X"0F",X"7D",X"6A",
		X"4E",X"4F",X"20",X"32",X"0F",X"7F",X"E2",X"00",X"04",X"22",X"12",X"30",X"80",X"00",X"41",X"44",
		X"4A",X"55",X"53",X"54",X"4D",X"45",X"4E",X"54",X"20",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",
		X"12",X"20",X"A0",X"00",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"0F",X"7E",X"BA",X"42",X"59",
		X"12",X"20",X"B0",X"00",X"0F",X"7E",X"E0",X"14",X"7E",X"F3",X"12",X"20",X"C0",X"00",X"41",X"4E",
		X"44",X"20",X"54",X"55",X"52",X"4E",X"49",X"4E",X"47",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",
		X"46",X"46",X"20",X"41",X"4E",X"44",X"20",X"4F",X"4E",X"00",X"20",X"46",X"41",X"43",X"54",X"4F",
		X"52",X"59",X"20",X"53",X"45",X"54",X"54",X"49",X"4E",X"47",X"53",X"20",X"00",X"04",X"99",X"12",
		X"21",X"80",X"00",X"0F",X"7E",X"BA",X"20",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"44",X"00",
		X"4F",X"50",X"45",X"4E",X"49",X"4E",X"47",X"20",X"46",X"52",X"4F",X"4E",X"54",X"20",X"44",X"4F",
		X"4F",X"52",X"00",X"12",X"20",X"B0",X"00",X"04",X"00",X"0F",X"7E",X"E0",X"12",X"20",X"B0",X"00",
		X"04",X"22",X"52",X"41",X"49",X"53",X"49",X"4E",X"47",X"20",X"54",X"41",X"42",X"4C",X"45",X"20",
		X"54",X"4F",X"50",X"00",X"04",X"99",X"5D",X"04",X"88",X"00",X"07",X"04",X"99",X"12",X"37",X"10",
		X"00",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"4D",X"45",X"4E",X"54",
		X"08",X"12",X"2D",X"C4",X"00",X"04",X"BB",X"0F",X"7F",X"A1",X"41",X"44",X"4A",X"55",X"53",X"54",
		X"4D",X"45",X"4E",X"54",X"12",X"2D",X"CE",X"00",X"55",X"53",X"45",X"20",X"54",X"48",X"52",X"55",
		X"53",X"54",X"20",X"41",X"4E",X"44",X"20",X"46",X"49",X"52",X"45",X"20",X"54",X"4F",X"20",X"43",
		X"48",X"41",X"4E",X"47",X"45",X"20",X"54",X"48",X"45",X"20",X"56",X"41",X"4C",X"55",X"45",X"12",
		X"11",X"B3",X"00",X"04",X"88",X"4D",X"4F",X"52",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",
		X"4D",X"45",X"4E",X"54",X"53",X"12",X"3D",X"DE",X"00",X"04",X"33",X"50",X"52",X"45",X"53",X"53",
		X"20",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",X"20",X"45",X"58",X"49",X"54",
		X"00",X"55",X"53",X"45",X"20",X"55",X"50",X"40",X"44",X"4F",X"57",X"4E",X"20",X"4C",X"45",X"56",
		X"45",X"52",X"20",X"54",X"4F",X"20",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"00",X"45",X"58",
		X"54",X"52",X"41",X"20",X"53",X"48",X"49",X"50",X"20",X"45",X"56",X"45",X"52",X"59",X"00",X"0F",
		X"7F",X"D7",X"31",X"0F",X"7F",X"E2",X"00",X"53",X"48",X"49",X"50",X"53",X"20",X"46",X"4F",X"52",
		X"20",X"00",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"47",X"41",X"4D",X"45",X"00",X"0F",
		X"7F",X"D7",X"32",X"0F",X"7F",X"E2",X"00",X"50",X"52",X"49",X"43",X"49",X"4E",X"47",X"20",X"53",
		X"45",X"4C",X"45",X"43",X"54",X"49",X"4F",X"4E",X"00",X"4C",X"45",X"46",X"54",X"0F",X"80",X"24",
		X"00",X"43",X"45",X"4E",X"54",X"45",X"52",X"0F",X"80",X"24",X"00",X"52",X"49",X"47",X"48",X"54",
		X"0F",X"80",X"24",X"00",X"20",X"53",X"4C",X"4F",X"54",X"20",X"55",X"4E",X"49",X"54",X"53",X"00",
		X"0F",X"80",X"67",X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"0F",X"80",X"67",X"42",X"4F",X"4E",
		X"55",X"53",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"4D",X"49",X"4E",X"49",X"4D",X"55",
		X"4D",X"20",X"55",X"4E",X"49",X"54",X"53",X"20",X"46",X"4F",X"52",X"20",X"41",X"4E",X"59",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"55",X"4E",X"49",X"54",X"53",X"20",X"52",X"45",X"51",
		X"55",X"49",X"52",X"45",X"44",X"20",X"46",X"4F",X"52",X"20",X"00",X"46",X"52",X"45",X"45",X"20",
		X"50",X"4C",X"41",X"59",X"00",X"4D",X"41",X"53",X"54",X"45",X"52",X"0F",X"80",X"96",X"43",X"4F",
		X"4E",X"54",X"52",X"4F",X"4C",X"00",X"20",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",X"54",
		X"59",X"20",X"00",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"0F",X"80",X"96",X"00",X"4D",X"41",
		X"58",X"49",X"4D",X"55",X"4D",X"0F",X"80",X"96",X"00",X"31",X"53",X"54",X"0F",X"80",X"C8",X"00",
		X"4C",X"41",X"53",X"54",X"0F",X"80",X"C8",X"00",X"20",X"57",X"41",X"56",X"45",X"20",X"4F",X"46",
		X"20",X"41",X"43",X"43",X"45",X"4C",X"45",X"52",X"41",X"54",X"45",X"44",X"20",X"44",X"49",X"46",
		X"46",X"49",X"43",X"55",X"4C",X"54",X"59",X"00",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",
		X"54",X"59",X"20",X"41",X"43",X"43",X"45",X"4C",X"45",X"52",X"41",X"54",X"49",X"4F",X"4E",X"20",
		X"52",X"41",X"54",X"45",X"00",X"49",X"4E",X"56",X"49",X"53",X"4F",X"20",X"54",X"49",X"4D",X"45",
		X"20",X"50",X"45",X"52",X"20",X"53",X"48",X"49",X"50",X"00",X"4D",X"45",X"4E",X"20",X"4E",X"45",
		X"45",X"44",X"45",X"44",X"20",X"54",X"4F",X"20",X"57",X"41",X"52",X"50",X"00",X"4C",X"41",X"53",
		X"54",X"20",X"57",X"41",X"56",X"45",X"20",X"57",X"41",X"52",X"50",X"20",X"41",X"4C",X"4C",X"4F",
		X"57",X"45",X"44",X"00",X"4C",X"45",X"54",X"54",X"45",X"52",X"53",X"20",X"46",X"4F",X"52",X"0F",
		X"81",X"53",X"00",X"20",X"48",X"49",X"47",X"48",X"45",X"53",X"54",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"20",X"4E",X"41",X"4D",X"45",X"00",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"0F",X"7E",
		X"BA",X"00",X"43",X"4C",X"45",X"41",X"52",X"0F",X"82",X"04",X"00",X"52",X"45",X"53",X"45",X"54",
		X"20",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"54",X"41",X"42",X"4C",
		X"45",X"00",X"41",X"55",X"54",X"4F",X"20",X"43",X"59",X"43",X"4C",X"45",X"00",X"53",X"45",X"54",
		X"20",X"41",X"54",X"54",X"52",X"41",X"43",X"54",X"20",X"4D",X"4F",X"44",X"45",X"20",X"4D",X"45",
		X"53",X"53",X"41",X"47",X"45",X"00",X"53",X"45",X"54",X"0F",X"81",X"53",X"00",X"15",X"10",X"00",
		X"0A",X"11",X"00",X"05",X"06",X"00",X"00",X"15",X"11",X"00",X"12",X"2F",X"10",X"00",X"04",X"99",
		X"0F",X"82",X"04",X"04",X"88",X"00",X"12",X"20",X"60",X"00",X"04",X"33",X"0F",X"82",X"04",X"43",
		X"4C",X"45",X"41",X"52",X"45",X"44",X"00",X"12",X"2A",X"40",X"00",X"04",X"88",X"48",X"49",X"47",
		X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",X"54",X"41",X"42",X"4C",X"45",X"20",X"52",X"45",
		X"53",X"45",X"54",X"00",X"20",X"42",X"4F",X"4F",X"4B",X"4B",X"45",X"45",X"50",X"49",X"4E",X"47",
		X"20",X"54",X"4F",X"54",X"41",X"4C",X"53",X"20",X"00",X"12",X"1C",X"60",X"00",X"50",X"41",X"49",
		X"44",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"12",X"6C",X"60",X"00",X"00",X"12",X"1C",
		X"70",X"00",X"45",X"58",X"54",X"52",X"41",X"20",X"53",X"48",X"49",X"50",X"53",X"12",X"6C",X"70",
		X"00",X"00",X"12",X"1C",X"80",X"00",X"50",X"4C",X"41",X"59",X"20",X"54",X"49",X"4D",X"45",X"20",
		X"49",X"4E",X"20",X"4D",X"49",X"4E",X"55",X"54",X"45",X"53",X"12",X"6C",X"80",X"00",X"00",X"12",
		X"1C",X"90",X"00",X"53",X"48",X"49",X"50",X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"44",X"12",
		X"6C",X"90",X"00",X"00",X"12",X"1C",X"A0",X"00",X"54",X"4F",X"54",X"41",X"4C",X"20",X"50",X"4C",
		X"41",X"59",X"53",X"12",X"6C",X"A0",X"00",X"00",X"12",X"1C",X"B0",X"00",X"57",X"41",X"52",X"50",
		X"53",X"12",X"6C",X"B0",X"00",X"00",X"12",X"1C",X"30",X"00",X"4C",X"45",X"46",X"54",X"0F",X"82",
		X"C9",X"12",X"6C",X"30",X"00",X"00",X"12",X"1C",X"40",X"00",X"43",X"45",X"4E",X"54",X"45",X"52",
		X"0F",X"82",X"C9",X"12",X"6C",X"40",X"00",X"00",X"12",X"1C",X"50",X"00",X"52",X"49",X"47",X"48",
		X"54",X"0F",X"82",X"C9",X"12",X"6C",X"50",X"00",X"00",X"20",X"53",X"4C",X"4F",X"54",X"20",X"43",
		X"4F",X"49",X"4E",X"53",X"00",X"04",X"33",X"12",X"3A",X"80",X"00",X"43",X"4F",X"4C",X"4F",X"52",
		X"20",X"52",X"41",X"4D",X"20",X"54",X"45",X"53",X"54",X"12",X"24",X"B0",X"00",X"56",X"45",X"52",
		X"54",X"49",X"43",X"41",X"4C",X"20",X"42",X"41",X"52",X"53",X"20",X"49",X"4E",X"44",X"49",X"43",
		X"41",X"54",X"45",X"20",X"45",X"52",X"52",X"4F",X"52",X"00",X"41",X"55",X"54",X"4F",X"20",X"55",
		X"50",X"00",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"00",X"52",X"49",X"47",X"48",X"54",X"20",
		X"43",X"4F",X"49",X"4E",X"00",X"48",X"49",X"47",X"48",X"20",X"53",X"43",X"4F",X"52",X"45",X"20",
		X"52",X"45",X"53",X"45",X"54",X"00",X"4C",X"45",X"46",X"54",X"20",X"43",X"4F",X"49",X"4E",X"00",
		X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",X"00",X"53",X"4C",X"41",X"4D",
		X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"00",X"46",X"49",X"52",X"45",X"14",X"83",X"C1",X"00",
		X"54",X"48",X"52",X"55",X"53",X"54",X"14",X"83",X"C1",X"00",X"53",X"4D",X"41",X"52",X"54",X"20",
		X"42",X"4F",X"4D",X"42",X"14",X"83",X"C1",X"00",X"48",X"59",X"50",X"45",X"52",X"53",X"50",X"41",
		X"43",X"45",X"14",X"83",X"C1",X"00",X"32",X"0F",X"83",X"90",X"00",X"31",X"0F",X"83",X"90",X"00",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"00",X"52",X"45",
		X"56",X"45",X"52",X"53",X"45",X"14",X"83",X"C1",X"00",X"44",X"4F",X"57",X"4E",X"14",X"83",X"C1",
		X"00",X"55",X"50",X"14",X"83",X"C1",X"00",X"49",X"4E",X"56",X"49",X"53",X"4F",X"14",X"83",X"C1",
		X"00",X"20",X"20",X"5B",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"09",X"10",X"5C",X"00",X"04",
		X"88",X"12",X"3A",X"1A",X"00",X"53",X"57",X"49",X"54",X"43",X"48",X"20",X"54",X"45",X"53",X"54",
		X"00",X"04",X"99",X"12",X"3E",X"50",X"00",X"41",X"4C",X"4C",X"20",X"52",X"4F",X"4D",X"53",X"20",
		X"4F",X"4B",X"12",X"36",X"90",X"00",X"04",X"33",X"52",X"41",X"4D",X"20",X"54",X"45",X"53",X"54",
		X"20",X"46",X"4F",X"4C",X"4C",X"4F",X"57",X"53",X"12",X"2E",X"A0",X"00",X"50",X"52",X"45",X"53",
		X"53",X"20",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"20",X"54",X"4F",X"20",X"45",X"58",X"49",
		X"54",X"00",X"20",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"53",X"20",X"44",X"45",
		X"54",X"45",X"43",X"54",X"45",X"44",X"00",X"04",X"99",X"12",X"2A",X"80",X"00",X"4E",X"4F",X"0F",
		X"84",X"22",X"00",X"04",X"99",X"12",X"21",X"80",X"00",X"4E",X"4F",X"20",X"43",X"4D",X"4F",X"53",
		X"0F",X"84",X"22",X"00",X"43",X"4D",X"4F",X"53",X"20",X"52",X"41",X"4D",X"0F",X"89",X"E3",X"00",
		X"04",X"22",X"12",X"36",X"80",X"00",X"0F",X"84",X"54",X"00",X"0F",X"84",X"60",X"12",X"28",X"90",
		X"00",X"4F",X"52",X"20",X"57",X"52",X"49",X"54",X"45",X"20",X"50",X"52",X"4F",X"54",X"45",X"43",
		X"54",X"20",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",X"04",X"99",X"0F",X"84",X"C1",X"14",X"84",
		X"92",X"00",X"04",X"00",X"0F",X"84",X"C1",X"04",X"99",X"12",X"17",X"B0",X"00",X"40",X"54",X"41",
		X"42",X"4C",X"45",X"20",X"54",X"4F",X"50",X"20",X"4D",X"55",X"53",X"54",X"20",X"42",X"45",X"20",
		X"52",X"41",X"49",X"53",X"45",X"44",X"20",X"46",X"4F",X"52",X"20",X"54",X"45",X"53",X"54",X"40",
		X"00",X"12",X"18",X"B0",X"00",X"40",X"46",X"52",X"4F",X"4E",X"54",X"20",X"44",X"4F",X"4F",X"52",
		X"20",X"4D",X"55",X"53",X"54",X"20",X"42",X"45",X"20",X"4F",X"50",X"45",X"4E",X"20",X"46",X"4F",
		X"52",X"20",X"54",X"45",X"53",X"54",X"40",X"00",X"04",X"99",X"12",X"3A",X"80",X"00",X"53",X"4F",
		X"55",X"4E",X"44",X"20",X"4C",X"49",X"4E",X"45",X"20",X"09",X"10",X"00",X"04",X"DD",X"46",X"49",
		X"52",X"45",X"42",X"4F",X"4D",X"42",X"45",X"52",X"40",X"32",X"35",X"30",X"20",X"20",X"20",X"46",
		X"49",X"52",X"45",X"42",X"41",X"4C",X"4C",X"40",X"31",X"30",X"30",X"00",X"04",X"FF",X"59",X"4C",
		X"4C",X"41",X"42",X"49",X"41",X"4E",X"20",X"53",X"50",X"41",X"43",X"45",X"20",X"47",X"55",X"50",
		X"50",X"59",X"40",X"32",X"30",X"30",X"00",X"04",X"88",X"50",X"48",X"52",X"45",X"44",X"40",X"32",
		X"30",X"30",X"04",X"FF",X"20",X"42",X"49",X"47",X"20",X"52",X"45",X"44",X"40",X"32",X"30",X"30",
		X"04",X"33",X"20",X"4D",X"55",X"4E",X"43",X"48",X"49",X"45",X"53",X"40",X"35",X"30",X"00",X"04",
		X"99",X"44",X"59",X"4E",X"41",X"4D",X"4F",X"40",X"32",X"30",X"30",X"20",X"20",X"20",X"53",X"50",
		X"41",X"43",X"45",X"20",X"48",X"55",X"4D",X"40",X"31",X"30",X"30",X"00",X"04",X"DD",X"42",X"4F",
		X"4D",X"42",X"45",X"52",X"40",X"32",X"35",X"30",X"00",X"04",X"33",X"42",X"41",X"49",X"54",X"45",
		X"52",X"40",X"32",X"30",X"30",X"00",X"04",X"22",X"50",X"4F",X"44",X"40",X"31",X"30",X"30",X"30",
		X"20",X"20",X"20",X"53",X"57",X"41",X"52",X"4D",X"45",X"52",X"40",X"31",X"35",X"30",X"00",X"04",
		X"44",X"4C",X"41",X"4E",X"44",X"45",X"52",X"40",X"31",X"35",X"30",X"00",X"04",X"CC",X"4D",X"55",
		X"54",X"41",X"4E",X"54",X"40",X"31",X"35",X"30",X"00",X"04",X"AA",X"07",X"53",X"54",X"41",X"52",
		X"47",X"41",X"54",X"45",X"20",X"20",X"20",X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",X"00",X"04",
		X"AA",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"31",X"00",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"3D",X"00",X"04",X"11",X"43",X"52",X"45",X"44",
		X"49",X"54",X"53",X"3F",X"3A",X"09",X"10",X"00",X"04",X"88",X"48",X"49",X"47",X"48",X"20",X"53",
		X"43",X"4F",X"52",X"45",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"3F",X"50",X"52",X"45",
		X"53",X"53",X"20",X"48",X"59",X"50",X"45",X"52",X"53",X"50",X"41",X"43",X"45",X"00",X"47",X"41",
		X"4D",X"45",X"20",X"53",X"45",X"43",X"52",X"45",X"54",X"53",X"3F",X"50",X"52",X"45",X"53",X"53",
		X"20",X"52",X"45",X"56",X"45",X"52",X"53",X"45",X"00",X"04",X"AA",X"09",X"10",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"53",X"54",X"41",X"52",X"54",X"00",X"04",X"FF",X"09",X"10",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"47",X"41",X"4D",X"45",X"00",X"04",X"11",X"09",X"10",
		X"20",X"53",X"48",X"49",X"50",X"53",X"00",X"10",X"20",X"53",X"4D",X"41",X"52",X"54",X"20",X"42",
		X"4F",X"4D",X"42",X"53",X"00",X"10",X"20",X"49",X"4E",X"56",X"49",X"53",X"4F",X"20",X"55",X"4E",
		X"49",X"54",X"53",X"00",X"04",X"AA",X"09",X"45",X"58",X"54",X"52",X"41",X"20",X"53",X"48",X"49",
		X"50",X"3C",X"20",X"53",X"4D",X"41",X"52",X"54",X"20",X"42",X"4F",X"4D",X"42",X"3C",X"20",X"49",
		X"4E",X"56",X"49",X"53",X"4F",X"20",X"54",X"49",X"4D",X"45",X"20",X"41",X"57",X"41",X"52",X"44",
		X"45",X"44",X"20",X"45",X"56",X"45",X"52",X"59",X"20",X"10",X"30",X"30",X"30",X"20",X"50",X"4F",
		X"49",X"4E",X"54",X"53",X"00",X"04",X"88",X"53",X"04",X"77",X"45",X"04",X"66",X"43",X"04",X"55",
		X"52",X"04",X"44",X"45",X"04",X"33",X"54",X"04",X"22",X"53",X"00",X"04",X"88",X"12",X"10",X"55",
		X"00",X"57",X"41",X"52",X"50",X"3F",X"08",X"20",X"52",X"45",X"53",X"43",X"55",X"45",X"20",X"09",
		X"11",X"20",X"48",X"55",X"4D",X"41",X"4E",X"4F",X"49",X"44",X"53",X"20",X"41",X"4E",X"44",X"20",
		X"43",X"41",X"52",X"52",X"59",X"20",X"54",X"48",X"45",X"4D",X"20",X"49",X"4E",X"54",X"4F",X"20",
		X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"12",X"22",X"5D",X"00",X"57",X"41",X"52",X"50",
		X"20",X"4E",X"4F",X"54",X"20",X"41",X"4C",X"4C",X"4F",X"57",X"45",X"44",X"20",X"41",X"46",X"54",
		X"45",X"52",X"20",X"57",X"41",X"56",X"45",X"20",X"10",X"12",X"22",X"63",X"00",X"46",X"4C",X"59",
		X"49",X"4E",X"47",X"20",X"42",X"41",X"43",X"4B",X"57",X"41",X"52",X"44",X"53",X"20",X"49",X"4E",
		X"54",X"4F",X"20",X"53",X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"49",X"4E",X"48",X"49",
		X"42",X"49",X"54",X"53",X"20",X"57",X"41",X"52",X"50",X"04",X"77",X"07",X"12",X"10",X"6F",X"00",
		X"49",X"4E",X"56",X"49",X"53",X"4F",X"3F",X"08",X"41",X"43",X"54",X"49",X"56",X"41",X"54",X"45",
		X"20",X"49",X"4E",X"56",X"49",X"53",X"4F",X"20",X"41",X"4E",X"54",X"49",X"4D",X"41",X"54",X"54",
		X"45",X"52",X"20",X"43",X"4C",X"4F",X"41",X"4B",X"49",X"4E",X"47",X"20",X"44",X"45",X"56",X"49",
		X"43",X"45",X"20",X"54",X"4F",X"20",X"44",X"49",X"53",X"41",X"50",X"50",X"45",X"41",X"52",X"12",
		X"24",X"77",X"00",X"41",X"4E",X"44",X"20",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"20",X"45",
		X"56",X"45",X"52",X"59",X"54",X"48",X"49",X"4E",X"47",X"20",X"49",X"4E",X"20",X"59",X"4F",X"55",
		X"52",X"20",X"50",X"41",X"54",X"48",X"12",X"23",X"7D",X"00",X"20",X"52",X"45",X"44",X"20",X"4C",
		X"49",X"4E",X"45",X"20",X"42",X"45",X"4C",X"4F",X"57",X"20",X"53",X"4D",X"41",X"52",X"54",X"20",
		X"42",X"4F",X"4D",X"42",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"20",X"53",X"48",X"4F",
		X"57",X"53",X"20",X"49",X"4E",X"56",X"49",X"53",X"4F",X"20",X"54",X"49",X"4D",X"45",X"20",X"4C",
		X"45",X"46",X"54",X"07",X"12",X"10",X"89",X"00",X"04",X"66",X"53",X"54",X"41",X"52",X"47",X"41",
		X"54",X"45",X"3F",X"12",X"3F",X"89",X"00",X"08",X"54",X"52",X"41",X"4E",X"53",X"50",X"4F",X"52",
		X"54",X"53",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"54",X"4F",X"20",X"48",X"55",X"4D",
		X"41",X"4E",X"4F",X"49",X"44",X"53",X"20",X"42",X"45",X"49",X"4E",X"47",X"12",X"3F",X"91",X"00",
		X"41",X"42",X"44",X"55",X"43",X"54",X"45",X"44",X"3D",X"3A",X"3A",X"4F",X"54",X"48",X"45",X"52",
		X"57",X"49",X"53",X"45",X"20",X"54",X"52",X"41",X"4E",X"53",X"50",X"4F",X"52",X"54",X"53",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"12",X"3F",X"97",X"00",X"54",X"4F",X"20",X"4F",X"50",X"50",
		X"4F",X"53",X"49",X"54",X"45",X"20",X"53",X"49",X"44",X"45",X"20",X"4F",X"46",X"20",X"50",X"4C",
		X"41",X"4E",X"45",X"54",X"07",X"12",X"10",X"B7",X"00",X"04",X"44",X"53",X"4D",X"41",X"52",X"54",
		X"20",X"42",X"4F",X"4D",X"42",X"3F",X"08",X"20",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"53",
		X"20",X"41",X"4C",X"4C",X"20",X"45",X"4E",X"45",X"4D",X"49",X"45",X"53",X"20",X"4F",X"4E",X"20",
		X"53",X"43",X"52",X"45",X"45",X"4E",X"07",X"12",X"10",X"A3",X"00",X"04",X"55",X"48",X"55",X"4D",
		X"41",X"4E",X"4F",X"49",X"44",X"53",X"3F",X"12",X"32",X"A3",X"00",X"08",X"50",X"4C",X"41",X"4E",
		X"45",X"54",X"20",X"45",X"58",X"50",X"4C",X"4F",X"44",X"45",X"53",X"20",X"57",X"48",X"45",X"4E",
		X"20",X"41",X"4C",X"4C",X"20",X"48",X"55",X"4D",X"41",X"4E",X"4F",X"49",X"44",X"53",X"20",X"4C",
		X"4F",X"53",X"54",X"12",X"32",X"AB",X"00",X"48",X"55",X"4D",X"41",X"4E",X"4F",X"49",X"44",X"53",
		X"20",X"52",X"45",X"53",X"54",X"4F",X"52",X"45",X"44",X"20",X"41",X"46",X"54",X"45",X"52",X"20",
		X"45",X"56",X"45",X"52",X"59",X"20",X"35",X"54",X"48",X"20",X"57",X"41",X"56",X"45",X"00",X"5B",
		X"43",X"5C",X"20",X"31",X"39",X"38",X"31",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",
		X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",
		X"3D",X"00",X"12",X"30",X"70",X"00",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"20",X"54",X"45",
		X"53",X"54",X"53",X"20",X"49",X"4E",X"44",X"49",X"43",X"41",X"54",X"45",X"3F",X"00",X"04",X"99",
		X"0F",X"89",X"72",X"12",X"3A",X"90",X"00",X"41",X"4C",X"4C",X"20",X"53",X"59",X"53",X"54",X"45",
		X"4D",X"53",X"20",X"47",X"4F",X"00",X"04",X"22",X"0F",X"89",X"72",X"12",X"40",X"90",X"00",X"00",
		X"12",X"40",X"80",X"00",X"04",X"22",X"00",X"0F",X"89",X"B0",X"52",X"4F",X"4D",X"0F",X"89",X"E3",
		X"10",X"00",X"0F",X"89",X"B0",X"52",X"41",X"4D",X"0F",X"89",X"E3",X"10",X"00",X"0F",X"89",X"A6",
		X"52",X"4F",X"4D",X"0F",X"89",X"E3",X"10",X"00",X"0F",X"89",X"A6",X"52",X"41",X"4D",X"0F",X"89",
		X"E3",X"10",X"00",X"20",X"45",X"52",X"52",X"4F",X"52",X"20",X"09",X"00",X"12",X"3F",X"70",X"00",
		X"04",X"DD",X"09",X"20",X"57",X"41",X"56",X"45",X"20",X"10",X"3F",X"00",X"0F",X"89",X"EC",X"04",
		X"AA",X"12",X"32",X"88",X"00",X"59",X"4C",X"4C",X"41",X"42",X"49",X"41",X"4E",X"20",X"44",X"4F",
		X"47",X"46",X"49",X"47",X"48",X"54",X"00",X"0F",X"89",X"EC",X"04",X"CC",X"12",X"2E",X"88",X"00",
		X"46",X"49",X"52",X"45",X"42",X"4F",X"4D",X"42",X"45",X"52",X"20",X"53",X"48",X"4F",X"57",X"44",
		X"4F",X"57",X"4E",X"00",X"04",X"55",X"32",X"30",X"30",X"30",X"3B",X"00",X"04",X"FF",X"12",X"37",
		X"27",X"00",X"20",X"48",X"55",X"4D",X"41",X"4E",X"4F",X"49",X"44",X"53",X"20",X"52",X"45",X"4D",
		X"41",X"49",X"4E",X"49",X"4E",X"47",X"3F",X"3A",X"09",X"10",X"00",X"04",X"88",X"12",X"38",X"27",
		X"00",X"50",X"4F",X"44",X"20",X"49",X"4E",X"54",X"45",X"52",X"53",X"45",X"43",X"54",X"49",X"4F",
		X"4E",X"20",X"40",X"20",X"30",X"3F",X"00",X"04",X"88",X"12",X"5D",X"27",X"00",X"0A",X"10",X"00",
		X"13",X"9C",X"DE",X"12",X"40",X"27",X"00",X"3E",X"20",X"20",X"53",X"43",X"41",X"4E",X"4E",X"45",
		X"52",X"20",X"20",X"3E",X"00",X"04",X"55",X"12",X"36",X"27",X"00",X"50",X"4C",X"41",X"4E",X"45",
		X"54",X"20",X"53",X"55",X"52",X"46",X"41",X"43",X"45",X"20",X"55",X"4E",X"53",X"54",X"41",X"42",
		X"4C",X"45",X"3B",X"00",X"04",X"55",X"12",X"38",X"27",X"00",X"41",X"4C",X"4C",X"20",X"4C",X"41",
		X"4E",X"44",X"45",X"52",X"53",X"20",X"44",X"45",X"53",X"54",X"52",X"4F",X"59",X"45",X"44",X"3B",
		X"00",X"04",X"77",X"12",X"30",X"27",X"00",X"09",X"0F",X"8A",X"E2",X"10",X"0F",X"8A",X"F1",X"45",
		X"4E",X"00",X"57",X"41",X"52",X"50",X"20",X"52",X"45",X"51",X"55",X"49",X"52",X"45",X"53",X"20",
		X"00",X"20",X"41",X"44",X"44",X"49",X"54",X"49",X"4F",X"4E",X"41",X"4C",X"20",X"4D",X"00",X"04",
		X"77",X"12",X"30",X"27",X"00",X"0F",X"8A",X"E2",X"31",X"0F",X"8A",X"F1",X"41",X"4E",X"00",X"04",
		X"11",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"09",X"10",X"00",X"04",X"AA",X"47",X"41",X"4D",
		X"45",X"20",X"4F",X"56",X"45",X"52",X"00",X"04",X"99",X"12",X"34",X"50",X"00",X"3D",X"3D",X"3D",
		X"57",X"41",X"52",X"50",X"20",X"54",X"4F",X"20",X"57",X"41",X"56",X"45",X"20",X"09",X"10",X"00",
		X"04",X"11",X"12",X"36",X"50",X"00",X"41",X"54",X"54",X"41",X"43",X"4B",X"20",X"57",X"41",X"56",
		X"45",X"20",X"09",X"10",X"12",X"3C",X"60",X"00",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",
		X"44",X"00",X"04",X"FF",X"12",X"38",X"90",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",X"58",
		X"20",X"20",X"11",X"00",X"24",X"2F",X"20",X"54",X"48",X"49",X"53",X"20",X"49",X"53",X"20",X"53",
		X"54",X"41",X"52",X"47",X"41",X"54",X"45",X"20",X"24",X"24",X"2F",X"20",X"44",X"45",X"53",X"49",
		X"47",X"4E",X"45",X"44",X"20",X"45",X"58",X"43",X"4C",X"55",X"53",X"49",X"56",X"45",X"4C",X"59",
		X"20",X"46",X"4F",X"52",X"20",X"24",X"2F",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",
		X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",
		X"20",X"24",X"2F",X"20",X"42",X"59",X"20",X"45",X"55",X"47",X"45",X"4E",X"45",X"20",X"50",X"2E",
		X"20",X"4A",X"41",X"52",X"56",X"49",X"53",X"20",X"41",X"4E",X"44",X"20",X"4C",X"41",X"57",X"52",
		X"45",X"4E",X"43",X"45",X"20",X"45",X"2E",X"20",X"44",X"45",X"4D",X"41",X"52",X"20",X"24",X"24",
		X"2F",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"31",
		X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",
		X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"20",X"24",X"2F",X"20",X"41",X"4C",
		X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"35",X"10",X"AF",X"4D",X"A7",X"4B",X"86",X"07",X"A7",X"4C",X"A6",X"4B",X"8E",X"8F",X"12",X"7E",
		X"00",X"A8",X"8E",X"9C",X"27",X"10",X"8E",X"BC",X"72",X"A6",X"84",X"E6",X"84",X"84",X"07",X"97",
		X"4F",X"A6",X"A4",X"84",X"07",X"91",X"4F",X"23",X"01",X"5C",X"A6",X"84",X"84",X"38",X"97",X"4F",
		X"A6",X"A4",X"84",X"38",X"91",X"4F",X"23",X"02",X"CB",X"08",X"A6",X"4C",X"85",X"01",X"26",X"10",
		X"A6",X"84",X"84",X"C0",X"97",X"4F",X"A6",X"A4",X"84",X"C0",X"91",X"4F",X"23",X"02",X"CB",X"40",
		X"E7",X"80",X"31",X"21",X"8C",X"9C",X"36",X"26",X"C0",X"6A",X"4C",X"26",X"AD",X"6E",X"D8",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
