library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_arith.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM is
	port (
		ROM_nCS :in  std_logic := '1';
		ROM_nOE :in  std_logic := '1';
		ROM_A   :in  std_logic_vector (16 downto 0) := (others => '0'); -- Address input
		ROM_D   :out std_logic_vector ( 7 downto 0)  -- Data output
	);
end entity;

architecture behavioral of ROM is
	type mem is array (0 to 131071) of std_logic_vector(7 downto 0);
	constant my_rom : mem := (
		x"C3",x"77",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"5F",x"16",x"00",x"19",x"C9",x"FF",x"FF",
		x"DF",x"EB",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"5E",x"23",x"56",x"23",x"C9",x"FF",x"FF",x"FF",
		x"E1",x"CF",x"D7",x"E9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"6E",x"0C",x"DD",x"66",x"0D",x"7E",x"23",
		x"DD",x"75",x"0C",x"DD",x"74",x"0D",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"08",x"D9",x"21",x"90",x"43",x"CB",x"C6",x"3A",x"00",x"60",
		x"32",x"91",x"43",x"D9",x"08",x"ED",x"45",x"31",x"00",x"44",x"3A",x"00",x"60",x"21",x"00",x"40",
		x"01",x"00",x"04",x"36",x"00",x"23",x"0B",x"78",x"B1",x"20",x"F8",x"CD",x"9F",x"00",x"CD",x"37",
		x"01",x"CD",x"9B",x"04",x"21",x"90",x"43",x"CB",x"46",x"28",x"FC",x"CB",x"86",x"18",x"EC",x"3A",
		x"91",x"43",x"B7",x"C8",x"FE",x"10",x"30",x"09",x"3D",x"21",x"AF",x"00",x"CF",x"D7",x"E9",x"77",
		x"00",x"0E",x"00",x"D6",x"10",x"CB",x"7F",x"28",x"03",x"0C",x"E6",x"7F",x"21",x"B2",x"06",x"CF",
		x"D7",x"7E",x"23",x"FD",x"21",x"00",x"40",x"B7",x"28",x"04",x"FD",x"21",x"B0",x"41",x"0D",x"28",
		x"44",x"7E",x"FE",x"FF",x"C8",x"23",x"DF",x"E5",x"6F",x"26",x"00",x"29",x"29",x"29",x"29",x"4D",
		x"44",x"29",x"09",x"4D",x"44",x"FD",x"E5",x"DD",x"E1",x"DD",x"09",x"DD",x"36",x"00",x"80",x"DD",
		x"73",x"0C",x"DD",x"72",x"0D",x"21",x"02",x"06",x"DF",x"DD",x"73",x"10",x"DD",x"72",x"11",x"DD",
		x"36",x"01",x"03",x"DD",x"36",x"2C",x"40",x"DD",x"36",x"2D",x"00",x"DD",x"36",x"0A",x"00",x"CD",
		x"CF",x"01",x"E1",x"18",x"BC",x"7E",x"FE",x"FF",x"C8",x"23",x"23",x"23",x"E5",x"6F",x"26",x"00",
		x"29",x"29",x"29",x"29",x"5D",x"54",x"29",x"19",x"EB",x"FD",x"E5",x"E1",x"19",x"06",x"30",x"36",
		x"00",x"23",x"10",x"FB",x"E1",x"18",x"DE",x"06",x"12",x"DD",x"21",x"00",x"40",x"C5",x"3E",x"12",
		x"90",x"32",x"92",x"43",x"DD",x"CB",x"00",x"7E",x"C4",x"54",x"01",x"11",x"30",x"00",x"DD",x"19",
		x"C1",x"10",x"EA",x"C9",x"DD",x"6E",x"14",x"DD",x"66",x"15",x"2B",x"DD",x"75",x"14",x"DD",x"74",
		x"15",x"7C",x"B5",x"CC",x"CF",x"01",x"DD",x"CB",x"00",x"5E",x"28",x"09",x"DD",x"36",x"02",x"00",
		x"DD",x"36",x"03",x"00",x"C9",x"DD",x"CB",x"00",x"56",x"28",x"15",x"DD",x"6E",x"28",x"DD",x"66",
		x"29",x"2B",x"DD",x"75",x"28",x"DD",x"74",x"29",x"7C",x"B5",x"20",x"04",x"DD",x"CB",x"00",x"96",
		x"DD",x"6E",x"02",x"DD",x"66",x"03",x"DD",x"5E",x"04",x"DD",x"56",x"05",x"19",x"DD",x"75",x"02",
		x"DD",x"74",x"03",x"DD",x"6E",x"06",x"DD",x"66",x"07",x"DD",x"5E",x"08",x"DD",x"56",x"09",x"19",
		x"DD",x"75",x"06",x"DD",x"74",x"07",x"DD",x"CB",x"00",x"76",x"C0",x"DD",x"6E",x"0E",x"DD",x"66",
		x"0F",x"2B",x"DD",x"75",x"0E",x"DD",x"74",x"0F",x"7D",x"B4",x"C0",x"CD",x"D1",x"03",x"C9",x"DD",
		x"CB",x"00",x"76",x"C2",x"35",x"04",x"DD",x"36",x"08",x"00",x"DD",x"36",x"09",x"00",x"DD",x"7E",
		x"00",x"E6",x"E6",x"DD",x"77",x"00",x"DD",x"6E",x"06",x"DD",x"66",x"07",x"DD",x"75",x"16",x"DD",
		x"74",x"17",x"DD",x"6E",x"2E",x"DD",x"66",x"2F",x"DD",x"75",x"14",x"DD",x"74",x"15",x"FF",x"FE",
		x"80",x"30",x"59",x"DD",x"CB",x"00",x"46",x"28",x"10",x"DD",x"6E",x"0C",x"DD",x"66",x"0D",x"2B",
		x"DD",x"75",x"0C",x"DD",x"74",x"0D",x"C3",x"AE",x"02",x"DD",x"CB",x"00",x"C6",x"47",x"E6",x"0F",
		x"FE",x"0C",x"20",x"06",x"DD",x"CB",x"00",x"DE",x"18",x"D4",x"21",x"B0",x"05",x"CF",x"DF",x"CB",
		x"38",x"CB",x"38",x"CB",x"38",x"CB",x"38",x"DD",x"7E",x"01",x"CB",x"2F",x"CB",x"2F",x"80",x"28",
		x"13",x"47",x"FE",x"08",x"38",x"08",x"DD",x"CB",x"01",x"46",x"20",x"08",x"06",x"07",x"CB",x"3A",
		x"CB",x"1B",x"10",x"FA",x"DD",x"73",x"06",x"DD",x"72",x"07",x"18",x"A2",x"FE",x"F0",x"38",x"27",
		x"E6",x"0F",x"21",x"FE",x"01",x"E5",x"E7",x"08",x"03",x"0D",x"03",x"1A",x"03",x"28",x"03",x"38",
		x"03",x"46",x"03",x"56",x"03",x"6D",x"03",x"72",x"03",x"77",x"03",x"7C",x"03",x"87",x"03",x"9B",
		x"03",x"A4",x"03",x"AD",x"03",x"B5",x"03",x"E6",x"7F",x"21",x"E0",x"05",x"CF",x"DF",x"DD",x"6E",
		x"2C",x"DD",x"66",x"2D",x"CD",x"17",x"04",x"06",x"06",x"CB",x"3C",x"CB",x"1D",x"10",x"FA",x"DD",
		x"75",x"14",x"DD",x"74",x"15",x"DD",x"75",x"2E",x"DD",x"74",x"2F",x"C3",x"FE",x"01",x"DD",x"6E",
		x"10",x"DD",x"66",x"11",x"DF",x"DD",x"73",x"02",x"DD",x"72",x"03",x"DD",x"75",x"12",x"DD",x"74",
		x"13",x"CD",x"D1",x"03",x"DD",x"CB",x"00",x"66",x"20",x"05",x"DD",x"CB",x"00",x"6E",x"C8",x"DD",
		x"6E",x"06",x"DD",x"66",x"07",x"DD",x"5E",x"17",x"DD",x"56",x"18",x"DD",x"4E",x"14",x"DD",x"46",
		x"15",x"CD",x"EB",x"02",x"DD",x"75",x"08",x"DD",x"74",x"09",x"C9",x"B7",x"ED",x"52",x"30",x"08",
		x"EB",x"21",x"00",x"00",x"B7",x"ED",x"52",x"37",x"F5",x"59",x"50",x"CD",x"F8",x"03",x"F1",x"D0",
		x"EB",x"21",x"00",x"00",x"B7",x"ED",x"52",x"C9",x"FF",x"DD",x"77",x"01",x"C9",x"FF",x"21",x"02",
		x"06",x"CF",x"D7",x"DD",x"75",x"10",x"DD",x"74",x"11",x"C9",x"DD",x"6E",x"0C",x"DD",x"66",x"0D",
		x"DF",x"DD",x"73",x"0C",x"DD",x"72",x"0D",x"C9",x"CD",x"C1",x"03",x"E5",x"CD",x"1A",x"03",x"EB",
		x"E1",x"73",x"23",x"72",x"DD",x"34",x"0A",x"C9",x"DD",x"35",x"0A",x"CD",x"C1",x"03",x"DF",x"DD",
		x"73",x"0C",x"DD",x"72",x"0D",x"C9",x"FF",x"DD",x"77",x"0B",x"E5",x"CD",x"C1",x"03",x"D1",x"73",
		x"23",x"72",x"DD",x"34",x"0A",x"C9",x"DD",x"35",x"0A",x"DD",x"35",x"0B",x"20",x"01",x"C9",x"CD",
		x"C1",x"03",x"DD",x"34",x"0A",x"DF",x"DD",x"73",x"0C",x"DD",x"72",x"0D",x"C9",x"DD",x"CB",x"00",
		x"E6",x"C9",x"DD",x"CB",x"00",x"EE",x"C9",x"DD",x"CB",x"00",x"AE",x"C9",x"FF",x"87",x"47",x"DD",
		x"7E",x"01",x"B0",x"DD",x"77",x"01",x"C9",x"DD",x"6E",x"0C",x"DD",x"66",x"0D",x"DF",x"DD",x"75",
		x"0C",x"DD",x"74",x"0D",x"DD",x"73",x"2C",x"DD",x"72",x"2D",x"C9",x"DD",x"7E",x"01",x"E6",x"03",
		x"DD",x"77",x"01",x"C9",x"DD",x"36",x"2C",x"40",x"DD",x"36",x"2D",x"00",x"C9",x"DD",x"CB",x"00",
		x"F6",x"E1",x"C3",x"35",x"04",x"E1",x"DD",x"E5",x"E1",x"06",x"20",x"36",x"00",x"23",x"10",x"FB",
		x"C9",x"DD",x"E5",x"E1",x"11",x"18",x"00",x"19",x"DD",x"7E",x"0A",x"87",x"5F",x"16",x"00",x"19",
		x"C9",x"DD",x"6E",x"12",x"DD",x"66",x"13",x"DF",x"4B",x"42",x"DD",x"73",x"0E",x"DD",x"72",x"0F",
		x"DF",x"DD",x"75",x"12",x"DD",x"74",x"13",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"EB",x"CD",x"EB",
		x"02",x"DD",x"75",x"04",x"DD",x"74",x"05",x"C9",x"F5",x"C5",x"EB",x"4D",x"44",x"21",x"00",x"00",
		x"3E",x"10",x"EB",x"29",x"EB",x"ED",x"6A",x"B7",x"ED",x"42",x"30",x"03",x"09",x"18",x"01",x"13",
		x"3D",x"20",x"EF",x"EB",x"C1",x"F1",x"C9",x"F5",x"C5",x"D5",x"4D",x"44",x"21",x"00",x"00",x"7A",
		x"B3",x"28",x"0E",x"CB",x"38",x"CB",x"19",x"30",x"01",x"19",x"EB",x"29",x"EB",x"79",x"B0",x"20",
		x"F2",x"D1",x"C1",x"F1",x"C9",x"FF",x"CB",x"7F",x"28",x"07",x"DD",x"CB",x"00",x"B6",x"C3",x"CF",
		x"01",x"DD",x"6E",x"0C",x"DD",x"66",x"0D",x"DF",x"DD",x"75",x"0C",x"DD",x"74",x"0D",x"DD",x"73",
		x"14",x"DD",x"72",x"15",x"CB",x"47",x"28",x"07",x"DF",x"DD",x"73",x"06",x"DD",x"72",x"07",x"CB",
		x"4F",x"28",x"07",x"DF",x"DD",x"73",x"08",x"DD",x"72",x"09",x"CB",x"57",x"28",x"07",x"DF",x"DD",
		x"73",x"02",x"DD",x"72",x"03",x"CB",x"5F",x"28",x"07",x"DF",x"DD",x"73",x"04",x"DD",x"72",x"05",
		x"CB",x"67",x"28",x"10",x"7E",x"DD",x"77",x"2A",x"23",x"DF",x"DD",x"73",x"28",x"DD",x"72",x"29",
		x"DD",x"CB",x"00",x"D6",x"DD",x"75",x"0C",x"DD",x"74",x"0D",x"C9",x"DD",x"21",x"B0",x"41",x"FD",
		x"21",x"60",x"43",x"06",x"03",x"C5",x"DD",x"E5",x"CD",x"F6",x"04",x"FD",x"71",x"07",x"11",x"50",
		x"FE",x"DD",x"19",x"CD",x"F6",x"04",x"FD",x"7E",x"07",x"B1",x"2F",x"FD",x"77",x"07",x"DD",x"E1",
		x"C1",x"11",x"90",x"00",x"DD",x"19",x"11",x"10",x"00",x"FD",x"19",x"10",x"D8",x"21",x"60",x"43",
		x"0E",x"00",x"CD",x"E6",x"04",x"21",x"70",x"43",x"0E",x"10",x"CD",x"E6",x"04",x"21",x"80",x"43",
		x"0E",x"80",x"CD",x"E6",x"04",x"C9",x"06",x"10",x"3E",x"10",x"90",x"ED",x"79",x"0C",x"7E",x"23",
		x"ED",x"79",x"0D",x"10",x"F3",x"C9",x"0E",x"00",x"DD",x"CB",x"00",x"7E",x"28",x"25",x"CB",x"C1",
		x"11",x"00",x"00",x"CD",x"8F",x"05",x"FD",x"75",x"00",x"FD",x"74",x"01",x"FD",x"77",x"08",x"DD",
		x"7E",x"01",x"E6",x"03",x"47",x"DD",x"CB",x"00",x"56",x"28",x"08",x"CB",x"D9",x"DD",x"7E",x"2A",
		x"FD",x"77",x"06",x"DD",x"CB",x"30",x"7E",x"28",x"28",x"CB",x"C9",x"11",x"30",x"00",x"CD",x"8F",
		x"05",x"FD",x"75",x"02",x"FD",x"74",x"03",x"FD",x"77",x"09",x"DD",x"7E",x"31",x"87",x"87",x"E6",
		x"0C",x"B0",x"47",x"DD",x"CB",x"30",x"56",x"28",x"08",x"CB",x"E1",x"DD",x"7E",x"58",x"FD",x"77",
		x"06",x"DD",x"CB",x"60",x"7E",x"28",x"34",x"CB",x"D1",x"11",x"60",x"00",x"CD",x"8F",x"05",x"FD",
		x"75",x"04",x"FD",x"74",x"05",x"FD",x"77",x"0A",x"DD",x"7E",x"61",x"87",x"87",x"87",x"87",x"E6",
		x"30",x"B0",x"47",x"DD",x"CB",x"60",x"56",x"28",x"12",x"CB",x"E9",x"11",x"88",x"00",x"DD",x"19",
		x"DD",x"7E",x"00",x"11",x"78",x"FF",x"DD",x"19",x"FD",x"77",x"06",x"FD",x"70",x"0E",x"C9",x"C5",
		x"DD",x"19",x"21",x"00",x"00",x"B7",x"ED",x"52",x"EB",x"DD",x"7E",x"03",x"DD",x"6E",x"06",x"DD",
		x"66",x"07",x"DD",x"19",x"06",x"04",x"CB",x"3F",x"CB",x"3C",x"CB",x"1D",x"10",x"F8",x"C1",x"C9",
		x"2B",x"B3",x"1D",x"A9",x"9F",x"9F",x"A9",x"96",x"35",x"8E",x"39",x"86",x"B1",x"7E",x"95",x"77",
		x"DE",x"70",x"89",x"6A",x"8E",x"64",x"E9",x"5E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"00",x"02",x"00",x"04",x"00",x"06",x"00",x"08",x"00",x"0C",x"00",x"10",x"00",x"18",x"00",
		x"20",x"00",x"30",x"00",x"40",x"00",x"60",x"00",x"80",x"00",x"C0",x"00",x"00",x"01",x"80",x"01",
		x"00",x"02",x"18",x"06",x"26",x"06",x"34",x"06",x"42",x"06",x"50",x"06",x"5E",x"06",x"6C",x"06",
		x"7A",x"06",x"88",x"06",x"96",x"06",x"A4",x"06",x"FF",x"FF",x"02",x"00",x"FF",x"FF",x"08",x"00",
		x"00",x"80",x"0A",x"00",x"00",x"00",x"FF",x"FF",x"02",x"00",x"FF",x"FF",x"08",x"00",x"00",x"80",
		x"14",x"00",x"00",x"00",x"01",x"00",x"02",x"00",x"FF",x"FF",x"3C",x"00",x"FF",x"FF",x"80",x"00",
		x"01",x"00",x"FF",x"FF",x"01",x"00",x"FF",x"FF",x"F0",x"00",x"00",x"80",x"F0",x"00",x"01",x"00",
		x"01",x"00",x"0A",x"00",x"00",x"F0",x"0A",x"00",x"00",x"80",x"14",x"00",x"01",x"00",x"FF",x"FF",
		x"02",x"00",x"FF",x"FF",x"14",x"00",x"00",x"60",x"32",x"00",x"00",x"00",x"00",x"80",x"02",x"00",
		x"FF",x"FF",x"08",x"00",x"00",x"80",x"1E",x"00",x"00",x"00",x"FF",x"FF",x"02",x"00",x"FF",x"FF",
		x"3C",x"00",x"00",x"80",x"B0",x"00",x"00",x"00",x"FF",x"FF",x"02",x"00",x"FF",x"FF",x"1E",x"00",
		x"00",x"80",x"60",x"00",x"00",x"00",x"00",x"40",x"04",x"00",x"FF",x"FF",x"60",x"00",x"00",x"80",
		x"3C",x"00",x"00",x"00",x"00",x"50",x"04",x"00",x"FF",x"FF",x"B0",x"00",x"00",x"80",x"A0",x"00",
		x"00",x"50",x"F2",x"06",x"3A",x"07",x"F0",x"06",x"8A",x"07",x"BE",x"07",x"D1",x"07",x"F8",x"07",
		x"50",x"08",x"8C",x"08",x"B6",x"08",x"87",x"17",x"00",x"09",x"F0",x"06",x"A2",x"09",x"FA",x"09",
		x"1E",x"0A",x"02",x"0B",x"F0",x"06",x"82",x"0C",x"38",x"0D",x"D7",x"13",x"0E",x"16",x"D7",x"16",
		x"44",x"0A",x"4F",x"18",x"E7",x"1A",x"A9",x"19",x"4F",x"1D",x"92",x"0A",x"CA",x"0A",x"1E",x"1E",
		x"00",x"FF",x"00",x"07",x"FA",x"06",x"08",x"1A",x"07",x"FF",x"F0",x"03",x"F1",x"03",x"FA",x"01",
		x"FB",x"40",x"00",x"20",x"80",x"24",x"27",x"30",x"34",x"37",x"40",x"44",x"47",x"50",x"54",x"57",
		x"60",x"64",x"80",x"F1",x"08",x"69",x"80",x"70",x"88",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"01",
		x"FB",x"40",x"00",x"21",x"80",x"25",x"28",x"31",x"35",x"38",x"41",x"45",x"48",x"51",x"55",x"58",
		x"61",x"65",x"80",x"F1",x"08",x"6A",x"80",x"71",x"86",x"FF",x"00",x"05",x"42",x"07",x"06",x"66",
		x"07",x"FF",x"FE",x"0F",x"05",x"00",x"00",x"10",x"00",x"FE",x"FF",x"FF",x"00",x"FF",x"0F",x"05",
		x"00",x"00",x"09",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"0F",x"20",x"00",x"00",x"05",x"F0",x"FF",
		x"FF",x"FF",x"00",x"F9",x"80",x"FF",x"FE",x"0F",x"05",x"00",x"00",x"12",x"00",x"FF",x"FF",x"FF",
		x"00",x"F9",x"0F",x"05",x"00",x"00",x"0B",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"0F",x"20",x"00",
		x"00",x"07",x"F0",x"FF",x"FF",x"FF",x"DD",x"F9",x"80",x"FF",x"01",x"05",x"92",x"07",x"06",x"A8",
		x"07",x"FF",x"F0",x"03",x"F1",x"05",x"FA",x"01",x"FB",x"10",x"00",x"F8",x"60",x"86",x"0C",x"84",
		x"50",x"86",x"0C",x"84",x"F2",x"92",x"07",x"FF",x"F0",x"03",x"F1",x"05",x"FA",x"01",x"FB",x"10",
		x"00",x"F8",x"61",x"86",x"0C",x"84",x"51",x"86",x"0C",x"84",x"F2",x"B1",x"07",x"FF",x"00",x"05",
		x"C3",x"07",x"FF",x"F8",x"50",x"82",x"54",x"57",x"60",x"64",x"67",x"82",x"F1",x"03",x"69",x"90",
		x"FF",x"01",x"07",x"D9",x"07",x"08",x"EA",x"07",x"FF",x"FB",x"1F",x"10",x"00",x"00",x"10",x"00",
		x"00",x"FF",x"FF",x"00",x"10",x"15",x"10",x"00",x"80",x"FF",x"FE",x"0F",x"10",x"00",x"00",x"05",
		x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"FF",x"00",x"07",x"00",x"08",x"08",x"28",x"08",x"FF",
		x"F0",x"03",x"F1",x"0C",x"FA",x"01",x"FB",x"30",x"00",x"70",x"84",x"6B",x"60",x"5B",x"82",x"5A",
		x"59",x"58",x"57",x"56",x"55",x"54",x"53",x"52",x"51",x"50",x"4B",x"4A",x"49",x"48",x"47",x"46",
		x"45",x"44",x"43",x"42",x"41",x"40",x"82",x"FF",x"F0",x"03",x"F1",x"0C",x"FA",x"01",x"FB",x"30",
		x"00",x"6B",x"84",x"6A",x"6B",x"5A",x"82",x"59",x"58",x"57",x"56",x"55",x"54",x"53",x"52",x"51",
		x"50",x"4B",x"4A",x"49",x"48",x"47",x"46",x"45",x"44",x"43",x"42",x"41",x"40",x"3B",x"82",x"FF",
		x"01",x"07",x"58",x"08",x"08",x"7C",x"08",x"FF",x"FE",x"0F",x"03",x"00",x"00",x"25",x"FF",x"FF",
		x"FF",x"FF",x"00",x"F2",x"0F",x"03",x"00",x"00",x"20",x"FF",x"FF",x"FF",x"FF",x"00",x"F0",x"0F",
		x"20",x"00",x"00",x"20",x"FC",x"FF",x"FF",x"FF",x"00",x"FB",x"80",x"FF",x"FE",x"0F",x"0A",x"00",
		x"00",x"00",x"00",x"20",x"00",x"00",x"FF",x"FF",x"FF",x"F9",x"80",x"FF",x"00",x"05",x"94",x"08",
		x"06",x"A5",x"08",x"FF",x"F5",x"03",x"FE",x"0F",x"06",x"00",x"00",x"03",x"C0",x"FF",x"DD",x"DD",
		x"00",x"FF",x"80",x"F6",x"FF",x"F5",x"03",x"FE",x"0F",x"06",x"00",x"00",x"03",x"D0",x"FF",x"DD",
		x"DD",x"00",x"FF",x"80",x"F6",x"FF",x"00",x"05",x"BE",x"08",x"06",x"D1",x"08",x"FF",x"FE",x"0F",
		x"10",x"00",x"00",x"02",x"E0",x"FF",x"DD",x"DD",x"00",x"EF",x"F0",x"03",x"F1",x"00",x"71",x"85",
		x"FF",x"FE",x"0F",x"03",x"00",x"00",x"04",x"00",x"00",x"DD",x"DD",x"FF",x"E0",x"0F",x"03",x"00",
		x"00",x"03",x"00",x"00",x"FF",x"FF",x"FF",x"E0",x"0F",x"03",x"00",x"00",x"02",x"00",x"00",x"FF",
		x"FF",x"FF",x"E0",x"0F",x"05",x"00",x"00",x"03",x"00",x"00",x"FF",x"FF",x"FF",x"E0",x"80",x"FF",
		x"00",x"00",x"0E",x"09",x"01",x"4A",x"09",x"02",x"82",x"09",x"03",x"92",x"09",x"FF",x"F0",x"00",
		x"F1",x"02",x"FA",x"01",x"FB",x"20",x"00",x"40",x"82",x"41",x"42",x"43",x"44",x"45",x"46",x"47",
		x"48",x"49",x"4A",x"4B",x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5A",x"59",
		x"58",x"57",x"56",x"55",x"54",x"53",x"52",x"51",x"50",x"4B",x"4A",x"49",x"48",x"47",x"46",x"45",
		x"44",x"43",x"42",x"41",x"40",x"82",x"F2",x"0E",x"09",x"FF",x"F0",x"00",x"F1",x"03",x"FA",x"01",
		x"FB",x"20",x"00",x"60",x"82",x"61",x"63",x"64",x"65",x"66",x"67",x"68",x"69",x"6A",x"6B",x"70",
		x"71",x"72",x"73",x"74",x"75",x"76",x"77",x"79",x"7A",x"79",x"78",x"77",x"76",x"75",x"74",x"73",
		x"72",x"71",x"70",x"6B",x"6A",x"69",x"68",x"67",x"66",x"65",x"64",x"63",x"62",x"82",x"F2",x"4A",
		x"09",x"FF",x"FE",x"0F",x"09",x"00",x"00",x"03",x"E0",x"FF",x"DD",x"DD",x"FF",x"FF",x"80",x"F2",
		x"82",x"09",x"FE",x"0F",x"09",x"00",x"00",x"05",x"E0",x"FF",x"DD",x"DD",x"FF",x"FF",x"80",x"F2",
		x"92",x"09",x"00",x"07",x"B0",x"09",x"08",x"C1",x"09",x"04",x"D4",x"09",x"05",x"E7",x"09",x"FF",
		x"F1",x"08",x"FB",x"10",x"00",x"65",x"83",x"63",x"61",x"63",x"82",x"65",x"80",x"67",x"69",x"86",
		x"FF",x"F1",x"08",x"FB",x"10",x"00",x"61",x"83",x"5B",x"82",x"59",x"83",x"5B",x"82",x"61",x"81",
		x"63",x"65",x"86",x"FF",x"F1",x"08",x"FB",x"10",x"00",x"0C",x"88",x"65",x"83",x"63",x"61",x"63",
		x"82",x"65",x"81",x"67",x"69",x"86",x"FF",x"F1",x"08",x"FB",x"10",x"00",x"0C",x"88",x"61",x"83",
		x"5B",x"59",x"5B",x"82",x"61",x"81",x"63",x"65",x"86",x"FF",x"00",x"05",x"02",x"0A",x"06",x"10",
		x"0A",x"FF",x"FE",x"0F",x"10",x"00",x"00",x"05",x"C0",x"FF",x"FF",x"FF",x"00",x"00",x"80",x"FF",
		x"FE",x"0F",x"09",x"00",x"00",x"04",x"C0",x"FF",x"FF",x"FF",x"00",x"00",x"80",x"FF",x"00",x"04",
		x"26",x"0A",x"08",x"35",x"0A",x"FF",x"F1",x"01",x"FB",x"30",x"00",x"F8",x"60",x"86",x"70",x"88",
		x"69",x"85",x"67",x"83",x"FF",x"F1",x"02",x"FB",x"30",x"00",x"F8",x"50",x"86",x"60",x"88",x"70",
		x"85",x"71",x"83",x"FF",x"00",x"00",x"4C",x"0A",x"01",x"73",x"0A",x"FF",x"F5",x"02",x"F1",x"08",
		x"FB",x"15",x"00",x"57",x"84",x"54",x"56",x"82",x"58",x"59",x"5B",x"61",x"63",x"65",x"67",x"83",
		x"69",x"82",x"F6",x"FE",x"1F",x"80",x"00",x"00",x"03",x"FC",x"FF",x"FF",x"FF",x"FE",x"FF",x"10",
		x"80",x"00",x"FF",x"FE",x"1F",x"0B",x"00",x"00",x"04",x"C0",x"FF",x"FF",x"FF",x"F0",x"FF",x"08",
		x"10",x"00",x"1F",x"20",x"00",x"00",x"02",x"40",x"00",x"FF",x"FF",x"FF",x"FF",x"05",x"09",x"00",
		x"80",x"FF",x"00",x"07",x"9A",x"0A",x"08",x"B9",x"0A",x"FF",x"FE",x"1F",x"0B",x"00",x"00",x"04",
		x"C0",x"FF",x"FF",x"FF",x"F0",x"FF",x"08",x"10",x"00",x"1F",x"40",x"00",x"00",x"02",x"40",x"00",
		x"FF",x"FF",x"FF",x"FF",x"05",x"40",x"00",x"80",x"FF",x"FE",x"1F",x"20",x"00",x"00",x"05",x"00",
		x"00",x"FF",x"FF",x"00",x"F8",x"10",x"20",x"00",x"80",x"FF",x"00",x"07",x"D2",x"0A",x"08",x"EC",
		x"0A",x"FF",x"F1",x"0C",x"FA",x"03",x"FB",x"40",x"00",x"20",x"80",x"24",x"27",x"30",x"34",x"37",
		x"40",x"44",x"47",x"50",x"54",x"57",x"60",x"64",x"67",x"70",x"82",x"FF",x"F1",x"0C",x"FA",x"03",
		x"FB",x"40",x"00",x"70",x"80",x"67",x"64",x"60",x"57",x"54",x"57",x"60",x"30",x"27",x"24",x"20",
		x"80",x"FF",x"00",x"00",x"13",x"0B",x"01",x"5C",x"0B",x"02",x"A5",x"0B",x"03",x"EE",x"0B",x"04",
		x"37",x"0C",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"20",x"00",x"54",x"86",x"57",x"0C",
		x"50",x"54",x"0C",x"49",x"50",x"0C",x"49",x"50",x"0C",x"49",x"0C",x"47",x"0C",x"52",x"55",x"0C",
		x"4B",x"52",x"0C",x"47",x"4B",x"0C",x"47",x"4B",x"0C",x"50",x"0C",x"52",x"0C",x"49",x"48",x"49",
		x"4B",x"50",x"4B",x"50",x"52",x"54",x"0C",x"57",x"59",x"0C",x"57",x"54",x"50",x"57",x"52",x"0C",
		x"55",x"54",x"52",x"50",x"4B",x"54",x"88",x"0C",x"50",x"0C",x"88",x"FF",x"F0",x"03",x"F1",x"00",
		x"FA",x"00",x"FB",x"20",x"00",x"44",x"86",x"47",x"0C",x"40",x"44",x"0C",x"39",x"40",x"0C",x"39",
		x"40",x"0C",x"39",x"0C",x"37",x"0C",x"42",x"45",x"0C",x"3B",x"42",x"0C",x"37",x"3B",x"0C",x"37",
		x"3B",x"0C",x"40",x"0C",x"42",x"0C",x"39",x"38",x"39",x"3B",x"40",x"3B",x"40",x"42",x"44",x"0C",
		x"47",x"49",x"0C",x"47",x"44",x"40",x"47",x"42",x"0C",x"45",x"44",x"42",x"40",x"3B",x"44",x"88",
		x"0C",x"40",x"0C",x"88",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"20",x"00",x"50",x"86",
		x"54",x"0C",x"49",x"50",x"0C",x"45",x"49",x"0C",x"45",x"49",x"0C",x"45",x"0C",x"44",x"0C",x"4B",
		x"52",x"0C",x"47",x"4B",x"0C",x"42",x"45",x"0C",x"42",x"47",x"0C",x"49",x"0C",x"4B",x"0C",x"45",
		x"44",x"45",x"47",x"49",x"48",x"49",x"4B",x"50",x"0C",x"54",x"55",x"0C",x"54",x"50",x"49",x"54",
		x"4B",x"0C",x"52",x"50",x"4B",x"49",x"47",x"50",x"88",x"0C",x"47",x"0C",x"88",x"FF",x"F0",x"03",
		x"F1",x"00",x"FA",x"00",x"FB",x"20",x"00",x"40",x"86",x"44",x"0C",x"39",x"40",x"0C",x"35",x"39",
		x"0C",x"39",x"35",x"0C",x"35",x"0C",x"34",x"0C",x"3B",x"42",x"0C",x"37",x"3B",x"0C",x"32",x"35",
		x"0C",x"32",x"37",x"0C",x"39",x"0C",x"3B",x"0C",x"35",x"34",x"35",x"37",x"39",x"38",x"39",x"3B",
		x"45",x"0C",x"44",x"45",x"0C",x"44",x"40",x"39",x"44",x"3B",x"0C",x"42",x"40",x"3B",x"39",x"37",
		x"40",x"88",x"0C",x"37",x"0C",x"88",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"20",x"00",
		x"24",x"86",x"0C",x"27",x"0C",x"24",x"24",x"27",x"0C",x"20",x"0C",x"24",x"0C",x"20",x"20",x"24",
		x"0C",x"22",x"0C",x"25",x"0C",x"22",x"22",x"25",x"0C",x"1B",x"0C",x"22",x"0C",x"1B",x"1B",x"22",
		x"0C",x"19",x"0C",x"17",x"0C",x"15",x"0C",x"14",x"0C",x"15",x"0C",x"17",x"0C",x"19",x"0C",x"1B",
		x"0C",x"20",x"0C",x"24",x"0C",x"1B",x"1B",x"22",x"0C",x"20",x"20",x"24",x"0C",x"20",x"88",x"0C",
		x"88",x"FF",x"01",x"00",x"90",x"0C",x"01",x"BD",x"0C",x"02",x"EA",x"0C",x"03",x"17",x"0D",x"FF",
		x"F0",x"01",x"F1",x"05",x"FA",x"00",x"FB",x"28",x"00",x"54",x"87",x"47",x"84",x"54",x"87",x"47",
		x"84",x"52",x"87",x"45",x"84",x"52",x"87",x"45",x"84",x"50",x"87",x"44",x"84",x"50",x"87",x"44",
		x"84",x"50",x"86",x"0C",x"84",x"4B",x"50",x"87",x"52",x"84",x"F2",x"AE",x"0D",x"F0",x"01",x"F1",
		x"05",x"FA",x"00",x"FB",x"28",x"00",x"50",x"87",x"44",x"84",x"50",x"87",x"44",x"84",x"4B",x"87",
		x"42",x"84",x"4B",x"87",x"42",x"84",x"47",x"87",x"40",x"84",x"47",x"87",x"40",x"84",x"47",x"86",
		x"0C",x"84",x"47",x"49",x"87",x"4B",x"84",x"F2",x"BA",x"0E",x"F0",x"01",x"F1",x"05",x"FA",x"00",
		x"FB",x"28",x"00",x"40",x"87",x"47",x"84",x"45",x"87",x"44",x"84",x"39",x"87",x"3B",x"84",x"40",
		x"87",x"42",x"84",x"37",x"87",x"39",x"84",x"3B",x"87",x"40",x"84",x"42",x"86",x"0C",x"84",x"42",
		x"44",x"87",x"45",x"84",x"F2",x"C7",x"0F",x"F0",x"01",x"F1",x"01",x"FA",x"00",x"FB",x"28",x"00",
		x"24",x"88",x"17",x"88",x"22",x"88",x"15",x"88",x"20",x"88",x"17",x"88",x"20",x"86",x"0C",x"84",
		x"1B",x"20",x"87",x"22",x"84",x"F2",x"D3",x"10",x"01",x"00",x"46",x"0D",x"01",x"5B",x"0D",x"02",
		x"73",x"0D",x"03",x"8B",x"0D",x"FF",x"F0",x"02",x"F1",x"08",x"FA",x"00",x"FB",x"30",x"00",x"55",
		x"88",x"54",x"52",x"50",x"49",x"8A",x"50",x"86",x"F2",x"87",x"11",x"F0",x"02",x"F1",x"08",x"FA",
		x"00",x"FB",x"30",x"00",x"0C",x"84",x"59",x"88",x"57",x"55",x"54",x"87",x"52",x"8A",x"57",x"86",
		x"F2",x"41",x"12",x"F0",x"02",x"F1",x"08",x"FA",x"00",x"FB",x"30",x"00",x"0C",x"86",x"60",x"88",
		x"5B",x"59",x"57",x"86",x"55",x"8A",x"57",x"86",x"F2",x"AF",x"12",x"F0",x"02",x"F1",x"07",x"FA",
		x"00",x"FB",x"30",x"00",x"17",x"88",x"15",x"14",x"12",x"10",x"8A",x"10",x"86",x"F2",x"21",x"13",
		x"01",x"00",x"AE",x"0D",x"01",x"BA",x"0E",x"02",x"C7",x"0F",x"03",x"D3",x"10",x"FF",x"F0",x"01",
		x"F1",x"05",x"FB",x"28",x"00",x"F3",x"DC",x"0D",x"F3",x"29",x"0E",x"F3",x"DC",x"0D",x"F3",x"37",
		x"0E",x"F3",x"3E",x"0E",x"F3",x"57",x"0E",x"F3",x"7C",x"0E",x"F3",x"95",x"0E",x"F3",x"3E",x"0E",
		x"F3",x"6A",x"0E",x"F3",x"7C",x"0E",x"F3",x"A7",x"0E",x"F2",x"AE",x"0D",x"54",x"87",x"53",x"84",
		x"54",x"87",x"53",x"84",x"54",x"86",x"50",x"0C",x"50",x"54",x"87",x"53",x"84",x"54",x"86",x"50",
		x"0C",x"50",x"0C",x"50",x"52",x"87",x"51",x"84",x"52",x"87",x"51",x"84",x"52",x"86",x"4B",x"0C",
		x"4B",x"52",x"87",x"51",x"84",x"52",x"86",x"4B",x"0C",x"4B",x"0C",x"4B",x"0C",x"88",x"50",x"4B",
		x"49",x"47",x"50",x"86",x"54",x"8A",x"0C",x"84",x"54",x"54",x"86",x"47",x"88",x"0C",x"84",x"54",
		x"52",x"86",x"45",x"88",x"0C",x"84",x"52",x"84",x"F4",x"50",x"88",x"4B",x"86",x"50",x"88",x"0C",
		x"84",x"4B",x"50",x"87",x"52",x"84",x"F4",x"50",x"88",x"50",x"4B",x"49",x"88",x"F4",x"54",x"87",
		x"53",x"84",x"54",x"87",x"53",x"84",x"54",x"86",x"4B",x"0C",x"4B",x"54",x"87",x"53",x"84",x"54",
		x"86",x"55",x"88",x"54",x"0C",x"86",x"F4",x"49",x"88",x"54",x"52",x"50",x"4B",x"86",x"50",x"88",
		x"49",x"88",x"0C",x"84",x"49",x"4B",x"87",x"50",x"84",x"F4",x"59",x"88",x"5B",x"60",x"86",x"5B",
		x"88",x"0C",x"84",x"59",x"89",x"0C",x"87",x"59",x"88",x"54",x"88",x"F4",x"52",x"87",x"51",x"84",
		x"52",x"87",x"51",x"84",x"52",x"86",x"49",x"0C",x"49",x"52",x"87",x"51",x"84",x"52",x"86",x"54",
		x"88",x"52",x"0C",x"86",x"F4",x"57",x"88",x"57",x"55",x"86",x"54",x"88",x"0C",x"84",x"52",x"89",
		x"0C",x"87",x"53",x"89",x"0C",x"86",x"F4",x"57",x"88",x"57",x"58",x"86",x"59",x"88",x"0C",x"86",
		x"5B",x"89",x"0C",x"84",x"4B",x"50",x"88",x"52",x"88",x"F4",x"F0",x"01",x"F1",x"05",x"FB",x"28",
		x"00",x"F3",x"E8",x"0E",x"F3",x"35",x"0F",x"F3",x"E8",x"0E",x"F3",x"43",x"0F",x"F3",x"4A",x"0F",
		x"F3",x"63",x"0F",x"F3",x"88",x"0F",x"F3",x"A1",x"0F",x"F3",x"4A",x"0F",x"F3",x"76",x"0F",x"F3",
		x"88",x"0F",x"F3",x"B3",x"0F",x"F2",x"BA",x"0E",x"50",x"87",x"4B",x"84",x"50",x"87",x"4B",x"84",
		x"50",x"86",x"49",x"0C",x"49",x"50",x"87",x"4B",x"84",x"50",x"86",x"47",x"0C",x"47",x"0C",x"47",
		x"4B",x"87",x"4A",x"84",x"4B",x"87",x"4A",x"84",x"4B",x"86",x"45",x"0C",x"45",x"4B",x"87",x"4A",
		x"84",x"4B",x"86",x"45",x"0C",x"45",x"0C",x"45",x"0C",x"88",x"49",x"47",x"45",x"44",x"47",x"86",
		x"50",x"8A",x"0C",x"84",x"50",x"50",x"86",x"44",x"88",x"0C",x"84",x"50",x"4B",x"86",x"42",x"88",
		x"0C",x"84",x"4B",x"84",x"F4",x"49",x"88",x"47",x"86",x"47",x"88",x"0C",x"84",x"47",x"49",x"87",
		x"4B",x"84",x"F4",x"47",x"88",x"47",x"47",x"45",x"88",x"F4",x"4B",x"87",x"4A",x"84",x"4B",x"87",
		x"4A",x"84",x"4B",x"86",x"48",x"0C",x"48",x"4B",x"87",x"4A",x"84",x"4B",x"86",x"50",x"88",x"4B",
		x"0C",x"86",x"F4",x"44",x"88",x"50",x"4B",x"49",x"47",x"86",x"49",x"88",x"44",x"0C",x"84",x"44",
		x"84",x"47",x"87",x"49",x"84",x"F4",x"54",x"88",x"57",x"59",x"86",x"57",x"88",x"0C",x"84",x"54",
		x"89",x"0C",x"87",x"54",x"88",x"49",x"88",x"F4",x"49",x"87",x"48",x"84",x"49",x"87",x"48",x"84",
		x"49",x"86",x"45",x"0C",x"45",x"49",x"87",x"48",x"84",x"49",x"86",x"50",x"88",x"49",x"0C",x"86",
		x"F4",x"54",x"88",x"54",x"52",x"86",x"50",x"88",x"0C",x"84",x"4B",x"89",x"0C",x"87",x"4A",x"89",
		x"0C",x"86",x"F4",x"52",x"88",x"52",x"54",x"86",x"55",x"88",x"0C",x"86",x"55",x"89",x"0C",x"84",
		x"47",x"84",x"49",x"88",x"4B",x"88",x"F4",x"F0",x"01",x"F1",x"00",x"FB",x"28",x"00",x"F3",x"F5",
		x"0F",x"F3",x"42",x"10",x"F3",x"F5",x"0F",x"F3",x"50",x"10",x"F3",x"57",x"10",x"F3",x"70",x"10",
		x"F3",x"94",x"10",x"F3",x"AD",x"10",x"F3",x"57",x"10",x"F3",x"82",x"10",x"F3",x"94",x"10",x"F3",
		x"BF",x"10",x"F2",x"C7",x"0F",x"44",x"87",x"43",x"84",x"44",x"87",x"43",x"84",x"44",x"86",x"40",
		x"0C",x"40",x"44",x"87",x"43",x"84",x"44",x"86",x"40",x"0C",x"40",x"0C",x"40",x"42",x"87",x"41",
		x"84",x"42",x"87",x"41",x"84",x"42",x"86",x"3B",x"0C",x"3B",x"42",x"87",x"41",x"84",x"42",x"86",
		x"3B",x"0C",x"3B",x"0C",x"3B",x"0C",x"88",x"40",x"3B",x"39",x"37",x"40",x"86",x"44",x"8A",x"0C",
		x"84",x"44",x"44",x"86",x"37",x"88",x"0C",x"84",x"44",x"42",x"86",x"45",x"88",x"0C",x"84",x"42",
		x"84",x"F4",x"40",x"88",x"3B",x"86",x"40",x"88",x"0C",x"84",x"3B",x"40",x"87",x"42",x"84",x"F4",
		x"40",x"88",x"40",x"3B",x"39",x"88",x"F4",x"44",x"87",x"43",x"84",x"44",x"87",x"43",x"84",x"44",
		x"86",x"3B",x"0C",x"3B",x"44",x"87",x"43",x"84",x"44",x"86",x"45",x"88",x"44",x"0C",x"86",x"F4",
		x"39",x"88",x"44",x"42",x"44",x"4B",x"86",x"40",x"88",x"39",x"0C",x"84",x"39",x"3B",x"87",x"40",
		x"84",x"F4",x"49",x"88",x"4B",x"50",x"86",x"4B",x"88",x"0C",x"84",x"49",x"89",x"0C",x"87",x"49",
		x"88",x"44",x"88",x"F4",x"42",x"87",x"41",x"84",x"42",x"87",x"41",x"84",x"42",x"86",x"49",x"0C",
		x"49",x"42",x"87",x"41",x"84",x"42",x"86",x"44",x"88",x"42",x"0C",x"86",x"F4",x"47",x"88",x"47",
		x"45",x"86",x"44",x"88",x"0C",x"84",x"42",x"89",x"0C",x"87",x"43",x"89",x"0C",x"86",x"F4",x"47",
		x"88",x"47",x"48",x"86",x"49",x"88",x"0C",x"86",x"4B",x"89",x"0C",x"84",x"3B",x"84",x"40",x"88",
		x"42",x"88",x"F4",x"F0",x"00",x"F1",x"01",x"FB",x"28",x"00",x"F3",x"01",x"11",x"F3",x"20",x"11",
		x"F3",x"01",x"11",x"F3",x"2D",x"11",x"F3",x"34",x"11",x"F3",x"3F",x"11",x"F3",x"55",x"11",x"F3",
		x"60",x"11",x"F3",x"34",x"11",x"F3",x"4A",x"11",x"F3",x"55",x"11",x"F3",x"6B",x"11",x"F2",x"D3",
		x"10",x"20",x"88",x"0C",x"17",x"0C",x"20",x"17",x"19",x"1B",x"19",x"0C",x"14",x"0C",x"19",x"14",
		x"15",x"17",x"20",x"0C",x"1B",x"0C",x"19",x"17",x"15",x"14",x"12",x"17",x"19",x"1B",x"88",x"F4",
		x"20",x"88",x"0C",x"89",x"0C",x"84",x"22",x"84",x"24",x"87",x"25",x"84",x"F4",x"20",x"88",x"20",
		x"1B",x"19",x"88",x"F4",x"24",x"88",x"0C",x"1B",x"0C",x"24",x"22",x"20",x"1B",x"88",x"F4",x"19",
		x"88",x"1B",x"20",x"1B",x"19",x"17",x"19",x"1B",x"88",x"F4",x"19",x"88",x"18",x"19",x"1B",x"20",
		x"0C",x"21",x"0C",x"88",x"F4",x"22",x"88",x"0C",x"19",x"0C",x"22",x"20",x"1B",x"19",x"88",x"F4",
		x"17",x"88",x"0C",x"1B",x"20",x"22",x"0C",x"23",x"0C",x"88",x"F4",x"17",x"89",x"17",x"86",x"1B",
		x"88",x"24",x"27",x"88",x"25",x"24",x"22",x"88",x"F4",x"01",x"00",x"87",x"11",x"01",x"41",x"12",
		x"02",x"AF",x"12",x"03",x"21",x"13",x"FF",x"F0",x"01",x"F1",x"00",x"FB",x"30",x"00",x"F3",x"A0",
		x"11",x"F3",x"B4",x"11",x"F3",x"A0",x"11",x"F3",x"C7",x"11",x"F3",x"E2",x"11",x"F2",x"87",x"11",
		x"40",x"86",x"42",x"44",x"47",x"45",x"44",x"45",x"47",x"45",x"44",x"45",x"4A",x"88",x"49",x"86",
		x"49",x"0C",x"86",x"F4",x"49",x"86",x"49",x"49",x"49",x"45",x"45",x"42",x"42",x"3A",x"3A",x"37",
		x"37",x"3A",x"42",x"40",x"0C",x"86",x"F4",x"52",x"86",x"52",x"52",x"52",x"49",x"49",x"45",x"45",
		x"42",x"45",x"49",x"50",x"88",x"49",x"86",x"45",x"0C",x"84",x"45",x"45",x"0C",x"45",x"86",x"0C",
		x"86",x"F4",x"39",x"88",x"40",x"47",x"89",x"45",x"86",x"44",x"45",x"40",x"39",x"40",x"84",x"0C",
		x"39",x"86",x"3A",x"40",x"3A",x"39",x"39",x"37",x"37",x"36",x"37",x"3A",x"47",x"8A",x"0C",x"3A",
		x"88",x"42",x"49",x"89",x"47",x"86",x"46",x"47",x"42",x"3A",x"42",x"84",x"0C",x"3A",x"86",x"40",
		x"42",x"44",x"42",x"42",x"40",x"40",x"42",x"44",x"40",x"49",x"8A",x"0C",x"88",x"40",x"50",x"0C",
		x"86",x"49",x"4A",x"49",x"88",x"4A",x"86",x"49",x"47",x"46",x"47",x"4A",x"88",x"0C",x"42",x"86",
		x"44",x"0C",x"42",x"44",x"0C",x"42",x"42",x"45",x"47",x"0C",x"45",x"47",x"8A",x"0C",x"0C",x"86",
		x"F4",x"F0",x"01",x"F1",x"00",x"FB",x"30",x"00",x"F3",x"5A",x"12",x"F3",x"6C",x"12",x"F3",x"5A",
		x"12",x"F3",x"74",x"12",x"F3",x"83",x"12",x"F2",x"41",x"12",x"0C",x"8A",x"35",x"86",x"0C",x"35",
		x"0C",x"35",x"0C",x"35",x"F5",x"08",x"0C",x"86",x"32",x"86",x"F6",x"F4",x"0C",x"86",x"34",x"0C",
		x"34",x"0C",x"86",x"F4",x"0C",x"86",x"34",x"0C",x"34",x"0C",x"84",x"40",x"40",x"0C",x"40",x"86",
		x"0C",x"86",x"F4",x"F5",x"08",x"0C",x"86",x"35",x"F6",x"F5",x"10",x"0C",x"32",x"F6",x"F5",x"04",
		x"0C",x"34",x"F6",x"F5",x"08",x"0C",x"35",x"F6",x"F5",x"04",x"0C",x"32",x"F6",x"3A",x"40",x"0C",
		x"3A",x"40",x"0C",x"3A",x"40",x"42",x"44",x"0C",x"42",x"44",x"8A",x"0C",x"0C",x"86",x"F4",x"F0",
		x"01",x"F1",x"00",x"FB",x"30",x"00",x"F3",x"C8",x"12",x"F3",x"D9",x"12",x"F3",x"C8",x"12",x"F3",
		x"E1",x"12",x"F3",x"F0",x"12",x"F2",x"AF",x"12",x"0C",x"8A",x"29",x"86",x"0C",x"29",x"F5",x"06",
		x"0C",x"29",x"F6",x"F5",x"04",x"0C",x"2A",x"F6",x"F4",x"0C",x"86",x"27",x"0C",x"27",x"0C",x"86",
		x"F4",x"0C",x"86",x"27",x"0C",x"27",x"0C",x"84",x"39",x"39",x"0C",x"39",x"86",x"0C",x"86",x"F4",
		x"F5",x"08",x"0C",x"86",x"29",x"F6",x"F5",x"08",x"0C",x"27",x"F6",x"F5",x"08",x"0C",x"2A",x"F6",
		x"F5",x"04",x"0C",x"27",x"F6",x"F5",x"08",x"0C",x"29",x"F6",x"F5",x"04",x"0C",x"27",x"F6",x"37",
		x"39",x"0C",x"37",x"39",x"0C",x"37",x"39",x"3A",x"40",x"0C",x"3A",x"40",x"8A",x"0C",x"0C",x"86",
		x"F4",x"F0",x"00",x"F1",x"00",x"FA",x"01",x"FB",x"30",x"00",x"F3",x"3C",x"13",x"F3",x"4F",x"13",
		x"F3",x"3C",x"13",x"F3",x"5E",x"13",x"F3",x"74",x"13",x"F2",x"21",x"13",x"10",x"86",x"12",x"14",
		x"15",x"88",x"10",x"10",x"09",x"12",x"09",x"12",x"86",x"12",x"15",x"19",x"1A",x"88",x"F4",x"15",
		x"88",x"1A",x"87",x"19",x"84",x"17",x"86",x"15",x"14",x"88",x"10",x"10",x"86",x"F4",x"12",x"88",
		x"1A",x"86",x"12",x"15",x"19",x"10",x"88",x"10",x"86",x"15",x"0C",x"84",x"15",x"15",x"0C",x"15",
		x"86",x"0C",x"86",x"F4",x"15",x"88",x"10",x"15",x"17",x"86",x"19",x"15",x"88",x"15",x"16",x"17",
		x"86",x"19",x"17",x"88",x"12",x"17",x"21",x"86",x"22",x"17",x"88",x"12",x"87",x"12",x"84",x"17",
		x"86",x"15",x"14",x"12",x"17",x"88",x"12",x"17",x"19",x"86",x"1A",x"17",x"88",x"12",x"0A",x"10",
		x"86",x"12",x"14",x"88",x"10",x"09",x"10",x"86",x"0A",x"09",x"88",x"05",x"09",x"07",x"86",x"09",
		x"07",x"09",x"0A",x"10",x"15",x"88",x"14",x"86",x"15",x"12",x"88",x"17",x"1A",x"86",x"17",x"14",
		x"12",x"0A",x"10",x"0C",x"0A",x"10",x"0C",x"0A",x"10",x"0A",x"10",x"0C",x"0A",x"10",x"8A",x"20",
		x"86",x"1A",x"17",x"14",x"10",x"86",x"F4",x"01",x"00",x"E5",x"13",x"01",x"1A",x"15",x"02",x"92",
		x"15",x"03",x"87",x"14",x"FF",x"F0",x"01",x"F1",x"05",x"FB",x"30",x"00",x"F3",x"0F",x"14",x"F3",
		x"2F",x"14",x"F3",x"2F",x"14",x"F0",x"02",x"F3",x"54",x"14",x"F3",x"6A",x"14",x"F3",x"54",x"14",
		x"F0",x"01",x"F1",x"08",x"F3",x"7D",x"14",x"F1",x"00",x"F3",x"2F",x"14",x"F2",x"E5",x"13",x"45",
		x"86",x"45",x"88",x"45",x"86",x"45",x"89",x"0C",x"86",x"45",x"45",x"45",x"45",x"43",x"89",x"0C",
		x"86",x"45",x"45",x"45",x"45",x"43",x"88",x"43",x"42",x"42",x"42",x"89",x"0C",x"86",x"F4",x"52",
		x"86",x"52",x"88",x"50",x"86",x"4A",x"88",x"0C",x"52",x"86",x"52",x"88",x"47",x"86",x"4A",x"88",
		x"0C",x"52",x"86",x"52",x"55",x"52",x"57",x"55",x"52",x"50",x"4A",x"4A",x"88",x"51",x"86",x"4A",
		x"88",x"0C",x"88",x"F4",x"53",x"86",x"53",x"84",x"53",x"87",x"51",x"86",x"53",x"53",x"84",x"53",
		x"87",x"51",x"86",x"53",x"88",x"48",x"8A",x"0C",x"88",x"F4",x"51",x"86",x"51",x"84",x"51",x"87",
		x"51",x"86",x"51",x"51",x"53",x"55",x"51",x"88",x"4A",x"8A",x"0C",x"88",x"F4",x"55",x"8A",x"57",
		x"88",x"57",x"55",x"8B",x"0C",x"88",x"F4",x"F0",x"00",x"F1",x"05",x"FA",x"01",x"FB",x"30",x"00",
		x"F3",x"AF",x"14",x"F3",x"CD",x"14",x"F3",x"CD",x"14",x"F3",x"ED",x"14",x"F3",x"00",x"15",x"F3",
		x"ED",x"14",x"F1",x"08",x"F3",x"13",x"15",x"F1",x"00",x"F3",x"CD",x"14",x"F2",x"87",x"14",x"F5",
		x"02",x"1A",x"86",x"2A",x"21",x"22",x"23",x"33",x"19",x"2A",x"F6",x"1A",x"2A",x"21",x"22",x"23",
		x"33",x"25",x"35",x"26",x"36",x"28",x"38",x"1A",x"1A",x"1A",x"1A",x"86",x"F4",x"F1",x"00",x"F5",
		x"02",x"0A",x"86",x"0A",x"11",x"12",x"13",x"13",x"19",x"1A",x"F6",x"0A",x"0A",x"11",x"12",x"13",
		x"13",x"15",x"15",x"16",x"16",x"18",x"18",x"1A",x"1A",x"1A",x"1A",x"86",x"F4",x"23",x"86",x"23",
		x"21",x"21",x"20",x"20",x"1A",x"1A",x"18",x"18",x"16",x"16",x"15",x"15",x"13",x"13",x"86",x"F4",
		x"11",x"86",x"11",x"10",x"10",x"0A",x"0A",x"08",x"08",x"0A",x"0A",x"10",x"10",x"11",x"11",x"12",
		x"12",x"86",x"F4",x"15",x"8A",x"10",x"15",x"15",x"8A",x"F4",x"F0",x"01",x"F1",x"05",x"FB",x"30",
		x"00",x"F3",x"40",x"15",x"F3",x"40",x"15",x"F3",x"40",x"15",x"F3",x"61",x"15",x"F3",x"72",x"15",
		x"F3",x"61",x"15",x"F1",x"08",x"F3",x"88",x"15",x"F1",x"05",x"F3",x"40",x"15",x"F2",x"1A",x"15",
		x"4A",x"86",x"4A",x"88",x"49",x"86",x"4A",x"89",x"0C",x"86",x"4A",x"4A",x"4A",x"49",x"86",x"45",
		x"89",x"0C",x"86",x"4A",x"4A",x"4A",x"49",x"45",x"88",x"45",x"45",x"45",x"45",x"89",x"0C",x"86",
		x"F4",x"4A",x"86",x"4A",x"4A",x"4A",x"88",x"0C",x"86",x"46",x"48",x"4A",x"4A",x"4A",x"8A",x"0C",
		x"88",x"F4",x"48",x"86",x"48",x"48",x"48",x"88",x"0C",x"86",x"48",x"48",x"51",x"88",x"50",x"86",
		x"48",x"88",x"0C",x"86",x"4A",x"45",x"86",x"F4",x"50",x"8A",x"53",x"88",x"53",x"50",x"8B",x"0C",
		x"88",x"F4",x"F0",x"01",x"F1",x"05",x"FA",x"00",x"FB",x"30",x"00",x"F3",x"BA",x"15",x"F3",x"BA",
		x"15",x"F3",x"BA",x"15",x"F3",x"DD",x"15",x"F3",x"EE",x"15",x"F3",x"DD",x"15",x"F1",x"08",x"F3",
		x"04",x"16",x"F1",x"05",x"F3",x"BA",x"15",x"F2",x"92",x"15",x"52",x"86",x"52",x"88",x"50",x"86",
		x"4A",x"47",x"4A",x"84",x"50",x"87",x"52",x"86",x"52",x"51",x"50",x"4A",x"89",x"0C",x"86",x"52",
		x"52",x"51",x"50",x"4A",x"88",x"4A",x"4A",x"4A",x"4A",x"89",x"0C",x"86",x"F4",x"46",x"86",x"46",
		x"46",x"46",x"88",x"0C",x"86",x"43",x"45",x"46",x"46",x"46",x"8A",x"0C",x"88",x"F4",x"45",x"86",
		x"45",x"45",x"45",x"88",x"0C",x"86",x"45",x"45",x"4A",x"88",x"48",x"86",x"45",x"88",x"0C",x"86",
		x"46",x"41",x"86",x"F4",x"49",x"8A",x"4A",x"88",x"4A",x"49",x"8B",x"0C",x"88",x"F4",x"00",x"00",
		x"22",x"16",x"01",x"42",x"16",x"02",x"62",x"16",x"03",x"82",x"16",x"04",x"9D",x"16",x"05",x"B9",
		x"16",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"1A",x"00",x"0C",x"89",x"47",x"8A",x"49",x"4B",x"50",
		x"86",x"F1",x"05",x"FB",x"34",x"00",x"49",x"86",x"4B",x"50",x"52",x"54",x"0C",x"84",x"50",x"0C",
		x"82",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"1A",x"00",x"0C",x"88",x"44",x"8A",x"45",x"47",x"49",
		x"88",x"F1",x"05",x"FB",x"34",x"00",x"39",x"86",x"3B",x"40",x"42",x"40",x"0C",x"84",x"40",x"0C",
		x"82",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"1A",x"00",x"0C",x"86",x"40",x"8A",x"42",x"44",x"45",
		x"89",x"F1",x"05",x"FB",x"34",x"00",x"35",x"86",x"37",x"39",x"3B",x"37",x"0C",x"84",x"37",x"0C",
		x"82",x"FF",x"F0",x"07",x"F1",x"00",x"FB",x"1A",x"00",x"0C",x"8C",x"0C",x"F1",x"01",x"FB",x"34",
		x"00",x"17",x"86",x"15",x"14",x"12",x"10",x"0C",x"84",x"10",x"0C",x"82",x"FF",x"F0",x"07",x"F1",
		x"00",x"FB",x"1A",x"00",x"0C",x"8C",x"0C",x"8C",x"F1",x"01",x"FB",x"34",x"00",x"27",x"86",x"25",
		x"24",x"22",x"20",x"0C",x"84",x"20",x"0C",x"82",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"1A",x"00",
		x"39",x"8A",x"3B",x"40",x"42",x"F1",x"05",x"FB",x"34",x"00",x"32",x"86",x"34",x"35",x"37",x"37",
		x"86",x"0C",x"84",x"34",x"0C",x"82",x"FF",x"00",x"00",x"EE",x"16",x"01",x"02",x"17",x"02",x"1B",
		x"17",x"03",x"32",x"17",x"04",x"46",x"17",x"05",x"5F",x"17",x"06",x"73",x"17",x"FF",x"F0",x"03",
		x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"54",x"54",x"52",x"52",x"49",x"4B",x"50",x"8A",x"0C",
		x"8F",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"0C",x"86",x"50",x"88",x"50",
		x"4B",x"4B",x"86",x"45",x"88",x"47",x"47",x"8A",x"0C",x"8F",x"FF",x"F0",x"03",x"F1",x"07",x"FB",
		x"30",x"00",x"0C",x"88",x"F5",x"04",x"47",x"88",x"F6",x"42",x"88",x"44",x"88",x"44",x"8A",x"0C",
		x"8F",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"44",x"44",x"42",x"42",x"40",
		x"3B",x"40",x"8A",x"0C",x"8F",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"0C",
		x"86",x"40",x"88",x"40",x"3B",x"3B",x"86",x"39",x"88",x"37",x"37",x"8A",x"0C",x"8F",x"FF",x"F0",
		x"03",x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"20",x"20",x"1B",x"1B",x"19",x"1B",x"20",x"8A",
		x"0C",x"8F",x"FF",x"F0",x"03",x"F1",x"07",x"FB",x"30",x"00",x"0C",x"88",x"15",x"15",x"14",x"14",
		x"12",x"14",x"17",x"8A",x"0C",x"8F",x"FF",x"00",x"00",x"95",x"17",x"01",x"E3",x"17",x"02",x"04",
		x"18",x"03",x"25",x"18",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"28",x"00",x"50",x"84",
		x"0C",x"50",x"54",x"57",x"0C",x"59",x"0C",x"60",x"0C",x"59",x"0C",x"57",x"0C",x"54",x"0C",x"49",
		x"0C",x"49",x"50",x"54",x"0C",x"57",x"0C",x"59",x"0C",x"57",x"0C",x"54",x"0C",x"50",x"0C",x"45",
		x"0C",x"45",x"49",x"50",x"0C",x"55",x"0C",x"57",x"0C",x"55",x"0C",x"50",x"0C",x"49",x"0C",x"47",
		x"0C",x"47",x"4B",x"52",x"0C",x"55",x"0C",x"57",x"0C",x"55",x"0C",x"52",x"0C",x"4B",x"0C",x"47",
		x"0C",x"8A",x"FF",x"F0",x"03",x"F1",x"09",x"FA",x"00",x"FB",x"28",x"00",x"47",x"8B",x"0C",x"86",
		x"47",x"49",x"8B",x"0C",x"86",x"44",x"40",x"8B",x"0C",x"86",x"3B",x"84",x"40",x"42",x"8B",x"0C",
		x"84",x"0C",x"8A",x"FF",x"F0",x"03",x"F1",x"09",x"FA",x"00",x"FB",x"28",x"00",x"40",x"8B",x"0C",
		x"86",x"40",x"39",x"8B",x"0C",x"86",x"39",x"35",x"8B",x"0C",x"86",x"34",x"84",x"35",x"37",x"8B",
		x"0C",x"84",x"0C",x"8A",x"FF",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"28",x"00",x"20",x"88",
		x"24",x"27",x"29",x"86",x"27",x"19",x"88",x"20",x"24",x"27",x"86",x"24",x"15",x"88",x"19",x"20",
		x"15",x"86",x"20",x"17",x"88",x"1B",x"22",x"25",x"86",x"22",x"17",x"84",x"0C",x"8A",x"FF",x"00",
		x"00",x"5D",x"18",x"01",x"BB",x"18",x"02",x"12",x"19",x"03",x"70",x"19",x"FF",x"F0",x"03",x"F1",
		x"09",x"FB",x"30",x"00",x"47",x"89",x"40",x"84",x"44",x"47",x"89",x"40",x"84",x"44",x"47",x"0C",
		x"47",x"0C",x"47",x"46",x"47",x"49",x"47",x"88",x"44",x"F1",x"00",x"59",x"84",x"58",x"59",x"86",
		x"5B",x"87",x"59",x"84",x"57",x"56",x"57",x"86",x"59",x"87",x"57",x"84",x"55",x"54",x"55",x"86",
		x"57",x"87",x"55",x"84",x"54",x"86",x"55",x"57",x"0C",x"59",x"84",x"58",x"59",x"86",x"5B",x"87",
		x"59",x"84",x"57",x"56",x"57",x"86",x"59",x"87",x"57",x"84",x"55",x"54",x"52",x"0C",x"5B",x"60",
		x"62",x"0C",x"60",x"86",x"0C",x"84",x"60",x"86",x"0C",x"86",x"FF",x"F0",x"03",x"F1",x"09",x"FB",
		x"30",x"00",x"44",x"89",x"37",x"84",x"40",x"44",x"89",x"37",x"84",x"40",x"44",x"0C",x"44",x"0C",
		x"44",x"43",x"44",x"45",x"44",x"88",x"40",x"F1",x"00",x"40",x"86",x"39",x"40",x"84",x"3B",x"39",
		x"86",x"3B",x"37",x"3B",x"84",x"39",x"37",x"86",x"39",x"35",x"39",x"84",x"37",x"35",x"86",x"0C",
		x"84",x"34",x"86",x"35",x"37",x"39",x"84",x"40",x"86",x"39",x"40",x"84",x"3B",x"39",x"86",x"3B",
		x"37",x"3B",x"84",x"39",x"37",x"86",x"39",x"35",x"3B",x"37",x"37",x"0C",x"84",x"37",x"86",x"0C",
		x"86",x"FF",x"F0",x"03",x"F1",x"09",x"FB",x"30",x"00",x"40",x"89",x"34",x"84",x"37",x"40",x"89",
		x"34",x"84",x"37",x"40",x"0C",x"40",x"0C",x"40",x"3B",x"40",x"42",x"40",x"88",x"37",x"F1",x"00",
		x"55",x"84",x"54",x"55",x"86",x"57",x"87",x"55",x"84",x"54",x"53",x"54",x"86",x"55",x"87",x"54",
		x"84",x"52",x"51",x"52",x"86",x"54",x"87",x"52",x"84",x"50",x"86",x"52",x"54",x"0C",x"55",x"84",
		x"54",x"55",x"86",x"57",x"87",x"55",x"84",x"54",x"53",x"54",x"86",x"55",x"87",x"54",x"84",x"52",
		x"50",x"4B",x"0C",x"57",x"59",x"5B",x"0C",x"57",x"86",x"0C",x"84",x"57",x"86",x"0C",x"86",x"FF",
		x"F0",x"03",x"F1",x"09",x"FB",x"30",x"00",x"37",x"89",x"30",x"84",x"34",x"37",x"89",x"30",x"84",
		x"34",x"37",x"0C",x"37",x"0C",x"37",x"36",x"37",x"39",x"37",x"88",x"34",x"F1",x"00",x"25",x"25",
		x"24",x"24",x"22",x"22",x"20",x"86",x"22",x"24",x"25",x"25",x"88",x"25",x"24",x"24",x"22",x"22",
		x"20",x"86",x"0C",x"84",x"20",x"86",x"0C",x"86",x"FF",x"00",x"00",x"BD",x"19",x"01",x"0A",x"1A",
		x"02",x"54",x"1A",x"03",x"99",x"1A",x"04",x"B3",x"1A",x"05",x"CD",x"1A",x"FF",x"F0",x"03",x"F1",
		x"08",x"FA",x"00",x"FB",x"30",x"00",x"40",x"86",x"40",x"88",x"47",x"45",x"86",x"44",x"42",x"40",
		x"47",x"88",x"45",x"44",x"42",x"86",x"42",x"42",x"88",x"49",x"47",x"86",x"45",x"44",x"42",x"49",
		x"47",x"88",x"45",x"44",x"44",x"86",x"47",x"88",x"4B",x"44",x"86",x"47",x"4B",x"45",x"49",x"88",
		x"50",x"45",x"86",x"49",x"50",x"52",x"52",x"0C",x"55",x"88",x"54",x"86",x"52",x"50",x"52",x"52",
		x"0C",x"89",x"52",x"86",x"50",x"4B",x"86",x"F2",x"BD",x"19",x"F0",x"03",x"F1",x"08",x"FA",x"00",
		x"FB",x"30",x"00",x"37",x"86",x"37",x"88",x"44",x"42",x"86",x"40",x"3B",x"37",x"44",x"88",x"42",
		x"40",x"3B",x"86",x"39",x"39",x"88",x"45",x"44",x"86",x"42",x"40",x"39",x"45",x"44",x"88",x"42",
		x"40",x"3B",x"86",x"44",x"88",x"47",x"3B",x"86",x"44",x"47",x"40",x"45",x"88",x"49",x"40",x"86",
		x"45",x"49",x"49",x"49",x"89",x"0C",x"8A",x"49",x"86",x"49",x"0C",x"89",x"4B",x"86",x"50",x"52",
		x"86",x"F2",x"0A",x"1A",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"30",x"00",x"F5",x"0D",x"20",
		x"86",x"F6",x"19",x"86",x"1B",x"20",x"86",x"F5",x"0D",x"22",x"86",x"F6",x"1B",x"86",x"20",x"22",
		x"86",x"F5",x"05",x"24",x"86",x"F6",x"20",x"86",x"22",x"24",x"86",x"F5",x"05",x"25",x"86",x"F6",
		x"22",x"86",x"24",x"25",x"22",x"22",x"0C",x"17",x"88",x"19",x"86",x"1B",x"20",x"22",x"22",x"0C",
		x"89",x"17",x"86",x"19",x"1B",x"86",x"F2",x"54",x"1A",x"F0",x"02",x"F1",x"0A",x"FB",x"30",x"00",
		x"30",x"8E",x"32",x"34",x"8C",x"35",x"37",x"86",x"37",x"0C",x"8B",x"37",x"86",x"37",x"0C",x"8B",
		x"F2",x"99",x"1A",x"F0",x"02",x"F1",x"0A",x"FB",x"30",x"00",x"34",x"8E",x"35",x"37",x"8C",x"39",
		x"3B",x"86",x"3B",x"0C",x"8B",x"3B",x"86",x"3B",x"0C",x"8B",x"F2",x"B3",x"1A",x"F0",x"02",x"F1",
		x"0A",x"FB",x"30",x"00",x"37",x"8E",x"39",x"3B",x"8C",x"40",x"42",x"86",x"42",x"0C",x"8B",x"42",
		x"86",x"42",x"0C",x"8B",x"F2",x"CD",x"1A",x"00",x"00",x"FE",x"1A",x"01",x"65",x"1B",x"02",x"24",
		x"1C",x"03",x"89",x"1C",x"04",x"DB",x"1C",x"05",x"F4",x"1C",x"06",x"0D",x"1D",x"FF",x"F0",x"03",
		x"F1",x"01",x"FA",x"00",x"FB",x"30",x"00",x"F5",x"04",x"50",x"88",x"F6",x"F5",x"04",x"4B",x"88",
		x"F6",x"F5",x"04",x"49",x"88",x"F6",x"0C",x"86",x"47",x"88",x"49",x"4B",x"50",x"86",x"F5",x"04",
		x"50",x"88",x"F6",x"F5",x"04",x"4B",x"88",x"F6",x"49",x"88",x"45",x"4B",x"47",x"50",x"49",x"52",
		x"52",x"55",x"55",x"88",x"F5",x"04",x"54",x"88",x"F6",x"F5",x"04",x"52",x"88",x"F6",x"F5",x"04",
		x"50",x"88",x"F6",x"4B",x"88",x"4B",x"4B",x"86",x"4B",x"50",x"52",x"86",x"F5",x"04",x"54",x"88",
		x"F6",x"F5",x"04",x"52",x"88",x"F6",x"50",x"88",x"49",x"52",x"4B",x"54",x"50",x"55",x"55",x"57",
		x"57",x"88",x"F2",x"FE",x"1A",x"F0",x"03",x"F1",x"00",x"FA",x"00",x"FB",x"30",x"00",x"F3",x"89",
		x"1B",x"F3",x"A2",x"1B",x"F3",x"89",x"1B",x"F3",x"B7",x"1B",x"F3",x"D7",x"1B",x"F3",x"F0",x"1B",
		x"F3",x"D7",x"1B",x"F3",x"06",x"1C",x"F2",x"65",x"1B",x"F5",x"03",x"0C",x"86",x"49",x"86",x"F6",
		x"50",x"84",x"4B",x"49",x"86",x"F5",x"03",x"0C",x"86",x"47",x"86",x"F6",x"4B",x"84",x"49",x"47",
		x"86",x"F4",x"F5",x"03",x"0C",x"86",x"45",x"86",x"F6",x"49",x"84",x"47",x"45",x"86",x"44",x"44",
		x"45",x"45",x"47",x"47",x"49",x"49",x"F4",x"0C",x"86",x"45",x"45",x"84",x"47",x"49",x"86",x"0C",
		x"47",x"47",x"84",x"49",x"4B",x"86",x"0C",x"49",x"49",x"84",x"4B",x"50",x"86",x"0C",x"4B",x"0C",
		x"4B",x"0C",x"52",x"0C",x"52",x"86",x"F4",x"F5",x"03",x"0C",x"86",x"50",x"86",x"F6",x"54",x"84",
		x"52",x"50",x"86",x"F5",x"03",x"0C",x"86",x"4B",x"86",x"F6",x"52",x"84",x"50",x"4B",x"86",x"F4",
		x"F5",x"03",x"0C",x"86",x"49",x"86",x"F6",x"50",x"84",x"4B",x"49",x"86",x"0C",x"47",x"0C",x"47",
		x"47",x"47",x"49",x"4B",x"86",x"F4",x"0C",x"86",x"49",x"49",x"84",x"4B",x"50",x"86",x"0C",x"4B",
		x"4B",x"84",x"50",x"52",x"86",x"0C",x"50",x"50",x"84",x"52",x"54",x"86",x"F5",x"04",x"0C",x"86",
		x"52",x"86",x"F6",x"F4",x"F0",x"03",x"F1",x"01",x"FA",x"00",x"FB",x"30",x"00",x"F5",x"04",x"45",
		x"88",x"F6",x"F5",x"04",x"44",x"88",x"F6",x"F5",x"04",x"42",x"88",x"F6",x"40",x"88",x"42",x"44",
		x"45",x"88",x"F5",x"04",x"45",x"88",x"F6",x"F5",x"04",x"44",x"88",x"F6",x"42",x"88",x"42",x"44",
		x"44",x"45",x"45",x"47",x"47",x"4B",x"4B",x"F5",x"04",x"49",x"88",x"F6",x"F5",x"04",x"47",x"88",
		x"F6",x"F5",x"04",x"45",x"88",x"F6",x"44",x"88",x"44",x"44",x"86",x"44",x"45",x"47",x"86",x"F5",
		x"04",x"49",x"88",x"F6",x"F5",x"04",x"47",x"88",x"F6",x"45",x"88",x"45",x"47",x"47",x"49",x"49",
		x"88",x"F5",x"04",x"4B",x"88",x"F6",x"F2",x"24",x"1C",x"F0",x"03",x"F1",x"01",x"FA",x"00",x"FB",
		x"30",x"00",x"F5",x"06",x"25",x"86",x"F6",x"27",x"86",x"25",x"86",x"F5",x"06",x"24",x"86",x"F6",
		x"25",x"86",x"24",x"86",x"F5",x"06",x"22",x"86",x"F6",x"24",x"86",x"22",x"20",x"20",x"22",x"22",
		x"24",x"24",x"25",x"25",x"F5",x"06",x"25",x"86",x"F6",x"27",x"86",x"25",x"86",x"F5",x"06",x"24",
		x"86",x"00",x"F6",x"25",x"86",x"24",x"22",x"22",x"20",x"22",x"24",x"24",x"22",x"24",x"25",x"25",
		x"24",x"25",x"86",x"F5",x"08",x"27",x"86",x"F6",x"F2",x"89",x"1C",x"F0",x"03",x"F1",x"09",x"FA",
		x"FF",x"FB",x"30",x"00",x"35",x"8C",x"34",x"32",x"30",x"35",x"34",x"32",x"8A",x"34",x"35",x"37",
		x"8C",x"F2",x"DB",x"1C",x"F0",x"03",x"F1",x"09",x"FA",x"00",x"FB",x"30",x"00",x"30",x"8C",x"2B",
		x"29",x"27",x"30",x"2B",x"29",x"8A",x"2B",x"30",x"32",x"8C",x"F2",x"F4",x"1C",x"F0",x"03",x"F1",
		x"00",x"FA",x"00",x"FB",x"30",x"00",x"F5",x"08",x"20",x"86",x"F6",x"F5",x"08",x"1B",x"86",x"F6",
		x"F5",x"08",x"19",x"86",x"F6",x"17",x"88",x"19",x"1B",x"86",x"17",x"19",x"86",x"1B",x"F5",x"08",
		x"20",x"86",x"F6",x"F5",x"08",x"1B",x"86",x"F6",x"F5",x"04",x"19",x"86",x"F6",x"F5",x"04",x"1B",
		x"86",x"F6",x"F5",x"04",x"20",x"86",x"F6",x"F5",x"08",x"22",x"86",x"F6",x"F2",x"0D",x"1D",x"00",
		x"00",x"66",x"1D",x"01",x"7C",x"1D",x"02",x"A2",x"1D",x"03",x"C7",x"1D",x"04",x"E3",x"1D",x"05",
		x"F1",x"1D",x"06",x"FF",x"1D",x"FF",x"F0",x"03",x"F1",x"08",x"FA",x"00",x"FB",x"28",x"00",x"F5",
		x"04",x"50",x"8B",x"F6",x"F5",x"04",x"52",x"8B",x"F6",x"F2",x"66",x"1D",x"F0",x"03",x"F1",x"08",
		x"FA",x"00",x"FB",x"28",x"00",x"0C",x"86",x"F5",x"03",x"54",x"8A",x"54",x"88",x"F6",x"54",x"8A",
		x"54",x"86",x"0C",x"86",x"F5",x"03",x"55",x"8A",x"55",x"88",x"F6",x"55",x"8A",x"55",x"86",x"F2",
		x"7C",x"1D",x"F0",x"03",x"F1",x"08",x"FA",x"00",x"FB",x"28",x"00",x"0C",x"88",x"F5",x"03",x"57",
		x"88",x"57",x"8A",x"F6",x"57",x"88",x"57",x"0C",x"88",x"F5",x"03",x"59",x"88",x"59",x"8A",x"F6",
		x"59",x"88",x"59",x"88",x"F2",x"A2",x"1D",x"F0",x"03",x"F1",x"08",x"FA",x"00",x"FB",x"28",x"00",
		x"0C",x"89",x"59",x"8B",x"59",x"59",x"59",x"89",x"0C",x"5B",x"8B",x"5B",x"5B",x"8B",x"5B",x"89",
		x"F2",x"C7",x"1D",x"F0",x"02",x"F1",x"03",x"FB",x"28",x"00",x"20",x"8F",x"22",x"8F",x"F2",x"E3",
		x"1D",x"F0",x"01",x"F1",x"03",x"FB",x"28",x"00",x"30",x"8F",x"32",x"8F",x"F2",x"F1",x"1D",x"F0",
		x"02",x"F1",x"08",x"FB",x"28",x"00",x"F5",x"04",x"40",x"86",x"44",x"47",x"49",x"47",x"44",x"F6",
		x"F5",x"04",x"42",x"86",x"45",x"49",x"4B",x"49",x"45",x"86",x"F6",x"F2",x"FF",x"1D",x"00",x"00",
		x"44",x"1E",x"01",x"64",x"1E",x"02",x"2C",x"1E",x"03",x"8C",x"1E",x"FF",x"F0",x"01",x"F1",x"07",
		x"FB",x"38",x"00",x"45",x"8A",x"F5",x"06",x"45",x"88",x"F6",x"47",x"8A",x"F5",x"06",x"47",x"88",
		x"F6",x"F2",x"2C",x"1E",x"F0",x"01",x"F1",x"07",x"FB",x"38",x"00",x"50",x"89",x"49",x"86",x"F5",
		x"06",x"50",x"86",x"49",x"86",x"F6",x"52",x"89",x"4B",x"86",x"F5",x"06",x"52",x"86",x"4B",x"86",
		x"F6",x"F2",x"44",x"1E",x"F0",x"01",x"F1",x"07",x"FB",x"38",x"00",x"0C",x"88",x"0C",x"84",x"F5",
		x"06",x"4B",x"86",x"47",x"86",x"F6",x"4B",x"86",x"47",x"84",x"0C",x"88",x"0C",x"84",x"F5",x"06",
		x"50",x"86",x"49",x"86",x"F6",x"50",x"86",x"49",x"84",x"F2",x"64",x"1E",x"F0",x"01",x"F1",x"01",
		x"FB",x"38",x"00",x"F5",x"02",x"15",x"86",x"15",x"19",x"19",x"20",x"20",x"19",x"19",x"86",x"F6",
		x"F5",x"02",x"17",x"86",x"17",x"1B",x"1B",x"22",x"22",x"1B",x"1B",x"86",x"F6",x"F2",x"8C",x"1E",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"45",x"0B",x"07",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"0D",x"44",x"0B",x"05",x"09",x"08",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"0E",x"10",x"11",x"45",x"03",x"07",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"12",x"13",x"11",x"44",x"0B",x"05",x"09",x"08",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"14",x"15",x"11",x"43",x"0B",x"05",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"16",x"17",x"11",x"45",x"03",x"04",x"09",x"6D",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"18",x"0F",x"11",x"42",x"0A",x"0A",x"0C",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"19",x"1A",x"1B",x"24",x"42",x"0A",x"0A",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"1C",x"1D",x"1E",x"25",x"42",x"0A",x"0A",x"04",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"1F",x"1D",x"1E",x"25",x"42",x"0A",x"0A",x"05",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"20",x"21",x"22",x"25",x"42",x"0A",x"0A",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"23",x"45",x"02",x"03",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"44",x"0B",x"0B",x"04",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"43",x"0B",x"0B",x"05",x"06",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"0A",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"0A",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3E",x"3F",x"40",x"41",x"4A",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3A",x"3B",x"3C",x"3D",x"49",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"36",x"37",x"38",x"39",x"4A",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"32",x"33",x"34",x"35",x"49",x"01",x"4B",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2E",x"2F",x"30",x"31",x"46",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2A",x"2B",x"2C",x"2D",x"48",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"26",x"27",x"28",x"29",x"47",x"01",x"4C",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"26",x"27",x"28",x"29",x"47",x"4B",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2A",x"2B",x"2C",x"2D",x"48",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2E",x"2F",x"30",x"31",x"46",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"32",x"33",x"34",x"35",x"4A",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"36",x"37",x"38",x"39",x"49",x"01",x"4C",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3A",x"3B",x"3C",x"3D",x"4A",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3E",x"3F",x"40",x"41",x"49",x"01",x"4B",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"80",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"82",x"83",x"84",x"85",x"86",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"8D",x"87",x"88",x"89",x"8A",x"8B",x"8C",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"8E",x"8F",x"90",x"91",x"92",x"C0",x"93",x"94",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"95",x"96",x"97",x"98",x"99",x"C1",x"9A",x"9B",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"9C",x"9D",x"9E",x"9F",x"A0",x"A1",x"A2",x"A3",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"A4",x"AA",x"A5",x"A6",x"A7",x"A8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"A9",x"AA",x"AA",x"AA",x"AB",x"AC",x"A8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"AD",x"AE",x"AA",x"AA",x"AA",x"AF",x"B0",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"B2",x"B3",x"AE",x"AA",x"AA",x"AA",x"B4",x"B5",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"B6",x"B7",x"B8",x"AE",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"BA",x"BB",x"AE",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"BC",x"BD",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"BE",x"BF",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F0",x"F9",x"F8",x"70",x"FC",x"F9",x"FC",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F1",x"70",x"FB",x"F8",x"F9",x"FB",x"F8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"FE",x"70",x"FB",x"FC",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F0",x"FA",x"70",x"FB",x"F9",x"FE",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F4",x"F5",x"F6",x"F8",x"F8",x"FC",x"FF",
		x"FF",x"01",x"01",x"C2",x"C3",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"CB",x"F7",x"FD",x"FF",
		x"FF",x"01",x"01",x"CC",x"CD",x"CE",x"CF",x"D0",x"D1",x"D2",x"D3",x"D4",x"D5",x"D6",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"D7",x"D8",x"D9",x"DA",x"DB",x"DC",x"DD",x"DE",x"DF",x"F8",x"FF",
		x"FF",x"01",x"01",x"01",x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E6",x"E7",x"E8",x"E9",x"FB",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"EA",x"EB",x"EC",x"ED",x"EE",x"EF",x"FA",x"70",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F4",x"6F",x"F6",x"FB",x"70",x"FA",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"FE",x"F9",x"F8",x"F9",x"FE",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"70",x"FB",x"F8",x"70",x"FC",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"F1",x"FA",x"F8",x"F9",x"FC",x"FA",x"FB",x"FE",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"8A",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"01",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"0A",x"0A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"8A",x"8A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"8A",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"55",x"54",x"54",x"54",x"54",x"54",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"56",x"57",x"57",x"57",x"58",x"58",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"5B",x"5A",x"5A",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"5E",x"5D",x"5C",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"5F",x"60",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"62",x"61",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"63",x"64",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"65",x"65",x"65",x"65",x"65",x"65",x"65",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"67",x"68",x"68",x"68",x"68",x"69",x"6A",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6C",x"6B",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6C",x"6B",x"53",x"52",x"51",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"45",x"0B",x"07",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"0D",x"44",x"0B",x"05",x"09",x"08",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"0E",x"10",x"11",x"45",x"03",x"07",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"12",x"13",x"11",x"44",x"0B",x"05",x"09",x"08",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"14",x"15",x"11",x"43",x"0B",x"05",x"08",x"09",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"16",x"17",x"11",x"45",x"03",x"04",x"09",x"6D",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"18",x"0F",x"11",x"42",x"0A",x"0A",x"0C",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"19",x"1A",x"1B",x"24",x"42",x"0A",x"0A",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"1C",x"1D",x"1E",x"25",x"42",x"0A",x"0A",x"04",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"1F",x"1D",x"1E",x"25",x"42",x"0A",x"0A",x"05",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"20",x"21",x"22",x"25",x"42",x"0A",x"0A",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"23",x"45",x"02",x"03",x"07",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"44",x"0B",x"0B",x"04",x"06",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6E",x"43",x"0B",x"0B",x"05",x"06",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"0A",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"0A",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"08",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"88",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3E",x"3F",x"40",x"41",x"4A",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3A",x"3B",x"3C",x"3D",x"49",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"36",x"37",x"38",x"39",x"4A",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"32",x"33",x"34",x"35",x"49",x"01",x"4B",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2E",x"2F",x"30",x"31",x"46",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2A",x"2B",x"2C",x"2D",x"48",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"26",x"27",x"28",x"29",x"47",x"01",x"4C",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"26",x"27",x"28",x"29",x"47",x"4B",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2A",x"2B",x"2C",x"2D",x"48",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"2E",x"2F",x"30",x"31",x"46",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"32",x"33",x"34",x"35",x"4A",x"4C",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"36",x"37",x"38",x"39",x"49",x"01",x"4C",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3A",x"3B",x"3C",x"3D",x"4A",x"01",x"01",x"FF",
		x"FF",x"01",x"71",x"72",x"73",x"74",x"75",x"76",x"3E",x"3F",x"40",x"41",x"49",x"01",x"4B",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"80",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"82",x"83",x"84",x"85",x"86",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"8D",x"87",x"88",x"89",x"8A",x"8B",x"8C",x"81",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"8E",x"8F",x"90",x"91",x"92",x"C0",x"93",x"94",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"95",x"96",x"97",x"98",x"99",x"C1",x"9A",x"9B",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"9C",x"9D",x"9E",x"9F",x"A0",x"A1",x"A2",x"A3",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"A4",x"AA",x"A5",x"A6",x"A7",x"A8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"A9",x"AA",x"AA",x"AA",x"AB",x"AC",x"A8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"AD",x"AE",x"AA",x"AA",x"AA",x"AF",x"B0",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"B2",x"B3",x"AE",x"AA",x"AA",x"AA",x"B4",x"B5",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"B6",x"B7",x"B8",x"AE",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"BA",x"BB",x"AE",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"BC",x"BD",x"AA",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"BE",x"BF",x"AA",x"AA",x"AA",x"B9",x"B1",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F0",x"F9",x"F8",x"70",x"FC",x"F9",x"FC",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F1",x"70",x"FB",x"F8",x"F9",x"FB",x"F8",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"FE",x"70",x"FB",x"FC",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F0",x"FA",x"70",x"FB",x"F9",x"FE",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F4",x"F5",x"F6",x"F8",x"F8",x"FC",x"FF",
		x"FF",x"01",x"01",x"C2",x"C3",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9",x"CA",x"CB",x"F7",x"FD",x"FF",
		x"FF",x"01",x"01",x"CC",x"CD",x"CE",x"CF",x"D0",x"D1",x"D2",x"D3",x"D4",x"D5",x"D6",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"D7",x"D8",x"D9",x"DA",x"DB",x"DC",x"DD",x"DE",x"DF",x"F8",x"FF",
		x"FF",x"01",x"01",x"01",x"E0",x"E1",x"E2",x"E3",x"E4",x"E5",x"E6",x"E7",x"E8",x"E9",x"FB",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"EA",x"EB",x"EC",x"ED",x"EE",x"EF",x"FA",x"70",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F4",x"6F",x"F6",x"FB",x"70",x"FA",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"FE",x"F9",x"F8",x"F9",x"FE",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"F2",x"F3",x"70",x"FB",x"F8",x"70",x"FC",x"FD",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"F1",x"FA",x"F8",x"F9",x"FC",x"FA",x"FB",x"FE",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"8A",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"01",x"0A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"08",x"08",x"08",x"08",x"0A",x"0A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"8A",x"8A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"8A",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"0A",
		x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"55",x"54",x"54",x"54",x"54",x"54",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"56",x"57",x"57",x"57",x"58",x"58",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"5B",x"5A",x"5A",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"59",x"59",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"5E",x"5D",x"5C",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"5F",x"60",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"62",x"61",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"63",x"64",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"65",x"65",x"65",x"65",x"65",x"65",x"65",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"67",x"68",x"68",x"68",x"68",x"69",x"6A",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6C",x"6B",x"53",x"52",x"51",x"FF",
		x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"6C",x"6B",x"53",x"52",x"51",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0A",x"0A",x"0A",x"0A",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"70",x"38",x"3C",x"7C",x"F0",x"00",x"00",x"00",x"40",x"E0",x"FC",x"7E",x"3E",
		x"F8",x"F0",x"7C",x"3C",x"38",x"70",x"00",x"00",x"7C",x"3E",x"7E",x"FC",x"E0",x"40",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"E0",x"20",x"18",
		x"08",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"C0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"1C",x"38",x"38",x"00",x"00",x"C0",x"E0",x"F0",x"38",x"1C",x"1C",
		x"38",x"38",x"1C",x"0F",x"07",x"03",x"00",x"00",x"1C",x"1C",x"38",x"F0",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"1F",x"38",x"70",x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"1C",x"0E",x"07",x"07",x"07",
		x"E0",x"E0",x"E0",x"70",x"38",x"1F",x"0F",x"07",x"07",x"07",x"07",x"0E",x"1C",x"F8",x"F0",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"1F",x"00",x"00",x"00",x"00",x"00",x"FE",x"FF",x"FF",
		x"1F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"05",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"1F",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"1F",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"1F",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
		x"00",x"00",x"00",x"03",x"07",x"0F",x"1F",x"1E",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"40",x"60",x"20",x"30",x"18",x"0C",
		x"18",x"30",x"30",x"60",x"60",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"06",x"06",x"06",x"04",x"04",x"00",x"18",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FA",x"FA",x"F2",x"E4",x"CC",x"18",x"E0",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"C0",x"E0",x"F1",x"F3",x"E7",x"0F",x"7F",x"FF",x"7A",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"20",x"BC",x"BF",x"BF",x"1F",x"07",x"01",x"C0",x"02",x"02",x"82",x"E2",x"E2",x"E2",x"E2",x"62",
		x"F0",x"F8",x"FE",x"7F",x"1F",x"0F",x"07",x"83",x"02",x"02",x"02",x"02",x"CA",x"8A",x"9A",x"3A",
		x"1F",x"07",x"00",x"00",x"80",x"00",x"70",x"F8",x"8A",x"0A",x"0A",x"3A",x"3A",x"7A",x"3A",x"1A",
		x"FC",x"00",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"0A",x"0A",x"02",x"02",x"82",x"C2",x"C2",x"02",
		x"80",x"00",x"00",x"00",x"00",x"08",x"18",x"38",x"3A",x"3A",x"FA",x"FA",x"FA",x"3A",x"0A",x"0A",
		x"7E",x"78",x"60",x"40",x"00",x"01",x"07",x"1F",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"8A",
		x"03",x"07",x"07",x"0F",x"0F",x"1F",x"1F",x"3E",x"C2",x"C2",x"C2",x"CA",x"8A",x"8A",x"0A",x"0A",
		x"38",x"62",x"0C",x"F8",x"F0",x"F0",x"E0",x"C0",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"F0",x"F0",x"F0",x"E0",x"E0",x"E0",x"C0",x"40",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
		x"00",x"00",x"80",x"00",x"00",x"00",x"01",x"03",x"1A",x"0A",x"0A",x"02",x"82",x"82",x"C2",x"C2",
		x"C0",x"8B",x"1B",x"7B",x"FF",x"FF",x"FF",x"FF",x"02",x"C2",x"C2",x"C2",x"82",x"82",x"82",x"1A",
		x"FF",x"FC",x"F1",x"C7",x"1F",x"01",x"00",x"00",x"1A",x"7A",x"FA",x"FA",x"FA",x"FA",x"1A",x"02",
		x"00",x"FF",x"00",x"FF",x"FF",x"F8",x"FC",x"FE",x"00",x"E0",x"18",x"CC",x"E4",x"12",x"FA",x"7A",
		x"FF",x"FE",x"FC",x"F8",x"FF",x"FA",x"F8",x"F1",x"3A",x"7A",x"FA",x"02",x"02",x"02",x"42",x"C2",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"03",x"07",x"07",x"07",x"03",x"07",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"07",x"07",x"05",x"00",x"00",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"0F",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"F0",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"1C",x"38",x"38",x"00",x"00",x"C0",x"E0",x"F0",x"38",x"1C",x"1C",
		x"38",x"38",x"1C",x"0F",x"07",x"03",x"00",x"00",x"1C",x"1C",x"38",x"F0",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"1F",x"38",x"70",x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"1C",x"0E",x"07",x"07",x"07",
		x"E0",x"E0",x"E0",x"70",x"38",x"1F",x"0F",x"07",x"07",x"07",x"07",x"0E",x"1C",x"F8",x"F0",x"E0",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3A",x"7E",x"7E",x"5C",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7E",x"7E",x"54",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7C",x"38",x"70",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"2E",x"7E",x"7E",x"74",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FE",x"FF",x"80",x"C0",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"00",x"7E",x"42",x"42",x"7E",x"00",x"00",x"00",x"00",x"02",x"7E",x"22",x"00",x"00",x"00",
		x"00",x"00",x"7A",x"4A",x"4A",x"6E",x"00",x"00",x"00",x"00",x"7E",x"52",x"42",x"66",x"00",x"00",
		x"00",x"00",x"04",x"1E",x"04",x"7C",x"00",x"00",x"00",x"00",x"5E",x"52",x"52",x"72",x"00",x"00",
		x"00",x"00",x"5E",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"7E",x"40",x"40",x"40",x"00",x"00",
		x"00",x"00",x"7E",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"7E",x"52",x"52",x"72",x"00",x"00",
		x"00",x"00",x"7E",x"50",x"50",x"7E",x"00",x"00",x"00",x"00",x"1E",x"12",x"12",x"7E",x"00",x"00",
		x"00",x"00",x"66",x"42",x"42",x"7E",x"00",x"00",x"00",x"00",x"7E",x"12",x"12",x"1E",x"00",x"00",
		x"00",x"00",x"42",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"40",x"50",x"50",x"7E",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"7F",x"00",x"00",x"00",x"00",x"00",x"FE",x"FF",x"FF",
		x"7F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"07",x"00",x"00",x"00",x"60",x"18",x"8C",x"C4",x"F2",
		x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"FA",x"FC",x"FC",x"F8",x"60",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"07",x"07",x"0F",x"3F",x"4F",x"00",x"00",x"00",x"AC",x"AC",x"AE",x"AE",x"AE",
		x"87",x"87",x"80",x"47",x"38",x"00",x"00",x"00",x"AC",x"AC",x"00",x"00",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"70",x"38",x"3C",x"7C",x"F0",x"00",x"00",x"00",x"40",x"E0",x"FC",x"7E",x"3E",
		x"F8",x"F0",x"7C",x"3C",x"38",x"70",x"00",x"00",x"7C",x"3E",x"7E",x"FC",x"E0",x"40",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"E0",x"20",x"18",
		x"08",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"C0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"1C",x"38",x"38",x"00",x"00",x"C0",x"E0",x"F0",x"38",x"1C",x"1C",
		x"38",x"38",x"1C",x"0F",x"07",x"03",x"00",x"00",x"1C",x"1C",x"38",x"F0",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"1F",x"38",x"70",x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"1C",x"0E",x"07",x"07",x"07",
		x"E0",x"E0",x"E0",x"70",x"38",x"1F",x"0F",x"07",x"07",x"07",x"07",x"0E",x"1C",x"F8",x"F0",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"1F",x"00",x"00",x"00",x"00",x"00",x"FE",x"FF",x"FF",
		x"1F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"05",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"1F",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"1F",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"1F",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",
		x"00",x"00",x"00",x"03",x"07",x"0F",x"1F",x"1E",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"40",x"60",x"20",x"30",x"18",x"0C",
		x"18",x"30",x"30",x"60",x"60",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"06",x"06",x"06",x"04",x"04",x"00",x"18",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FA",x"FA",x"F2",x"E4",x"CC",x"18",x"E0",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"C0",x"E0",x"F1",x"F3",x"E7",x"0F",x"7F",x"FF",x"7A",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",x"FA",
		x"20",x"BC",x"BF",x"BF",x"1F",x"07",x"01",x"C0",x"02",x"02",x"82",x"E2",x"E2",x"E2",x"E2",x"62",
		x"F0",x"F8",x"FE",x"7F",x"1F",x"0F",x"07",x"83",x"02",x"02",x"02",x"02",x"CA",x"8A",x"9A",x"3A",
		x"1F",x"07",x"00",x"00",x"80",x"00",x"70",x"F8",x"8A",x"0A",x"0A",x"3A",x"3A",x"7A",x"3A",x"1A",
		x"FC",x"00",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"0A",x"0A",x"02",x"02",x"82",x"C2",x"C2",x"02",
		x"80",x"00",x"00",x"00",x"00",x"08",x"18",x"38",x"3A",x"3A",x"FA",x"FA",x"FA",x"3A",x"0A",x"0A",
		x"7E",x"78",x"60",x"40",x"00",x"01",x"07",x"1F",x"0A",x"0A",x"0A",x"0A",x"0A",x"8A",x"8A",x"8A",
		x"03",x"07",x"07",x"0F",x"0F",x"1F",x"1F",x"3E",x"C2",x"C2",x"C2",x"CA",x"8A",x"8A",x"0A",x"0A",
		x"38",x"62",x"0C",x"F8",x"F0",x"F0",x"E0",x"C0",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
		x"F0",x"F0",x"F0",x"E0",x"E0",x"E0",x"C0",x"40",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
		x"00",x"00",x"80",x"00",x"00",x"00",x"01",x"03",x"1A",x"0A",x"0A",x"02",x"82",x"82",x"C2",x"C2",
		x"C0",x"8B",x"1B",x"7B",x"FF",x"FF",x"FF",x"FF",x"02",x"C2",x"C2",x"C2",x"82",x"82",x"82",x"1A",
		x"FF",x"FC",x"F1",x"C7",x"1F",x"01",x"00",x"00",x"1A",x"7A",x"FA",x"FA",x"FA",x"FA",x"1A",x"02",
		x"00",x"FF",x"00",x"FF",x"FF",x"F8",x"FC",x"FE",x"00",x"E0",x"18",x"CC",x"E4",x"12",x"FA",x"7A",
		x"FF",x"FE",x"FC",x"F8",x"FF",x"FA",x"F8",x"F1",x"3A",x"7A",x"FA",x"02",x"02",x"02",x"42",x"C2",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"C0",x"E0",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"78",x"38",x"18",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"78",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"F9",x"F8",
		x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FB",x"F9",x"78",x"38",x"18",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"00",x"00",x"03",x"07",x"07",x"07",x"03",x"07",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"07",x"07",x"05",x"00",x"00",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"0F",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"F0",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0F",x"1C",x"38",x"38",x"00",x"00",x"C0",x"E0",x"F0",x"38",x"1C",x"1C",
		x"38",x"38",x"1C",x"0F",x"07",x"03",x"00",x"00",x"1C",x"1C",x"38",x"F0",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"1F",x"38",x"70",x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"1C",x"0E",x"07",x"07",x"07",
		x"E0",x"E0",x"E0",x"70",x"38",x"1F",x"0F",x"07",x"07",x"07",x"07",x"0E",x"1C",x"F8",x"F0",x"E0",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3A",x"7E",x"7E",x"5C",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7E",x"7E",x"54",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7C",x"38",x"70",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"2E",x"7E",x"7E",x"74",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FE",x"FF",x"80",x"C0",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"00",x"7E",x"42",x"42",x"7E",x"00",x"00",x"00",x"00",x"02",x"7E",x"22",x"00",x"00",x"00",
		x"00",x"00",x"7A",x"4A",x"4A",x"6E",x"00",x"00",x"00",x"00",x"7E",x"52",x"42",x"66",x"00",x"00",
		x"00",x"00",x"04",x"1E",x"04",x"7C",x"00",x"00",x"00",x"00",x"5E",x"52",x"52",x"72",x"00",x"00",
		x"00",x"00",x"5E",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"7E",x"40",x"40",x"40",x"00",x"00",
		x"00",x"00",x"7E",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"7E",x"52",x"52",x"72",x"00",x"00",
		x"00",x"00",x"7E",x"50",x"50",x"7E",x"00",x"00",x"00",x"00",x"1E",x"12",x"12",x"7E",x"00",x"00",
		x"00",x"00",x"66",x"42",x"42",x"7E",x"00",x"00",x"00",x"00",x"7E",x"12",x"12",x"1E",x"00",x"00",
		x"00",x"00",x"42",x"52",x"52",x"7E",x"00",x"00",x"00",x"00",x"40",x"50",x"50",x"7E",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"7F",x"00",x"00",x"00",x"00",x"00",x"FE",x"FF",x"FF",
		x"7F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"07",x"00",x"00",x"00",x"60",x"18",x"8C",x"C4",x"F2",
		x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"FA",x"FC",x"FC",x"F8",x"60",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"30",x"1C",x"06",x"C2",x"F1",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FC",x"70",x"00",x"00",
		x"00",x"00",x"00",x"07",x"07",x"0F",x"3F",x"4F",x"00",x"00",x"00",x"AC",x"AC",x"AE",x"AE",x"AE",
		x"87",x"87",x"80",x"47",x"38",x"00",x"00",x"00",x"AC",x"AC",x"00",x"00",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"13",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"0F",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"70",x"38",x"3F",x"63",x"E3",x"00",x"00",x"0E",x"0E",x"1E",x"12",x"90",x"90",
		x"FF",x"E3",x"63",x"3F",x"38",x"70",x"00",x"00",x"92",x"90",x"90",x"12",x"1E",x"0E",x"0C",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"CF",x"CF",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F3",x"F3",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"00",x"00",x"00",x"00",x"00",x"02",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",
		x"0B",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"E0",x"20",x"C0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"00",x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",
		x"30",x"30",x"18",x"0C",x"07",x"03",x"00",x"00",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"60",x"C0",x"C0",x"C0",x"E0",x"F0",x"18",x"0C",x"06",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"60",x"30",x"18",x"0F",x"07",x"03",x"03",x"03",x"06",x"0C",x"18",x"F0",x"E0",
		x"20",x"00",x"24",x"00",x"00",x"A7",x"30",x"40",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",
		x"78",x"70",x"07",x"28",x"80",x"20",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"21",x"01",x"00",x"AC",x"54",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"A8",x"01",x"01",x"20",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"20",x"00",x"14",x"21",x"83",x"24",x"10",x"38",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"58",x"A9",x"51",x"00",x"08",x"40",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"27",x"13",x"08",x"04",x"03",x"00",x"00",x"00",x"26",x"26",x"26",x"26",x"26",x"26",x"26",x"26",
		x"00",x"00",x"03",x"04",x"08",x"13",x"27",x"26",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"C8",x"90",x"20",x"40",x"80",x"00",x"00",x"00",
		x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"00",x"00",x"80",x"40",x"20",x"90",x"C8",x"C8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"0E",x"02",x"00",x"00",x"00",x"00",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"30",x"38",x"1C",x"20",x"20",x"30",x"30",x"33",x"3F",x"F8",x"00",
		x"00",x"0F",x"3C",x"78",x"38",x"10",x"40",x"40",x"E0",x"F0",x"F0",x"78",x"38",x"1B",x"09",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"F9",x"F9",x"F1",x"E3",x"C2",x"06",x"1C",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"81",x"81",x"81",x"C1",x"C1",x"E1",x"E1",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E1",x"F1",x"F1",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"C0",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F8",x"09",x"09",x"01",x"01",x"01",x"01",x"01",x"01",
		x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"1F",x"1F",x"0F",x"0F",x"07",x"07",x"03",x"03",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"01",x"01",x"00",x"00",x"00",x"80",x"80",x"80",x"F9",x"F9",x"F9",x"79",x"79",x"39",x"19",x"19",
		x"3E",x"1C",x"08",x"00",x"04",x"0E",x"7F",x"FF",x"79",x"79",x"39",x"19",x"01",x"01",x"01",x"81",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"C1",x"E1",x"F1",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"1F",x"03",x"00",x"00",x"20",x"78",x"7E",x"3F",x"E1",x"E1",x"61",x"01",x"01",x"01",x"01",x"81",
		x"0F",x"07",x"01",x"80",x"E0",x"F0",x"F8",x"7C",x"E1",x"E1",x"C1",x"C1",x"09",x"09",x"19",x"39",
		x"00",x"00",x"01",x"00",x"00",x"E0",x"80",x"00",x"09",x"89",x"89",x"B9",x"39",x"79",x"39",x"19",
		x"00",x"FE",x"FF",x"FF",x"00",x"00",x"00",x"7F",x"01",x"01",x"01",x"81",x"01",x"01",x"01",x"E1",
		x"7F",x"F8",x"F8",x"F8",x"38",x"F0",x"E0",x"C0",x"B9",x"39",x"F9",x"F9",x"F9",x"39",x"09",x"09",
		x"80",x"07",x"1F",x"3F",x"FF",x"FE",x"F8",x"60",x"09",x"89",x"81",x"81",x"81",x"01",x"01",x"09",
		x"0C",x"38",x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"C0",x"81",x"03",x"07",x"0F",x"0F",x"1F",x"3F",x"81",x"81",x"81",x"81",x"81",x"89",x"89",x"89",
		x"00",x"0F",x"0F",x"1F",x"1F",x"1F",x"30",x"00",x"01",x"01",x"C1",x"C1",x"C1",x"C1",x"C1",x"41",
		x"0C",x"3E",x"7F",x"FF",x"FF",x"7F",x"3E",x"1C",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"41",x"41",x"41",x"D9",
		x"00",x"00",x"01",x"01",x"03",x"01",x"00",x"00",x"19",x"79",x"F9",x"F9",x"F9",x"F9",x"19",x"01",
		x"FF",x"00",x"00",x"E0",x"C0",x"C0",x"C0",x"C0",x"F0",x"1C",x"06",x"02",x"03",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"00",x"00",x"03",x"07",x"07",x"07",x"03",x"07",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"07",x"07",x"05",x"00",x"00",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0E",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"70",
		x"0E",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"70",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"00",x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",
		x"30",x"30",x"18",x"0C",x"07",x"03",x"00",x"00",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"60",x"C0",x"C0",x"C0",x"E0",x"F0",x"18",x"0C",x"06",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"60",x"30",x"18",x"0F",x"07",x"03",x"03",x"03",x"06",x"0C",x"18",x"F0",x"E0",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3A",x"7E",x"7E",x"5C",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7E",x"7E",x"54",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7C",x"38",x"70",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"2E",x"7E",x"7E",x"74",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"03",x"03",x"03",x"03",x"03",x"03",x"01",x"00",x"7F",x"3F",x"03",x"03",x"03",x"03",x"03",x"03",
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",
		x"78",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"50",x"00",x"00",x"00",x"60",x"F8",x"7C",x"3C",x"0E",
		x"29",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"28",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"10",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"64",x"94",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"08",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"07",x"00",x"07",x"00",x"07",x"00",x"00",x"00",x"FC",x"50",x"FE",x"50",x"FE",
		x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"50",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"70",x"38",x"3F",x"63",x"E3",x"00",x"00",x"0E",x"0E",x"1E",x"12",x"90",x"90",
		x"FF",x"E3",x"63",x"3F",x"38",x"70",x"00",x"00",x"92",x"90",x"90",x"12",x"1E",x"0E",x"0C",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"CF",x"CF",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F3",x"F3",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"00",x"00",x"00",x"00",x"00",x"02",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",
		x"0B",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"E0",x"20",x"C0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"00",x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",
		x"30",x"30",x"18",x"0C",x"07",x"03",x"00",x"00",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"60",x"C0",x"C0",x"C0",x"E0",x"F0",x"18",x"0C",x"06",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"60",x"30",x"18",x"0F",x"07",x"03",x"03",x"03",x"06",x"0C",x"18",x"F0",x"E0",
		x"20",x"00",x"24",x"00",x"00",x"A7",x"30",x"40",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",
		x"78",x"70",x"07",x"28",x"80",x"20",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"21",x"01",x"00",x"AC",x"54",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"A8",x"01",x"01",x"20",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"20",x"00",x"14",x"21",x"83",x"24",x"10",x"38",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"58",x"A9",x"51",x"00",x"08",x"40",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"27",x"13",x"08",x"04",x"03",x"00",x"00",x"00",x"26",x"26",x"26",x"26",x"26",x"26",x"26",x"26",
		x"00",x"00",x"03",x"04",x"08",x"13",x"27",x"26",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"C8",x"90",x"20",x"40",x"80",x"00",x"00",x"00",
		x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"00",x"00",x"80",x"40",x"20",x"90",x"C8",x"C8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"0E",x"02",x"00",x"00",x"00",x"00",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"30",x"38",x"1C",x"20",x"20",x"30",x"30",x"33",x"3F",x"F8",x"00",
		x"00",x"0F",x"3C",x"78",x"38",x"10",x"40",x"40",x"E0",x"F0",x"F0",x"78",x"38",x"1B",x"09",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"F9",x"F9",x"F1",x"E3",x"C2",x"06",x"1C",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"81",x"81",x"81",x"C1",x"C1",x"E1",x"E1",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E1",x"F1",x"F1",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"C0",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F8",x"09",x"09",x"01",x"01",x"01",x"01",x"01",x"01",
		x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"1F",x"1F",x"0F",x"0F",x"07",x"07",x"03",x"03",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"01",x"01",x"00",x"00",x"00",x"80",x"80",x"80",x"F9",x"F9",x"F9",x"79",x"79",x"39",x"19",x"19",
		x"3E",x"1C",x"08",x"00",x"04",x"0E",x"7F",x"FF",x"79",x"79",x"39",x"19",x"01",x"01",x"01",x"81",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"C1",x"E1",x"F1",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"1F",x"03",x"00",x"00",x"20",x"78",x"7E",x"3F",x"E1",x"E1",x"61",x"01",x"01",x"01",x"01",x"81",
		x"0F",x"07",x"01",x"80",x"E0",x"F0",x"F8",x"7C",x"E1",x"E1",x"C1",x"C1",x"09",x"09",x"19",x"39",
		x"00",x"00",x"01",x"00",x"00",x"E0",x"80",x"00",x"09",x"89",x"89",x"B9",x"39",x"79",x"39",x"19",
		x"00",x"FE",x"FF",x"FF",x"00",x"00",x"00",x"7F",x"01",x"01",x"01",x"81",x"01",x"01",x"01",x"E1",
		x"7F",x"F8",x"F8",x"F8",x"38",x"F0",x"E0",x"C0",x"B9",x"39",x"F9",x"F9",x"F9",x"39",x"09",x"09",
		x"80",x"07",x"1F",x"3F",x"FF",x"FE",x"F8",x"60",x"09",x"89",x"81",x"81",x"81",x"01",x"01",x"09",
		x"0C",x"38",x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"C0",x"81",x"03",x"07",x"0F",x"0F",x"1F",x"3F",x"81",x"81",x"81",x"81",x"81",x"89",x"89",x"89",
		x"00",x"0F",x"0F",x"1F",x"1F",x"1F",x"30",x"00",x"01",x"01",x"C1",x"C1",x"C1",x"C1",x"C1",x"41",
		x"0C",x"3E",x"7F",x"FF",x"FF",x"7F",x"3E",x"1C",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"41",x"41",x"41",x"D9",
		x"00",x"00",x"01",x"01",x"03",x"01",x"00",x"00",x"19",x"79",x"F9",x"F9",x"F9",x"F9",x"19",x"01",
		x"FF",x"00",x"00",x"E0",x"C0",x"C0",x"C0",x"C0",x"F0",x"1C",x"06",x"02",x"03",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"66",x"66",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",x"E6",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FE",
		x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"FF",x"FF",x"FF",x"80",x"FF",x"FF",x"E0",x"E0",x"E7",x"E7",x"E6",
		x"66",x"E6",x"E6",x"06",x"06",x"FE",x"FE",x"FF",x"00",x"FE",x"FE",x"06",x"06",x"E6",x"E6",x"E6",
		x"E6",x"E7",x"E7",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"E7",x"E7",x"E6",
		x"E6",x"E7",x"E7",x"E0",x"E0",x"E7",x"E7",x"E7",x"66",x"E6",x"E6",x"06",x"06",x"E6",x"E6",x"E6",
		x"00",x"00",x"03",x"07",x"07",x"07",x"03",x"07",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",
		x"07",x"07",x"03",x"07",x"07",x"05",x"00",x"00",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0E",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"70",
		x"0E",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"70",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"07",x"0C",x"18",x"30",x"30",x"00",x"00",x"C0",x"E0",x"30",x"18",x"0C",x"0C",
		x"30",x"30",x"18",x"0C",x"07",x"03",x"00",x"00",x"0C",x"0C",x"18",x"30",x"E0",x"C0",x"00",x"00",
		x"07",x"0F",x"18",x"30",x"60",x"C0",x"C0",x"C0",x"E0",x"F0",x"18",x"0C",x"06",x"03",x"03",x"03",
		x"C0",x"C0",x"C0",x"60",x"30",x"18",x"0F",x"07",x"03",x"03",x"03",x"06",x"0C",x"18",x"F0",x"E0",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3A",x"7E",x"7E",x"5C",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7E",x"7E",x"54",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"3E",x"7C",x"38",x"70",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"1F",x"3F",x"3F",x"3E",x"1F",x"3F",x"00",x"00",x"00",x"2E",x"7E",x"7E",x"74",x"00",
		x"3F",x"3E",x"1D",x"3F",x"3F",x"2E",x"00",x"00",x"0A",x"14",x"0A",x"14",x"00",x"00",x"00",x"00",
		x"03",x"03",x"03",x"03",x"03",x"03",x"01",x"00",x"7F",x"3F",x"03",x"03",x"03",x"03",x"03",x"03",
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",
		x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",
		x"78",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"50",x"00",x"00",x"00",x"60",x"F8",x"7C",x"3C",x"0E",
		x"29",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"28",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"10",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"64",x"94",x"00",x"00",x"70",x"FC",x"FE",x"3E",x"0F",x"07",
		x"08",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"80",x"E0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"07",x"00",x"07",x"00",x"07",x"00",x"00",x"00",x"FC",x"50",x"FE",x"50",x"FE",
		x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"50",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"02",x"03",x"0F",x"00",x"00",x"30",x"70",x"E0",x"ED",x"6F",x"6F",
		x"07",x"0F",x"03",x"02",x"00",x"00",x"00",x"00",x"7C",x"6F",x"6F",x"ED",x"E0",x"70",x"30",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF",
		x"CC",x"CC",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"F3",x"F3",x"F3",x"F3",x"03",x"03",x"FF",x"FF",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"33",x"33",x"F3",x"F3",x"03",x"03",x"FF",x"FF",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"03",x"03",x"F3",x"F3",x"33",x"33",
		x"FF",x"FF",x"03",x"03",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"FF",x"FF",x"C0",x"C0",x"CF",x"CF",x"CC",x"CC",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",x"C0",x"C0",x"CF",x"CF",x"CF",x"CF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"38",
		x"0C",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"18",x"C0",x"E0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",
		x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"00",x"00",x"C0",x"20",x"10",x"08",x"04",x"04",
		x"20",x"20",x"10",x"08",x"04",x"03",x"00",x"00",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",x"00",
		x"07",x"08",x"10",x"20",x"40",x"80",x"80",x"80",x"E0",x"10",x"08",x"04",x"02",x"01",x"01",x"01",
		x"80",x"80",x"80",x"40",x"20",x"10",x"08",x"07",x"01",x"01",x"01",x"02",x"04",x"08",x"10",x"E0",
		x"20",x"00",x"00",x"80",x"28",x"A8",x"5C",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"2F",x"AF",x"08",x"00",x"24",x"00",x"20",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"08",x"81",x"03",x"50",x"00",x"27",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"07",x"57",x"03",x"83",x"09",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"40",x"09",x"03",x"50",x"A8",x"43",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"27",x"17",x"27",x"83",x"21",x"14",x"00",x"20",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"C0",x"C2",x"C1",x"C0",x"C0",x"C0",x"C1",x"C2",x"03",x"0B",x"13",x"A3",x"43",x"A3",x"13",x"0B",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"1B",
		x"C0",x"DF",x"DF",x"C6",x"C6",x"C0",x"C0",x"C0",x"1B",x"FB",x"FB",x"1B",x"1B",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"CF",x"DF",x"DD",x"FF",x"FF",x"FF",x"FF",x"03",x"1B",x"9B",x"9B",
		x"D9",x"D8",x"D8",x"DC",x"DE",x"CE",x"C0",x"C0",x"DB",x"FB",x"FB",x"7B",x"3B",x"1B",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"DC",x"DF",x"DF",x"FF",x"FF",x"FF",x"FF",x"03",x"F3",x"FB",x"FB",
		x"DB",x"DB",x"DB",x"D8",x"D8",x"D8",x"C0",x"C0",x"3B",x"1B",x"1B",x"3B",x"7B",x"73",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"DF",x"DF",x"FF",x"FF",x"FF",x"FF",x"03",x"63",x"FB",x"FB",
		x"DC",x"CE",x"C7",x"C3",x"C1",x"C0",x"C0",x"C0",x"63",x"63",x"63",x"E3",x"E3",x"E3",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C1",x"DB",x"DB",x"FF",x"FF",x"FF",x"FF",x"03",x"F3",x"FB",x"BB",
		x"DB",x"DB",x"DB",x"DB",x"DF",x"DF",x"C0",x"C0",x"1B",x"1B",x"1B",x"3B",x"7B",x"73",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"2B",x"14",x"0B",x"04",x"03",x"00",x"00",x"00",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"00",x"00",x"03",x"04",x"0B",x"14",x"2B",x"2A",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"A8",x"50",x"A0",x"40",x"80",x"00",x"00",x"00",
		x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"00",x"00",x"80",x"40",x"A0",x"50",x"A8",x"A8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"18",x"10",x"00",x"20",x"20",
		x"06",x"07",x"03",x"03",x"03",x"03",x"02",x"02",x"58",x"DE",x"C3",x"01",x"03",x"1F",x"D8",x"00",
		x"00",x"0F",x"24",x"C0",x"C0",x"63",x"3F",x"1E",x"00",x"00",x"01",x"00",x"C0",x"E3",x"15",x"04",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"F0",x"F0",x"F0",x"F0",x"F8",x"00",x"00",x"FF",x"01",x"01",x"01",x"03",x"02",x"06",x"1C",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F9",x"79",x"79",x"79",x"39",x"39",x"19",x"19",
		x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"3F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"01",x"01",x"00",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"C1",x"E1",x"E1",x"F1",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"3E",x"1C",x"09",x"03",x"03",x"01",x"00",x"C0",x"79",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"79",
		x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"39",x"19",x"09",x"01",x"01",x"01",x"01",x"81",
		x"1F",x"83",x"80",x"80",x"20",x"78",x"7E",x"3F",x"E1",x"E1",x"61",x"01",x"01",x"01",x"01",x"81",
		x"0F",x"07",x"01",x"80",x"E0",x"F0",x"F8",x"7C",x"E1",x"E1",x"C1",x"C1",x"01",x"01",x"19",x"39",
		x"00",x"00",x"01",x"00",x"00",x"E0",x"80",x"00",x"01",x"81",x"81",x"81",x"39",x"79",x"39",x"19",
		x"00",x"FE",x"FF",x"FF",x"00",x"00",x"00",x"7F",x"09",x"09",x"01",x"81",x"01",x"01",x"01",x"E1",
		x"7F",x"F8",x"F8",x"F8",x"38",x"F0",x"E0",x"C0",x"81",x"01",x"01",x"01",x"19",x"39",x"09",x"09",
		x"80",x"07",x"1F",x"3F",x"FF",x"FE",x"F8",x"60",x"09",x"89",x"89",x"89",x"89",x"09",x"09",x"01",
		x"0C",x"38",x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"01",x"01",x"01",x"09",x"09",x"09",x"09",x"09",
		x"C0",x"81",x"03",x"07",x"0F",x"0F",x"1F",x"3F",x"89",x"89",x"89",x"89",x"89",x"81",x"81",x"81",
		x"00",x"0F",x"0F",x"1F",x"1F",x"1F",x"30",x"00",x"01",x"01",x"C1",x"C1",x"C1",x"C1",x"C1",x"41",
		x"0C",x"3E",x"7F",x"FF",x"FF",x"7F",x"3E",x"1C",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"C7",x"84",x"04",x"04",x"00",x"00",x"00",x"00",x"E1",x"01",x"01",x"01",x"41",x"41",x"41",x"C1",
		x"00",x"00",x"00",x"06",x"1C",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"1C",x"06",x"C2",x"E3",x"F1",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F4",x"F9",x"F9",x"F9",x"E1",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"00",x"00",x"00",x"07",x"04",x"07",x"00",x"07",x"00",x"00",x"00",x"C0",x"40",x"C0",x"00",x"C0",
		x"04",x"07",x"00",x"07",x"05",x"05",x"00",x"00",x"40",x"C0",x"00",x"40",x"40",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"06",x"0C",x"08",x"00",x"00",x"00",x"00",x"C0",x"60",x"30",x"10",
		x"08",x"0C",x"06",x"03",x"00",x"00",x"00",x"00",x"10",x"30",x"60",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"00",x"00",x"C0",x"20",x"10",x"08",x"04",x"04",
		x"20",x"20",x"10",x"08",x"04",x"03",x"00",x"00",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",x"00",
		x"07",x"08",x"10",x"20",x"40",x"80",x"80",x"80",x"E0",x"10",x"08",x"04",x"02",x"01",x"01",x"01",
		x"80",x"80",x"80",x"40",x"20",x"10",x"08",x"07",x"01",x"01",x"01",x"02",x"04",x"08",x"10",x"E0",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"74",x"54",x"5C",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"7C",x"54",x"54",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"7C",x"10",x"70",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"5C",x"54",x"74",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"FF",x"FF",x"FF",x"FF",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",
		x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"FF",x"81",x"FF",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"83",x"FF",x"A3",x"81",x"81",x"FF",
		x"FF",x"81",x"FB",x"CB",x"CB",x"EF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"C3",x"E7",x"81",x"FF",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"08",x"1C",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"2F",x"00",x"00",x"00",x"00",x"E0",x"70",x"38",x"8C",
		x"57",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"C4",x"E0",x"F0",x"F0",x"60",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"13",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"2F",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"07",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"04",x"01",x"03",x"00",x"00",x"00",x"50",x"FC",x"50",x"FE",x"FE",
		x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"02",x"03",x"0F",x"00",x"00",x"30",x"70",x"E0",x"ED",x"6F",x"6F",
		x"07",x"0F",x"03",x"02",x"00",x"00",x"00",x"00",x"7C",x"6F",x"6F",x"ED",x"E0",x"70",x"30",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF",
		x"CC",x"CC",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"F3",x"F3",x"F3",x"F3",x"03",x"03",x"FF",x"FF",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"33",x"33",x"F3",x"F3",x"03",x"03",x"FF",x"FF",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"03",x"03",x"F3",x"F3",x"33",x"33",
		x"FF",x"FF",x"03",x"03",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"FF",x"FF",x"C0",x"C0",x"CF",x"CF",x"CC",x"CC",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",x"C0",x"C0",x"CF",x"CF",x"CF",x"CF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"C6",x"7C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"C6",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"7C",x"C2",x"82",x"86",x"7C",x"38",x"00",x"00",x"02",x"02",x"FE",x"FE",x"42",x"02",x"00",
		x"62",x"F2",x"BA",x"9A",x"9E",x"CE",x"46",x"00",x"8C",x"DE",x"F2",x"B2",x"92",x"86",x"04",x"00",
		x"08",x"FE",x"FE",x"C8",x"68",x"38",x"18",x"00",x"9C",x"BE",x"A2",x"A2",x"A2",x"E6",x"E4",x"00",
		x"0C",x"9E",x"92",x"92",x"D2",x"7E",x"3C",x"00",x"C0",x"E0",x"B0",x"9E",x"8E",x"C0",x"C0",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"6C",x"00",x"78",x"FC",x"96",x"92",x"92",x"F2",x"60",x"00",
		x"7C",x"82",x"AA",x"AA",x"BA",x"82",x"7C",x"00",x"7C",x"82",x"BA",x"AA",x"BE",x"82",x"7C",x"00",
		x"2E",x"2E",x"3A",x"3A",x"00",x"20",x"7E",x"7E",x"00",x"00",x"00",x"E0",x"C0",x"00",x"00",x"00",
		x"20",x"00",x"70",x"50",x"50",x"7E",x"7E",x"00",x"00",x"00",x"00",x"F0",x"FA",x"FA",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"C8",x"88",x"C8",x"7E",x"3E",x"00",
		x"6C",x"FE",x"92",x"92",x"92",x"FE",x"FE",x"00",x"44",x"C6",x"82",x"82",x"C6",x"7C",x"38",x"00",
		x"38",x"7C",x"C6",x"82",x"82",x"FE",x"FE",x"00",x"00",x"82",x"92",x"92",x"92",x"FE",x"FE",x"00",
		x"80",x"90",x"90",x"90",x"90",x"FE",x"FE",x"00",x"9E",x"9E",x"92",x"82",x"C6",x"7C",x"38",x"00",
		x"FE",x"FE",x"10",x"10",x"10",x"FE",x"FE",x"00",x"00",x"82",x"82",x"FE",x"FE",x"82",x"82",x"00",
		x"FC",x"FE",x"02",x"02",x"02",x"06",x"04",x"00",x"82",x"C6",x"6E",x"3C",x"18",x"FE",x"FE",x"00",
		x"00",x"02",x"02",x"02",x"02",x"FE",x"FE",x"00",x"FE",x"FE",x"70",x"38",x"70",x"FE",x"FE",x"00",
		x"FE",x"FE",x"1C",x"38",x"70",x"FE",x"FE",x"00",x"7C",x"FE",x"82",x"82",x"82",x"FE",x"7C",x"00",
		x"70",x"88",x"88",x"88",x"88",x"FE",x"FE",x"00",x"7A",x"FC",x"8E",x"8A",x"82",x"FE",x"7C",x"00",
		x"72",x"F6",x"9E",x"8C",x"88",x"FE",x"FE",x"00",x"4C",x"DE",x"92",x"92",x"92",x"F6",x"64",x"00",
		x"00",x"80",x"80",x"FE",x"FE",x"80",x"80",x"00",x"FC",x"FE",x"02",x"02",x"02",x"FE",x"FC",x"00",
		x"F0",x"F8",x"1C",x"0E",x"1C",x"F8",x"F0",x"00",x"FC",x"FE",x"1C",x"38",x"1C",x"FE",x"FC",x"00",
		x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"C0",x"F0",x"1E",x"1E",x"F0",x"C0",x"00",
		x"C2",x"E2",x"F2",x"BA",x"9E",x"8E",x"86",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"38",
		x"0C",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"18",x"C0",x"E0",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",
		x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"00",x"00",x"C0",x"20",x"10",x"08",x"04",x"04",
		x"20",x"20",x"10",x"08",x"04",x"03",x"00",x"00",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",x"00",
		x"07",x"08",x"10",x"20",x"40",x"80",x"80",x"80",x"E0",x"10",x"08",x"04",x"02",x"01",x"01",x"01",
		x"80",x"80",x"80",x"40",x"20",x"10",x"08",x"07",x"01",x"01",x"01",x"02",x"04",x"08",x"10",x"E0",
		x"20",x"00",x"00",x"80",x"28",x"A8",x"5C",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"2F",x"AF",x"08",x"00",x"24",x"00",x"20",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"08",x"81",x"03",x"50",x"00",x"27",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"07",x"57",x"03",x"83",x"09",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"40",x"09",x"03",x"50",x"A8",x"43",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"27",x"17",x"27",x"83",x"21",x"14",x"00",x"20",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"C0",x"C2",x"C1",x"C0",x"C0",x"C0",x"C1",x"C2",x"03",x"0B",x"13",x"A3",x"43",x"A3",x"13",x"0B",
		x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"1B",
		x"C0",x"DF",x"DF",x"C6",x"C6",x"C0",x"C0",x"C0",x"1B",x"FB",x"FB",x"1B",x"1B",x"03",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"CF",x"DF",x"DD",x"FF",x"FF",x"FF",x"FF",x"03",x"1B",x"9B",x"9B",
		x"D9",x"D8",x"D8",x"DC",x"DE",x"CE",x"C0",x"C0",x"DB",x"FB",x"FB",x"7B",x"3B",x"1B",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"DC",x"DF",x"DF",x"FF",x"FF",x"FF",x"FF",x"03",x"F3",x"FB",x"FB",
		x"DB",x"DB",x"DB",x"D8",x"D8",x"D8",x"C0",x"C0",x"3B",x"1B",x"1B",x"3B",x"7B",x"73",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"DF",x"DF",x"FF",x"FF",x"FF",x"FF",x"03",x"63",x"FB",x"FB",
		x"DC",x"CE",x"C7",x"C3",x"C1",x"C0",x"C0",x"C0",x"63",x"63",x"63",x"E3",x"E3",x"E3",x"03",x"03",
		x"FF",x"FF",x"FF",x"FF",x"C0",x"C1",x"DB",x"DB",x"FF",x"FF",x"FF",x"FF",x"03",x"F3",x"FB",x"BB",
		x"DB",x"DB",x"DB",x"DB",x"DF",x"DF",x"C0",x"C0",x"1B",x"1B",x"1B",x"3B",x"7B",x"73",x"03",x"03",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"2B",x"14",x"0B",x"04",x"03",x"00",x"00",x"00",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",
		x"00",x"00",x"03",x"04",x"0B",x"14",x"2B",x"2A",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"A8",x"50",x"A0",x"40",x"80",x"00",x"00",x"00",
		x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"00",x"00",x"80",x"40",x"A0",x"50",x"A8",x"A8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"18",x"10",x"00",x"20",x"20",
		x"06",x"07",x"03",x"03",x"03",x"03",x"02",x"02",x"58",x"DE",x"C3",x"01",x"03",x"1F",x"D8",x"00",
		x"00",x"0F",x"24",x"C0",x"C0",x"63",x"3F",x"1E",x"00",x"00",x"01",x"00",x"C0",x"E3",x"15",x"04",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"F0",x"F0",x"F0",x"F0",x"F8",x"00",x"00",x"FF",x"01",x"01",x"01",x"03",x"02",x"06",x"1C",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F9",x"79",x"79",x"79",x"39",x"39",x"19",x"19",
		x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"3F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"07",x"07",x"03",x"03",x"01",x"01",x"01",x"00",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"C1",x"E1",x"E1",x"F1",x"F9",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",
		x"3E",x"1C",x"09",x"03",x"03",x"01",x"00",x"C0",x"79",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"79",
		x"E0",x"F0",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"39",x"19",x"09",x"01",x"01",x"01",x"01",x"81",
		x"1F",x"83",x"80",x"80",x"20",x"78",x"7E",x"3F",x"E1",x"E1",x"61",x"01",x"01",x"01",x"01",x"81",
		x"0F",x"07",x"01",x"80",x"E0",x"F0",x"F8",x"7C",x"E1",x"E1",x"C1",x"C1",x"01",x"01",x"19",x"39",
		x"00",x"00",x"01",x"00",x"00",x"E0",x"80",x"00",x"01",x"81",x"81",x"81",x"39",x"79",x"39",x"19",
		x"00",x"FE",x"FF",x"FF",x"00",x"00",x"00",x"7F",x"09",x"09",x"01",x"81",x"01",x"01",x"01",x"E1",
		x"7F",x"F8",x"F8",x"F8",x"38",x"F0",x"E0",x"C0",x"81",x"01",x"01",x"01",x"19",x"39",x"09",x"09",
		x"80",x"07",x"1F",x"3F",x"FF",x"FE",x"F8",x"60",x"09",x"89",x"89",x"89",x"89",x"09",x"09",x"01",
		x"0C",x"38",x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"01",x"01",x"01",x"09",x"09",x"09",x"09",x"09",
		x"C0",x"81",x"03",x"07",x"0F",x"0F",x"1F",x"3F",x"89",x"89",x"89",x"89",x"89",x"81",x"81",x"81",
		x"00",x"0F",x"0F",x"1F",x"1F",x"1F",x"30",x"00",x"01",x"01",x"C1",x"C1",x"C1",x"C1",x"C1",x"41",
		x"0C",x"3E",x"7F",x"FF",x"FF",x"7F",x"3E",x"1C",x"19",x"09",x"09",x"01",x"01",x"01",x"01",x"01",
		x"C7",x"84",x"04",x"04",x"00",x"00",x"00",x"00",x"E1",x"01",x"01",x"01",x"41",x"41",x"41",x"C1",
		x"00",x"00",x"00",x"06",x"1C",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"1C",x"06",x"C2",x"E3",x"F1",x"F9",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F4",x"F9",x"F9",x"F9",x"E1",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"14",x"14",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"95",
		x"7F",x"00",x"FF",x"00",x"FF",x"00",x"00",x"7F",x"FE",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FE",
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",
		x"95",x"94",x"97",x"90",x"9F",x"80",x"80",x"FF",x"FF",x"80",x"9F",x"90",x"97",x"94",x"94",x"95",
		x"95",x"15",x"F5",x"05",x"FD",x"01",x"01",x"FF",x"FF",x"01",x"FD",x"05",x"F5",x"15",x"15",x"95",
		x"95",x"14",x"D7",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"14",x"14",x"95",
		x"95",x"94",x"97",x"90",x"97",x"90",x"94",x"95",x"95",x"15",x"F5",x"15",x"F5",x"15",x"15",x"95",
		x"00",x"00",x"00",x"07",x"04",x"07",x"00",x"07",x"00",x"00",x"00",x"C0",x"40",x"C0",x"00",x"C0",
		x"04",x"07",x"00",x"07",x"05",x"05",x"00",x"00",x"40",x"C0",x"00",x"40",x"40",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"06",x"0C",x"08",x"00",x"00",x"00",x"00",x"C0",x"60",x"30",x"10",
		x"08",x"0C",x"06",x"03",x"00",x"00",x"00",x"00",x"10",x"30",x"60",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"04",x"08",x"10",x"20",x"20",x"00",x"00",x"C0",x"20",x"10",x"08",x"04",x"04",
		x"20",x"20",x"10",x"08",x"04",x"03",x"00",x"00",x"04",x"04",x"08",x"10",x"20",x"C0",x"00",x"00",
		x"07",x"08",x"10",x"20",x"40",x"80",x"80",x"80",x"E0",x"10",x"08",x"04",x"02",x"01",x"01",x"01",
		x"80",x"80",x"80",x"40",x"20",x"10",x"08",x"07",x"01",x"01",x"01",x"02",x"04",x"08",x"10",x"E0",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"74",x"54",x"5C",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"7C",x"54",x"54",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"7C",x"10",x"70",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"3E",x"22",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00",x"5C",x"54",x"74",x"00",
		x"22",x"3E",x"00",x"3A",x"2A",x"2E",x"00",x"00",x"00",x"14",x"08",x"14",x"00",x"00",x"00",x"00",
		x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"FF",x"FF",x"FF",x"FF",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",
		x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"FF",x"81",x"FF",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"83",x"FF",x"A3",x"81",x"81",x"FF",
		x"FF",x"81",x"FB",x"CB",x"CB",x"EF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"C3",x"E7",x"81",x"FF",
		x"FF",x"81",x"85",x"9F",x"85",x"FD",x"81",x"FF",x"FF",x"81",x"DF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"DF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"C1",x"C1",x"C1",x"81",x"FF",
		x"FF",x"81",x"FF",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"D3",x"D3",x"F3",x"81",x"FF",
		x"FF",x"81",x"FF",x"D1",x"D1",x"FF",x"81",x"FF",x"FF",x"81",x"9F",x"93",x"93",x"FF",x"81",x"FF",
		x"FF",x"81",x"E7",x"C3",x"C3",x"FF",x"81",x"FF",x"FF",x"81",x"FF",x"93",x"93",x"9F",x"81",x"FF",
		x"FF",x"81",x"C3",x"D3",x"D3",x"FF",x"81",x"FF",x"FF",x"81",x"C1",x"D1",x"D1",x"FF",x"81",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"08",x"1C",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"2F",x"00",x"00",x"00",x"00",x"E0",x"70",x"38",x"8C",
		x"57",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"C4",x"E0",x"F0",x"F0",x"60",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"13",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"2F",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"07",x"00",x"00",x"40",x"E0",x"F8",x"3C",x"0E",x"86",
		x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"E3",x"F3",x"F0",x"F8",x"F8",x"70",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"04",x"01",x"03",x"00",x"00",x"00",x"50",x"FC",x"50",x"FE",x"FE",
		x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"30",x"FC",x"FE",x"FE",x"FF",
		x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FC",x"30",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FB",x"BF",x"BB",x"FE",x"EF",x"FB",x"E9",x"FE",x"FF",x"ED",x"AA",x"FA",x"FA",x"EF",x"B3",x"FF",
		x"BF",x"F2",x"AF",x"EB",x"EE",x"FA",x"F9",x"00",x"BA",x"FE",x"AB",x"EF",x"BF",x"FE",x"FF",x"00",
		x"BB",x"FA",x"FE",x"AB",x"FF",x"EF",x"DA",x"EB",x"BC",x"EA",x"7F",x"BB",x"BF",x"BE",x"EF",x"EB",
		x"BD",x"3A",x"BE",x"EB",x"EE",x"FF",x"A0",x"00",x"BA",x"FF",x"EF",x"EE",x"BF",x"A3",x"01",x"00",
		x"C0",x"00",x"00",x"80",x"C0",x"80",x"80",x"80",x"00",x"01",x"00",x"01",x"06",x"05",x"00",x"00",
		x"80",x"00",x"00",x"80",x"80",x"80",x"C0",x"F4",x"01",x"01",x"07",x"00",x"00",x"06",x"07",x"0D",
		x"80",x"80",x"C0",x"00",x"80",x"80",x"C0",x"C0",x"0B",x"37",x"3A",x"CE",x"3F",x"05",x"03",x"BF",
		x"80",x"80",x"00",x"01",x"80",x"80",x"80",x"80",x"0A",x"7B",x"6F",x"4F",x"B6",x"FD",x"2B",x"01",
		x"38",x"68",x"5C",x"BC",x"EC",x"AE",x"4E",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F6",x"76",x"73",x"D3",x"D9",x"F9",x"B8",x"B0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"80",x"00",x"80",x"80",x"C0",x"80",x"80",x"01",x"01",x"0E",x"04",x"03",x"00",x"01",x"00",
		x"C0",x"C0",x"E0",x"C0",x"C0",x"80",x"80",x"80",x"00",x"03",x"07",x"02",x"05",x"01",x"00",x"03",
		x"FE",x"F8",x"7C",x"B8",x"90",x"80",x"C1",x"1A",x"7F",x"FF",x"7F",x"3F",x"1F",x"D9",x"E2",x"F1",
		x"37",x"5F",x"BD",x"FF",x"5F",x"13",x"F0",x"FE",x"F9",x"BE",x"FF",x"E4",x"D9",x"F3",x"E7",x"37",
		x"F4",x"F0",x"E5",x"EA",x"DF",x"FC",x"FE",x"BB",x"FB",x"F4",x"E3",x"F3",x"FB",x"1F",x"3F",x"9F",
		x"07",x"EF",x"CD",x"A3",x"F3",x"F8",x"FC",x"F4",x"EE",x"D8",x"B8",x"B1",x"6D",x"7A",x"FD",x"FF",
		x"FB",x"BF",x"BB",x"FE",x"EF",x"FB",x"E9",x"FE",x"FF",x"ED",x"AA",x"FA",x"FA",x"EF",x"B3",x"FF",
		x"BF",x"F2",x"AF",x"EB",x"EE",x"BA",x"B9",x"BF",x"BA",x"FE",x"AB",x"EF",x"BF",x"FE",x"FB",x"AA",
		x"BF",x"EE",x"AA",x"EF",x"3B",x"9F",x"FA",x"B9",x"FA",x"7F",x"FA",x"E8",x"FA",x"BF",x"FF",x"FB",
		x"EE",x"EE",x"F3",x"BF",x"CE",x"AB",x"EE",x"BE",x"EF",x"CA",x"EE",x"FF",x"BE",x"FB",x"BF",x"FB",
		x"77",x"8D",x"87",x"CD",x"C6",x"E4",x"AC",x"F8",x"FC",x"E8",x"61",x"01",x"00",x"01",x"00",x"01",
		x"F0",x"D0",x"E0",x"E0",x"C0",x"80",x"40",x"80",x"01",x"03",x"03",x"03",x"00",x"03",x"07",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"06",x"06",x"36",x"36",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"04",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"00",x"80",x"FF",x"FF",x"C0",x"40",x"80",x"FF",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"C0",x"40",x"80",x"FF",x"FF",x"C0",x"40",
		x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"80",x"FF",x"FF",x"C0",x"40",x"80",x"FF",x"FF",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"FF",x"FF",x"FC",x"FE",x"FE",x"E0",x"C0",x"C0",
		x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",
		x"F0",x"E0",x"00",x"3F",x"3F",x"3F",x"3F",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F8",x"F0",x"00",
		x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"C0",x"C0",x"D8",x"FC",x"FE",x"FE",x"E0",x"C0",
		x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"C0",x"C0",x"C0",x"D0",x"F0",x"F0",x"F0",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"07",x"07",x"00",x"3F",x"3F",x"00",x"00",x"00",x"FF",x"FF",x"00",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"3F",x"FF",x"C0",x"40",x"80",x"FF",x"FF",x"C0",x"40",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"80",x"FF",x"FF",x"C0",x"40",x"80",x"FF",x"FF",
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"C0",x"40",x"80",x"FF",x"FF",x"C0",x"40",x"80",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"C0",x"40",x"80",x"FF",x"FF",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"40",x"80",x"FF",x"FF",x"FF",x"FF",x"80",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"80",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"FF",x"7F",x"37",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"80",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"80",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"03",x"03",x"03",x"01",x"01",x"01",x"00",x"00",x"BF",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"7F",x"7F",x"7F",x"3F",x"3B",x"07",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2F",x"27",x"37",x"17",x"17",x"07",x"07",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"05",x"06",x"02",x"02",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"80",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"80",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"3F",x"3F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F7",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"25",x"10",x"A5",x"01",x"00",x"11",x"00",x"08",x"BF",x"52",x"29",x"06",x"F0",x"36",x"5C",x"23",
		x"A0",x"82",x"10",x"09",x"80",x"00",x"22",x"04",x"55",x"02",x"58",x"82",x"40",x"21",x"0A",x"26",
		x"FF",x"91",x"00",x"4A",x"91",x"00",x"10",x"50",x"FF",x"C4",x"4D",x"84",x"02",x"00",x"AC",x"00",
		x"81",x"72",x"1C",x"27",x"54",x"11",x"00",x"28",x"8C",x"08",x"80",x"A2",x"C4",x"74",x"9F",x"83",
		x"FF",x"30",x"0A",x"31",x"00",x"B8",x"15",x"80",x"FF",x"94",x"20",x"52",x"22",x"10",x"14",x"40",
		x"54",x"11",x"49",x"10",x"00",x"14",x"30",x"30",x"B1",x"10",x"40",x"90",x"0A",x"15",x"20",x"30",
		x"FF",x"99",x"52",x"04",x"1C",x"30",x"10",x"2A",x"28",x"14",x"00",x"44",x"40",x"08",x"00",x"20",
		x"14",x"82",x"08",x"92",x"70",x"19",x"10",x"90",x"80",x"24",x"04",x"90",x"50",x"08",x"00",x"62",
		x"00",x"02",x"00",x"0A",x"24",x"80",x"00",x"80",x"20",x"12",x"4A",x"28",x"8C",x"12",x"9A",x"43",
		x"01",x"08",x"12",x"00",x"A0",x"00",x"00",x"01",x"00",x"3A",x"80",x"10",x"53",x"02",x"29",x"0B",
		x"88",x"41",x"28",x"10",x"48",x"4D",x"02",x"08",x"84",x"04",x"80",x"00",x"0C",x"84",x"80",x"05",
		x"85",x"08",x"50",x"00",x"48",x"40",x"09",x"50",x"80",x"C0",x"A4",x"00",x"0C",x"04",x"0A",x"14",
		x"D0",x"30",x"5E",x"43",x"00",x"00",x"10",x"18",x"42",x"04",x"40",x"41",x"A8",x"70",x"08",x"4F",
		x"40",x"8A",x"10",x"14",x"21",x"B1",x"04",x"30",x"03",x"D0",x"80",x"42",x"24",x"40",x"40",x"21",
		x"14",x"10",x"00",x"90",x"04",x"D0",x"09",x"30",x"20",x"02",x"80",x"50",x"02",x"00",x"42",x"10",
		x"F0",x"72",x"34",x"77",x"09",x"12",x"91",x"30",x"10",x"08",x"80",x"02",x"80",x"18",x"00",x"48",
		x"08",x"00",x"20",x"00",x"44",x"80",x"00",x"02",x"80",x"02",x"44",x"20",x"52",x"00",x"09",x"83",
		x"00",x"00",x"00",x"08",x"20",x"00",x"82",x"80",x"00",x"44",x"00",x"02",x"0A",x"10",x"81",x"06",
		x"64",x"88",x"04",x"40",x"08",x"48",x"04",x"02",x"09",x"86",x"01",x"54",x"80",x"04",x"44",x"82",
		x"48",x"88",x"01",x"00",x"4A",x"04",x"49",x"80",x"A4",x"10",x"0D",x"84",x"94",x"20",x"04",x"84",
		x"90",x"4C",x"20",x"30",x"18",x"04",x"93",x"10",x"28",x"30",x"40",x"61",x"02",x"60",x"20",x"14",
		x"00",x"30",x"04",x"38",x"14",x"00",x"80",x"58",x"C0",x"60",x"22",x"14",x"A0",x"26",x"42",x"23",
		x"80",x"18",x"10",x"24",x"28",x"81",x"09",x"42",x"80",x"05",x"0A",x"1B",x"99",x"1B",x"D9",x"FC",
		x"01",x"02",x"29",x"07",x"84",x"04",x"23",x"01",x"7E",x"73",x"68",x"BC",x"4E",x"39",x"B4",x"DE",
		x"21",x"10",x"00",x"00",x"84",x"00",x"40",x"08",x"25",x"00",x"12",x"44",x"10",x"21",x"04",x"00",
		x"00",x"00",x"02",x"00",x"24",x"01",x"00",x"40",x"89",x"08",x"02",x"20",x"05",x"01",x"04",x"50",
		x"20",x"80",x"40",x"00",x"23",x"08",x"84",x"18",x"A5",x"00",x"14",x"82",x"00",x"84",x"04",x"00",
		x"02",x"20",x"00",x"20",x"00",x"C2",x"08",x"02",x"88",x"40",x"0D",x"00",x"80",x"46",x"01",x"01",
		x"00",x"98",x"52",x"20",x"00",x"92",x"18",x"09",x"B0",x"00",x"40",x"64",x"02",x"20",x"D0",x"08",
		x"14",x"10",x"26",x"41",x"90",x"08",x"10",x"08",x"24",x"22",x"60",x"11",x"80",x"E1",x"4A",x"A1",
		x"A4",x"0A",x"04",x"83",x"03",x"44",x"0E",x"03",x"F0",x"EE",x"3C",x"B0",x"EC",x"58",x"F6",x"BD",
		x"81",x"8E",x"81",x"43",x"34",x"0D",x"87",x"03",x"C7",x"EE",x"38",x"E0",x"DE",x"FC",x"C8",x"B7",
		x"02",x"00",x"80",x"10",x"00",x"00",x"80",x"00",x"12",x"00",x"00",x"00",x"21",x"10",x"04",x"01",
		x"00",x"00",x"02",x"20",x"00",x"00",x"00",x"44",x"10",x"00",x"08",x"02",x"00",x"41",x"04",x"00",
		x"04",x"A4",x"00",x"02",x"11",x"04",x"00",x"20",x"48",x"22",x"84",x"90",x"04",x"11",x"94",x"08",
		x"0A",x"02",x"80",x"24",x"00",x"20",x"40",x"09",x"00",x"34",x"46",x"00",x"8A",x"54",x"89",x"61",
		x"90",x"B2",x"00",x"14",x"88",x"01",x"10",x"12",x"20",x"10",x"2E",x"A8",x"44",x"46",x"22",x"21",
		x"00",x"A0",x"90",x"0C",x"14",x"13",x"04",x"30",x"10",x"21",x"B4",x"01",x"21",x"40",x"22",x"24",
		x"84",x"03",x"01",x"24",x"71",x"8F",x"0B",x"CA",x"3C",x"38",x"8B",x"D6",x"EC",x"7D",x"AB",x"EE",
		x"07",x"43",x"31",x"0C",x"87",x"03",x"23",x"86",x"F0",x"D8",x"B7",x"F8",x"EC",x"D6",x"90",x"78",
		x"00",x"80",x"00",x"00",x"00",x"80",x"08",x"00",x"01",x"12",x"80",x"01",x"24",x"82",x"08",x"01",
		x"80",x"00",x"00",x"08",x"42",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"01",x"00",x"00",x"08",
		x"02",x"08",x"51",x"00",x"2A",x"02",x"00",x"90",x"64",x"02",x"14",x"20",x"86",x"08",x"81",x"14",
		x"00",x"02",x"40",x"0C",x"80",x"01",x"04",x"19",x"62",x"01",x"82",x"0A",x"84",x"10",x"05",x"92",
		x"15",x"A2",x"10",x"01",x"70",x"10",x"A0",x"01",x"A0",x"00",x"46",x"60",x"A0",x"08",x"31",x"20",
		x"14",x"40",x"10",x"00",x"00",x"11",x"72",x"08",x"28",x"12",x"24",x"80",x"2A",x"21",x"51",x"29",
		x"50",x"A1",x"00",x"50",x"89",x"21",x"02",x"50",x"F5",x"78",x"B8",x"74",x"8E",x"30",x"F3",x"EE",
		x"80",x"18",x"21",x"80",x"51",x"21",x"12",x"62",x"14",x"30",x"F0",x"E4",x"CA",x"BD",x"FA",x"A0",
		x"00",x"80",x"00",x"80",x"00",x"02",x"80",x"00",x"24",x"00",x"00",x"02",x"00",x"08",x"00",x"41",
		x"04",x"20",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"02",x"10",x"08",x"01",x"01",x"04",
		x"04",x"40",x"08",x"20",x"01",x"40",x"02",x"00",x"00",x"10",x"82",x"00",x"00",x"04",x"42",x"00",
		x"08",x"00",x"00",x"00",x"20",x"00",x"02",x"00",x"40",x"02",x"88",x"00",x"00",x"11",x"02",x"80",
		x"0A",x"90",x"01",x"80",x"50",x"00",x"00",x"22",x"23",x"10",x"22",x"04",x"48",x"A3",x"00",x"08",
		x"41",x"14",x"02",x"00",x"10",x"20",x"02",x"04",x"52",x"10",x"22",x"02",x"95",x"00",x"04",x"0A",
		x"86",x"A0",x"50",x"93",x"A7",x"01",x"00",x"56",x"FF",x"3E",x"FC",x"78",x"6B",x"B6",x"F8",x"7C",
		x"03",x"01",x"A0",x"40",x"10",x"04",x"11",x"A1",x"38",x"FB",x"D6",x"3C",x"78",x"FB",x"D7",x"7E",
		x"FB",x"FF",x"FB",x"FE",x"EF",x"FB",x"E9",x"FE",x"FF",x"ED",x"AA",x"FA",x"FE",x"EF",x"B7",x"FF",
		x"FF",x"F2",x"EF",x"EB",x"EE",x"FA",x"F9",x"FF",x"BA",x"FE",x"AF",x"EF",x"BB",x"FE",x"FB",x"AA",
		x"FF",x"EE",x"EA",x"EF",x"FB",x"FF",x"FA",x"F9",x"FA",x"7F",x"FA",x"EB",x"FA",x"BF",x"FF",x"FB",
		x"EE",x"EE",x"F3",x"FF",x"CE",x"EB",x"EE",x"FE",x"EF",x"CA",x"EE",x"FF",x"BE",x"FB",x"BF",x"FB",
		x"BB",x"FA",x"FE",x"EB",x"FF",x"FF",x"FA",x"EB",x"BC",x"EA",x"7F",x"BB",x"BF",x"BE",x"EF",x"EB",
		x"BD",x"FE",x"BE",x"EB",x"EE",x"FF",x"BA",x"EE",x"BA",x"FF",x"EF",x"EE",x"BB",x"AF",x"EA",x"FA",
		x"FB",x"BF",x"FB",x"FE",x"EF",x"FB",x"E9",x"FE",x"FF",x"ED",x"AA",x"FA",x"FA",x"EF",x"B3",x"FF",
		x"BF",x"F2",x"EF",x"EB",x"EE",x"FA",x"FB",x"E0",x"BA",x"FE",x"AB",x"EF",x"BF",x"FE",x"FB",x"00",
		x"AF",x"4C",x"6B",x"B6",x"9D",x"C7",x"CB",x"3C",x"2D",x"16",x"AC",x"1F",x"8E",x"E8",x"5E",x"2D",
		x"56",x"B8",x"1F",x"74",x"38",x"8E",x"37",x"09",x"98",x"3E",x"6B",x"9E",x"26",x"74",x"DB",x"1E",
		x"03",x"07",x"08",x"10",x"0F",x"47",x"0A",x"3C",x"FC",x"68",x"BE",x"9D",x"C2",x"26",x"7B",x"8E",
		x"5F",x"0E",x"11",x"BB",x"7E",x"2C",x"55",x"BF",x"04",x"EF",x"DA",x"2D",x"0E",x"F4",x"86",x"67",
		x"AF",x"76",x"B8",x"1D",x"47",x"61",x"0C",x"15",x"BE",x"C4",x"62",x"F9",x"62",x"86",x"FB",x"B6",
		x"88",x"6E",x"11",x"BB",x"7E",x"25",x"07",x"3B",x"45",x"E8",x"B2",x"3C",x"DA",x"F4",x"86",x"77",
		x"33",x"C4",x"6B",x"B6",x"9D",x"47",x"CB",x"3C",x"2D",x"16",x"AD",x"1F",x"8E",x"E8",x"5E",x"2D",
		x"56",x"B8",x"1F",x"74",x"38",x"8E",x"37",x"09",x"98",x"3E",x"6B",x"9E",x"26",x"74",x"DB",x"1E",
		x"29",x"D4",x"6B",x"B7",x"1E",x"35",x"EB",x"3F",x"3D",x"96",x"E4",x"28",x"1C",x"C0",x"78",x"C8",
		x"58",x"B6",x"1E",x"70",x"6C",x"FF",x"74",x"09",x"F2",x"30",x"C0",x"B0",x"7C",x"70",x"DF",x"16",
		x"00",x"00",x"00",x"02",x"02",x"08",x"07",x"00",x"00",x"00",x"00",x"40",x"00",x"80",x"60",x"B0",
		x"00",x"07",x"08",x"02",x"04",x"01",x"02",x"00",x"A0",x"10",x"50",x"A0",x"40",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"00",x"24",x"13",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"05",x"38",x"02",x"05",x"02",x"08",x"10",x"80",x"00",x"80",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"04",x"1C",x"1C",x"1C",x"00",x"00",
		x"00",x"00",x"04",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"04",x"1C",x"1C",x"1C",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"EF",x"AF",x"AF",x"AF",x"3F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"7F",x"2F",x"2F",x"2F",x"AF",x"BF",x"BF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"05",x"05",x"01",x"08",x"08",x"0A",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"02",x"08",x"08",x"09",x"09",x"09",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",
		x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"FF",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"FF",
		x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",
		x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"FF",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"FF",
		x"FF",x"7F",x"33",x"19",x"0C",x"06",x"03",x"01",x"FF",x"FF",x"33",x"99",x"CC",x"66",x"33",x"99",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CC",x"66",x"33",x"19",x"0C",x"06",x"03",x"01",
		x"FF",x"FF",x"33",x"99",x"CC",x"66",x"33",x"99",x"FF",x"FF",x"33",x"99",x"CC",x"66",x"33",x"99",
		x"CC",x"66",x"33",x"99",x"CC",x"66",x"33",x"FF",x"CC",x"66",x"33",x"99",x"CC",x"66",x"33",x"FF",
		x"FF",x"FF",x"33",x"FF",x"CC",x"CC",x"CC",x"FF",x"FF",x"FF",x"33",x"FF",x"CC",x"CC",x"CC",x"FF",
		x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",
		x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",
		x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",x"CC",x"CC",x"CC",x"FF",
		x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
		x"AA",x"AA",x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"AA",x"00",x"00",x"00",x"00",x"00",x"00",
		x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
		x"AA",x"AA",x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"AA",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"92",x"92",x"92",x"92",x"92",x"FF",x"FF",x"FF",x"49",x"49",x"49",x"49",x"49",
		x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
		x"FF",x"FF",x"FF",x"FF",x"3F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"14",x"1F",x"00",x"11",x"0A",x"04",x"1F",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"1F",x"04",x"55",x"5F",x"55",x"55",x"55",x"55",
		x"55",x"55",x"55",x"00",x"00",x"00",x"00",x"00",x"5F",x"55",x"55",x"10",x"1F",x"10",x"10",x"00",
		x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
		x"92",x"92",x"92",x"92",x"92",x"FF",x"FF",x"FF",x"49",x"49",x"49",x"49",x"49",x"FF",x"FF",x"FF",
		x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
		x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"47",x"44",x"44",x"44",x"44",x"44",
		x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"C0",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",
		x"00",x"00",x"7E",x"7E",x"7E",x"7F",x"7E",x"7E",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",
		x"7F",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"C4",x"C4",x"C4",x"C4",x"C0",x"00",x"00",x"00",
		x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"47",x"44",x"44",x"44",x"44",x"44",
		x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F3",x"B3",x"F3",x"B3",x"FF",x"B3",x"F3",x"F3",x"33",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",x"38",x"38",x"38",x"3F",x"F8",x"38",x"38",x"38",
		x"FF",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",x"F8",x"38",x"38",x"3F",x"F8",x"38",x"38",x"38",
		x"FF",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",x"F8",x"38",x"38",x"3F",x"F8",x"38",x"38",x"38",
		x"FF",x"B3",x"F3",x"B3",x"FF",x"B3",x"F3",x"B3",x"FF",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",
		x"FF",x"B3",x"F3",x"B3",x"FF",x"B3",x"F3",x"B3",x"FF",x"33",x"33",x"33",x"FF",x"33",x"33",x"33",
		x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"EF",x"8F",x"1F",x"3F",x"3F",x"7F",x"FF",x"7F",
		x"80",x"82",x"C1",x"83",x"81",x"00",x"8B",x"19",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"7F",x"7F",x"7E",x"7E",x"7C",x"79",x"73",x"BF",x"7F",x"3F",x"3F",x"FF",x"DF",x"DF",x"9F",
		x"4F",x"7E",x"78",x"74",x"60",x"78",x"70",x"64",x"9F",x"0F",x"1F",x"3F",x"3F",x"1F",x"0F",x"27",
		x"1C",x"3A",x"3C",x"3C",x"7C",x"3E",x"3C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"34",x"3C",x"3E",x"3C",x"3C",x"34",x"7E",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"0C",x"0C",x"1C",
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"0A",x"3E",x"9E",x"8E",x"1F",x"FE",x"AF",x"9F",x"BF",
		x"00",x"00",x"00",x"00",x"43",x"C7",x"C7",x"CF",x"00",x"00",x"00",x"0C",x"1E",x"7E",x"FE",x"BE",
		x"CF",x"DF",x"47",x"43",x"40",x"21",x"47",x"7F",x"BE",x"BE",x"CE",x"9F",x"BE",x"BE",x"9E",x"9E",
		x"76",x"66",x"EF",x"EF",x"FF",x"FF",x"FF",x"FC",x"37",x"73",x"79",x"7C",x"7E",x"FE",x"FE",x"FC",
		x"F0",x"FC",x"FE",x"FF",x"FE",x"FF",x"7F",x"7F",x"00",x"0E",x"3F",x"7F",x"3F",x"1F",x"3F",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"02",x"06",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0E",x"0E",x"0E",x"06",x"02",x"00",x"01",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"BF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"0F",x"03",x"01",x"00",x"01",x"00",x"01",
		x"3F",x"9F",x"8E",x"9F",x"BF",x"BF",x"9F",x"FF",x"8E",x"1E",x"9E",x"5E",x"3E",x"BE",x"FE",x"FE",
		x"D7",x"DB",x"DB",x"F3",x"DB",x"B3",x"CB",x"DB",x"FC",x"FE",x"FC",x"FC",x"FE",x"FF",x"FF",x"FF",
		x"7F",x"7F",x"7C",x"7F",x"7F",x"7F",x"7F",x"7F",x"3F",x"2F",x"37",x"1F",x"B7",x"B7",x"3F",x"9B",
		x"7F",x"7F",x"3F",x"3F",x"1F",x"00",x"00",x"03",x"BF",x"1F",x"8E",x"80",x"00",x"2C",x"FE",x"E6",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"0B",x"0F",x"1F",x"3F",x"3F",x"03",x"FC",x"F0",
		x"01",x"03",x"03",x"03",x"03",x"01",x"01",x"01",x"8F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F4",x"F0",x"F0",x"F0",x"F0",x"F8",x"FC",x"FC",x"0E",x"0E",x"04",x"00",x"00",x"00",x"00",x"01",
		x"FE",x"FF",x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"02",x"EC",x"FE",x"3F",x"1F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"30",x"30",x"38",x"3C",x"38",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"30",
		x"30",x"30",x"38",x"38",x"BD",x"FD",x"FD",x"FD",x"78",x"78",x"78",x"F8",x"F8",x"F8",x"FC",x"FC",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"0F",x"3F",x"3F",x"5F",x"5F",x"FF",
		x"00",x"01",x"01",x"03",x"03",x"07",x"1F",x"7F",x"EF",x"EF",x"FF",x"FF",x"FF",x"EF",x"FF",x"E7",
		x"3F",x"7F",x"71",x"70",x"60",x"28",x"2E",x"7D",x"FE",x"FE",x"FF",x"0F",x"03",x"01",x"00",x"00",
		x"7D",x"6F",x"67",x"73",x"73",x"7D",x"7C",x"7E",x"C1",x"C1",x"E1",x"C1",x"E1",x"F9",x"F9",x"FC",
		x"38",x"30",x"30",x"30",x"20",x"20",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"C0",x"C0",x"80",x"00",x"00",x"00",x"03",x"03",x"03",x"03",x"0D",x"1D",x"0D",x"19",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FB",x"FB",x"FF",x"7F",x"7F",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7F",x"7F",x"3F",x"3F",x"20",x"10",x"08",
		x"F2",x"F1",x"F8",x"FE",x"FE",x"F7",x"F7",x"FF",x"07",x"07",x"0F",x"0E",x"2E",x"2E",x"7F",x"7E",
		x"FF",x"FB",x"FB",x"FD",x"FF",x"05",x"06",x"06",x"FF",x"FF",x"FF",x"FF",x"1F",x"4F",x"AB",x"FF",
		x"FD",x"FD",x"FE",x"FE",x"FE",x"FF",x"FF",x"7F",x"F8",x"F8",x"F8",x"F8",x"F0",x"70",x"70",x"60",
		x"7E",x"78",x"E0",x"80",x"C0",x"80",x"C0",x"80",x"18",x"70",x"80",x"00",x"00",x"00",x"01",x"01",
		x"00",x"00",x"00",x"00",x"07",x"3F",x"7F",x"3F",x"01",x"0F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"3F",x"7F",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"77",x"13",x"3F",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"E7",x"E7",x"E3",x"E1",x"E1",
		x"FF",x"3F",x"0D",x"81",x"41",x"47",x"CF",x"CF",x"E1",x"E0",x"F3",x"A7",x"33",x"3F",x"7F",x"FF",
		x"76",x"66",x"62",x"63",x"71",x"78",x"7F",x"7F",x"1C",x"1C",x"08",x"80",x"20",x"28",x"F8",x"F0",
		x"7F",x"7F",x"7F",x"3F",x"3F",x"3F",x"3F",x"1F",x"F8",x"F8",x"80",x"E0",x"E0",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"16",x"1E",x"0A",x"15",x"0B",x"1F",x"2B",x"1F",
		x"02",x"07",x"0F",x"0F",x"0F",x"3F",x"3F",x"3F",x"17",x"2F",x"1B",x"2F",x"3F",x"3F",x"7F",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"03",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"06",x"03",x"C1",x"70",x"1C",x"07",x"01",x"00",x"61",x"01",x"F0",x"00",x"00",x"00",x"80",x"78",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"F0",x"1E",x"03",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"81",x"E1",x"1D",x"03",
		x"E9",x"FF",x"EF",x"CE",x"C8",x"C0",x"C0",x"C0",x"FF",x"F9",x"80",x"00",x"00",x"00",x"00",x"02",
		x"C0",x"C0",x"80",x"81",x"82",x"1D",x"52",x"6A",x"0F",x"04",x"6A",x"4A",x"15",x"5A",x"AD",x"DA",
		x"DF",x"EF",x"7F",x"1F",x"0F",x"07",x"03",x"01",x"FD",x"FB",x"FF",x"FD",x"FD",x"FB",x"FF",x"FD",
		x"C1",x"F8",x"5E",x"A7",x"2B",x"55",x"6D",x"92",x"FF",x"FF",x"FB",x"FE",x"FE",x"FC",x"FD",x"FF",
		x"FC",x"FE",x"FE",x"FF",x"F6",x"FD",x"F4",x"F4",x"DF",x"DF",x"DF",x"DF",x"BF",x"9F",x"BF",x"BF",
		x"F0",x"F2",x"F5",x"E8",x"E2",x"F3",x"7B",x"7B",x"BF",x"9F",x"9F",x"5F",x"EF",x"6E",x"6E",x"B6",
		x"9F",x"9F",x"8F",x"8F",x"BF",x"9F",x"BF",x"9F",x"F0",x"F0",x"F8",x"F4",x"F0",x"F8",x"FC",x"F8",
		x"9F",x"BF",x"BE",x"9E",x"82",x"FF",x"FE",x"FE",x"E8",x"F0",x"F0",x"73",x"E7",x"F7",x"F3",x"FB",
		x"37",x"6E",x"6E",x"7C",x"5C",x"FE",x"FE",x"FD",x"FF",x"7F",x"F7",x"FF",x"FD",x"FF",x"FF",x"FF",
		x"F9",x"F9",x"FB",x"F9",x"FB",x"F3",x"F7",x"EF",x"FD",x"FF",x"EF",x"FF",x"FF",x"F7",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"02",x"14",x"03",x"4A",
		x"00",x"01",x"01",x"03",x"09",x"00",x"05",x"50",x"22",x"28",x"22",x"64",x"20",x"89",x"A2",x"CA",
		x"85",x"10",x"44",x"A5",x"0C",x"44",x"91",x"00",x"3F",x"7F",x"1F",x"1F",x"4F",x"57",x"63",x"41",
		x"24",x"84",x"84",x"A9",x"04",x"A0",x"62",x"24",x"42",x"14",x"84",x"05",x"08",x"44",x"C4",x"69",
		x"7B",x"7B",x"79",x"BD",x"FD",x"DF",x"DF",x"C3",x"36",x"17",x"0E",x"9B",x"03",x"87",x"87",x"83",
		x"F7",x"73",x"BB",x"3B",x"BB",x"1D",x"4F",x"97",x"01",x"80",x"D0",x"F6",x"F7",x"FF",x"FF",x"FF",
		x"7F",x"7F",x"7F",x"FF",x"87",x"E7",x"E7",x"E7",x"F8",x"F8",x"F8",x"FC",x"FE",x"FC",x"F8",x"E1",
		x"F3",x"F9",x"68",x"84",x"C0",x"F0",x"E0",x"FF",x"E3",x"CF",x"87",x"C3",x"49",x"26",x"27",x"83",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"04",x"06",x"10",x"15",
		x"00",x"00",x"01",x"05",x"05",x"05",x"15",x"56",x"54",x"5E",x"14",x"44",x"54",x"72",x"55",x"55",
		x"52",x"85",x"52",x"22",x"4B",x"C4",x"40",x"54",x"50",x"12",x"15",x"80",x"15",x"98",x"25",x"92",
		x"24",x"41",x"44",x"82",x"54",x"44",x"44",x"8A",x"80",x"0C",x"45",x"94",x"90",x"91",x"44",x"81",
		x"91",x"07",x"63",x"07",x"13",x"A3",x"27",x"47",x"74",x"F4",x"F5",x"3B",x"9F",x"99",x"98",x"D8",
		x"47",x"93",x"23",x"8B",x"23",x"21",x"2D",x"43",x"DE",x"FE",x"DE",x"FC",x"FC",x"FC",x"FF",x"FF",
		x"FE",x"FE",x"FF",x"F8",x"FE",x"FF",x"FF",x"FF",x"43",x"33",x"38",x"3F",x"3F",x"3F",x"07",x"0F",
		x"FC",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF",x"9F",x"9F",x"87",x"9D",x"85",x"8D",x"BD",x"99",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"05",x"0D",x"15",
		x"00",x"00",x"00",x"05",x"0C",x"1E",x"3E",x"3F",x"11",x"4C",x"05",x"C7",x"61",x"11",x"54",x"D5",
		x"51",x"5D",x"55",x"75",x"75",x"56",x"55",x"91",x"55",x"35",x"55",x"55",x"57",x"55",x"54",x"5D",
		x"55",x"45",x"0D",x"15",x"55",x"51",x"56",x"75",x"15",x"50",x"B5",x"C5",x"47",x"55",x"55",x"5D",
		x"0D",x"51",x"01",x"09",x"83",x"21",x"29",x"20",x"FF",x"DF",x"DF",x"DF",x"FF",x"FF",x"EF",x"EE",
		x"42",x"92",x"06",x"24",x"00",x"88",x"20",x"A2",x"E4",x"69",x"6C",x"7E",x"76",x"B6",x"B7",x"17",
		x"F3",x"E3",x"C3",x"E3",x"E3",x"83",x"01",x"01",x"85",x"83",x"81",x"83",x"87",x"9F",x"C3",x"C1",
		x"00",x"90",x"C0",x"C0",x"F4",x"F0",x"F0",x"DC",x"E1",x"E1",x"FD",x"F9",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"5F",
		x"00",x"01",x"03",x"07",x"0F",x"1F",x"3B",x"7B",x"DB",x"D9",x"FC",x"3E",x"3E",x"5A",x"DA",x"DA",
		x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF",x"FF",x"C6",x"D5",x"CD",x"C9",x"D4",x"C5",x"CA",x"CE",
		x"EF",x"DF",x"5F",x"7F",x"DF",x"DD",x"DD",x"DC",x"85",x"89",x"85",x"8E",x"8D",x"C5",x"E1",x"F1",
		x"0A",x"41",x"53",x"02",x"24",x"82",x"02",x"52",x"27",x"17",x"11",x"58",x"01",x"94",x"20",x"02",
		x"40",x"88",x"42",x"62",x"40",x"08",x"90",x"42",x"90",x"31",x"10",x"90",x"16",x"03",x"42",x"12",
		x"DF",x"5F",x"50",x"40",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"C3",x"FC",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"05",x"0D",x"15",x"37",x"3E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"25",x"3D",x"1D",x"0D",x"07",x"03",x"01",
		x"FB",x"FB",x"7B",x"7D",x"5D",x"59",x"5B",x"DB",x"B7",x"BF",x"B7",x"B7",x"BD",x"BD",x"DF",x"DF",
		x"FB",x"DA",x"DE",x"FA",x"EB",x"BB",x"AF",x"AB",x"DE",x"DE",x"DD",x"FD",x"FD",x"7D",x"7F",x"7F",
		x"DD",x"ED",x"DD",x"D9",x"DB",x"53",x"57",x"5E",x"F5",x"F1",x"E1",x"FA",x"F5",x"F3",x"F0",x"F1",
		x"7E",x"5F",x"4F",x"5B",x"5D",x"DE",x"DD",x"FB",x"F9",x"78",x"5C",x"7D",x"F4",x"FD",x"F1",x"71",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"EB",x"7F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"6F",x"6F",x"6B",x"6B",x"EE",x"FE",x"FF",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"00",
		x"D7",x"D6",x"D6",x"DE",x"FF",x"F7",x"F7",x"D5",x"59",x"79",x"79",x"E1",x"C6",x"C5",x"C1",x"40",
		x"C4",x"C4",x"C1",x"C4",x"C1",x"C9",x"41",x"01",x"51",x"19",x"59",x"15",x"74",x"40",x"16",x"54",
		x"1C",x"0D",x"03",x"01",x"00",x"00",x"00",x"00",x"D5",x"54",x"13",x"7D",x"D5",x"45",x"34",x"0D",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"03",x"01",x"00",x"00",x"00",x"00",x"00",
		x"51",x"1D",x"75",x"D5",x"56",x"57",x"55",x"55",x"65",x"53",x"17",x"13",x"5B",x"57",x"57",x"D7",
		x"65",x"11",x"15",x"55",x"15",x"14",x"0D",x"01",x"46",x"5D",x"54",x"55",x"B8",x"58",x"58",x"52",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B8",x"54",x"48",x"58",x"05",x"08",x"06",x"02",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"24",x"82",x"2A",x"02",x"49",x"9A",x"21",x"22",x"21",x"08",x"88",x"1B",x"48",x"4C",x"49",x"28",
		x"AA",x"02",x"22",x"08",x"02",x"04",x"01",x"00",x"40",x"08",x"B0",x"62",x"28",x"28",x"88",x"26",
		x"59",x"49",x"7B",x"68",x"C8",x"48",x"E0",x"C4",x"FE",x"FE",x"7E",x"FF",x"7E",x"7F",x"3E",x"0F",
		x"A5",x"C9",x"DD",x"DF",x"CF",x"87",x"8F",x"DF",x"06",x"3F",x"FF",x"FD",x"FC",x"FE",x"7E",x"FE",
		x"DD",x"D9",x"D9",x"D8",x"DC",x"DC",x"D8",x"CC",x"FF",x"FF",x"DF",x"FF",x"FE",x"FE",x"DE",x"EE",
		x"88",x"9C",x"C8",x"CC",x"E4",x"E4",x"E0",x"E8",x"E5",x"FC",x"4E",x"5C",x"EE",x"5E",x"CE",x"DE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"FF",x"00",x"00",x"30",x"30",x"3B",x"1B",x"FD",x"FD",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"10",x"20",x"28",x"FF",x"FF",x"FF",x"FF",x"00",x"40",x"30",x"3B",x"FD",x"FD",x"FD",x"FD",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"02",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"E0",x"FC",x"E7",x"FF",x"E6",x"FF",x"E7",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"00",x"00",x"00",
		x"01",x"00",x"03",x"87",x"0F",x"3F",x"FF",x"FF",x"F0",x"FC",x"FD",x"FE",x"FE",x"FE",x"FE",x"FE",
		x"04",x"03",x"3F",x"FF",x"FF",x"FF",x"7E",x"1C",x"80",x"FF",x"3F",x"FF",x"3F",x"F8",x"8C",x"8F",
		x"04",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"8F",x"8F",x"FF",x"FF",x"8F",x"8F",
		x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
		x"FF",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"FF",
		x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"F8",x"04",x"04",x"0F",
		x"FE",x"FF",x"FF",x"F7",x"FB",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",
		x"00",x"40",x"F0",x"FA",x"FE",x"00",x"3F",x"FF",x"00",x"0A",x"77",x"BF",x"FC",x"01",x"FF",x"3F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"F3",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF",x"F9",x"F9",x"FF",
		x"00",x"00",x"80",x"60",x"00",x"E0",x"98",x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FC",x"FB",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"D0",x"F4",x"FB",x"FF",x"FF",x"FF",
		x"20",x"FF",x"20",x"00",x"00",x"00",x"00",x"00",x"1F",x"FF",x"1F",x"03",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"01",x"00",x"FD",x"FD",x"FC",x"FC",x"F8",x"F8",x"F0",x"30",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"03",x"0F",x"0F",x"03",x"23",x"2F",x"FD",x"FD",x"FD",x"FC",x"FC",x"FC",x"F8",x"F0",
		x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"01",x"03",
		x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"02",x"FF",x"E7",x"C0",x"40",x"40",x"40",x"40",x"C0",
		x"01",x"07",x"1F",x"3F",x"7F",x"FF",x"FF",x"FE",x"80",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"00",
		x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"0E",x"FF",x"FE",x"FE",x"FE",x"00",x"00",x"03",x"0E",x"F8",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"70",x"F8",
		x"FF",x"FF",x"00",x"00",x"00",x"FC",x"04",x"04",x"FF",x"FF",x"8F",x"8F",x"FF",x"07",x"07",x"07",
		x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"E0",x"E0",x"FF",x"7F",x"00",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"55",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"57",
		x"55",x"55",x"55",x"55",x"D5",x"D5",x"7F",x"7F",x"57",x"57",x"57",x"57",x"57",x"56",x"FE",x"FE",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FB",x"07",x"1F",x"1F",x"07",x"07",x"1F",x"DF",
		x"8F",x"8F",x"0F",x"0F",x"0F",x"0E",x"0E",x"0E",x"FF",x"F8",x"C0",x"C6",x"C6",x"06",x"3E",x"3C",
		x"D0",x"10",x"50",x"10",x"50",x"10",x"50",x"10",x"01",x"03",x"02",x"03",x"00",x"03",x"02",x"03",
		x"50",x"1F",x"D0",x"50",x"D0",x"50",x"D0",x"41",x"00",x"FF",x"00",x"00",x"00",x"7C",x"7F",x"FF",
		x"00",x"F7",x"17",x"F7",x"07",x"F7",x"17",x"F7",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"07",x"FF",x"07",x"07",x"07",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F8",x"F0",x"F8",x"FC",x"F8",x"F8",x"F0",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F8",x"FC",x"F8",x"FC",x"FC",x"FE",x"FC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"07",x"0F",x"0F",x"1F",x"7F",x"3F",x"8F",x"E3",
		x"0F",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FE",x"FF",x"7F",x"1F",x"0F",x"03",x"00",
		x"FC",x"F8",x"F0",x"E0",x"C0",x"E0",x"F0",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FC",x"7E",x"3F",x"8F",x"E3",x"F9",x"FC",x"FE",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"78",
		x"3F",x"38",x"38",x"7F",x"70",x"70",x"7F",x"38",x"FC",x"7C",x"7C",x"FC",x"7C",x"7C",x"FC",x"7C",
		x"38",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"7C",x"FC",x"F8",x"70",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"03",
		x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"0F",x"0E",x"2E",x"6E",x"EE",x"EE",x"EE",x"EF",x"EF",
		x"1F",x"3F",x"7F",x"E1",x"E1",x"FF",x"E1",x"E1",x"EF",x"EE",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",
		x"00",x"01",x"11",x"01",x"0F",x"8F",x"0E",x"7C",x"38",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",
		x"0E",x"EF",x"6F",x"61",x"1D",x"0D",x"8C",x"8F",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"38",x"BC",
		x"FE",x"FF",x"00",x"01",x"00",x"01",x"00",x"01",x"07",x"8F",x"3F",x"BC",x"18",x"B8",x"38",x"98",
		x"00",x"01",x"00",x"01",x"00",x"01",x"FE",x"FF",x"38",x"B8",x"18",x"BC",x"3F",x"8F",x"07",x"FF",
		x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"07",x"FF",x"3F",x"07",x"00",x"02",x"02",x"3F",x"FF",x"FF",x"FF",x"FF",x"FE",
		x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"0E",x"00",x"00",x"03",x"FF",x"0F",x"03",x"00",
		x"FF",x"7B",x"7B",x"7B",x"7B",x"7B",x"7B",x"00",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
		x"00",x"07",x"3F",x"FF",x"FF",x"FC",x"FC",x"38",x"1F",x"E0",x"F7",x"F7",x"F7",x"00",x"00",x"00",
		x"00",x"F3",x"E7",x"8F",x"FF",x"FE",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",
		x"FF",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"00",x"FC",x"F8",x"F1",x"07",x"3F",x"1F",
		x"00",x"FF",x"FE",x"F8",x"F0",x"00",x"F0",x"00",x"00",x"00",x"00",x"1F",x"01",x"3E",x"7E",x"FD",
		x"F1",x"03",x"F3",x"F7",x"F7",x"F7",x"F7",x"F3",x"FB",x"F7",x"EF",x"DF",x"DE",x"FC",x"F9",x"F3",
		x"00",x"00",x"00",x"3F",x"21",x"00",x"30",x"30",x"0F",x"00",x"00",x"7C",x"44",x"00",x"60",x"60",
		x"30",x"B0",x"B0",x"30",x"30",x"FF",x"FF",x"0E",x"60",x"60",x"60",x"60",x"60",x"FF",x"FF",x"1C",
		x"FF",x"7F",x"7F",x"7F",x"7F",x"3F",x"BF",x"DF",x"BE",x"86",x"F6",x"F6",x"F0",x"FF",x"FF",x"FF",
		x"DF",x"CF",x"CF",x"CF",x"CF",x"F7",x"F7",x"37",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"C4",x"84",
		x"50",x"D0",x"50",x"D0",x"50",x"DF",x"10",x"50",x"7F",x"7D",x"00",x"00",x"00",x"FF",x"00",x"03",
		x"10",x"50",x"10",x"50",x"10",x"50",x"00",x"7F",x"02",x"03",x"00",x"03",x"02",x"00",x"01",x"FF",
		x"FF",x"FF",x"07",x"07",x"07",x"FF",x"05",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"B5",x"20",x"00",
		x"14",x"F0",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"F4",x"F8",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"83",x"81",x"80",x"80",x"80",x"00",x"00",x"00",x"E7",x"C6",x"C6",x"63",x"31",x"38",x"3C",x"3E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0E",x"0C",x"0C",x"0E",x"0E",x"FF",x"7F",x"7F",x"1C",x"18",x"18",x"1C",x"1C",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"37",x"36",x"35",x"37",x"37",x"F7",x"F7",x"FF",x"0F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7B",x"3B",x"07",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"E5",x"E4",x"3F",x"36",x"F8",x"F0",x"C0",x"30",x"00",x"00",
		x"F0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"1C",x"78",x"F4",x"F8",x"F8",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"AA",x"15",x"AA",x"54",x"AA",x"51",x"A8",x"54",x"A2",x"45",x"AA",x"50",x"8A",x"44",x"A2",x"55",
		x"2A",x"50",x"A2",x"40",x"AA",x"50",x"28",x"00",x"AA",x"54",x"AA",x"45",x"A8",x"54",x"AA",x"00",
		x"A2",x"50",x"AA",x"01",x"AA",x"41",x"0A",x"41",x"A0",x"40",x"2A",x"01",x"0A",x"10",x"AA",x"41",
		x"A8",x"00",x"A8",x"41",x"AA",x"55",x"20",x"00",x"8A",x"55",x"AA",x"40",x"AA",x"00",x"00",x"00",
		x"BF",x"FF",x"FF",x"7F",x"BF",x"7F",x"FF",x"7F",x"FD",x"FC",x"FE",x"F0",x"E9",x"E2",x"FF",x"FE",
		x"FF",x"FF",x"FF",x"7F",x"FF",x"7F",x"BF",x"5F",x"C8",x"82",x"D0",x"FB",x"FE",x"D1",x"E0",x"D2",
		x"FF",x"7E",x"BD",x"FE",x"FE",x"7F",x"BF",x"7F",x"E4",x"08",x"45",x"31",x"40",x"9A",x"F4",x"40",
		x"FF",x"7E",x"FC",x"F8",x"FD",x"7E",x"FF",x"7F",x"B5",x"04",x"90",x"B0",x"49",x"02",x"04",x"FE",
		x"C7",x"97",x"A3",x"43",x"13",x"51",x"B1",x"11",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"09",x"89",x"8C",x"2C",x"26",x"06",x"47",x"4F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"BF",x"7F",x"FF",x"7F",x"FF",x"7F",x"FF",x"7F",x"FC",x"FA",x"D1",x"E3",x"F8",x"F9",x"FC",x"EE",
		x"BF",x"7F",x"BF",x"7F",x"BF",x"7F",x"FF",x"7F",x"FD",x"E8",x"E0",x"F9",x"F2",x"FA",x"FE",x"F8",
		x"01",x"06",x"83",x"47",x"6F",x"7F",x"3E",x"E5",x"80",x"00",x"00",x"C0",x"E0",x"26",x"19",x"0C",
		x"C8",x"A0",x"42",x"00",x"20",x"AC",x"0F",x"01",x"06",x"41",x"00",x"1B",x"26",x"08",x"18",x"C0",
		x"0A",x"0F",x"1A",x"15",x"20",x"03",x"01",x"44",x"04",x"0B",x"1C",x"0C",x"04",x"60",x"C0",x"20",
		x"D0",x"10",x"32",x"5C",x"0C",x"05",x"02",x"0A",x"11",x"26",x"47",x"4E",x"92",x"05",x"02",x"00",
		x"AA",x"15",x"AA",x"54",x"AA",x"51",x"A8",x"54",x"A2",x"45",x"AA",x"50",x"8A",x"44",x"A2",x"55",
		x"2A",x"50",x"A2",x"40",x"AA",x"00",x"28",x"15",x"AA",x"54",x"AA",x"45",x"A8",x"54",x"A2",x"00",
		x"AA",x"44",x"AA",x"45",x"2A",x"15",x"AA",x"11",x"AA",x"55",x"AA",x"40",x"AA",x"15",x"AA",x"51",
		x"AA",x"44",x"A2",x"15",x"8A",x"01",x"AA",x"14",x"AA",x"40",x"AA",x"55",x"AA",x"51",x"AA",x"51",
		x"88",x"72",x"78",x"32",x"B9",x"1B",x"D3",x"07",x"03",x"17",x"9E",x"FC",x"FE",x"F8",x"FF",x"FC",
		x"8F",x"6F",x"BF",x"5F",x"BF",x"7F",x"BF",x"7F",x"FC",x"F8",x"F8",x"F0",x"FE",x"F8",x"F0",x"F8",
		x"01",x"03",x"01",x"00",x"01",x"03",x"03",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"01",x"03",x"07",x"01",x"01",x"09",x"09",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"38",x"00",x"38",x"00",x"38",x"00",x"00",x"00",x"3F",x"3F",x"BF",x"BF",x"7F",x"3F",
		x"38",x"00",x"38",x"00",x"38",x"00",x"38",x"00",x"3F",x"BF",x"BF",x"7F",x"3F",x"3F",x"BF",x"BF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"38",x"00",x"38",x"00",x"38",x"00",x"38",x"3F",x"7F",x"3F",x"3F",x"BF",x"BF",x"7F",x"3F",x"3F",
		x"1F",x"1F",x"1E",x"1F",x"1E",x"17",x"17",x"16",x"BF",x"80",x"EF",x"EF",x"EF",x"E0",x"80",x"C0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"1F",x"FF",x"FF",x"FF",x"3F",x"00",x"00",x"FF",x"FF",x"FF",x"BF",x"DF",x"FF",x"0F",x"00",
		x"04",x"17",x"16",x"1F",x"17",x"1F",x"1E",x"16",x"40",x"E0",x"E7",x"E3",x"EF",x"EF",x"E0",x"C0",
		x"00",x"1E",x"16",x"17",x"17",x"17",x"1F",x"13",x"40",x"C0",x"E0",x"EF",x"EF",x"EF",x"6F",x"3F",
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"3D",x"3F",x"FF",x"FF",x"FF",x"F7",x"EF",x"FF",
		x"07",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",
		x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"3F",x"BF",x"BF",x"7F",x"3F",x"3F",x"BF",x"BF",
		x"38",x"00",x"38",x"00",x"38",x"00",x"38",x"00",x"7F",x"3F",x"3F",x"BF",x"BF",x"7F",x"3F",x"3F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"38",x"00",x"38",x"00",x"38",x"00",x"38",x"00",x"BF",x"BF",x"7F",x"3F",x"3F",x"BF",x"BF",x"7F",
		x"38",x"00",x"38",x"00",x"38",x"00",x"38",x"00",x"3F",x"3F",x"BF",x"BF",x"7F",x"3F",x"3F",x"BF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"03",x"07",x"07",x"07",x"0F",x"0F",
		x"7C",x"44",x"FC",x"C4",x"FF",x"FF",x"E7",x"FF",x"BF",x"7F",x"00",x"BF",x"BF",x"BF",x"FF",x"FF",
		x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"FF",x"C0",x"80",x"BF",x"BF",x"BF",x"FF",x"FF",
		x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7F",x"FF",x"FF",x"FF",x"7F",x"37",x"0F",
		x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"FF",x"C0",x"80",x"BF",x"BF",x"BF",x"FF",x"FF",
		x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"FF",x"C0",x"80",x"BF",x"BF",x"BF",x"FF",x"FF",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"03",x"03",x"01",x"01",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"7F",x"7F",x"7F",x"3F",x"3F",x"0F",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"1F",x"1F",x"07",x"07",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"07",x"03",x"03",x"00",x"00",
		x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"FF",x"C0",x"80",x"BF",x"BF",x"BF",x"FF",x"FF",
		x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"E7",x"FF",x"FF",x"C0",x"80",x"BF",x"BF",x"BF",x"80",x"00",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",
		x"C0",x"00",x"00",x"00",x"07",x"03",x"03",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"03",x"01",x"03",x"01",x"03",x"01",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"08",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"24",x"90",x"84",x"11",x"80",x"10",x"02",x"00",x"BF",x"06",x"00",x"2A",x"C2",x"3B",x"08",x"03",
		x"20",x"86",x"11",x"21",x"02",x"00",x"B0",x"05",x"01",x"0A",x"00",x"03",x"40",x"10",x"02",x"63",
		x"FF",x"12",x"08",x"00",x"10",x"02",x"80",x"10",x"FF",x"8C",x"04",x"A6",x"00",x"40",x"84",x"25",
		x"C0",x"60",x"1C",x"17",x"11",x"10",x"00",x"A4",x"84",x"00",x"C0",x"84",x"C4",x"74",x"94",x"A7",
		x"DF",x"10",x"50",x"14",x"00",x"10",x"10",x"80",x"D7",x"10",x"00",x"18",x"20",x"10",x"91",x"50",
		x"34",x"11",x"00",x"12",x"10",x"10",x"80",x"10",x"10",x"14",x"40",x"30",x"00",x"14",x"00",x"91",
		x"FF",x"10",x"12",x"10",x"15",x"90",x"10",x"22",x"28",x"00",x"08",x"40",x"00",x"00",x"00",x"04",
		x"11",x"10",x"48",x"12",x"10",x"14",x"10",x"30",x"00",x"20",x"04",x"A0",x"10",x"00",x"00",x"28",
		x"00",x"82",x"04",x"0A",x"20",x"80",x"00",x"00",x"28",x"42",x"6A",x"08",x"A4",x"02",x"92",x"41",
		x"20",x"0A",x"82",x"00",x"20",x"01",x"00",x"21",x"10",x"2A",x"A9",x"00",x"52",x"12",x"09",x"0D",
		x"88",x"44",x"68",x"10",x"48",x"0C",x"0A",x"0A",x"84",x"04",x"90",x"01",x"04",x"84",x"80",x"44",
		x"80",x"08",x"44",x"00",x"08",x"52",x"08",x"C0",x"82",x"C0",x"A4",x"00",x"2C",x"04",x"02",x"05",
		x"D1",x"70",x"1C",x"03",x"02",x"08",x"10",x"90",x"40",x"00",x"44",x"40",x"C0",x"70",x"0C",x"47",
		x"20",x"80",x"10",x"54",x"03",x"10",x"08",x"10",x"81",x"44",x"00",x"40",x"00",x"40",x"C8",x"00",
		x"90",x"10",x"22",x"10",x"90",x"90",x"24",x"30",x"00",x"04",x"00",x"01",x"20",x"00",x"00",x"00",
		x"D0",x"70",x"1C",x"37",x"81",x"10",x"18",x"50",x"04",x"90",x"00",x"00",x"C4",x"01",x"00",x"60",
		x"00",x"80",x"20",x"00",x"14",x"80",x"00",x"00",x"90",x"00",x"45",x"20",x"42",x"84",x"09",x"81",
		x"00",x"82",x"00",x"00",x"20",x"00",x"22",x"80",x"10",x"04",x"02",x"02",x"00",x"10",x"03",x"04",
		x"46",x"88",x"40",x"40",x"08",x"48",x"04",x"00",x"08",x"94",x"01",x"04",x"80",x"85",x"44",x"80",
		x"C8",x"89",x"08",x"00",x"4A",x"00",x"49",x"08",x"AC",x"10",x"0C",x"86",x"84",x"00",x"44",x"8C",
		x"90",x"40",x"30",x"10",x"18",x"44",x"12",x"11",x"A0",x"21",x"00",x"20",x"20",x"20",x"20",x"02",
		x"08",x"10",x"00",x"18",x"91",x"00",x"84",x"10",x"80",x"60",x"20",x"10",x"20",x"24",x"0A",x"21",
		x"10",x"18",x"91",x"00",x"08",x"01",x"25",x"00",x"20",x"05",x"4A",x"5F",x"3B",x"3F",x"DF",x"FF",
		x"01",x"04",x"0D",x"87",x"03",x"0C",x"03",x"01",x"7F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"04",x"90",x"00",x"00",x"00",x"11",x"40",x"00",x"24",x"02",x"52",x"01",x"10",x"09",x"04",x"02",
		x"04",x"00",x"80",x"80",x"84",x"00",x"10",x"40",x"88",x"00",x"42",x"04",x"04",x"01",x"26",x"40",
		x"A0",x"80",x"40",x"00",x"21",x"08",x"05",x"08",x"86",x"00",x"04",x"88",x"00",x"85",x"04",x"00",
		x"22",x"20",x"00",x"22",x"00",x"42",x"00",x"43",x"88",x"04",x"04",x"20",x"80",x"04",x"03",x"01",
		x"20",x"90",x"50",x"21",x"08",x"10",x"08",x"08",x"20",x"20",x"42",x"20",x"00",x"20",x"40",x"18",
		x"14",x"10",x"22",x"01",x"10",x"00",x"54",x"00",x"20",x"22",x"A2",x"00",x"80",x"A0",x"68",x"A1",
		x"86",x"0B",x"04",x"93",x"01",x"04",x"07",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",
		x"41",x"87",x"01",x"53",x"14",x"0C",x"87",x"23",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"00",x"00",x"10",x"00",x"00",x"A0",x"04",x"02",x"00",x"80",x"02",x"09",x"10",x"00",x"03",
		x"00",x"00",x"02",x"20",x"80",x"00",x"01",x"40",x"00",x"00",x"28",x"02",x"00",x"08",x"04",x"02",
		x"05",x"20",x"04",x"02",x"10",x"04",x"10",x"00",x"40",x"01",x"84",x"D0",x"0C",x"10",x"84",x"08",
		x"08",x"06",x"80",x"34",x"00",x"00",x"44",x"88",x"22",x"24",x"04",x"01",x"C2",x"54",x"90",x"21",
		x"90",x"98",x"00",x"14",x"42",x"01",x"14",x"00",x"29",x"90",x"28",x"28",x"46",x"12",x"22",x"A5",
		x"00",x"90",x"50",x"05",x"10",x"12",x"08",x"90",x"10",x"20",x"26",x"00",x"21",x"44",x"00",x"60",
		x"14",x"03",x"83",x"00",x"51",x"0F",x"27",x"88",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"07",x"43",x"11",x"8C",x"07",x"0B",x"03",x"84",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"40",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"20",x"12",x"00",x"03",x"2C",x"80",x"08",x"01",
		x"00",x"04",x"00",x"08",x"40",x"00",x"00",x"80",x"02",x"00",x"10",x"04",x"00",x"00",x"40",x"09",
		x"02",x"88",x"43",x"00",x"2A",x"00",x"10",x"91",x"24",x"12",x"14",x"20",x"04",x"08",x"85",x"14",
		x"00",x"02",x"40",x"08",x"00",x"01",x"84",x"10",x"40",x"11",x"82",x"0A",x"84",x"22",x"05",x"D0",
		x"50",x"82",x"14",x"00",x"50",x"51",x"20",x"08",x"A4",x"20",x"40",x"00",x"A0",x"04",x"30",x"20",
		x"10",x"00",x"14",x"40",x"00",x"10",x"50",x"40",x"28",x"84",x"04",x"00",x"A3",x"20",x"45",x"88",
		x"91",x"A5",x"00",x"10",x"A0",x"25",x"00",x"13",x"FF",x"3F",x"FF",x"FF",x"9F",x"3F",x"7F",x"BF",
		x"81",x"12",x"A1",x"00",x"51",x"09",x"52",x"22",x"1F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"BF",
		x"00",x"84",x"00",x"00",x"00",x"02",x"80",x"00",x"21",x"00",x"04",x"22",x"01",x"00",x"00",x"41",
		x"00",x"20",x"00",x"08",x"00",x"82",x"00",x"00",x"08",x"01",x"02",x"00",x"08",x"01",x"10",x"04",
		x"80",x"44",x"08",x"00",x"00",x"50",x"42",x"01",x"02",x"10",x"80",x"44",x"00",x"04",x"50",x"01",
		x"08",x"00",x"00",x"84",x"00",x"00",x"00",x"40",x"00",x"02",x"A0",x"00",x"00",x"55",x"00",x"81",
		x"42",x"90",x"01",x"08",x"50",x"20",x"02",x"22",x"26",x"00",x"20",x"95",x"08",x"A2",x"04",x"28",
		x"00",x"90",x"02",x"04",x"10",x"80",x"08",x"04",x"42",x"19",x"22",x"04",x"B5",x"00",x"01",x"2A",
		x"82",x"22",x"40",x"01",x"A7",x"09",x"80",x"42",x"FF",x"7F",x"7F",x"FF",x"FF",x"BF",x"FF",x"7F",
		x"03",x"01",x"08",x"50",x"40",x"00",x"13",x"81",x"3F",x"FF",x"FF",x"7F",x"7F",x"FF",x"9F",x"3F",
		x"EA",x"D5",x"EA",x"D4",x"EA",x"F1",x"E8",x"D4",x"A2",x"45",x"AA",x"50",x"8A",x"44",x"A2",x"55",
		x"EA",x"D0",x"E2",x"C0",x"EA",x"E0",x"E8",x"D5",x"AA",x"54",x"AA",x"41",x"A8",x"54",x"A2",x"00",
		x"AA",x"C4",x"EA",x"C5",x"EA",x"95",x"AA",x"91",x"AA",x"55",x"AA",x"40",x"AA",x"15",x"AA",x"51",
		x"EA",x"C4",x"82",x"D5",x"8A",x"81",x"CA",x"D4",x"AA",x"40",x"AA",x"55",x"AA",x"51",x"AA",x"51",
		x"AA",x"D0",x"EA",x"E1",x"AA",x"E5",x"EA",x"C1",x"A8",x"40",x"2A",x"11",x"AA",x"14",x"AA",x"41",
		x"A8",x"D0",x"AA",x"C1",x"EA",x"D5",x"AA",x"C4",x"AA",x"55",x"AA",x"44",x"AA",x"21",x"CA",x"20",
		x"AA",x"95",x"EA",x"D4",x"AA",x"D1",x"E8",x"D4",x"A2",x"45",x"AA",x"50",x"8A",x"44",x"A2",x"55",
		x"AA",x"D0",x"E2",x"C0",x"EA",x"D0",x"EA",x"E0",x"AA",x"54",x"AA",x"45",x"A8",x"54",x"AA",x"00",
		x"AF",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FE",x"FC",x"FF",x"FE",x"F8",x"FE",x"FD",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FE",x"FF",x"FE",x"FE",x"FC",x"FF",x"FE",
		x"03",x"1F",x"0F",x"13",x"0F",x"07",x"0F",x"3F",x"FC",x"F8",x"FE",x"FF",x"FE",x"FE",x"FF",x"FE",
		x"5F",x"1F",x"1F",x"BF",x"7F",x"BF",x"5F",x"BF",x"FC",x"FF",x"FA",x"FD",x"FE",x"FC",x"FE",x"FF",
		x"3F",x"7F",x"BF",x"1F",x"4F",x"3F",x"1F",x"3F",x"FE",x"FC",x"FE",x"FF",x"FE",x"FE",x"FF",x"FE",
		x"CF",x"7F",x"1F",x"BF",x"7F",x"BF",x"7F",x"BF",x"FD",x"F8",x"F2",x"FC",x"FA",x"FC",x"FE",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FE",x"FD",x"FF",x"FE",x"F8",x"FE",x"FD",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FE",x"FF",x"FE",x"FE",x"FC",x"FF",x"FE",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FE",x"E4",x"F8",x"FC",x"F0",x"F8",x"E8",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"F8",x"C4",x"F0",x"FC",x"F0",x"FF",x"FE",
		x"00",x"00",x"00",x"02",x"03",x"0B",x"07",x"05",x"00",x"00",x"00",x"40",x"80",x"C0",x"E0",x"F0",
		x"03",x"07",x"0A",x"03",x"06",x"01",x"02",x"00",x"E0",x"F0",x"F0",x"E0",x"C0",x"40",x"80",x"00",
		x"00",x"00",x"00",x"00",x"02",x"0C",x"26",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"2F",x"1F",x"3F",x"17",x"0F",x"17",x"0A",x"14",x"80",x"00",x"80",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"7F",x"7B",x"63",x"6B",x"63",x"7F",x"7F",x"01",x"7F",x"7B",x"63",x"6B",x"63",x"7F",x"7F",
		x"01",x"7F",x"7B",x"63",x"6B",x"63",x"7F",x"7F",x"01",x"7F",x"7B",x"63",x"6B",x"63",x"7F",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"10",x"50",x"50",x"50",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"D0",x"D0",x"D0",x"50",x"40",x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FA",x"FA",x"FE",x"F7",x"F7",x"F5",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FD",x"FD",x"F7",x"F7",x"F6",x"F6",x"F6",
		x"EE",x"EB",x"EB",x"FB",x"FF",x"FB",x"EB",x"EF",x"DF",x"FF",x"DF",x"DF",x"5F",x"7F",x"6F",x"7F",
		x"EF",x"EF",x"EB",x"EA",x"FA",x"FA",x"FE",x"FF",x"5F",x"7F",x"EF",x"EF",x"AF",x"EF",x"DF",x"F7",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"FF",
		x"00",x"00",x"00",x"06",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"66",x"00",x"99",x"00",x"66",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"19",x"00",x"06",x"00",x"01",x"00",x"00",
		x"00",x"00",x"00",x"66",x"00",x"99",x"00",x"66",x"00",x"00",x"00",x"66",x"00",x"99",x"00",x"66",
		x"00",x"99",x"00",x"66",x"00",x"99",x"00",x"00",x"00",x"99",x"00",x"66",x"00",x"99",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"EE",x"EE",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"EE",x"EE",x"FF",
		x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",
		x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",
		x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",x"FF",x"EE",x"EE",x"FF",
		x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
		x"55",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"55",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
		x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
		x"55",x"55",x"7F",x"7F",x"3F",x"3F",x"1F",x"00",x"55",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
		x"00",x"00",x"92",x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"49",x"49",x"49",x"49",x"49",x"49",
		x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
		x"00",x"00",x"80",x"80",x"C0",x"C0",x"E0",x"E0",x"00",x"1F",x"06",x"0C",x"1F",x"00",x"1F",x"14",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"1F",x"04",x"AE",x"BF",x"AA",x"BF",x"BF",x"BF",
		x"AA",x"AA",x"AA",x"FF",x"7F",x"3F",x"1F",x"00",x"BF",x"AA",x"BA",x"FF",x"FF",x"FF",x"FF",x"00",
		x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
		x"92",x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"49",x"49",x"49",x"49",x"49",x"49",x"00",x"00",
		x"FF",x"00",x"00",x"00",x"BB",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"B8",x"00",x"00",x"00",
		x"BB",x"00",x"00",x"00",x"BB",x"00",x"00",x"00",x"B8",x"00",x"03",x"00",x"B8",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"00",x"00",x"00",x"3B",x"00",x"00",x"00",
		x"0F",x"0F",x"7E",x"7E",x"7E",x"7F",x"7E",x"7E",x"3B",x"00",x"00",x"00",x"3B",x"00",x"00",x"00",
		x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"3B",x"00",x"00",x"00",x"3B",x"00",x"00",x"00",
		x"7F",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"3B",x"00",x"00",x"00",x"3F",x"FF",x"FF",x"FF",
		x"BB",x"00",x"00",x"00",x"BB",x"00",x"00",x"00",x"B8",x"00",x"03",x"00",x"B8",x"00",x"00",x"00",
		x"BB",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"B8",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",
		x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",
		x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",
		x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"FF",x"CC",x"CC",x"FF",x"CC",x"CC",x"FF",
		x"00",x"66",x"3F",x"19",x"0F",x"06",x"03",x"01",x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"66",x"3F",x"19",x"0F",x"06",x"03",x"00",
		x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",
		x"FF",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"00",x"FF",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"00",
		x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",
		x"CC",x"C0",x"C0",x"80",x"C0",x"C0",x"C0",x"80",x"CC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",x"00",x"66",x"FF",x"99",x"FF",x"66",x"FF",x"99",
		x"CC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CF",x"08",x"08",x"08",x"0F",x"08",x"08",x"08",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"0F",x"08",x"08",x"08",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"0F",x"08",x"08",x"08",
		x"C0",x"80",x"C0",x"80",x"C0",x"80",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C0",x"80",x"C0",x"80",x"C0",x"80",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"10",x"70",x"E0",x"C0",x"C0",x"80",x"00",x"80",
		x"7F",x"7D",x"3E",x"7C",x"7E",x"FF",x"74",x"E6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"03",x"01",x"01",x"03",x"01",x"03",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"01",x"03",x"01",x"03",x"03",x"01",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"52",x"FC",x"FF",x"FF",x"FF",x"FF",x"01",x"0B",x"47",x"EF",x"C7",x"F7",x"FB",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FF",x"F7",x"EF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"01",x"03",x"06",x"0C",x"40",x"80",x"C0",x"C0",x"00",x"20",x"20",x"60",
		x"30",x"41",x"47",x"4B",x"5F",x"47",x"4F",x"5B",x"64",x"FA",x"FE",x"FE",x"FF",x"FF",x"FF",x"DF",
		x"E3",x"C5",x"C3",x"C3",x"83",x"C1",x"C3",x"C7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"CB",x"C3",x"C1",x"C3",x"C3",x"CB",x"81",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"07",x"1F",x"FF",x"00",x"00",x"00",x"3E",x"FE",x"FE",x"FE",x"FE",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"00",x"00",x"00",x"00",x"03",x"1F",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"0B",x"0B",
		x"00",x"00",x"00",x"3C",x"FB",x"F7",x"F6",x"F4",x"45",x"69",x"75",x"E8",x"05",x"54",x"E2",x"C4",
		x"00",x"00",x"00",x"00",x"02",x"23",x"3A",x"33",x"00",x"00",x"06",x"03",x"01",x"01",x"01",x"41",
		x"33",x"21",x"F8",x"BC",x"FF",x"DE",x"F8",x"C0",x"41",x"49",x"B9",x"F8",x"F1",x"73",x"7B",x"7F",
		x"49",x"39",x"30",x"10",x"00",x"00",x"00",x"03",x"CF",x"8F",x"87",x"83",x"81",x"01",x"01",x"03",
		x"1F",x"33",x"71",x"F8",x"F9",x"F8",x"F8",x"F8",x"FF",x"F1",x"C0",x"80",x"C0",x"E0",x"C0",x"E0",
		x"00",x"00",x"00",x"00",x"01",x"03",x"0F",x"1D",x"01",x"07",x"17",x"77",x"F7",x"D5",x"55",x"55",
		x"7D",x"C0",x"80",x"7F",x"FE",x"FE",x"FA",x"FC",x"50",x"00",x"00",x"01",x"03",x"05",x"08",x"08",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"00",x"00",
		x"00",x"00",x"00",x"F0",x"FE",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"80",x"F0",x"F8",
		x"03",x"07",x"07",x"06",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"0B",x"19",x"19",x"1D",x"10",x"39",x"F9",x"F8",x"F9",x"FD",x"FD",x"FC",
		x"E0",x"E0",x"01",x"01",x"01",x"01",x"00",x"00",x"84",x"82",x"02",x"82",x"C2",x"82",x"A2",x"C0",
		x"80",x"C0",x"C0",x"C0",x"C0",x"80",x"80",x"80",x"80",x"F1",x"FD",x"FF",x"FF",x"7F",x"7F",x"7F",
		x"C4",x"61",x"71",x"61",x"43",x"42",x"61",x"00",x"7F",x"F5",x"FB",x"AB",x"DF",x"DF",x"1F",x"1D",
		x"28",x"25",x"24",x"0C",x"24",x"4C",x"34",x"24",x"3F",x"15",x"5F",x"2F",x"37",x"3F",x"1F",x"5D",
		x"F8",x"E0",x"F3",x"F0",x"F8",x"F0",x"D0",x"F8",x"C0",x"D0",x"C8",x"E0",x"48",x"48",x"C0",x"64",
		x"F8",x"F8",x"F0",x"F0",x"F0",x"FF",x"FF",x"FC",x"40",x"E0",x"71",x"7F",x"FF",x"D3",x"01",x"19",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"08",x"18",x"30",x"20",x"7C",x"03",x"0F",
		x"00",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"70",x"00",x"00",x"00",x"00",x"00",x"C0",x"02",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"00",x"01",x"03",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"03",x"01",x"00",x"00",x"00",x"00",x"10",
		x"7F",x"3D",x"9D",x"CD",x"CD",x"05",x"C1",x"C1",x"F0",x"F8",x"FC",x"7E",x"3E",x"0E",x"0F",x"0F",
		x"C1",x"C9",x"C1",x"C0",x"40",x"00",x"00",x"00",x"07",x"07",x"07",x"07",x"07",x"07",x"03",x"03",
		x"18",x"19",x"1D",x"8F",x"BF",x"9D",x"98",x"BC",x"FE",x"FF",x"FD",x"F9",x"F9",x"F9",x"F1",x"F9",
		x"9D",x"9F",x"8F",x"9F",x"BF",x"1F",x"0F",x"1F",x"F9",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"80",x"C0",x"C0",x"C0",x"F8",x"FC",x"FC",x"7F",x"7C",x"35",x"3D",x"18",x"37",x"2E",x"0B",
		x"FC",x"E7",x"8F",x"CF",x"DF",x"FF",x"FF",x"FE",x"13",x"15",x"EF",x"DD",x"EF",x"FF",x"9F",x"1F",
		x"C0",x"80",x"80",x"87",x"8F",x"C7",x"C1",x"A0",x"01",x"01",x"00",x"70",x"30",x"B8",x"B0",x"F8",
		x"80",x"B0",x"D8",x"CC",x"8C",x"C2",x"80",x"C0",x"38",x"38",x"1C",x"18",x"00",x"00",x"00",x"00",
		x"C5",x"C7",x"CD",x"C3",x"DF",x"DF",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"7F",x"7F",x"3F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FC",x"FC",x"FC",x"FC",x"F2",x"E2",x"F2",x"E6",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"82",x"86",x"84",x"80",x"40",x"40",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"40",x"00",x"00",x"00",x"00",x"08",
		x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"08",x"08",x"00",x"11",x"11",x"11",x"00",x"01",
		x"00",x"04",x"04",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"30",x"14",x"00",
		x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"80",x"07",x"07",x"07",x"07",x"0F",x"8F",x"8F",x"9F",
		x"81",x"87",x"1F",x"7F",x"00",x"00",x"00",x"00",x"E7",x"8F",x"7F",x"FF",x"1F",x"03",x"04",x"1A",
		x"67",x"B3",x"94",x"88",x"CB",x"C1",x"80",x"C0",x"FF",x"FD",x"FF",x"FF",x"FF",x"F9",x"CF",x"09",
		x"C0",x"80",x"00",x"00",x"1F",x"1F",x"1F",x"1F",x"87",x"04",x"00",x"80",x"E8",x"EC",x"C0",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"FD",x"32",x"83",x"C1",x"18",x"98",x"18",x"1C",x"1E",x"1E",
		x"00",x"C0",x"F2",x"7E",x"BE",x"B8",x"30",x"30",x"1E",x"1F",x"0C",x"58",x"CC",x"C0",x"81",x"01",
		x"C9",x"D9",x"DD",x"DC",x"EE",x"D7",x"C0",x"D0",x"60",x"60",x"B0",x"78",x"C0",x"C0",x"06",x"0C",
		x"C0",x"F8",x"E0",x"E8",x"E0",x"E0",x"C8",x"E8",x"06",x"06",x"70",x"1C",x"1C",x"0C",x"0C",x"0C",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"E9",x"E1",x"F5",x"EA",x"F4",x"E0",x"D4",x"E0",
		x"FD",x"F8",x"F0",x"F0",x"F0",x"C0",x"C0",x"C0",x"E8",x"D0",x"E4",x"D0",x"C0",x"C0",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"02",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"C6",x"0C",x"00",x"02",x"0A",x"2A",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"01",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"02",x"52",x"52",x"56",x"D6",x"D3",x"6E",x"EE",x"EE",x"EE",x"AA",x"AA",x"AA",x"AA",
		x"F3",x"F7",x"F7",x"1F",x"03",x"00",x"00",x"00",x"AA",x"AA",x"AA",x"AA",x"AA",x"FA",x"1E",x"00",
		x"16",x"00",x"10",x"11",x"17",x"1F",x"0F",x"0F",x"00",x"06",x"7F",x"FF",x"FF",x"FF",x"FF",x"FD",
		x"07",x"07",x"03",x"02",x"05",x"02",x"2D",x"95",x"F0",x"FB",x"95",x"B5",x"EA",x"A5",x"52",x"25",
		x"20",x"10",x"80",x"E0",x"F0",x"F8",x"FC",x"FE",x"03",x"07",x"03",x"03",x"03",x"05",x"01",x"03",
		x"3E",x"07",x"A1",x"58",x"D4",x"AA",x"92",x"6D",x"00",x"00",x"04",x"01",x"01",x"03",x"02",x"00",
		x"83",x"81",x"01",x"00",x"89",x"82",x"8B",x"8B",x"66",x"66",x"26",x"23",x"41",x"E3",x"C0",x"40",
		x"8F",x"0D",x"8A",x"97",x"1D",x"0C",x"84",x"84",x"41",x"61",x"60",x"E3",x"31",x"B1",x"93",x"4D",
		x"60",x"70",x"78",x"7C",x"44",x"64",x"40",x"E2",x"0C",x"0E",x"06",x"0A",x"0E",x"06",x"02",x"06",
		x"E1",x"C1",x"C1",x"E1",x"FD",x"80",x"81",x"81",x"16",x"0E",x"0C",x"88",x"18",x"08",x"0C",x"04",
		x"08",x"11",x"11",x"03",x"23",x"01",x"01",x"02",x"00",x"80",x"08",x"00",x"02",x"00",x"00",x"00",
		x"06",x"06",x"04",x"06",x"04",x"0C",x"08",x"10",x"02",x"00",x"10",x"00",x"00",x"08",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"05",x"0D",x"0B",x"3C",x"35",
		x"00",x"00",x"02",x"04",x"06",x"1F",x"3A",x"2F",x"DD",x"D7",x"DD",x"9B",x"DF",x"76",x"5D",x"35",
		x"7A",x"EF",x"BB",x"5A",x"F3",x"BB",x"6E",x"FF",x"C0",x"80",x"E0",x"E0",x"B0",x"A8",x"9C",x"BE",
		x"DB",x"7B",x"7B",x"56",x"FB",x"5F",x"9D",x"DB",x"BD",x"EB",x"7B",x"FA",x"F7",x"BB",x"3B",x"96",
		x"84",x"84",x"86",x"42",x"02",x"20",x"20",x"3C",x"CF",x"EF",x"F7",x"67",x"FF",x"78",x"78",x"7C",
		x"0C",x"8E",x"46",x"C4",x"44",x"E2",x"B0",x"68",x"FE",x"7F",x"2F",x"09",x"08",x"00",x"00",x"00",
		x"80",x"80",x"80",x"00",x"78",x"18",x"98",x"98",x"07",x"07",x"07",x"03",x"01",x"03",x"07",x"1E",
		x"0C",x"06",x"97",x"7B",x"3F",x"0F",x"1F",x"00",x"1C",x"30",x"78",x"3C",x"B6",x"D9",x"D8",x"7C",
		x"80",x"00",x"A0",x"80",x"40",x"A0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"90",x"40",x"20",x"80",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"02",x"03",x"09",x"0F",x"2A",
		x"00",x"00",x"02",x"02",x"0A",x"1A",x"2A",x"29",x"2B",x"A1",x"EB",x"BB",x"AB",x"8D",x"AA",x"AA",
		x"AD",x"7A",x"AD",x"DD",x"B4",x"3B",x"BF",x"AB",x"AF",x"ED",x"EA",x"7F",x"EA",x"67",x"DA",x"6D",
		x"DB",x"BE",x"BB",x"7D",x"AB",x"BB",x"BB",x"75",x"7F",x"F3",x"BA",x"6B",x"6F",x"6E",x"BB",x"7E",
		x"6E",x"FA",x"9E",x"FA",x"EC",x"5C",x"DA",x"BA",x"8B",x"0B",x"0A",x"C4",x"60",x"66",x"67",x"27",
		x"BA",x"6C",x"DE",x"76",x"DD",x"DF",x"D3",x"BD",x"21",x"01",x"21",x"03",x"03",x"03",x"00",x"00",
		x"01",x"41",x"20",x"37",x"11",x"18",x"08",x"08",x"BC",x"EC",x"E7",x"E0",x"E0",x"C0",x"F8",x"F0",
		x"0F",x"0C",x"07",x"03",x"83",x"83",x"03",x"03",x"60",x"60",x"78",x"62",x"FA",x"F2",x"C2",x"E6",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"02",x"0A",
		x"00",x"00",x"01",x"02",x"03",x"01",x"01",x"40",x"2E",x"33",x"FA",x"38",x"9E",x"EE",x"AB",x"2A",
		x"AE",x"A2",x"AA",x"8A",x"8A",x"A9",x"AA",x"6E",x"AA",x"CA",x"AA",x"AA",x"A8",x"AA",x"AB",x"A2",
		x"AA",x"BA",x"F2",x"EA",x"AA",x"AE",x"A9",x"8A",x"EA",x"AF",x"4A",x"3A",x"B8",x"AA",x"AA",x"A2",
		x"F3",x"AF",x"FF",x"F7",x"7D",x"DE",x"D6",x"DF",x"0C",x"2E",x"2E",x"26",x"86",x"82",x"92",x"91",
		x"BD",x"6D",x"F9",x"DB",x"FF",x"77",x"DF",x"5D",x"1B",x"D6",x"D3",x"81",x"A9",x"69",x"48",x"E8",
		x"0F",x"1F",x"3F",x"1F",x"1F",x"7F",x"FF",x"FF",x"7A",x"7C",x"7E",x"7C",x"78",x"60",x"BC",x"BE",
		x"FF",x"6F",x"3F",x"3F",x"0B",x"0F",x"0F",x"23",x"9E",x"9E",x"82",x"C6",x"80",x"C0",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",
		x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"26",x"03",x"C1",x"C1",x"A5",x"25",x"25",
		x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"39",x"2A",x"32",x"36",x"2B",x"3A",x"35",x"31",
		x"10",x"20",x"A0",x"80",x"20",x"22",x"22",x"23",x"7A",x"76",x"7A",x"71",x"72",x"3A",x"1E",x"0E",
		x"F5",x"BE",x"AC",x"FD",x"DB",x"7D",x"FD",x"AD",x"D8",x"E8",x"EE",x"A7",x"FE",x"6B",x"DF",x"FD",
		x"BF",x"77",x"BD",x"9D",x"BF",x"F7",x"6F",x"BD",x"6F",x"CE",x"EF",x"6F",x"E9",x"FC",x"BD",x"ED",
		x"20",x"A0",x"AF",x"BF",x"FC",x"F6",x"FA",x"EF",x"80",x"80",x"80",x"80",x"80",x"C0",x"40",x"40",
		x"F5",x"FE",x"F5",x"FA",x"FD",x"FE",x"F5",x"FB",x"40",x"C0",x"3C",x"D7",x"4A",x"10",x"A8",x"44",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"0A",x"08",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"31",x"3A",x"32",x"12",x"02",x"00",x"00",x"00",
		x"04",x"04",x"84",x"82",x"A2",x"A6",x"A4",x"24",x"48",x"40",x"48",x"48",x"42",x"42",x"20",x"20",
		x"04",x"25",x"21",x"05",x"14",x"44",x"50",x"54",x"21",x"21",x"22",x"02",x"02",x"82",x"80",x"80",
		x"22",x"12",x"22",x"26",x"24",x"AC",x"A8",x"A1",x"0A",x"0E",x"1E",x"05",x"0A",x"0C",x"0F",x"0E",
		x"81",x"A0",x"B0",x"A4",x"A2",x"21",x"22",x"04",x"06",x"87",x"A3",x"82",x"0B",x"02",x"0E",x"8E",
		x"FF",x"FE",x"FB",x"FD",x"FF",x"FF",x"FD",x"FF",x"AA",x"E8",x"54",x"A4",x"78",x"C2",x"28",x"D4",
		x"FE",x"FB",x"FF",x"FD",x"FF",x"FF",x"FB",x"FE",x"B0",x"C8",x"32",x"60",x"D4",x"68",x"D0",x"A8",
		x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"90",x"90",x"94",x"94",x"11",x"01",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"28",x"29",x"29",x"21",x"00",x"08",x"08",x"2A",x"A6",x"86",x"86",x"1E",x"39",x"3A",x"3E",x"BF",
		x"3B",x"3B",x"3E",x"3B",x"3E",x"36",x"3E",x"1E",x"AE",x"E6",x"A6",x"EA",x"8B",x"BF",x"E9",x"AB",
		x"03",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"2A",x"AB",x"EC",x"82",x"2A",x"3A",x"0B",x"02",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"AE",x"E2",x"8A",x"2A",x"A9",x"A8",x"AA",x"AA",x"9A",x"AC",x"E8",x"EC",x"A4",x"A8",x"A8",x"28",
		x"9A",x"EE",x"EA",x"AA",x"6A",x"0B",x"02",x"06",x"B9",x"A2",x"AB",x"AA",x"47",x"A7",x"A7",x"AD",
		x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"47",x"AB",x"B7",x"27",x"1A",x"07",x"01",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"DB",x"7D",x"D5",x"FD",x"B6",x"65",x"DE",x"DD",x"DE",x"F7",x"77",x"E4",x"B7",x"B3",x"B6",x"D7",
		x"55",x"7D",x"1D",x"17",x"0D",x"03",x"02",x"00",x"BF",x"F7",x"4F",x"9D",x"D7",x"D7",x"77",x"D9",
		x"A6",x"B6",x"94",x"97",x"37",x"B7",x"1F",x"3B",x"3B",x"27",x"AD",x"16",x"8D",x"9D",x"C7",x"F2",
		x"5A",x"36",x"22",x"20",x"30",x"78",x"F0",x"20",x"F9",x"C8",x"1C",x"2A",x"1F",x"1B",x"FD",x"3D",
		x"E2",x"76",x"66",x"67",x"33",x"A3",x"67",x"F3",x"38",x"1E",x"AC",x"0C",x"0D",x"19",x"31",x"1D",
		x"F7",x"63",x"37",x"33",x"5B",x"9B",x"1F",x"97",x"1A",x"03",x"B1",x"AB",x"11",x"A5",x"33",x"2D",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"FF",x"00",x"00",x"30",x"30",x"3B",x"1B",x"FC",x"FC",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F7",x"FD",x"01",x"27",x"00",x"40",x"30",x"3B",x"ED",x"E0",x"E0",x"E0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"60",x"3C",x"A7",x"83",x"00",x"03",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"00",x"00",x"00",
		x"01",x"00",x"03",x"87",x"0F",x"3F",x"FF",x"FF",x"F0",x"FC",x"01",x"00",x"80",x"80",x"80",x"80",
		x"04",x"03",x"3E",x"FE",x"FE",x"3E",x"00",x"00",x"80",x"FF",x"20",x"00",x"00",x"FF",x"8C",x"8F",
		x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"8F",x"8F",x"FF",x"FF",x"07",x"07",
		x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"08",x"C4",x"04",x"0F",
		x"FE",x"FF",x"07",x"07",x"03",x"00",x"00",x"00",x"7F",x"FF",x"FD",x"FD",x"FD",x"0D",x"01",x"07",
		x"FF",x"FF",x"0F",x"07",x"07",x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"01",x"FF",x"3F",
		x"FF",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"0F",x"FF",x"9F",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"04",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"3F",x"1B",x"14",x"10",x"10",x"30",
		x"20",x"FF",x"20",x"00",x"00",x"00",x"00",x"00",x"1F",x"FF",x"1F",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"3F",x"07",x"00",x"00",x"00",x"FC",x"FC",x"FD",x"FD",x"E3",x"C3",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"07",x"01",x"FD",x"F7",x"F7",x"FD",x"01",x"00",x"FC",x"FC",x"FC",x"FD",x"E1",x"E1",x"C3",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"3F",x"A7",x"BF",x"A7",x"B8",x"22",
		x"00",x"07",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"02",x"FE",x"FD",x"FB",x"F7",x"EF",x"DC",x"BC",
		x"FF",x"3F",x"07",x"80",x"C0",x"E0",x"01",x"F9",x"80",x"80",x"80",x"FE",x"FD",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"03",x"09",
		x"00",x"00",x"FF",x"FF",x"FF",x"F8",x"F8",x"F8",x"07",x"07",x"07",x"07",x"07",x"F8",x"88",x"88",
		x"FC",x"86",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"F8",x"F8",x"60",x"60",x"3F",x"80",x"FF",x"FF",
		x"00",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"55",x"00",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"50",
		x"55",x"55",x"55",x"55",x"D5",x"55",x"80",x"80",x"50",x"50",x"50",x"50",x"50",x"51",x"01",x"01",
		x"00",x"FF",x"FF",x"F8",x"F0",x"F8",x"FF",x"03",x"04",x"F8",x"EF",x"EF",x"FB",x"FB",x"EF",x"EF",
		x"73",x"73",x"F3",x"F3",x"F3",x"F2",x"F2",x"F2",x"FB",x"F8",x"CF",x"CF",x"CF",x"7F",x"7F",x"7F",
		x"5F",x"1F",x"5E",x"1F",x"5F",x"1F",x"5E",x"1F",x"EF",x"FC",x"2C",x"FC",x"EF",x"FC",x"2C",x"FC",
		x"5F",x"1F",x"1F",x"18",x"1F",x"1E",x"1F",x"01",x"EF",x"FF",x"FF",x"FF",x"83",x"7C",x"8E",x"84",
		x"FF",x"08",x"08",x"08",x"F8",x"08",x"08",x"08",x"FE",x"FE",x"FC",x"FC",x"FC",x"F8",x"F8",x"F8",
		x"F8",x"F8",x"F8",x"18",x"F8",x"00",x"00",x"00",x"F8",x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1E",x"1E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"07",x"0F",x"03",x"10",x"78",x"3C",x"8E",x"E3",
		x"0F",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FE",x"FF",x"7F",x"1F",x"0F",x"03",x"00",
		x"FF",x"FE",x"FD",x"FB",x"33",x"19",x"0C",x"06",x"7F",x"F9",x"F9",x"FF",x"F3",x"F3",x"FF",x"79",
		x"83",x"41",x"20",x"80",x"E0",x"F8",x"FC",x"FE",x"39",x"9F",x"CC",x"64",x"33",x"19",x"0C",x"06",
		x"CF",x"D8",x"D8",x"9F",x"B0",x"B0",x"9F",x"D8",x"8D",x"0D",x"0D",x"8D",x"0D",x"0D",x"8D",x"0D",
		x"D8",x"CF",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"0D",x"8D",x"0B",x"87",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"87",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"FF",x"C3",x"C3",x"FF",x"C3",x"C3",x"FF",
		x"FF",x"FF",x"FF",x"87",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"FF",x"C3",x"C2",x"FC",x"C0",x"C0",
		x"FF",x"FF",x"E1",x"E1",x"FE",x"E0",x"E0",x"F0",x"ED",x"CD",x"8D",x"0D",x"0D",x"0D",x"0F",x"0F",
		x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"0F",x"0D",x"0C",x"0C",x"0E",x"0E",x"0E",x"0E",
		x"F3",x"F3",x"F3",x"9F",x"9F",x"9F",x"FF",x"FF",x"FE",x"FD",x"FB",x"F7",x"EF",x"DF",x"BF",x"3C",
		x"FF",x"1F",x"9F",x"9F",x"E3",x"F3",x"73",x"72",x"9F",x"CF",x"E7",x"F3",x"F9",x"FC",x"FE",x"7F",
		x"01",x"01",x"FF",x"FF",x"87",x"FF",x"FF",x"FF",x"80",x"81",x"B3",x"A3",x"83",x"A3",x"A3",x"83",
		x"FF",x"FF",x"87",x"FF",x"FF",x"01",x"01",x"01",x"A3",x"A3",x"81",x"A0",x"B3",x"81",x"80",x"FC",
		x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0",x"E0",
		x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
		x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"7F",x"3F",x"0F",x"0F",x"1F",x"1F",x"3F",x"3F",
		x"1E",x"1E",x"1E",x"1E",x"1F",x"1F",x"1E",x"1E",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",x"7F",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"07",x"FF",x"07",x"00",x"00",x"00",x"00",x"3E",x"FE",x"FE",x"FE",x"7E",x"00",
		x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"FF",x"03",x"00",x"00",
		x"FF",x"7B",x"7B",x"00",x"00",x"00",x"00",x"7B",x"82",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",
		x"F0",x"07",x"3F",x"FC",x"FC",x"FF",x"3F",x"07",x"1F",x"E0",x"F7",x"00",x"00",x"F7",x"F7",x"E0",
		x"00",x"F2",x"E7",x"0F",x"1F",x"0D",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",
		x"FF",x"00",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"00",x"FC",x"00",x"01",x"E7",x"FF",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"F0",x"00",x"F0",x"00",x"00",x"1F",x"00",x"00",x"3F",x"7F",x"FF",
		x"F1",x"03",x"F3",x"F7",x"87",x"87",x"87",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",
		x"00",x"00",x"FF",x"C0",x"C0",x"00",x"4F",x"4F",x"0F",x"00",x"FF",x"83",x"83",x"00",x"9F",x"9F",
		x"0F",x"8F",x"8F",x"8F",x"8F",x"00",x"00",x"F1",x"9F",x"9F",x"9F",x"9F",x"9F",x"00",x"00",x"E3",
		x"B2",x"52",x"53",x"43",x"63",x"33",x"33",x"13",x"7F",x"7F",x"CF",x"CF",x"CF",x"FB",x"FB",x"EF",
		x"13",x"23",x"23",x"23",x"23",x"03",x"03",x"C3",x"EF",x"FB",x"FB",x"EF",x"EF",x"F8",x"C4",x"84",
		x"1F",x"1F",x"1F",x"18",x"1F",x"1F",x"1F",x"5F",x"8E",x"86",x"FF",x"FF",x"FF",x"FF",x"EF",x"FC",
		x"1E",x"5F",x"1F",x"5F",x"1E",x"5F",x"00",x"7F",x"2C",x"FC",x"EF",x"FC",x"2C",x"FC",x"01",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"F8",x"02",x"07",x"E0",x"E0",x"E0",x"C0",x"C0",x"CA",x"DF",x"FF",
		x"0B",x"07",x"0F",x"3F",x"1F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"DE",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"73",x"71",x"70",x"00",x"00",x"00",x"00",x"00",x"F8",x"F1",x"F1",x"78",x"3C",x"3E",x"3F",x"3F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"81",x"F3",x"F3",x"81",x"F1",x"00",x"00",x"FF",x"02",x"E7",x"E7",x"02",x"E3",x"00",x"00",x"FF",
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"C2",x"C1",x"07",x"C7",x"03",x"02",x"FF",x"0F",x"7D",x"FD",x"FD",x"FD",x"FD",x"1D",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"04",x"08",x"00",x"00",x"00",x"00",x"00",
		x"DF",x"DF",x"C0",x"C0",x"C0",x"C1",x"C2",x"C3",x"3F",x"3F",x"07",x"0F",x"3F",x"CF",x"FF",x"FF",
		x"0F",x"07",x"1F",x"0F",x"3F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"7F",x"3F",x"3F",x"1F",x"1F",x"3F",x"2F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"1B",x"07",x"07",x"03",x"05",x"00",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"03",x"03",x"07",x"0F",x"07",x"0F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"1F",x"2F",x"1F",x"3F",x"5F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"7F",x"1F",x"2F",x"0F",x"17",x"1F",x"0F",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"07",x"0F",x"0B",x"07",x"03",x"05",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"67",x"02",
		x"FE",x"FF",x"FA",x"FF",x"EE",x"FD",x"FB",x"FD",x"AF",x"77",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",
		x"FD",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"BF",x"7F",x"5F",x"17",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"0F",x"07",x"03",x"05",x"01",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"AF",x"D7",x"EF",x"DF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"EE",x"C5",x"A0",x"00",x"FF",x"FF",x"FF",x"3F",x"9F",x"3F",x"0F",x"06",
		x"DF",x"BF",x"EF",x"FF",x"AB",x"F7",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"EF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"F7",x"F3",x"D7",x"DB",x"77",x"77",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"EF",x"FF",x"EF",x"F7",x"EF",x"F7",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F3",x"E9",x"F7",x"F9",x"F3",x"FF",x"EF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"FF",x"BF",x"DF",x"BF",x"FF",x"FF",x"DF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"DF",x"FF",x"5F",x"FF",x"FF",x"AF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"F7",x"FF",x"F7",x"DF",x"F7",x"EF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"04",x"40",x"54",x"01",x"10",x"26",x"16",x"01",x"08",x"12",x"55",x"07",x"25",x"11",x"4C",x"00",
		x"C0",x"0D",x"58",x"15",x"11",x"05",x"86",x"00",x"45",x"29",x"54",x"10",x"42",x"01",x"00",x"00",
		x"4C",x"05",x"01",x"54",x"00",x"14",x"A5",x"14",x"4B",x"15",x"80",x"54",x"E0",x"45",x"10",x"14",
		x"42",x"D5",x"43",x"14",x"11",x"00",x"C0",x"00",x"65",x"00",x"10",x"15",x"40",x"41",x"00",x"00",
		x"76",x"DA",x"F6",x"EC",x"68",x"F6",x"7C",x"F1",x"B5",x"08",x"D0",x"10",x"88",x"20",x"42",x"08",
		x"48",x"F8",x"ED",x"DA",x"79",x"ED",x"7F",x"A2",x"00",x"02",x"00",x"10",x"02",x"40",x"00",x"42",
		x"78",x"E8",x"74",x"F2",x"78",x"E0",x"76",x"B9",x"46",x"00",x"05",x"6E",x"7F",x"06",x"27",x"00",
		x"70",x"D8",x"F0",x"C1",x"70",x"E4",x"60",x"F1",x"00",x"0C",x"85",x"D7",x"76",x"5F",x"03",x"13",
		x"84",x"D4",x"8A",x"CA",x"9A",x"1D",x"B4",x"55",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"6D",x"A5",x"4A",x"CA",x"84",x"71",x"6E",x"AC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7E",x"F5",x"FE",x"F9",x"76",x"BD",x"79",x"FC",x"84",x"12",x"08",x"07",x"8B",x"40",x"81",x"80",
		x"76",x"B8",x"5E",x"B9",x"3C",x"F9",x"76",x"FA",x"09",x"C0",x"00",x"03",x"A1",x"8B",x"40",x"90",
		x"FF",x"FD",x"7E",x"3D",x"58",x"DE",x"EA",x"A5",x"71",x"F3",x"FB",x"BF",x"7F",x"1F",x"17",x"0B",
		x"C9",x"3B",x"7F",x"FF",x"FF",x"7F",x"02",x"01",x"BC",x"FF",x"FF",x"F6",x"FC",x"FC",x"F6",x"0F",
		x"0B",x"84",x"90",x"15",x"B0",x"FE",x"FF",x"BC",x"07",x"82",x"A0",x"E8",x"FC",x"DD",x"5D",x"7F",
		x"E8",x"18",x"DF",x"DF",x"0F",x"07",x"01",x"9B",x"0E",x"A5",x"FE",x"FA",x"D0",x"84",x"C2",x"E0",
		x"04",x"40",x"54",x"01",x"10",x"26",x"16",x"01",x"08",x"12",x"55",x"07",x"25",x"11",x"4C",x"00",
		x"C0",x"0D",x"58",x"15",x"11",x"55",x"C6",x"40",x"45",x"29",x"54",x"10",x"42",x"01",x"0C",x"D5",
		x"40",x"11",x"55",x"10",x"C4",x"60",x"05",x"46",x"05",x"80",x"05",x"17",x"05",x"40",x"00",x"04",
		x"11",x"11",x"0C",x"40",x"31",x"54",x"11",x"41",x"10",x"35",x"11",x"00",x"41",x"04",x"40",x"04",
		x"F2",x"9C",x"61",x"36",x"33",x"DB",x"53",x"87",x"D7",x"BE",x"F8",x"F8",x"F0",x"A0",x"E0",x"90",
		x"7E",x"AF",x"5D",x"BE",x"7F",x"FE",x"FC",x"F5",x"D4",x"80",x"00",x"90",x"40",x"01",x"20",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FF",x"4A",x"A0",x"D4",x"94",x"08",x"40",x"E4",x"30",
		x"FC",x"FE",x"FC",x"F8",x"F9",x"F9",x"C9",x"C9",x"50",x"08",x"04",x"44",x"12",x"80",x"20",x"48",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FF",x"FF",x"BF",x"BF",x"BF",x"3F",x"80",x"BF",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"BF",x"BF",x"3F",x"80",x"BF",x"BF",x"BF",x"3F",
		x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",
		x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",
		x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"40",x"A0",x"34",x"44",x"A8",x"30",x"3A",x"60",
		x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"C9",x"50",x"10",x"A8",x"34",x"60",x"10",x"08",x"50",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FF",x"80",x"BF",x"BF",x"BF",x"3F",x"80",x"BF",x"BF",
		x"E7",x"E0",x"E1",x"E0",x"E1",x"E8",x"E8",x"E9",x"BF",x"BF",x"83",x"01",x"01",x"1F",x"7F",x"3F",
		x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FB",x"E8",x"E9",x"E0",x"E8",x"E0",x"E1",x"E9",x"BF",x"1F",x"0F",x"0F",x"01",x"01",x"1F",x"3F",
		x"FC",x"E0",x"E9",x"E8",x"E8",x"E8",x"E0",x"EC",x"3F",x"3F",x"1F",x"0F",x"0F",x"0F",x"8F",x"BF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",
		x"E3",x"E3",x"E3",x"E3",x"E3",x"E3",x"E3",x"FB",x"BF",x"BF",x"3F",x"80",x"BF",x"BF",x"BF",x"3F",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"80",x"BF",x"BF",x"BF",x"3F",x"80",x"BF",x"BF",
		x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"BF",x"3F",x"80",x"BF",x"BF",x"BF",x"3F",x"80",
		x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"BF",x"BF",x"BF",x"3F",x"80",x"BF",x"BF",x"BF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"FC",x"FC",x"F8",x"F8",x"F8",x"F0",x"F0",
		x"FB",x"FB",x"7B",x"7B",x"44",x"44",x"5C",x"44",x"3F",x"80",x"BF",x"3F",x"3F",x"3F",x"00",x"00",
		x"5C",x"44",x"5C",x"44",x"5C",x"44",x"5C",x"44",x"00",x"BF",x"BF",x"BF",x"3F",x"3F",x"00",x"00",
		x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"E0",x"E0",x"E0",x"C0",x"C0",x"C0",x"80",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"80",x"00",x"00",x"00",x"80",x"C8",x"F0",
		x"5C",x"44",x"5C",x"44",x"5C",x"44",x"5C",x"44",x"00",x"BF",x"BF",x"BF",x"3F",x"3F",x"00",x"00",
		x"5C",x"44",x"5C",x"44",x"5C",x"44",x"5C",x"44",x"00",x"BF",x"BF",x"BF",x"3F",x"3F",x"00",x"00",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"FC",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",x"FF",x"40",x"30",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"80",x"80",x"C0",x"C4",x"F8",x"F8",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D0",x"D8",x"C8",x"E8",x"E8",x"F8",x"F8",x"F8",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"FC",x"FA",x"F9",x"FD",x"FD",x"FF",x"FF",
		x"5C",x"44",x"5C",x"44",x"5C",x"44",x"5C",x"44",x"00",x"BF",x"BF",x"BF",x"3F",x"3F",x"00",x"00",
		x"5C",x"44",x"5C",x"44",x"5C",x"44",x"5C",x"44",x"00",x"BF",x"BF",x"BF",x"3F",x"3F",x"7F",x"FF",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"36",x"F6",x"F6",x"FE",x"FF",x"FF",x"FD",x"FE",x"48",x"A8",x"58",x"54",x"08",x"A8",x"E0",x"C0",
		x"FE",x"FF",x"FF",x"FE",x"FF",x"FF",x"FE",x"FF",x"54",x"8C",x"84",x"94",x"52",x"A8",x"26",x"54",
		x"CE",x"CE",x"F6",x"36",x"36",x"36",x"36",x"36",x"20",x"82",x"56",x"44",x"40",x"A8",x"50",x"44",
		x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"A0",x"F0",x"24",x"B0",x"78",x"A8",x"28",x"54",
		x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"48",x"A0",x"50",x"50",x"28",x"A8",x"64",x"58",
		x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"10",x"A8",x"20",x"78",x"70",x"B8",x"34",x"54",
		x"25",x"10",x"A4",x"01",x"00",x"11",x"00",x"08",x"BF",x"52",x"01",x"02",x"D0",x"32",x"0C",x"23",
		x"20",x"82",x"10",x"09",x"80",x"00",x"20",x"04",x"41",x"02",x"48",x"02",x"40",x"21",x"02",x"26",
		x"FF",x"11",x"00",x"48",x"91",x"00",x"00",x"50",x"FF",x"84",x"4C",x"84",x"02",x"00",x"A4",x"00",
		x"81",x"70",x"1C",x"27",x"54",x"10",x"00",x"28",x"8C",x"00",x"80",x"A2",x"C4",x"74",x"9E",x"83",
		x"DF",x"30",x"08",x"11",x"00",x"B0",x"14",x"80",x"D7",x"94",x"20",x"12",x"20",x"10",x"14",x"40",
		x"54",x"11",x"08",x"10",x"00",x"14",x"10",x"30",x"B1",x"10",x"40",x"90",x"08",x"15",x"00",x"30",
		x"FF",x"18",x"52",x"04",x"14",x"10",x"10",x"2A",x"28",x"04",x"00",x"44",x"40",x"00",x"00",x"20",
		x"10",x"02",x"08",x"92",x"30",x"18",x"10",x"90",x"00",x"24",x"04",x"90",x"10",x"00",x"00",x"62",
		x"00",x"02",x"00",x"0A",x"24",x"80",x"00",x"80",x"20",x"12",x"4A",x"28",x"8C",x"12",x"9A",x"43",
		x"01",x"08",x"12",x"00",x"A0",x"00",x"00",x"01",x"00",x"3A",x"80",x"10",x"53",x"02",x"29",x"0B",
		x"88",x"41",x"28",x"10",x"48",x"4D",x"02",x"08",x"84",x"04",x"80",x"00",x"0C",x"84",x"80",x"05",
		x"85",x"08",x"50",x"00",x"48",x"40",x"09",x"50",x"80",x"C0",x"A4",x"00",x"0C",x"04",x"0A",x"14",
		x"D0",x"30",x"1E",x"43",x"00",x"00",x"10",x"18",x"40",x"04",x"40",x"41",x"A0",x"70",x"08",x"47",
		x"40",x"88",x"10",x"14",x"21",x"91",x"04",x"30",x"03",x"D0",x"00",x"40",x"24",x"40",x"40",x"01",
		x"10",x"10",x"00",x"90",x"04",x"90",x"01",x"30",x"00",x"02",x"00",x"40",x"00",x"00",x"02",x"10",
		x"D0",x"70",x"34",x"37",x"01",x"12",x"90",x"30",x"00",x"08",x"00",x"02",x"80",x"10",x"00",x"48",
		x"08",x"00",x"20",x"00",x"44",x"80",x"00",x"02",x"80",x"02",x"44",x"20",x"52",x"00",x"09",x"83",
		x"00",x"00",x"00",x"08",x"20",x"00",x"82",x"80",x"00",x"44",x"00",x"02",x"02",x"10",x"81",x"06",
		x"64",x"88",x"04",x"40",x"08",x"48",x"04",x"02",x"08",x"86",x"01",x"44",x"80",x"04",x"44",x"80",
		x"48",x"88",x"00",x"00",x"4A",x"04",x"49",x"80",x"A4",x"10",x"0D",x"84",x"84",x"20",x"04",x"84",
		x"90",x"44",x"20",x"30",x"18",x"04",x"13",x"10",x"28",x"20",x"40",x"60",x"02",x"20",x"20",x"10",
		x"00",x"30",x"04",x"18",x"10",x"00",x"80",x"50",x"80",x"60",x"20",x"14",x"20",x"24",x"42",x"23",
		x"80",x"18",x"10",x"24",x"28",x"00",x"08",x"40",x"80",x"00",x"40",x"40",x"22",x"24",x"06",x"03",
		x"00",x"06",x"04",x"00",x"87",x"00",x"20",x"00",x"01",x"CC",x"97",x"43",x"B1",x"C6",x"4B",x"21",
		x"21",x"10",x"00",x"00",x"84",x"00",x"40",x"08",x"25",x"00",x"12",x"44",x"10",x"21",x"04",x"00",
		x"00",x"00",x"02",x"00",x"24",x"01",x"00",x"40",x"89",x"08",x"02",x"20",x"05",x"01",x"04",x"50",
		x"20",x"80",x"40",x"00",x"23",x"08",x"84",x"18",x"A4",x"00",x"14",x"82",x"00",x"84",x"04",x"00",
		x"02",x"20",x"00",x"20",x"00",x"C2",x"08",x"02",x"88",x"40",x"05",x"00",x"80",x"46",x"01",x"01",
		x"00",x"98",x"50",x"20",x"00",x"92",x"18",x"09",x"B0",x"00",x"40",x"60",x"02",x"20",x"50",x"08",
		x"14",x"10",x"22",x"41",x"10",x"08",x"10",x"00",x"20",x"22",x"60",x"01",x"80",x"E0",x"4A",x"A1",
		x"A0",x"01",x"00",x"80",x"02",x"40",x"00",x"00",x"8F",x"11",x"C3",x"4F",x"13",x"27",x"09",x"42",
		x"00",x"89",x"80",x"40",x"00",x"00",x"80",x"00",x"38",x"11",x"C7",x"1F",x"21",x"03",x"37",x"48",
		x"02",x"00",x"80",x"10",x"00",x"00",x"80",x"00",x"12",x"00",x"00",x"00",x"21",x"10",x"04",x"01",
		x"00",x"00",x"02",x"20",x"00",x"00",x"00",x"44",x"00",x"00",x"08",x"02",x"00",x"41",x"04",x"00",
		x"04",x"A4",x"00",x"02",x"10",x"04",x"00",x"20",x"40",x"22",x"84",x"90",x"04",x"10",x"94",x"08",
		x"0A",x"02",x"80",x"24",x"00",x"20",x"40",x"09",x"00",x"24",x"46",x"00",x"82",x"54",x"88",x"21",
		x"90",x"B2",x"00",x"14",x"88",x"01",x"10",x"12",x"20",x"10",x"2A",x"28",x"44",x"46",x"22",x"21",
		x"00",x"80",x"90",x"0C",x"14",x"13",x"00",x"30",x"10",x"20",x"B4",x"01",x"21",x"40",x"22",x"20",
		x"80",x"00",x"00",x"24",x"60",x"00",x"08",x"C0",x"83",x"C7",x"74",x"29",x"13",x"82",x"54",x"11",
		x"00",x"40",x"00",x"00",x"80",x"00",x"20",x"82",x"0F",x"27",x"48",x"07",x"13",x"29",x"6F",x"87",
		x"00",x"80",x"00",x"00",x"00",x"80",x"08",x"00",x"01",x"12",x"80",x"01",x"24",x"82",x"08",x"01",
		x"80",x"00",x"00",x"08",x"42",x"00",x"00",x"00",x"00",x"04",x"00",x"04",x"01",x"00",x"00",x"08",
		x"02",x"08",x"51",x"00",x"2A",x"02",x"00",x"90",x"64",x"02",x"14",x"20",x"86",x"08",x"81",x"14",
		x"00",x"02",x"40",x"0C",x"80",x"01",x"04",x"19",x"62",x"01",x"82",x"0A",x"84",x"10",x"05",x"92",
		x"14",x"A2",x"10",x"01",x"70",x"10",x"A0",x"01",x"A0",x"00",x"44",x"20",x"A0",x"08",x"30",x"20",
		x"14",x"40",x"10",x"00",x"00",x"11",x"70",x"08",x"28",x"12",x"04",x"80",x"2A",x"21",x"51",x"08",
		x"50",x"A0",x"00",x"50",x"89",x"20",x"02",x"52",x"0A",x"47",x"47",x"8B",x"11",x"0F",x"8C",x"51",
		x"81",x"18",x"20",x"80",x"50",x"20",x"10",x"60",x"0B",x"CF",x"8F",x"1B",x"35",x"42",x"05",x"1F",
		x"00",x"80",x"00",x"80",x"00",x"02",x"80",x"00",x"24",x"00",x"00",x"02",x"00",x"08",x"00",x"41",
		x"04",x"20",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"02",x"10",x"08",x"01",x"01",x"04",
		x"04",x"40",x"08",x"20",x"01",x"40",x"02",x"00",x"00",x"10",x"82",x"00",x"00",x"04",x"42",x"00",
		x"08",x"00",x"00",x"00",x"20",x"00",x"02",x"00",x"40",x"02",x"88",x"00",x"00",x"11",x"02",x"80",
		x"0A",x"90",x"01",x"80",x"50",x"00",x"00",x"22",x"23",x"10",x"22",x"04",x"48",x"A3",x"00",x"08",
		x"41",x"14",x"02",x"00",x"10",x"20",x"02",x"04",x"52",x"10",x"22",x"02",x"95",x"00",x"04",x"0A",
		x"84",x"20",x"40",x"92",x"A0",x"00",x"00",x"50",x"00",x"01",x"03",x"87",x"94",x"09",x"07",x"03",
		x"00",x"00",x"A0",x"40",x"00",x"04",x"10",x"A0",x"07",x"04",x"29",x"43",x"07",x"04",x"08",x"41",
		x"E4",x"C0",x"E4",x"C1",x"D0",x"E6",x"F6",x"C1",x"08",x"12",x"55",x"07",x"21",x"11",x"48",x"00",
		x"C0",x"CD",x"F8",x"D5",x"D1",x"F5",x"C6",x"C0",x"45",x"29",x"50",x"10",x"46",x"01",x"0C",x"D5",
		x"80",x"91",x"D5",x"D0",x"C4",x"80",x"85",x"86",x"05",x"80",x"05",x"14",x"05",x"40",x"00",x"04",
		x"D1",x"D1",x"8C",x"C0",x"B1",x"94",x"91",x"C1",x"10",x"35",x"11",x"00",x"41",x"04",x"40",x"04",
		x"C4",x"85",x"C1",x"F4",x"80",x"80",x"E5",x"D4",x"43",x"15",x"80",x"44",x"40",x"41",x"10",x"14",
		x"C2",x"C1",x"C1",x"94",x"D1",x"80",x"C5",x"D1",x"45",x"00",x"10",x"11",x"44",x"50",x"15",x"05",
		x"84",x"C0",x"D4",x"81",x"90",x"E6",x"D6",x"81",x"08",x"12",x"55",x"07",x"25",x"11",x"4C",x"00",
		x"C0",x"CD",x"D8",x"95",x"D1",x"85",x"C4",x"E0",x"45",x"29",x"54",x"10",x"42",x"01",x"04",x"00",
		x"80",x"13",x"94",x"49",x"62",x"38",x"34",x"C3",x"D0",x"E9",x"50",x"E0",x"70",x"13",x"A0",x"D0",
		x"A9",x"47",x"E0",x"8B",x"C7",x"71",x"C8",x"F6",x"61",x"C0",x"94",x"61",x"D8",x"89",x"24",x"E1",
		x"00",x"08",x"07",x"03",x"00",x"40",x"05",x"03",x"01",x"93",x"40",x"62",x"3D",x"D8",x"84",x"70",
		x"10",x"11",x"0E",x"04",x"01",x"13",x"0A",x"00",x"F9",x"10",x"21",x"D0",x"F1",x"09",x"78",x"98",
		x"10",x"09",x"07",x"02",x"08",x"5E",x"13",x"2A",x"40",x"39",x"9D",x"06",x"9C",x"79",x"04",x"48",
		x"C7",x"71",x"0E",x"04",x"01",x"1A",x"78",x"84",x"BA",x"15",x"40",x"C1",x"21",x"09",x"78",x"88",
		x"CC",x"3B",x"94",x"49",x"62",x"B8",x"34",x"C3",x"D0",x"E8",x"50",x"E0",x"71",x"10",x"A0",x"D0",
		x"A9",x"47",x"E0",x"8B",x"C7",x"71",x"C8",x"F6",x"61",x"C0",x"94",x"60",x"D8",x"89",x"24",x"E1",
		x"D6",x"2B",x"94",x"48",x"E1",x"CA",x"14",x"C0",x"C0",x"68",x"01",x"D3",x"E1",x"37",x"83",x"27",
		x"A7",x"49",x"E1",x"8F",x"93",x"00",x"8B",x"F6",x"05",x"CB",x"0F",x"45",x"83",x"83",x"20",x"E8",
		x"FF",x"FF",x"FF",x"FD",x"FD",x"F7",x"F8",x"FF",x"FF",x"FF",x"CF",x"AF",x"CB",x"47",x"83",x"47",
		x"FF",x"F8",x"F7",x"FD",x"FB",x"FE",x"FD",x"FF",x"43",x"E3",x"A3",x"47",x"87",x"CF",x"DB",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"DA",x"EC",x"FF",x"FF",x"FF",x"FF",x"FF",x"5F",x"7F",x"1F",
		x"FE",x"FA",x"C7",x"FD",x"FA",x"FD",x"F6",x"EF",x"3F",x"1F",x"1F",x"1F",x"3F",x"3F",x"7F",x"DF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FE",x"82",x"BA",x"AA",x"B2",x"A2",x"BE",x"80",x"FE",x"82",x"BA",x"AA",x"B2",x"A2",x"BE",x"80",
		x"FE",x"82",x"BA",x"AA",x"B2",x"A2",x"BE",x"80",x"FE",x"82",x"BA",x"AA",x"B2",x"A2",x"BE",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"82",x"12",x"52",x"50",x"50",x"C0",x"C1",x"85",x"D6",x"F3",x"D5",x"D2",x"56",x"77",x"6D",x"7A",
		x"85",x"D5",x"D3",x"D2",x"52",x"42",x"42",x"43",x"5D",x"74",x"EC",x"E9",x"AC",x"EC",x"DB",x"F6",
		x"4E",x"0B",x"2B",x"79",x"F7",x"49",x"4B",x"6F",x"FB",x"FB",x"FA",x"FA",x"7E",x"77",x"67",x"75",
		x"6F",x"2F",x"AB",x"A2",x"92",x"B2",x"16",x"77",x"5D",x"7D",x"ED",x"F7",x"B7",x"F6",x"F6",x"F6",
		x"51",x"54",x"54",x"44",x"40",x"44",x"54",x"50",x"20",x"01",x"25",x"25",x"A1",x"81",x"91",x"85",
		x"50",x"50",x"54",x"55",x"45",x"45",x"41",x"40",x"A4",x"84",x"14",x"15",x"51",x"10",x"21",x"08",
		x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",
		x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",
		x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",
		x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",x"33",x"00",x"00",x"33",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"F0",x"FE",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"66",x"00",x"99",x"00",x"E6",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"F9",x"F0",x"FE",x"FC",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"00",x"66",x"00",x"99",x"00",x"66",x"FF",x"FF",x"00",x"66",x"00",x"99",x"00",x"66",
		x"00",x"99",x"00",x"66",x"00",x"99",x"00",x"FF",x"00",x"99",x"00",x"66",x"00",x"99",x"00",x"FF",
		x"FF",x"FF",x"00",x"00",x"11",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"11",x"00",x"00",x"00",
		x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",
		x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",
		x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",x"11",x"00",x"00",x"00",
		x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
		x"55",x"55",x"AA",x"AA",x"55",x"55",x"AA",x"FF",x"55",x"55",x"AA",x"AA",x"55",x"55",x"AA",x"FF",
		x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
		x"55",x"55",x"AA",x"AA",x"D5",x"D5",x"EA",x"FF",x"55",x"55",x"AA",x"AA",x"55",x"55",x"AA",x"FF",
		x"FF",x"FF",x"6D",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"B6",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"0A",x"04",x"1F",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"C0",x"E0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"FF",x"FF",x"AE",x"BF",x"AA",x"BF",x"BF",x"BF",
		x"AA",x"AA",x"AA",x"00",x"80",x"C0",x"E0",x"FF",x"BF",x"AA",x"BA",x"10",x"1F",x"10",x"10",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FF",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"FF",x"FF",x"FF",x"C3",x"C3",x"C2",x"C3",x"C3",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"C2",x"C3",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"FF",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
		x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",
		x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",
		x"FF",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"33",x"33",x"31",x"33",x"33",x"73",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"30",x"30",x"30",x"30",x"37",x"30",x"30",x"30",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"30",x"30",x"30",x"30",x"37",x"30",x"30",x"30",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"30",x"30",x"30",x"30",x"37",x"30",x"30",x"30",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"01",x"DC",x"F8",x"F8",x"7E",x"78",x"3C",x"32",x"C0",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FA",x"F0",x"28",x"F2",x"53",x"E4",x"47",x"D7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"48",x"A0",x"14",x"D2",x"8A",x"28",x"20",x"50",
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"D4",x"A0",x"84",x"58",x"D0",x"80",x"A4",x"58",
		x"FF",x"FF",x"BF",x"77",x"78",x"ED",x"73",x"F9",x"FF",x"FF",x"BF",x"9E",x"3F",x"9E",x"4E",x"A5",
		x"73",x"A1",x"53",x"0C",x"C6",x"17",x"4A",x"54",x"CC",x"C6",x"B7",x"E2",x"A5",x"42",x"37",x"16",
		x"0F",x"55",x"93",x"39",x"9C",x"11",x"38",x"74",x"69",x"C2",x"EC",x"8A",x"D4",x"78",x"F4",x"7E",
		x"B0",x"38",x"14",x"38",x"9E",x"1C",x"48",x"02",x"3D",x"5C",x"BA",x"1E",x"2D",x"87",x"0E",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"F0",x"E2",x"01",x"03",x"07",x"07",x"87",x"2F",x"2F",x"7F",
		x"CF",x"BF",x"BF",x"BF",x"BE",x"BE",x"BC",x"BC",x"6B",x"F5",x"E1",x"C1",x"00",x"00",x"00",x"00",
		x"DF",x"FF",x"BF",x"FF",x"BF",x"FF",x"BF",x"FF",x"DC",x"EE",x"FB",x"7D",x"EE",x"DF",x"FA",x"EE",
		x"FF",x"BF",x"BF",x"FF",x"BF",x"F7",x"BE",x"BF",x"7D",x"DA",x"E6",x"BD",x"F7",x"FE",x"39",x"9F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"2A",x"FF",x"FF",x"FF",x"FF",x"EF",x"AB",x"AB",x"AF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"0F",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F0",x"F6",x"92",
		x"FF",x"FF",x"FE",x"FC",x"FB",x"F7",x"F6",x"FE",x"70",x"70",x"79",x"F4",x"78",x"78",x"78",x"78",
		x"FF",x"FF",x"FF",x"FF",x"BC",x"1C",x"05",x"0C",x"FF",x"FF",x"F9",x"FC",x"78",x"38",x"30",x"50",
		x"0C",x"1E",x"07",x"03",x"30",x"41",x"27",x"1F",x"FC",x"D4",x"34",x"67",x"4E",x"CC",x"E4",x"E0",
		x"BE",x"9E",x"1C",x"1C",x"0C",x"18",x"18",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"40",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"FF",x"FE",x"F1",x"E1",x"81",x"01",x"01",x"01",
		x"F0",x"C3",x"84",x"00",x"00",x"FC",x"FA",x"FC",x"00",x"80",x"00",x"00",x"00",x"04",x"08",x"0C",
		x"2A",x"6A",x"6A",x"6A",x"2A",x"2A",x"2A",x"00",x"BF",x"BF",x"BF",x"FF",x"FF",x"FC",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"08",
		x"03",x"07",x"07",x"06",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"EC",x"E4",x"0E",x"05",x"02",x"00",x"00",x"00",x"1A",x"4D",x"9D",x"0C",x"10",x"38",x"1D",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"0E",x"02",x"00",x"00",x"00",x"00",x"00",
		x"CB",x"2E",x"17",x"AE",x"0C",x"05",x"06",x"39",x"F0",x"EA",x"64",x"F4",x"E0",x"60",x"A0",x"62",
		x"93",x"0A",x"89",x"08",x"1B",x"38",x"99",x"19",x"82",x"EA",x"A2",x"92",x"48",x"C0",x"C0",x"A2",
		x"00",x"00",x"07",x"0F",x"07",x"0F",x"2F",x"07",x"C0",x"D0",x"C8",x"E0",x"C8",x"C8",x"C0",x"E4",
		x"07",x"07",x"0E",x"0F",x"0F",x"01",x"00",x"00",x"C0",x"E0",x"F1",x"F9",x"FC",x"D2",x"01",x"19",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F2",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F3",x"E0",x"C0",x"C0",x"80",x"80",x"0F",
		x"FF",x"FC",x"FC",x"FC",x"FD",x"FE",x"FE",x"FE",x"70",x"00",x"00",x"02",x"1C",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"0E",x"07",x"03",x"00",x"01",x"03",x"06",
		x"00",x"00",x"08",x"00",x"00",x"10",x"10",x"10",x"0D",x"8E",x"C6",x"37",x"0E",x"0F",x"0C",x"1E",
		x"00",x"20",x"98",x"E8",x"F1",x"19",x"CD",x"C9",x"00",x"00",x"00",x"00",x"00",x"30",x"31",x"21",
		x"91",x"31",x"39",x"38",x"9D",x"0D",x"14",x"04",x"41",x"79",x"71",x"F1",x"E0",x"E0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0A",x"02",x"27",x"68",x"71",x"E4",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"7F",x"FC",x"FA",x"10",x"22",x"10",x"10",x"60",x"F8",
		x"FC",x"FE",x"D1",x"B0",x"A0",x"E0",x"E0",x"D8",x"00",x"00",x"80",x"00",x"00",x"20",x"20",x"70",
		x"F8",x"DC",x"BC",x"AE",x"EE",x"A2",x"E0",x"A0",x"30",x"38",x"1C",x"18",x"00",x"00",x"00",x"00",
		x"BD",x"F7",x"FD",x"B3",x"FE",x"FE",x"40",x"00",x"DF",x"FA",x"FF",x"FD",x"EF",x"36",x"00",x"00",
		x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"40",x"44",x"65",x"63",x"A3",x"B7",x"BF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BE",x"BC",x"B8",x"F0",x"E0",x"E0",x"F0",x"F0",
		x"10",x"50",x"F8",x"FE",x"FE",x"CF",x"8F",x"07",x"0E",x"0C",x"0C",x"1C",x"38",x"38",x"78",x"79",
		x"01",x"03",x"07",x"03",x"00",x"04",x"06",x"06",x"D0",x"F0",x"E0",x"F0",x"F0",x"0F",x"03",x"01",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"80",x"83",x"87",
		x"81",x"87",x"1F",x"FE",x"C0",x"80",x"C0",x"00",x"FB",x"F1",x"80",x"00",x"00",x"00",x"01",x"01",
		x"00",x"00",x"00",x"00",x"04",x"0E",x"87",x"CF",x"01",x"0F",x"7F",x"1F",x"0B",x"02",x"30",x"A6",
		x"CF",x"8F",x"0F",x"13",x"1F",x"17",x"17",x"17",x"18",x"BB",x"F4",x"7C",x"96",x"FA",x"FE",x"FF",
		x"FE",x"EE",x"DC",x"FC",x"F0",x"49",x"02",x"CD",x"6C",x"26",x"FB",x"59",x"D8",x"D4",x"96",x"90",
		x"FF",x"3E",x"1E",x"1E",x"AE",x"AC",x"37",x"BF",x"90",x"12",x"04",x"1B",x"4D",x"41",x"00",x"00",
		x"A9",x"A9",x"A5",x"BC",x"9A",x"AB",x"BF",x"AF",x"20",x"20",x"90",x"08",x"C0",x"C0",x"E6",x"4C",
		x"BC",x"84",x"9C",x"D6",x"DE",x"DE",x"F6",x"F6",x"06",x"04",x"60",x"18",x"18",x"08",x"08",x"08",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"07",x"0F",x"0E",x"0F",x"3F",x"3D",x"3E",x"00",x"00",x"00",x"20",x"38",x"3C",x"7C",x"78",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"06",x"03",x"81",x"E0",x"F8",x"FE",x"FF",x"FF",x"61",x"04",x"FC",x"00",x"00",x"00",x"00",x"E0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
		x"00",x"00",x"00",x"E0",x"FC",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"E1",x"FD",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"07",x"07",x"03",x"02",x"05",x"02",x"2D",x"95",x"FF",x"EB",x"95",x"B5",x"EA",x"A5",x"52",x"25",
		x"DF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"E4",x"C0",x"AA",x"E2",x"C4",x"A0",x"E2",
		x"FF",x"FF",x"BB",x"5C",x"D6",x"AB",x"92",x"6D",x"C1",x"C7",x"E7",x"4B",x"A1",x"CB",x"E2",x"7A",
		x"57",x"79",x"E9",x"68",x"6D",x"6A",x"6F",x"5F",x"B8",x"A8",x"D0",x"6C",x"DE",x"2C",x"1F",x"5F",
		x"6F",x"6D",x"4A",x"77",x"DE",x"C4",x"E1",x"F1",x"9E",x"3E",x"4F",x"AC",x"52",x"D7",x"71",x"3B",
		x"7E",x"6E",x"77",x"73",x"53",x"73",x"5B",x"71",x"0C",x"08",x"04",x"00",x"0C",x"02",x"02",x"84",
		x"68",x"18",x"0D",x"2D",x"01",x"7E",x"7E",x"7E",x"94",x"8C",x"8C",x"8B",x"9F",x"63",x"77",x"73",
		x"3F",x"7E",x"6E",x"7C",x"7C",x"FE",x"FE",x"FC",x"38",x"3C",x"32",x"78",x"70",x"68",x"42",x"E8",
		x"F8",x"FC",x"FD",x"FF",x"FF",x"FD",x"FE",x"FF",x"94",x"A4",x"48",x"B0",x"CA",x"F0",x"A8",x"52",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FD",x"FD",x"EB",x"FC",x"B5",
		x"FF",x"FE",x"FE",x"FC",x"F6",x"FF",x"FA",x"AF",x"DD",x"D7",x"DD",x"9B",x"DF",x"76",x"5D",x"35",
		x"7A",x"EF",x"BB",x"5A",x"F3",x"BB",x"6E",x"FF",x"F0",x"A0",x"F0",x"E0",x"B8",x"AC",x"9E",x"BE",
		x"DB",x"7B",x"7B",x"56",x"FB",x"5F",x"9D",x"DB",x"BD",x"EB",x"7B",x"FA",x"F7",x"BB",x"3B",x"96",
		x"F0",x"F8",x"F8",x"78",x"18",x"2C",x"20",x"FC",x"88",x"88",x"C0",x"40",x"C0",x"61",x"60",x"7C",
		x"F8",x"FD",x"7D",x"FF",x"5F",x"FF",x"BF",x"6F",x"FE",x"1C",x"88",x"88",x"C9",x"E1",x"E7",x"F7",
		x"7F",x"7F",x"7F",x"7F",x"78",x"91",x"40",x"53",x"CB",x"D3",x"EB",x"E3",x"09",x"7F",x"BF",x"FF",
		x"81",x"81",x"01",x"01",x"81",x"80",x"D0",x"C0",x"FF",x"F3",x"E1",x"F1",x"F8",x"7E",x"3F",x"1F",
		x"7E",x"FF",x"5F",x"7B",x"BE",x"5F",x"3F",x"FF",x"D0",x"A8",x"D4",x"68",x"D2",x"B0",x"24",x"D0",
		x"6F",x"BE",x"DF",x"7D",x"FF",x"FB",x"FF",x"7D",x"A8",x"D0",x"72",x"A8",x"52",x"F0",x"68",x"A4",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FE",x"FB",x"F9",x"EB",x"EA",
		x"FF",x"FF",x"FE",x"FA",x"FA",x"EA",x"E8",x"A9",x"A9",x"A1",x"E9",x"A9",x"8B",x"89",x"A2",x"AA",
		x"AD",x"7A",x"AD",x"DD",x"B4",x"3B",x"BF",x"AB",x"AF",x"ED",x"EA",x"7F",x"EA",x"67",x"DA",x"6D",
		x"DB",x"BE",x"BB",x"7D",x"AB",x"BB",x"BB",x"75",x"7F",x"F3",x"BA",x"6B",x"6F",x"6E",x"BB",x"7E",
		x"60",x"F8",x"9C",x"F8",x"EE",x"5F",x"D9",x"B9",x"79",x"39",x"3A",x"14",x"30",x"54",x"54",x"9E",
		x"B9",x"6F",x"DD",x"75",x"DC",x"DE",x"D2",x"BC",x"B9",x"98",x"B8",x"9A",x"93",x"B3",x"30",x"30",
		x"CD",x"99",x"48",x"43",x"A7",x"A0",x"B2",x"32",x"4F",x"1F",x"9C",x"1E",x"1C",x"98",x"A4",x"9C",
		x"93",x"03",x"58",x"4C",x"AC",x"AC",x"24",x"54",x"06",x"66",x"E1",x"C6",x"43",x"43",x"43",x"66",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F2",x"E8",
		x"FF",x"FF",x"FE",x"F8",x"F0",x"E0",x"C0",x"F0",x"EE",x"92",x"0A",x"60",x"96",x"0A",x"0B",x"08",
		x"AE",x"A2",x"A2",x"8A",x"8A",x"A8",x"AA",x"6E",x"AA",x"CA",x"AA",x"A2",x"A8",x"AA",x"AB",x"A2",
		x"8A",x"BA",x"72",x"E2",x"AA",x"AE",x"A8",x"0A",x"AA",x"AE",x"4A",x"32",x"98",x"AA",x"AA",x"A2",
		x"F2",x"AE",x"FE",x"F6",x"7C",x"DE",x"D6",x"DF",x"C2",x"E1",x"E1",x"E9",x"49",x"45",x"54",x"75",
		x"BD",x"6D",x"F9",x"DB",x"FF",x"77",x"DF",x"5D",x"5A",x"B6",x"B7",x"F7",x"8B",x"5B",x"7A",x"FE",
		x"00",x"00",x"80",x"88",x"98",x"F8",x"F0",x"80",x"FA",x"FC",x"DE",x"FC",x"F8",x"E0",x"7C",x"7E",
		x"E1",x"69",x"7D",x"FD",x"D9",x"DF",x"DF",x"73",x"7E",x"7E",x"7E",x"3E",x"70",x"38",x"78",x"7C",
		x"FE",x"FF",x"FF",x"FB",x"FE",x"FF",x"FF",x"FF",x"D0",x"A8",x"D4",x"68",x"D2",x"B0",x"24",x"D0",
		x"FF",x"FE",x"FF",x"FD",x"FF",x"FB",x"FF",x"FD",x"A8",x"D0",x"72",x"A8",x"52",x"F0",x"68",x"A4",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
		x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"D2",x"83",x"12",x"15",x"12",x"45",x"67",x"33",x"3B",x"3B",
		x"02",x"03",x"03",x"02",x"02",x"00",x"10",x"68",x"19",x"0A",x"12",x"16",x"0B",x"1A",x"14",x"11",
		x"54",x"50",x"D8",x"F5",x"DB",x"9F",x"9B",x"13",x"3A",x"36",x"38",x"11",x"12",x"8A",x"CA",x"C6",
		x"F5",x"BE",x"AC",x"FD",x"DB",x"7D",x"FD",x"AD",x"D7",x"EB",x"EF",x"A7",x"FE",x"6B",x"DF",x"FD",
		x"BF",x"77",x"BD",x"9D",x"BF",x"F7",x"6F",x"BD",x"6F",x"CE",x"EF",x"6F",x"E9",x"FC",x"BD",x"ED",
		x"20",x"A8",x"AF",x"B0",x"03",x"09",x"05",x"10",x"7F",x"7E",x"7C",x"79",x"79",x"3B",x"B9",x"B9",
		x"0A",x"01",x"0A",x"05",x"02",x"01",x"0A",x"04",x"BB",x"79",x"FD",x"2B",x"B5",x"EF",x"57",x"BB",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"FA",x"F2",x"EA",x"C8",x"C0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"C1",x"C1",x"E3",x"F2",x"F8",x"FC",x"FE",
		x"01",x"03",x"85",x"BA",x"CE",x"9B",x"D3",x"0A",x"59",x"B0",x"12",x"A3",x"D1",x"B0",x"39",x"3A",
		x"40",x"B3",x"A5",x"D5",x"8A",x"E7",x"42",x"6C",x"AB",x"F1",x"B5",x"5C",x"5B",x"63",x"65",x"72",
		x"31",x"B9",x"21",x"3B",x"D5",x"4A",x"31",x"08",x"CA",x"4E",x"82",x"05",x"22",x"88",x"C6",x"A2",
		x"44",x"6C",x"11",x"45",x"13",x"55",x"16",x"93",x"52",x"61",x"21",x"40",x"49",x"80",x"82",x"C2",
		x"00",x"01",x"04",x"02",x"00",x"00",x"02",x"00",x"55",x"17",x"AB",x"5B",x"87",x"3D",x"D7",x"2B",
		x"01",x"04",x"00",x"02",x"00",x"00",x"04",x"01",x"4F",x"37",x"CD",x"9F",x"2B",x"97",x"2F",x"57",
		x"04",x"80",x"F0",x"F8",x"FC",x"FC",x"FF",x"FF",x"73",x"7B",x"D2",x"98",x"1B",x"13",x"03",x"82",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"F8",x"FC",x"FC",x"FE",x"FF",x"FF",
		x"C3",x"9C",x"2C",x"60",x"00",x"88",x"88",x"08",x"A0",x"80",x"82",x"1E",x"19",x"0A",x"06",x"83",
		x"19",x"0B",x"1E",x"0B",x"1E",x"02",x"8A",x"E2",x"82",x"E0",x"A0",x"E8",x"88",x"1C",x"E8",x"AA",
		x"F2",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"2A",x"8B",x"E8",x"82",x"AA",x"FA",x"F9",x"FA",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"AA",x"E2",x"8A",x"08",x"A8",x"AA",x"AB",x"2A",x"9A",x"2C",x"EA",x"EC",x"A6",x"8E",x"AC",x"AC",
		x"BA",x"EA",x"EA",x"AA",x"AA",x"EB",x"F2",x"FE",x"B9",x"A2",x"A9",x"AA",x"44",x"A2",x"87",x"AD",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"47",x"AB",x"B6",x"A7",x"FA",x"F7",x"F9",x"FD",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"DB",x"7D",x"D5",x"FD",x"B6",x"65",x"DE",x"DD",x"DE",x"F7",x"77",x"E4",x"B7",x"B3",x"B6",x"D7",
		x"55",x"FD",x"DD",x"F7",x"FD",x"FB",x"FE",x"FF",x"BF",x"F7",x"4F",x"9D",x"D7",x"D7",x"77",x"D9",
		x"9A",x"BA",x"8F",x"97",x"25",x"AE",x"04",x"32",x"C5",x"D9",x"91",x"08",x"F1",x"A0",x"79",x"04",
		x"4D",x"BB",x"2A",x"84",x"39",x"D6",x"3D",x"95",x"1F",x"50",x"22",x"D7",x"63",x"E5",x"81",x"C1",
		x"3F",x"2E",x"3C",x"3F",x"0B",x"18",x"15",x"02",x"C4",x"E0",x"70",x"92",x"D1",x"63",x"AD",x"91",
		x"4C",x"5A",x"AF",x"A2",x"20",x"62",x"36",x"7D",x"1F",x"8F",x"FF",x"A7",x"5F",x"EB",x"7D",x"F3",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"E1",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FE",x"F0",x"00",x"0F",x"FF",x"FF",x"FF",x"FF",x"3F",x"3B",x"18",x"E1",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"E0",x"C0",x"C0",x"F7",x"01",x"FD",x"17",x"FF",x"7F",x"3F",x"38",x"FC",x"FD",x"FD",x"FC",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"87",x"C3",x"40",x"40",x"C0",x"C3",x"40",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"FF",x"FF",x"FC",x"FF",x"FF",x"FF",
		x"F0",x"E0",x"C3",x"07",x"0F",x"3F",x"FF",x"FF",x"0F",x"03",x"FC",x"FE",x"FE",x"FE",x"80",x"80",
		x"E0",x"80",x"3F",x"FF",x"00",x"C0",x"FC",x"F8",x"7F",x"00",x"1F",x"E0",x"20",x"07",x"04",x"07",
		x"F8",x"F8",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"07",x"07",x"07",x"07",x"07",x"07",x"8F",x"88",
		x"FF",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",
		x"00",x"00",x"F8",x"F0",x"F8",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"F8",x"00",x"00",x"00",
		x"FF",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"00",x"08",x"C4",x"04",x"0D",
		x"00",x"03",x"FF",x"F7",x"FB",x"01",x"00",x"00",x"7D",x"FD",x"E3",x"03",x"03",x"F0",x"FC",x"7C",
		x"1F",x"4F",x"FE",x"06",x"07",x"00",x"3F",x"C0",x"40",x"0F",x"7F",x"FF",x"FC",x"01",x"FF",x"00",
		x"C0",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"C0",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"03",x"27",x"EF",x"FE",x"0F",x"FF",x"9F",x"0F",x"56",x"C9",x"9A",x"E1",x"E8",x"92",x"68",x"C1",
		x"03",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"A8",x"CD",x"CE",x"EE",x"0C",x"0C",x"0C",x"0C",
		x"DF",x"00",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"01",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"07",x"C0",x"F8",x"FF",x"FF",x"FF",x"F0",x"F0",x"F1",x"61",x"1B",x"3B",x"CF",x"CF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"17",x"01",x"FD",x"F7",x"F0",x"FC",x"C0",x"C7",x"E0",x"E0",x"E0",x"E1",x"1D",x"1D",x"3B",x"CF",
		x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",x"43",x"41",x"7F",x"E7",x"FF",x"E7",x"F8",x"E2",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"82",x"FE",x"FD",x"FB",x"F7",x"EF",x"DC",x"BC",
		x"03",x"C0",x"F8",x"FF",x"FF",x"FF",x"0F",x"FF",x"80",x"00",x"00",x"FE",x"FD",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"03",x"81",
		x"00",x"00",x"FF",x"FF",x"FF",x"F8",x"F8",x"F8",x"F8",x"F8",x"00",x"00",x"00",x"FF",x"8F",x"8F",
		x"FC",x"86",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"FC",x"F8",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"00",x"00",x"FF",x"F8",x"F0",x"F8",x"FF",x"FF",x"07",
		x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"07",x"06",x"04",x"04",x"04",x"05",x"05",x"05",
		x"00",x"FF",x"FF",x"F8",x"F0",x"F8",x"FF",x"FB",x"3F",x"FF",x"F0",x"F0",x"FC",x"FC",x"F0",x"F0",
		x"7B",x"7B",x"FB",x"FB",x"FB",x"FA",x"FA",x"FA",x"FC",x"F8",x"CF",x"CF",x"CF",x"7F",x"7F",x"7F",
		x"C0",x"03",x"46",x"03",x"40",x"03",x"46",x"03",x"01",x"C0",x"00",x"C0",x"00",x"C0",x"00",x"C0",
		x"40",x"00",x"C0",x"40",x"C0",x"40",x"C1",x"41",x"00",x"00",x"00",x"00",x"00",x"7C",x"FE",x"FC",
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F1",x"F1",x"F3",x"F3",x"E3",x"E7",x"E7",x"E7",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"CE",x"8E",x"8E",x"8E",x"8E",x"8E",
		x"9F",x"9F",x"9F",x"9D",x"1E",x"1F",x"1F",x"1F",x"8E",x"4B",x"1E",x"8F",x"0D",x"5E",x"9F",x"0E",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1E",x"1E",x"A7",x"F3",x"A1",x"E4",x"C8",x"EC",x"DC",x"7C",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"F8",x"F8",x"FF",x"FF",x"EF",x"9F",x"7F",x"3F",x"0F",x"03",
		x"F0",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"80",x"E0",x"F0",x"FC",x"FF",
		x"FF",x"FE",x"FD",x"FB",x"F3",x"F9",x"FC",x"FE",x"7F",x"F9",x"F9",x"FF",x"F3",x"F3",x"FF",x"79",
		x"FF",x"7F",x"3F",x"0F",x"03",x"01",x"00",x"00",x"39",x"9F",x"CC",x"E4",x"F3",x"F9",x"FC",x"7E",
		x"FF",x"F8",x"F8",x"FF",x"F0",x"F0",x"FF",x"F8",x"85",x"05",x"05",x"85",x"05",x"05",x"85",x"05",
		x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"05",x"85",x"83",x"87",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"87",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"FF",x"C3",x"C3",x"FF",x"C3",x"C3",x"FF",
		x"FF",x"FF",x"FF",x"87",x"87",x"FF",x"87",x"87",x"FF",x"FF",x"FF",x"C3",x"C3",x"FF",x"C3",x"C3",
		x"FF",x"FF",x"E1",x"E1",x"FF",x"E1",x"E1",x"FF",x"E9",x"E9",x"E9",x"E9",x"EB",x"EB",x"EB",x"EB",
		x"FF",x"FF",x"FF",x"E1",x"E1",x"FF",x"E1",x"E1",x"EB",x"EB",x"EB",x"EB",x"E9",x"ED",x"ED",x"ED",
		x"F3",x"F3",x"E3",x"9F",x"9F",x"1F",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",
		x"FF",x"9F",x"9F",x"9F",x"F3",x"F3",x"F3",x"FE",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"7F",
		x"FF",x"FF",x"01",x"79",x"81",x"79",x"01",x"01",x"80",x"81",x"B3",x"A0",x"80",x"A0",x"A0",x"80",
		x"01",x"79",x"81",x"79",x"01",x"01",x"FF",x"FF",x"A0",x"A0",x"80",x"A0",x"B3",x"81",x"80",x"FC",
		x"00",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"8E",x"8E",x"8E",x"8E",x"8E",x"9E",x"9C",x"9C",
		x"00",x"00",x"00",x"00",x"FE",x"FF",x"00",x"00",x"9C",x"9C",x"9C",x"9C",x"9C",x"1C",x"1C",x"1C",
		x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"7C",x"2A",x"04",x"09",x"14",x"1E",x"3C",x"39",
		x"1E",x"1E",x"1E",x"1E",x"1F",x"1F",x"1E",x"1E",x"36",x"7D",x"7C",x"F1",x"E4",x"EA",x"74",x"F9",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"F8",x"C7",x"FF",x"F8",x"FF",x"FF",x"F0",x"00",x"3E",x"FE",x"FE",x"00",x"80",x"FC",
		x"FF",x"FF",x"FF",x"FF",x"FC",x"FF",x"FF",x"FF",x"FC",x"FF",x"FC",x"F3",x"3F",x"FC",x"FF",x"FF",
		x"F0",x"7B",x"00",x"7B",x"7B",x"00",x"00",x"7B",x"7E",x"FF",x"00",x"FF",x"FF",x"00",x"00",x"FF",
		x"F0",x"C7",x"3C",x"FF",x"FC",x"03",x"C3",x"FF",x"1F",x"E0",x"00",x"F7",x"00",x"F7",x"F7",x"FF",
		x"00",x"F1",x"06",x"8E",x"E6",x"03",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"FF",
		x"FF",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"F8",x"01",x"E7",x"FF",x"E3",
		x"00",x"FF",x"00",x"00",x"00",x"F0",x"00",x"F0",x"00",x"00",x"1F",x"00",x"00",x"3F",x"7F",x"FF",
		x"F1",x"03",x"F3",x"07",x"77",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"3E",x"3C",
		x"00",x"00",x"FF",x"FF",x"E1",x"00",x"7F",x"7F",x"0F",x"00",x"FF",x"FF",x"C7",x"00",x"FF",x"FF",
		x"3F",x"BF",x"BF",x"BF",x"BF",x"00",x"00",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"E3",
		x"FA",x"7A",x"7B",x"7B",x"7B",x"3B",x"BB",x"DB",x"7F",x"7F",x"CF",x"CF",x"CF",x"F8",x"F8",x"E0",
		x"DB",x"EB",x"EB",x"EB",x"EB",x"03",x"03",x"C3",x"E0",x"F8",x"F8",x"E0",x"E0",x"F8",x"C4",x"84",
		x"41",x"C0",x"40",x"C0",x"40",x"C0",x"00",x"43",x"8E",x"04",x"00",x"00",x"00",x"00",x"00",x"C0",
		x"06",x"43",x"00",x"43",x"06",x"43",x"00",x"7F",x"00",x"C0",x"00",x"C0",x"00",x"C0",x"01",x"FF",
		x"00",x"00",x"F8",x"18",x"F8",x"00",x"FA",x"0D",x"1C",x"1C",x"1C",x"38",x"38",x"7A",x"FF",x"EF",
		x"0A",x"0F",x"FE",x"3F",x"1F",x"7D",x"FE",x"FF",x"1E",x"57",x"E9",x"E4",x"A1",x"F0",x"55",x"2A",
		x"1E",x"1E",x"18",x"3E",x"7F",x"BE",x"F6",x"EF",x"FA",x"78",x"75",x"3C",x"5A",x"91",x"2A",x"04",
		x"6F",x"F6",x"C7",x"AB",x"F2",x"6C",x"E8",x"C5",x"0A",x"9C",x"07",x"22",x"85",x"42",x"00",x"68",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"F0",x"F0",x"F0",x"70",x"70",x"F0",x"F8",x"FE",x"18",x"31",x"31",x"18",x"0C",x"06",x"3F",x"3F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"81",x"F3",x"F3",x"81",x"F1",x"00",x"00",x"FF",x"02",x"E7",x"E7",x"02",x"E3",x"00",x"00",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"07",x"C6",x"C5",x"07",x"C7",x"04",x"07",x"FF",x"0D",x"7F",x"FF",x"E3",x"01",x"00",x"E0",x"FE",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"E0",x"E0",x"FF",x"FF",x"3F",x"00",x"02",x"02",x"00",x"09",x"FB",x"F7",x"D3",x"06",x"07",x"AB",
		x"CB",x"FF",x"FF",x"FF",x"FF",x"DF",x"AF",x"3D",x"C5",x"E1",x"C2",x"61",x"A9",x"C4",x"D0",x"B2",
		x"C5",x"F0",x"F8",x"D0",x"58",x"E9",x"F0",x"E3",x"FC",x"BA",x"1D",x"2C",x"2A",x"44",x"C6",x"E0",
		x"F1",x"B9",x"A8",x"D0",x"89",x"EC",x"BD",x"EF",x"92",x"E0",x"50",x"80",x"24",x"00",x"60",x"28",
		x"FD",x"F7",x"FF",x"FE",x"FB",x"FF",x"FE",x"FF",x"91",x"60",x"B4",x"C0",x"11",x"C8",x"F4",x"A2",
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"58",x"C4",x"B9",x"D0",x"EC",x"C9",x"BA",x"ED",
		x"FF",x"FC",x"FE",x"FE",x"FF",x"FE",x"FF",x"FF",x"EA",x"FC",x"E9",x"7A",x"1C",x"DA",x"1D",x"4C",
		x"FF",x"FE",x"FF",x"FD",x"FF",x"FB",x"FE",x"FD",x"89",x"86",x"EA",x"90",x"55",x"E2",x"B0",x"C9",
		x"FD",x"FE",x"FD",x"FA",x"FC",x"FE",x"FC",x"FB",x"6A",x"88",x"24",x"91",x"04",x"8A",x"C8",x"85",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D0",x"45",x"D8",x"B5",x"EA",x"FE",x"FF",x"FF",
		x"B0",x"04",x"A0",x"68",x"80",x"20",x"A1",x"94",x"07",x"47",x"66",x"2F",x"65",x"EE",x"C7",x"B6",
		x"41",x"03",x"95",x"97",x"4F",x"9F",x"15",x"BE",x"C7",x"CB",x"C1",x"AD",x"D2",x"68",x"91",x"C8",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"FE",x"FB",x"FE",x"FF",x"FD",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C8",x"E2",x"94",x"F1",x"68",x"AA",x"D0",x"E5",x"8D",x"07",x"8F",x"5A",x"1C",x"39",x"0A",x"3E",
		x"40",x"D8",x"88",x"5D",x"BF",x"BF",x"FF",x"FF",x"74",x"BD",x"FE",x"FD",x"FE",x"FB",x"FF",x"FF",
		x"1F",x"1F",x"8B",x"57",x"03",x"03",x"85",x"16",x"54",x"88",x"C1",x"90",x"60",x"80",x"12",x"A0",
		x"8E",x"1E",x"BF",x"36",x"7F",x"5F",x"3E",x"2B",x"08",x"80",x"54",x"82",x"C8",x"94",x"E4",x"B0",
		x"C7",x"6F",x"CF",x"87",x"43",x"83",x"88",x"23",x"7A",x"DC",x"F5",x"EA",x"FD",x"78",x"D0",x"01",
		x"87",x"06",x"17",x"B7",x"3F",x"F7",x"F6",x"3F",x"54",x"A0",x"D4",x"A1",x"43",x"97",x"87",x"57",
		x"07",x"0B",x"17",x"8E",x"1F",x"0F",x"1F",x"2E",x"AA",x"40",x"94",x"A0",x"48",x"B0",x"04",x"A1",
		x"9F",x"1F",x"8E",x"1F",x"0F",x"07",x"0B",x"07",x"50",x"84",x"D0",x"84",x"40",x"A9",x"C0",x"70",
		x"4F",x"0F",x"8F",x"07",x"07",x"03",x"83",x"02",x"A8",x"58",x"D2",x"E0",x"B4",x"E0",x"48",x"B0",
		x"00",x"81",x"43",x"01",x"03",x"87",x"03",x"07",x"F9",x"C0",x"AA",x"A8",x"D2",x"48",x"E4",x"98",
		x"88",x"28",x"41",x"EA",x"30",x"7C",x"39",x"7C",x"0A",x"1D",x"0E",x"1E",x"3A",x"1C",x"3D",x"52",
		x"28",x"BC",x"1A",x"3C",x"9E",x"6E",x"14",x"88",x"1C",x"9F",x"3C",x"1E",x"3D",x"1E",x"8F",x"0E",
		x"87",x"8B",x"47",x"AF",x"27",x"4F",x"E3",x"45",x"A8",x"62",x"E4",x"56",x"CC",x"98",x"F4",x"F8",
		x"73",x"E9",x"74",x"30",x"70",x"1A",x"90",x"42",x"DA",x"ED",x"FA",x"D4",x"52",x"28",x"80",x"20",
		x"43",x"61",x"23",x"71",x"28",x"70",x"E4",x"38",x"F7",x"E2",x"F9",x"F0",x"F9",x"EB",x"B7",x"55",
		x"70",x"65",x"B4",x"7B",x"51",x"28",x"38",x"11",x"2E",x"1D",x"1D",x"4C",x"08",x"A0",x"00",x"00",
		x"DA",x"E3",x"C2",x"ED",x"D2",x"CB",x"90",x"FD",x"00",x"24",x"08",x"05",x"04",x"02",x"00",x"40",
		x"B8",x"FC",x"F3",x"7B",x"E7",x"7B",x"2F",x"0F",x"C0",x"A0",x"02",x"40",x"A0",x"50",x"94",x"EA",
		x"00",x"24",x"88",x"0D",x"1A",x"8C",x"5E",x"1D",x"8D",x"47",x"16",x"0D",x"06",x"0F",x"16",x"0C",
		x"0E",x"9D",x"0D",x"1E",x"88",x"2C",x"04",x"80",x"5E",x"36",x"3D",x"66",x"73",x"C1",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"00",x"32",x"00",x"B0",x"3E",x"00",x"32",x"00",x"9E",x"3E",x"01",x"32",x"00",x"B8",x"31",
		x"00",x"90",x"C3",x"20",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"F5",x"3E",x"00",x"32",x"00",x"B0",x"F1",x"C3",x"C0",x"01",
		x"00",x"10",x"00",x"20",x"00",x"30",x"00",x"50",x"00",x"40",x"80",x"8F",x"00",x"8F",x"80",x"8E",
		x"00",x"8E",x"80",x"8D",x"05",x"00",x"20",x"20",x"20",x"20",x"40",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"05",x"00",x"00",x"00",x"00",x"00",x"20",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"05",x"FF",x"40",
		x"40",x"40",x"40",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C3",x"AD",x"01",x"C3",x"18",x"07",x"C3",x"92",x"01",x"C3",x"64",x"08",x"C3",x"50",x"08",x"C3",
		x"1D",x"0B",x"C3",x"41",x"0B",x"C3",x"21",x"0A",x"C3",x"FD",x"09",x"C3",x"82",x"0A",x"C3",x"98",
		x"0A",x"C3",x"EE",x"09",x"C3",x"AC",x"0B",x"C3",x"18",x"06",x"C3",x"B0",x"0B",x"C3",x"E4",x"0B",
		x"C3",x"F2",x"0B",x"C3",x"01",x"0C",x"C3",x"42",x"0C",x"C3",x"4C",x"0C",x"C3",x"0F",x"60",x"C3",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CD",x"C7",x"03",x"CD",x"20",x"07",x"31",x"00",x"90",x"21",x"00",x"80",x"01",x"00",x"08",x"CD",
		x"50",x"08",x"21",x"00",x"88",x"01",x"F6",x"07",x"CD",x"50",x"08",x"21",x"00",x"90",x"01",x"FF",
		x"03",x"CD",x"5A",x"08",x"21",x"00",x"94",x"01",x"FF",x"03",x"CD",x"50",x"08",x"21",x"20",x"98",
		x"01",x"60",x"00",x"CD",x"50",x"08",x"21",x"00",x"9C",x"01",x"00",x"01",x"CD",x"50",x"08",x"21",
		x"00",x"9A",x"01",x"C8",x"00",x"CD",x"50",x"08",x"3E",x"01",x"32",x"00",x"87",x"3E",x"01",x"32",
		x"01",x"87",x"3A",x"04",x"B0",x"32",x"13",x"80",x"3A",x"05",x"B0",x"32",x"14",x"80",x"CD",x"B9",
		x"02",x"CD",x"08",x"09",x"CD",x"18",x"06",x"3E",x"01",x"32",x"8C",x"80",x"21",x"01",x"00",x"22",
		x"22",x"80",x"3E",x"00",x"32",x"00",x"B0",x"3E",x"FF",x"32",x"02",x"80",x"31",x"00",x"90",x"3E",
		x"00",x"32",x"03",x"80",x"21",x"84",x"00",x"CD",x"68",x"03",x"C3",x"05",x"02",x"3E",x"00",x"32",
		x"00",x"B0",x"3E",x"00",x"32",x"03",x"80",x"21",x"90",x"00",x"CD",x"68",x"03",x"C3",x"05",x"02",
		x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"CD",x"9F",x"02",x"31",x"00",x"90",x"00",x"00",
		x"00",x"CD",x"58",x"09",x"CD",x"AB",x"09",x"CD",x"1B",x"60",x"CD",x"12",x"60",x"CD",x"82",x"03",
		x"CD",x"2F",x"06",x"CD",x"D9",x"5F",x"CD",x"BD",x"02",x"CD",x"64",x"08",x"CD",x"E2",x"09",x"3A",
		x"77",x"80",x"B7",x"20",x"05",x"CD",x"65",x"03",x"18",x"0B",x"3E",x"00",x"32",x"03",x"80",x"21",
		x"84",x"00",x"CD",x"68",x"03",x"3A",x"03",x"80",x"B7",x"C2",x"47",x"02",x"3E",x"FF",x"32",x"02",
		x"80",x"3E",x"00",x"32",x"00",x"B0",x"3E",x"01",x"32",x"00",x"B0",x"06",x"05",x"0E",x"00",x"21",
		x"0E",x"80",x"7E",x"E6",x"30",x"C2",x"2E",x"02",x"7E",x"E6",x"C0",x"C2",x"35",x"02",x"23",x"0C",
		x"10",x"F0",x"C3",x"16",x"02",x"3E",x"00",x"32",x"00",x"B0",x"32",x"02",x"80",x"79",x"32",x"00",
		x"80",x"7E",x"E6",x"80",x"CA",x"68",x"02",x"2A",x"00",x"80",x"29",x"11",x"04",x"80",x"19",x"5E",
		x"23",x"56",x"EB",x"F9",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"3E",x"00",x"32",x"00",x"B0",
		x"3E",x"01",x"32",x"00",x"B0",x"F1",x"ED",x"45",x"36",x"80",x"2A",x"00",x"80",x"29",x"11",x"7A",
		x"00",x"19",x"5E",x"23",x"56",x"EB",x"F9",x"2A",x"00",x"80",x"29",x"11",x"70",x"00",x"19",x"5E",
		x"23",x"56",x"EB",x"3E",x"00",x"32",x"00",x"B0",x"3E",x"01",x"32",x"00",x"B0",x"E9",x"3E",x"00",
		x"32",x"00",x"B0",x"2A",x"00",x"80",x"11",x"0E",x"80",x"19",x"CB",x"BE",x"C3",x"05",x"02",x"3A",
		x"02",x"80",x"FE",x"FF",x"C8",x"2A",x"00",x"80",x"29",x"11",x"04",x"80",x"19",x"EB",x"21",x"00",
		x"00",x"39",x"23",x"23",x"EB",x"73",x"23",x"72",x"C9",x"CD",x"D0",x"5F",x"C9",x"3A",x"02",x"B0",
		x"E6",x"01",x"C2",x"D0",x"02",x"DD",x"21",x"15",x"80",x"26",x"00",x"CD",x"EE",x"02",x"18",x"05",
		x"3E",x"01",x"32",x"15",x"80",x"3A",x"02",x"B0",x"E6",x"02",x"C2",x"E8",x"02",x"DD",x"21",x"82",
		x"80",x"26",x"01",x"CD",x"EE",x"02",x"18",x"05",x"3E",x"01",x"32",x"82",x"80",x"C9",x"DD",x"7E",
		x"00",x"FE",x"00",x"28",x"6F",x"3A",x"17",x"80",x"32",x"90",x"80",x"7C",x"FE",x"00",x"28",x"17",
		x"3A",x"84",x"80",x"FE",x"FF",x"20",x"10",x"3A",x"85",x"80",x"3C",x"32",x"85",x"80",x"FE",x"02",
		x"38",x"4E",x"3E",x"00",x"32",x"85",x"80",x"DD",x"46",x"01",x"3A",x"17",x"80",x"FE",x"99",x"D2",
		x"33",x"03",x"3A",x"17",x"80",x"C6",x"01",x"27",x"32",x"17",x"80",x"05",x"78",x"FE",x"00",x"20",
		x"E9",x"18",x"07",x"3A",x"87",x"80",x"80",x"32",x"87",x"80",x"DD",x"36",x"00",x"00",x"3A",x"70",
		x"80",x"B7",x"C0",x"CD",x"F0",x"00",x"3E",x"10",x"CD",x"FC",x"00",x"3A",x"81",x"80",x"B7",x"28",
		x"07",x"3A",x"90",x"80",x"FE",x"01",x"20",x"0C",x"3E",x"00",x"32",x"03",x"80",x"C3",x"C6",x"00",
		x"DD",x"36",x"00",x"00",x"C9",x"21",x"9D",x"00",x"11",x"0E",x"80",x"46",x"23",x"7E",x"FE",x"FF",
		x"28",x"08",x"23",x"7E",x"12",x"13",x"10",x"FA",x"18",x"07",x"23",x"1A",x"B6",x"12",x"13",x"10",
		x"F9",x"C9",x"F5",x"C5",x"E5",x"21",x"18",x"80",x"3A",x"27",x"80",x"47",x"3A",x"70",x"80",x"B7",
		x"C2",x"98",x"03",x"3A",x"7A",x"80",x"18",x"0A",x"3A",x"00",x"B0",x"CB",x"40",x"28",x"03",x"C3",
		x"E0",x"0F",x"01",x"00",x"05",x"1F",x"30",x"15",x"CB",x"16",x"F5",x"7E",x"FE",x"03",x"28",x"07",
		x"F1",x"23",x"30",x"0B",x"34",x"18",x"09",x"F1",x"23",x"36",x"FF",x"18",x"03",x"71",x"23",x"71",
		x"23",x"10",x"E2",x"E1",x"C1",x"F1",x"C9",x"3E",x"00",x"32",x"8F",x"80",x"CD",x"18",x"06",x"3E",
		x"01",x"32",x"8C",x"80",x"CD",x"AB",x"09",x"21",x"20",x"98",x"01",x"60",x"00",x"CD",x"CC",x"00",
		x"21",x"00",x"90",x"01",x"00",x"04",x"CD",x"CC",x"00",x"21",x"00",x"94",x"01",x"00",x"04",x"CD",
		x"CC",x"00",x"21",x"62",x"C6",x"11",x"C0",x"9C",x"01",x"40",x"00",x"ED",x"B0",x"CD",x"CF",x"00",
		x"B8",x"C5",x"16",x"CD",x"CF",x"00",x"A2",x"C6",x"08",x"FD",x"21",x"56",x"C3",x"FD",x"6E",x"00",
		x"FD",x"66",x"01",x"AF",x"4F",x"57",x"5F",x"06",x"08",x"7E",x"0F",x"30",x"07",x"1C",x"20",x"04",
		x"14",x"20",x"01",x"0C",x"C3",x"10",x"1F",x"E6",x"10",x"C2",x"39",x"05",x"10",x"EC",x"23",x"FD",
		x"7E",x"02",x"BD",x"20",x"E2",x"FD",x"7E",x"03",x"BC",x"20",x"DC",x"CD",x"6C",x"05",x"FD",x"7E",
		x"0C",x"FD",x"A6",x"0D",x"FE",x"FF",x"28",x"07",x"11",x"0C",x"00",x"FD",x"19",x"18",x"BE",x"FD",
		x"21",x"94",x"C3",x"FD",x"6E",x"00",x"FD",x"66",x"01",x"C3",x"20",x"1F",x"E6",x"10",x"C2",x"39",
		x"05",x"3E",x"FF",x"AE",x"77",x"23",x"7D",x"FD",x"BE",x"02",x"20",x"ED",x"7C",x"FD",x"BE",x"03",
		x"20",x"E7",x"FD",x"6E",x"00",x"FD",x"66",x"01",x"11",x"00",x"00",x"D9",x"11",x"00",x"00",x"D9",
		x"06",x"08",x"7E",x"0F",x"30",x"03",x"13",x"18",x"03",x"D9",x"13",x"D9",x"10",x"F5",x"23",x"FD",
		x"7E",x"02",x"BD",x"20",x"EB",x"C3",x"20",x"3F",x"BC",x"20",x"E5",x"FD",x"6E",x"00",x"FD",x"66",
		x"01",x"C3",x"30",x"1F",x"E6",x"10",x"C2",x"39",x"05",x"3E",x"FF",x"AE",x"77",x"23",x"7D",x"FD",
		x"BE",x"02",x"20",x"ED",x"7C",x"FD",x"BE",x"03",x"20",x"E7",x"FD",x"6E",x"00",x"FD",x"66",x"01",
		x"06",x"08",x"7E",x"0F",x"30",x"03",x"13",x"18",x"03",x"D9",x"13",x"D9",x"10",x"F5",x"23",x"FD",
		x"7E",x"02",x"BD",x"20",x"EB",x"C3",x"30",x"3F",x"BC",x"20",x"E5",x"FD",x"4E",x"04",x"FD",x"46",
		x"05",x"D9",x"7B",x"D9",x"BB",x"20",x"06",x"D9",x"7A",x"D9",x"BA",x"28",x"06",x"FD",x"4E",x"06",
		x"FD",x"46",x"07",x"C5",x"DD",x"E1",x"C3",x"E0",x"1F",x"C3",x"C0",x"1F",x"FD",x"19",x"FD",x"7E",
		x"00",x"FD",x"A6",x"01",x"FE",x"FF",x"C2",x"53",x"04",x"21",x"6C",x"84",x"01",x"28",x"00",x"CD",
		x"CC",x"00",x"CD",x"8B",x"05",x"3E",x"01",x"32",x"15",x"80",x"06",x"04",x"C3",x"40",x"1F",x"E6",
		x"10",x"C2",x"39",x"05",x"21",x"FF",x"FF",x"C3",x"40",x"3F",x"20",x"FB",x"10",x"EE",x"C9",x"F5",
		x"3E",x"FF",x"3D",x"FE",x"00",x"20",x"FB",x"F1",x"C9",x"21",x"6C",x"84",x"01",x"28",x"00",x"CD",
		x"CC",x"00",x"DD",x"21",x"48",x"C6",x"CD",x"D2",x"00",x"C3",x"50",x"1F",x"E6",x"10",x"C2",x"56",
		x"05",x"3E",x"00",x"32",x"15",x"80",x"3A",x"15",x"80",x"B7",x"C2",x"65",x"05",x"3A",x"00",x"B0",
		x"E6",x"10",x"C2",x"6B",x"05",x"CD",x"8B",x"05",x"C3",x"49",x"05",x"C9",x"FD",x"6E",x"04",x"FD",
		x"66",x"05",x"B7",x"FD",x"4E",x"06",x"FD",x"46",x"07",x"ED",x"52",x"CA",x"84",x"05",x"FD",x"4E",
		x"08",x"FD",x"46",x"09",x"C5",x"DD",x"E1",x"CD",x"D2",x"00",x"C9",x"DD",x"21",x"81",x"84",x"FD",
		x"21",x"00",x"B0",x"11",x"14",x"00",x"21",x"E4",x"C5",x"06",x"05",x"C5",x"D5",x"E5",x"DD",x"E5",
		x"11",x"6C",x"84",x"01",x"14",x"00",x"ED",x"B0",x"C3",x"F7",x"1F",x"B7",x"CA",x"B9",x"05",x"CD",
		x"CE",x"05",x"DD",x"21",x"6C",x"84",x"CD",x"D2",x"00",x"DD",x"E1",x"E1",x"D1",x"C1",x"78",x"FE",
		x"03",x"C2",x"C6",x"05",x"FD",x"23",x"FD",x"23",x"19",x"DD",x"23",x"10",x"CE",x"C9",x"C5",x"DD",
		x"E5",x"DD",x"21",x"6E",x"84",x"FD",x"E5",x"C1",x"79",x"FE",x"02",x"C2",x"E3",x"05",x"06",x"04",
		x"C3",x"E5",x"05",x"06",x"08",x"FD",x"7E",x"00",x"B7",x"1F",x"D2",x"F4",x"05",x"DD",x"36",x"00",
		x"31",x"C3",x"F8",x"05",x"C3",x"80",x"1F",x"00",x"DD",x"23",x"DD",x"23",x"10",x"EA",x"DD",x"E1",
		x"C1",x"C9",x"DD",x"7E",x"00",x"FD",x"BE",x"00",x"CA",x"16",x"06",x"FD",x"7E",x"00",x"DD",x"77",
		x"00",x"3E",x"01",x"C3",x"17",x"06",x"AF",x"C9",x"11",x"00",x"8C",x"21",x"00",x"D5",x"01",x"00",
		x"01",x"ED",x"B0",x"11",x"00",x"88",x"21",x"1A",x"0F",x"01",x"70",x"00",x"ED",x"B0",x"C9",x"C5",
		x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"DD",x"21",x"00",x"88",x"DD",x"7E",x"00",x"FE",x"FF",x"CA",
		x"A8",x"06",x"DD",x"CB",x"00",x"7E",x"C2",x"95",x"06",x"DD",x"7E",x"03",x"DD",x"BE",x"07",x"28",
		x"03",x"D2",x"9D",x"06",x"DD",x"36",x"07",x"00",x"DD",x"66",x"02",x"DD",x"6E",x"01",x"16",x"00",
		x"DD",x"5E",x"08",x"19",x"E5",x"23",x"23",x"0E",x"00",x"23",x"7E",x"FE",x"FF",x"28",x"05",x"DD",
		x"4E",x"08",x"0C",x"0C",x"DD",x"71",x"08",x"E1",x"FD",x"21",x"00",x"00",x"11",x"10",x"00",x"DD",
		x"7E",x"00",x"E6",x"7F",x"FE",x"00",x"28",x"05",x"FD",x"19",x"3D",x"18",x"F7",x"11",x"00",x"8C",
		x"FD",x"19",x"CD",x"B0",x"06",x"11",x"0A",x"00",x"DD",x"19",x"C3",x"3A",x"06",x"DD",x"34",x"07",
		x"11",x"0A",x"00",x"DD",x"19",x"C3",x"3A",x"06",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",
		x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"7E",x"32",x"72",x"88",x"23",x"7E",x"32",x"73",x"88",
		x"DD",x"7E",x"05",x"87",x"11",x"00",x"00",x"5F",x"FD",x"19",x"FD",x"E5",x"DD",x"4E",x"06",x"0D",
		x"11",x"02",x"00",x"DD",x"7E",x"04",x"FE",x"01",x"28",x"03",x"11",x"FE",x"FF",x"21",x"74",x"88",
		x"79",x"FE",x"00",x"28",x"0F",x"FD",x"7E",x"00",x"77",x"23",x"FD",x"7E",x"01",x"77",x"23",x"FD",
		x"19",x"0D",x"18",x"EC",x"FD",x"E1",x"21",x"72",x"88",x"DD",x"4E",x"06",x"79",x"FE",x"00",x"28",
		x"0F",x"7E",x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77",x"01",x"23",x"FD",x"19",x"0D",x"18",x"EC",
		x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",x"3A",x"70",x"80",x"B7",x"C2",x"8E",x"02",x"C9",
		x"DD",x"21",x"00",x"90",x"FD",x"21",x"00",x"94",x"01",x"00",x"00",x"78",x"FE",x"10",x"28",x"3A",
		x"79",x"FE",x"10",x"20",x"0A",x"04",x"0E",x"00",x"11",x"20",x"00",x"DD",x"19",x"FD",x"19",x"DD",
		x"36",x"00",x"5C",x"DD",x"36",x"01",x"5D",x"DD",x"36",x"20",x"5E",x"DD",x"36",x"21",x"5F",x"FD",
		x"36",x"00",x"05",x"FD",x"36",x"01",x"05",x"FD",x"36",x"20",x"05",x"FD",x"36",x"21",x"05",x"DD",
		x"23",x"DD",x"23",x"FD",x"23",x"FD",x"23",x"0C",x"18",x"C1",x"06",x"00",x"21",x"FF",x"FF",x"C3",
		x"90",x"1F",x"CB",x"67",x"20",x"0C",x"2B",x"7C",x"B5",x"20",x"F4",x"04",x"78",x"FE",x"03",x"38",
		x"EB",x"C9",x"16",x"FF",x"15",x"7A",x"20",x"FC",x"C3",x"A0",x"1F",x"CB",x"67",x"28",x"F3",x"16",
		x"FF",x"15",x"7A",x"20",x"FC",x"C3",x"B0",x"1F",x"CB",x"67",x"20",x"F3",x"04",x"78",x"FE",x"03",
		x"38",x"E0",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"36",x"00",x"23",x"0B",x"79",x"B0",x"C2",x"50",x"08",x"C9",x"36",x"00",x"23",x"0B",x"79",x"B0",
		x"C2",x"5A",x"08",x"C9",x"D5",x"E5",x"2A",x"24",x"80",x"5D",x"54",x"19",x"19",x"E5",x"2A",x"22",
		x"80",x"5D",x"54",x"CB",x"23",x"CB",x"12",x"19",x"22",x"22",x"80",x"E1",x"ED",x"5A",x"22",x"24",
		x"80",x"E1",x"D1",x"C9",x"07",x"11",x"54",x"05",x"2E",x"05",x"54",x"05",x"FF",x"FF",x"09",x"11",
		x"45",x"05",x"2E",x"05",x"45",x"05",x"FF",x"FF",x"0B",x"11",x"48",x"05",x"2E",x"05",x"48",x"05",
		x"FF",x"FF",x"0D",x"11",x"4B",x"05",x"2E",x"05",x"4B",x"05",x"FF",x"FF",x"0F",x"11",x"41",x"05",
		x"2E",x"05",x"41",x"05",x"FF",x"FF",x"11",x"11",x"4E",x"05",x"2E",x"05",x"4E",x"05",x"FF",x"FF",
		x"13",x"11",x"4C",x"05",x"2E",x"05",x"4C",x"05",x"FF",x"FF",x"15",x"11",x"54",x"05",x"2E",x"05",
		x"54",x"05",x"FF",x"FF",x"17",x"11",x"44",x"05",x"2E",x"05",x"44",x"05",x"FF",x"FF",x"19",x"11",
		x"2E",x"05",x"2E",x"05",x"2E",x"05",x"FF",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"10",x"00",
		x"00",x"00",x"03",x"00",x"00",x"00",x"05",x"00",x"00",x"00",x"10",x"00",x"00",x"00",x"05",x"00",
		x"00",x"00",x"10",x"00",x"00",x"00",x"05",x"00",x"21",x"00",x"B0",x"06",x"10",x"36",x"00",x"23",
		x"10",x"FB",x"21",x"84",x"08",x"11",x"32",x"81",x"01",x"64",x"00",x"ED",x"B0",x"11",x"00",x"81",
		x"06",x"0A",x"0E",x"04",x"CD",x"45",x"09",x"ED",x"A0",x"79",x"B7",x"20",x"FA",x"10",x"F3",x"CD",
		x"45",x"09",x"11",x"E2",x"80",x"01",x"04",x"00",x"ED",x"B0",x"21",x"28",x"81",x"06",x"0A",x"36",
		x"01",x"23",x"10",x"FB",x"C9",x"C5",x"D5",x"3A",x"14",x"80",x"E6",x"07",x"21",x"E8",x"08",x"01",
		x"04",x"00",x"CD",x"F6",x"00",x"D1",x"C1",x"C9",x"DD",x"21",x"78",x"98",x"FD",x"21",x"20",x"98",
		x"21",x"00",x"85",x"06",x"0C",x"0E",x"03",x"78",x"FE",x"00",x"28",x"11",x"23",x"7E",x"2B",x"CB",
		x"6F",x"20",x"05",x"CD",x"82",x"09",x"18",x"EF",x"CD",x"96",x"09",x"18",x"EA",x"79",x"32",x"00",
		x"9A",x"C9",x"05",x"C5",x"D5",x"DD",x"E5",x"D1",x"01",x"08",x"00",x"ED",x"B0",x"11",x"F8",x"FF",
		x"B7",x"DD",x"19",x"D1",x"C1",x"C9",x"0C",x"05",x"C5",x"D5",x"FD",x"E5",x"D1",x"01",x"08",x"00",
		x"ED",x"B0",x"11",x"08",x"00",x"B7",x"FD",x"19",x"D1",x"C1",x"C9",x"21",x"40",x"8C",x"11",x"40",
		x"9C",x"01",x"10",x"00",x"ED",x"B0",x"21",x"A0",x"8C",x"11",x"A0",x"9C",x"01",x"60",x"00",x"ED",
		x"B0",x"3A",x"8C",x"80",x"B7",x"C8",x"FE",x"02",x"28",x"12",x"3E",x"00",x"32",x"8C",x"80",x"21",
		x"00",x"8C",x"11",x"00",x"9C",x"01",x"A0",x"00",x"ED",x"B0",x"18",x"05",x"3E",x"00",x"32",x"8C",
		x"80",x"C9",x"2A",x"6E",x"80",x"7D",x"B4",x"28",x"04",x"2B",x"22",x"6E",x"80",x"C9",x"F5",x"ED",
		x"43",x"6E",x"80",x"ED",x"4B",x"6E",x"80",x"79",x"B0",x"20",x"F8",x"F1",x"C9",x"F5",x"C5",x"D5",
		x"E5",x"DD",x"E5",x"FD",x"E5",x"CD",x"8A",x"0B",x"C5",x"E1",x"4E",x"23",x"46",x"23",x"C5",x"DD",
		x"E1",x"CD",x"21",x"0A",x"3D",x"C2",x"0A",x"0A",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",
		x"C9",x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"CD",x"82",x"0A",x"E5",x"DD",x"7E",x"05",
		x"3D",x"CB",x"2F",x"16",x"00",x"5F",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"19",x"E5",x"D1",x"E1",
		x"0E",x"00",x"DD",x"46",x"05",x"78",x"3D",x"20",x"02",x"0E",x"0F",x"CD",x"59",x"0A",x"10",x"F5",
		x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",x"C9",x"1A",x"CB",x"40",x"C2",x"67",x"0A",x"E6",
		x"F0",x"0F",x"0F",x"0F",x"0F",x"18",x"02",x"E6",x"0F",x"CD",x"07",x"0B",x"77",x"D5",x"11",x"00",
		x"04",x"19",x"DD",x"7E",x"04",x"77",x"11",x"E0",x"FB",x"19",x"D1",x"CB",x"40",x"CA",x"81",x"0A",
		x"1B",x"C9",x"F5",x"DD",x"46",x"01",x"21",x"00",x"94",x"11",x"E0",x"FF",x"04",x"19",x"10",x"FD",
		x"06",x"00",x"DD",x"4E",x"00",x"09",x"F1",x"C9",x"F5",x"C5",x"D5",x"FD",x"E5",x"CB",x"38",x"CB",
		x"38",x"CB",x"38",x"CB",x"39",x"CB",x"39",x"CB",x"39",x"FD",x"21",x"C7",x"0A",x"16",x"00",x"CB",
		x"20",x"58",x"FD",x"19",x"FD",x"5E",x"00",x"FD",x"56",x"01",x"21",x"00",x"94",x"19",x"06",x"00",
		x"09",x"FD",x"E1",x"D1",x"C1",x"F1",x"C9",x"E0",x"FF",x"C0",x"FF",x"A0",x"FF",x"80",x"FF",x"60",
		x"FF",x"40",x"FF",x"20",x"FF",x"00",x"FF",x"E0",x"FE",x"C0",x"FE",x"A0",x"FE",x"80",x"FE",x"60",
		x"FE",x"40",x"FE",x"20",x"FE",x"00",x"FE",x"E0",x"FD",x"C0",x"FD",x"A0",x"FD",x"80",x"FD",x"60",
		x"FD",x"40",x"FD",x"20",x"FD",x"00",x"FD",x"E0",x"FC",x"C0",x"FC",x"A0",x"FC",x"80",x"FC",x"60",
		x"FC",x"40",x"FC",x"20",x"FC",x"00",x"FC",x"B7",x"20",x"07",x"B9",x"20",x"04",x"3E",x"00",x"18",
		x"0B",x"0E",x"0F",x"C6",x"30",x"FE",x"3A",x"DA",x"1C",x"0B",x"C6",x"07",x"C9",x"F5",x"C5",x"D5",
		x"E5",x"DD",x"E5",x"FD",x"E5",x"CD",x"8A",x"0B",x"C5",x"E1",x"4E",x"23",x"46",x"23",x"C5",x"DD",
		x"E1",x"CD",x"41",x"0B",x"3D",x"C2",x"2A",x"0B",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",
		x"C9",x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"CD",x"82",x"0A",x"DD",x"23",x"DD",x"23",
		x"DD",x"5E",x"00",x"DD",x"56",x"01",x"3E",x"FF",x"BA",x"CA",x"65",x"0B",x"CD",x"D3",x"5F",x"CD",
		x"9F",x"0B",x"C3",x"4C",x"0B",x"BB",x"CA",x"81",x"0B",x"7B",x"DD",x"23",x"DD",x"23",x"DD",x"5E",
		x"00",x"DD",x"56",x"01",x"CD",x"D3",x"5F",x"CD",x"9F",x"0B",x"3D",x"C2",x"77",x"0B",x"C3",x"4C",
		x"0B",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",x"C9",x"21",x"0E",x"00",x"39",x"5E",x"23",
		x"56",x"E5",x"EB",x"4E",x"23",x"46",x"23",x"7E",x"23",x"EB",x"E1",x"72",x"2B",x"73",x"C9",x"73",
		x"C5",x"01",x"00",x"04",x"09",x"72",x"01",x"E0",x"FB",x"09",x"C1",x"C9",x"CD",x"1E",x"60",x"C9",
		x"87",x"16",x"00",x"5F",x"19",x"5E",x"23",x"56",x"EB",x"E9",x"C5",x"D5",x"E5",x"DD",x"E5",x"DD",
		x"21",x"00",x"94",x"21",x"00",x"90",x"5F",x"16",x"00",x"19",x"DD",x"19",x"11",x"20",x"00",x"06",
		x"20",x"36",x"00",x"DD",x"36",x"00",x"0A",x"DD",x"19",x"19",x"05",x"C2",x"D1",x"0B",x"DD",x"E1",
		x"E1",x"D1",x"C1",x"C9",x"F5",x"C5",x"78",x"CD",x"BA",x"0B",x"3C",x"0D",x"C2",x"E7",x"0B",x"C1",
		x"F1",x"C9",x"DD",x"21",x"12",x"C8",x"CD",x"D2",x"00",x"DD",x"21",x"22",x"C8",x"CD",x"D5",x"00",
		x"C9",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"11",x"8A",x"0F",x"29",x"19",x"5E",x"23",x"56",x"26",
		x"00",x"6F",x"19",x"7E",x"DD",x"77",x"02",x"DD",x"36",x"03",x"05",x"3A",x"AC",x"81",x"16",x"00",
		x"5F",x"21",x"A8",x"0F",x"19",x"7E",x"FD",x"77",x"04",x"FD",x"36",x"05",x"05",x"DD",x"7E",x"04",
		x"C6",x"10",x"FD",x"77",x"06",x"DD",x"7E",x"05",x"FD",x"77",x"07",x"FD",x"E1",x"DD",x"E1",x"E1",
		x"D1",x"C9",x"B7",x"CA",x"4B",x"0C",x"09",x"3D",x"C2",x"46",x"0C",x"C9",x"B7",x"CA",x"55",x"0C",
		x"09",x"3D",x"C2",x"50",x"0C",x"5E",x"23",x"56",x"EB",x"C9",x"3A",x"00",x"B0",x"E6",x"20",x"CA",
		x"92",x"0C",x"3A",x"02",x"B0",x"E6",x"04",x"C2",x"62",x"0C",x"3A",x"00",x"B0",x"E6",x"20",x"CA",
		x"92",x"0C",x"3A",x"02",x"B0",x"E6",x"04",x"C2",x"7D",x"0C",x"C3",x"6A",x"0C",x"06",x"FF",x"3E",
		x"1C",x"3D",x"C2",x"81",x"0C",x"10",x"F8",x"3A",x"02",x"B0",x"E6",x"04",x"C2",x"92",x"0C",x"C3",
		x"6A",x"0C",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"00",x"FF",x"02",x"FF",x"04",x"FF",x"06",x"FF",x"08",x"FF",x"0A",x"FF",x"0C",x"FF",x"0F",
		x"CC",x"0F",x"AA",x"0F",x"88",x"0F",x"66",x"0F",x"44",x"0F",x"22",x"0F",x"00",x"0F",x"02",x"0F",
		x"04",x"0F",x"06",x"0F",x"08",x"0F",x"0A",x"0F",x"0C",x"0F",x"0F",x"0F",x"0F",x"0C",x"0F",x"0A",
		x"0F",x"08",x"0F",x"06",x"0F",x"04",x"0F",x"02",x"0F",x"00",x"2F",x"00",x"4F",x"00",x"6F",x"00",
		x"8F",x"00",x"AF",x"00",x"CF",x"00",x"FF",x"FF",x"0F",x"00",x"2F",x"00",x"4F",x"00",x"6F",x"00",
		x"8F",x"00",x"AF",x"00",x"CF",x"00",x"FF",x"00",x"FC",x"00",x"FA",x"00",x"F8",x"00",x"F6",x"00",
		x"F4",x"00",x"F2",x"00",x"F0",x"00",x"F0",x"02",x"F0",x"04",x"F0",x"06",x"F0",x"08",x"F0",x"0A",
		x"F0",x"0C",x"F0",x"0F",x"C0",x"0F",x"A0",x"0F",x"80",x"0F",x"60",x"0F",x"40",x"0F",x"20",x"0F",
		x"00",x"0F",x"02",x"0F",x"04",x"0F",x"06",x"0F",x"08",x"0F",x"0A",x"0F",x"0C",x"0F",x"0F",x"0F",
		x"0F",x"0C",x"0F",x"0A",x"0F",x"08",x"0F",x"06",x"0F",x"04",x"0F",x"02",x"FF",x"FF",x"00",x"0F",
		x"22",x"0F",x"44",x"0F",x"66",x"0F",x"88",x"0F",x"AA",x"0F",x"CC",x"0F",x"EE",x"0F",x"FF",x"FF",
		x"0F",x"00",x"2F",x"02",x"4F",x"04",x"6F",x"06",x"8F",x"08",x"AF",x"0A",x"CF",x"0C",x"EF",x"0E",
		x"FF",x"FF",x"0F",x"0F",x"2F",x"0F",x"4F",x"0F",x"6F",x"0F",x"8F",x"0F",x"AF",x"0F",x"CF",x"0F",
		x"EF",x"0F",x"FF",x"FF",x"F0",x"00",x"F2",x"02",x"F4",x"04",x"F6",x"06",x"F8",x"08",x"FA",x"0A",
		x"FC",x"0C",x"FE",x"0E",x"FF",x"FF",x"F0",x"0F",x"F2",x"0F",x"F4",x"0F",x"F6",x"0F",x"F8",x"0F",
		x"FA",x"0F",x"FC",x"0F",x"FE",x"0F",x"FF",x"FF",x"FF",x"00",x"FF",x"02",x"FF",x"04",x"FF",x"06",
		x"FF",x"08",x"FF",x"0A",x"FF",x"0C",x"FF",x"0E",x"FF",x"FF",x"FF",x"0F",x"EE",x"0E",x"DD",x"0D",
		x"CC",x"0C",x"BB",x"0B",x"AA",x"0A",x"99",x"09",x"88",x"08",x"FF",x"FF",x"0F",x"00",x"00",x"00",
		x"9F",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"0F",x"00",x"00",x"0F",x"00",x"00",x"00",
		x"9F",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"0F",x"00",x"00",x"0F",x"00",x"00",x"00",
		x"9F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"0F",x"00",x"00",x"00",x"0F",x"00",x"00",x"FF",x"00",
		x"00",x"00",x"9F",x"00",x"00",x"00",x"0F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"08",x"00",x"FF",x"FF",x"0F",x"0F",x"00",x"00",x"0F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0C",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"0D",x"00",x"0B",x"00",x"09",x"00",x"07",x"00",x"05",x"00",x"03",x"00",x"01",x"00",
		x"00",x"00",x"00",x"FF",x"CC",x"00",x"88",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"0F",x"FF",x"FF",x"00",x"0F",x"22",x"0F",x"44",x"0F",x"66",x"0F",x"88",x"0F",x"AA",x"0F",
		x"CC",x"0F",x"FF",x"0F",x"FF",x"FF",x"FF",x"00",x"FF",x"02",x"FF",x"04",x"FF",x"06",x"FF",x"08",
		x"FF",x"0A",x"FF",x"0C",x"FF",x"0F",x"FF",x"FF",x"0F",x"00",x"2F",x"02",x"4F",x"04",x"6F",x"06",
		x"8F",x"08",x"AF",x"0A",x"CF",x"0C",x"FF",x"0F",x"FF",x"FF",x"99",x"00",x"AA",x"00",x"BB",x"00",
		x"CC",x"00",x"DD",x"00",x"EE",x"00",x"FF",x"00",x"FF",x"FF",x"84",x"D0",x"0F",x"03",x"01",x"05",
		x"03",x"02",x"00",x"00",x"8A",x"00",x"00",x"04",x"01",x"01",x"06",x"00",x"00",x"00",x"8B",x"0A",
		x"0F",x"01",x"07",x"07",x"07",x"01",x"00",x"00",x"0C",x"C4",x"0E",x"02",x"01",x"07",x"01",x"00",
		x"00",x"00",x"0D",x"1C",x"0E",x"01",x"01",x"01",x"01",x"02",x"00",x"00",x"0D",x"46",x"0E",x"01",
		x"01",x"02",x"01",x"02",x"00",x"00",x"0D",x"70",x"0E",x"01",x"01",x"03",x"01",x"02",x"00",x"00",
		x"0D",x"9A",x"0E",x"04",x"01",x"04",x"01",x"02",x"00",x"00",x"0E",x"48",x"0D",x"02",x"07",x"07",
		x"07",x"04",x"00",x"00",x"0F",x"00",x"0D",x"02",x"07",x"07",x"07",x"02",x"00",x"00",x"04",x"BB",
		x"0F",x"03",x"01",x"01",x"01",x"03",x"00",x"00",x"FF",x"FF",x"92",x"0F",x"9A",x"0F",x"9D",x"0F",
		x"9F",x"0F",x"00",x"70",x"71",x"72",x"74",x"76",x"78",x"7A",x"77",x"79",x"7B",x"71",x"73",x"70",
		x"71",x"72",x"74",x"76",x"78",x"7A",x"7A",x"7A",x"00",x"7C",x"7D",x"7E",x"7F",x"FF",x"00",x"FB",
		x"00",x"F8",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"00",x"0C",x"00",x"08",
		x"00",x"04",x"00",x"00",x"00",x"04",x"00",x"08",x"00",x"0C",x"00",x"FF",x"FF",x"FF",x"FF",x"00",
		x"B0",x"0F",x"80",x"0F",x"50",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"3A",x"13",x"80",x"CB",x"77",x"C2",x"EE",x"0F",x"3A",x"01",x"B0",x"C3",x"A2",x"03",x"3A",x"00",
		x"B0",x"C3",x"A2",x"03",x"00",x"00",x"00",x"00",x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C9",x"00",
		x"3A",x"8E",x"80",x"FE",x"00",x"28",x"0B",x"3A",x"28",x"80",x"CB",x"97",x"32",x"28",x"80",x"C3",
		x"C3",x"00",x"DD",x"21",x"28",x"80",x"DD",x"CB",x"00",x"56",x"C2",x"DD",x"12",x"DD",x"CB",x"00",
		x"7E",x"28",x"42",x"DD",x"36",x"02",x"00",x"2A",x"36",x"80",x"2B",x"22",x"36",x"80",x"7C",x"B5",
		x"20",x"14",x"CD",x"F9",x"2F",x"CD",x"E6",x"2F",x"DD",x"CB",x"00",x"BE",x"DD",x"CB",x"00",x"B6",
		x"DD",x"36",x"02",x"00",x"18",x"1F",x"7C",x"B7",x"20",x"1B",x"7D",x"FE",x"39",x"30",x"16",x"E6",
		x"03",x"FE",x"00",x"20",x"10",x"DD",x"CB",x"00",x"76",x"28",x"06",x"DD",x"CB",x"00",x"B6",x"18",
		x"04",x"DD",x"CB",x"00",x"F6",x"DD",x"7E",x"19",x"DD",x"34",x"23",x"CB",x"5F",x"20",x"04",x"DD",
		x"36",x"23",x"00",x"E6",x"0A",x"28",x"0A",x"DD",x"7E",x"0B",x"FE",x"FF",x"28",x"03",x"C3",x"72",
		x"12",x"3A",x"3F",x"80",x"FE",x"00",x"28",x"17",x"3A",x"20",x"80",x"FE",x"03",x"C2",x"CE",x"12",
		x"DD",x"36",x"17",x"00",x"DD",x"36",x"0B",x"00",x"DD",x"36",x"1C",x"00",x"C3",x"72",x"12",x"DD",
		x"CB",x"00",x"4E",x"C2",x"D2",x"10",x"CD",x"DD",x"1A",x"7C",x"B5",x"20",x"1F",x"ED",x"5B",x"40",
		x"80",x"7A",x"B3",x"28",x"17",x"CB",x"5A",x"28",x"05",x"3E",x"11",x"CD",x"FD",x"1B",x"01",x"10",
		x"00",x"CD",x"E4",x"00",x"3A",x"53",x"84",x"F6",x"C0",x"32",x"53",x"84",x"DD",x"74",x"18",x"DD",
		x"75",x"19",x"CD",x"70",x"18",x"CD",x"B7",x"17",x"DD",x"7E",x"12",x"FE",x"FF",x"C2",x"25",x"12",
		x"2A",x"42",x"80",x"7C",x"B5",x"20",x"0A",x"2A",x"31",x"80",x"7C",x"B5",x"20",x"03",x"C3",x"38",
		x"11",x"DD",x"CB",x"00",x"46",x"C2",x"52",x"11",x"3A",x"20",x"80",x"FE",x"03",x"C2",x"1D",x"11",
		x"CD",x"73",x"17",x"3E",x"12",x"CD",x"FD",x"1B",x"DD",x"36",x"0B",x"00",x"DD",x"36",x"1C",x"00",
		x"DD",x"CB",x"19",x"5E",x"28",x"07",x"DD",x"CB",x"00",x"C6",x"C3",x"72",x"12",x"3A",x"41",x"80",
		x"CB",x"5F",x"28",x"11",x"DD",x"CB",x"00",x"46",x"20",x"0B",x"CD",x"73",x"17",x"DD",x"36",x"17",
		x"08",x"DD",x"CB",x"00",x"C6",x"C3",x"A7",x"11",x"3A",x"20",x"80",x"FE",x"03",x"20",x"10",x"3E",
		x"12",x"CD",x"FD",x"1B",x"DD",x"36",x"0B",x"00",x"DD",x"36",x"1C",x"00",x"C3",x"72",x"12",x"C3",
		x"A7",x"11",x"3A",x"20",x"80",x"FE",x"03",x"C2",x"77",x"11",x"CD",x"73",x"17",x"3E",x"12",x"CD",
		x"FD",x"1B",x"DD",x"36",x"0B",x"00",x"DD",x"36",x"1C",x"00",x"DD",x"CB",x"19",x"4E",x"28",x"07",
		x"DD",x"CB",x"00",x"86",x"C3",x"72",x"12",x"3A",x"41",x"80",x"CB",x"4F",x"28",x"11",x"DD",x"CB",
		x"00",x"46",x"28",x"0B",x"CD",x"73",x"17",x"DD",x"36",x"17",x"00",x"DD",x"CB",x"00",x"86",x"2A",
		x"42",x"80",x"CB",x"7C",x"20",x"04",x"7C",x"B5",x"20",x"0A",x"21",x"00",x"00",x"22",x"42",x"80",
		x"DD",x"CB",x"00",x"86",x"C3",x"A7",x"11",x"3A",x"41",x"80",x"CB",x"5F",x"28",x"12",x"2A",x"42",
		x"80",x"7C",x"B5",x"20",x"0B",x"21",x"00",x"00",x"22",x"31",x"80",x"22",x"38",x"80",x"18",x"1E",
		x"CD",x"E3",x"18",x"DD",x"CB",x"00",x"46",x"20",x"0C",x"2A",x"5A",x"80",x"11",x"0A",x"00",x"19",
		x"22",x"31",x"80",x"18",x"09",x"2A",x"5A",x"80",x"CD",x"D9",x"18",x"22",x"31",x"80",x"CD",x"9A",
		x"18",x"2A",x"42",x"80",x"ED",x"5B",x"31",x"80",x"3A",x"1C",x"80",x"FE",x"00",x"20",x"09",x"3A",
		x"1E",x"80",x"FE",x"00",x"20",x"09",x"18",x"0C",x"B7",x"CB",x"2A",x"CB",x"1B",x"18",x"05",x"B7",
		x"CB",x"23",x"CB",x"12",x"19",x"CB",x"7C",x"20",x"09",x"7C",x"B5",x"28",x"05",x"22",x"42",x"80",
		x"18",x"10",x"DD",x"CB",x"00",x"46",x"28",x"0A",x"21",x"00",x"00",x"22",x"42",x"80",x"DD",x"CB",
		x"00",x"86",x"C3",x"72",x"12",x"DD",x"CB",x"00",x"46",x"C2",x"4F",x"12",x"3A",x"20",x"80",x"FE",
		x"03",x"20",x"06",x"CD",x"73",x"17",x"CD",x"0D",x"17",x"3A",x"20",x"80",x"FE",x"FF",x"20",x"03",
		x"CD",x"33",x"17",x"3A",x"20",x"80",x"B7",x"20",x"03",x"CD",x"53",x"17",x"C3",x"1D",x"11",x"3A",
		x"20",x"80",x"FE",x"03",x"20",x"06",x"CD",x"73",x"17",x"CD",x"0D",x"17",x"3A",x"20",x"80",x"FE",
		x"FF",x"20",x"03",x"CD",x"33",x"17",x"3A",x"20",x"80",x"B7",x"20",x"03",x"CD",x"53",x"17",x"C3",
		x"77",x"11",x"DD",x"CB",x"00",x"9E",x"CD",x"8E",x"15",x"DD",x"CB",x"00",x"5E",x"20",x"03",x"CD",
		x"B4",x"14",x"CD",x"51",x"19",x"DD",x"CB",x"00",x"8E",x"3A",x"02",x"85",x"DD",x"BE",x"03",x"20",
		x"0C",x"3A",x"03",x"85",x"DD",x"BE",x"04",x"20",x"04",x"DD",x"CB",x"00",x"CE",x"DD",x"CB",x"00",
		x"7E",x"28",x"04",x"DD",x"36",x"02",x"0E",x"CD",x"F4",x"16",x"3A",x"3A",x"80",x"FE",x"FF",x"28",
		x"1A",x"FE",x"00",x"20",x"0F",x"3A",x"35",x"80",x"3C",x"32",x"35",x"80",x"CD",x"B7",x"17",x"CD",
		x"FC",x"17",x"18",x"07",x"3A",x"3A",x"80",x"3D",x"32",x"3A",x"80",x"C3",x"C3",x"00",x"3E",x"19",
		x"32",x"00",x"85",x"3A",x"3F",x"80",x"3D",x"32",x"3F",x"80",x"C3",x"C3",x"00",x"3A",x"95",x"80",
		x"FE",x"FF",x"28",x"06",x"CD",x"70",x"13",x"C3",x"6D",x"13",x"DD",x"21",x"5E",x"80",x"FD",x"21",
		x"00",x"85",x"3A",x"5F",x"80",x"FE",x"FF",x"28",x"2C",x"3E",x"01",x"CD",x"FC",x"00",x"3E",x"14",
		x"CD",x"FC",x"00",x"DD",x"36",x"00",x"00",x"DD",x"36",x"01",x"FF",x"FD",x"36",x"00",x"A4",x"FD",
		x"36",x"01",x"20",x"FD",x"7E",x"02",x"D6",x"08",x"FD",x"77",x"02",x"FD",x"7E",x"03",x"D6",x"08",
		x"FD",x"77",x"03",x"18",x"48",x"DD",x"7E",x"00",x"FE",x"40",x"D2",x"41",x"13",x"DD",x"34",x"00",
		x"DD",x"7E",x"00",x"FE",x"40",x"D2",x"41",x"13",x"E6",x"0F",x"20",x"31",x"FD",x"34",x"00",x"18",
		x"2C",x"21",x"00",x"00",x"22",x"00",x"85",x"3A",x"88",x"80",x"FE",x"00",x"20",x"1F",x"3A",x"8E",
		x"80",x"FE",x"00",x"20",x"18",x"3E",x"00",x"32",x"95",x"80",x"3A",x"70",x"80",x"FE",x"00",x"20",
		x"07",x"3E",x"01",x"32",x"78",x"80",x"18",x"05",x"3E",x"01",x"32",x"77",x"80",x"C3",x"C3",x"00",
		x"DD",x"21",x"95",x"80",x"DD",x"7E",x"00",x"E6",x"0F",x"FE",x"0F",x"28",x"0A",x"FE",x"07",x"28",
		x"06",x"CD",x"2D",x"14",x"C3",x"2C",x"14",x"21",x"00",x"00",x"22",x"31",x"80",x"CD",x"DD",x"1A",
		x"CB",x"5D",x"28",x"0C",x"DD",x"36",x"00",x"FF",x"3E",x"A7",x"CD",x"FC",x"00",x"C3",x"2C",x"14",
		x"DD",x"7E",x"00",x"FE",x"0F",x"28",x"27",x"DD",x"36",x"00",x"0F",x"2A",x"AA",x"14",x"DD",x"75",
		x"01",x"DD",x"74",x"02",x"DD",x"36",x"03",x"00",x"3A",x"03",x"85",x"DD",x"77",x"04",x"DD",x"36",
		x"05",x"00",x"DD",x"36",x"06",x"00",x"DD",x"36",x"07",x"00",x"DD",x"36",x"08",x"00",x"2A",x"9A",
		x"80",x"11",x"0A",x"00",x"19",x"22",x"9A",x"80",x"ED",x"5B",x"98",x"80",x"19",x"22",x"98",x"80",
		x"DD",x"34",x"07",x"DD",x"7E",x"07",x"FE",x"05",x"38",x"30",x"DD",x"36",x"07",x"00",x"FD",x"21",
		x"AA",x"14",x"16",x"00",x"DD",x"5E",x"08",x"FD",x"19",x"FD",x"7E",x"00",x"FE",x"FF",x"20",x"08",
		x"FD",x"21",x"AA",x"14",x"DD",x"36",x"08",x"00",x"DD",x"34",x"08",x"DD",x"34",x"08",x"FD",x"7E",
		x"00",x"DD",x"77",x"01",x"FD",x"7E",x"01",x"DD",x"77",x"02",x"3A",x"96",x"80",x"32",x"00",x"85",
		x"3A",x"97",x"80",x"32",x"01",x"85",x"3A",x"99",x"80",x"32",x"03",x"85",x"C9",x"DD",x"7E",x"00",
		x"FE",x"03",x"28",x"1F",x"3E",x"01",x"32",x"8D",x"80",x"DD",x"36",x"00",x"03",x"DD",x"36",x"07",
		x"00",x"DD",x"36",x"08",x"00",x"DD",x"36",x"09",x"00",x"3E",x"01",x"CD",x"FC",x"00",x"3E",x"27",
		x"CD",x"FC",x"00",x"DD",x"7E",x"07",x"FE",x"3C",x"38",x"07",x"DD",x"36",x"00",x"07",x"C3",x"9F",
		x"14",x"DD",x"7E",x"09",x"FE",x"03",x"38",x"2B",x"DD",x"36",x"09",x"00",x"FD",x"21",x"A0",x"14",
		x"16",x"00",x"DD",x"5E",x"08",x"B7",x"FD",x"19",x"FD",x"7E",x"00",x"FE",x"FF",x"20",x"08",x"FD",
		x"21",x"A0",x"14",x"DD",x"36",x"08",x"00",x"FD",x"7E",x"00",x"32",x"00",x"85",x"FD",x"7E",x"01",
		x"32",x"01",x"85",x"DD",x"34",x"07",x"DD",x"34",x"08",x"DD",x"34",x"08",x"DD",x"34",x"09",x"C9",
		x"28",x"C0",x"28",x"80",x"28",x"00",x"28",x"40",x"FF",x"FF",x"48",x"00",x"49",x"00",x"4A",x"00",
		x"4B",x"00",x"FF",x"FF",x"E5",x"D5",x"2A",x"2F",x"80",x"ED",x"5B",x"31",x"80",x"7A",x"B3",x"20",
		x"48",x"3A",x"41",x"80",x"CB",x"5F",x"28",x"41",x"7C",x"B5",x"20",x"11",x"3A",x"29",x"80",x"FE",
		x"1B",x"38",x"06",x"FE",x"23",x"30",x"02",x"18",x"5A",x"3E",x"18",x"18",x"56",x"CB",x"7C",x"20",
		x"14",x"DD",x"34",x"22",x"3A",x"4A",x"80",x"FE",x"04",x"DA",x"4B",x"15",x"DD",x"36",x"22",x"00",
		x"CD",x"4E",x"15",x"18",x"4B",x"DD",x"34",x"22",x"3A",x"4A",x"80",x"FE",x"04",x"DA",x"4B",x"15",
		x"DD",x"36",x"22",x"00",x"CD",x"6E",x"15",x"18",x"37",x"CB",x"7A",x"28",x"14",x"7C",x"B5",x"20",
		x"04",x"3E",x"23",x"18",x"1E",x"CB",x"7C",x"20",x"04",x"3E",x"25",x"18",x"16",x"3E",x"27",x"18",
		x"12",x"7C",x"B5",x"20",x"04",x"3E",x"24",x"18",x"0A",x"CB",x"7C",x"20",x"04",x"3E",x"26",x"18",
		x"02",x"3E",x"28",x"32",x"29",x"80",x"32",x"00",x"85",x"3E",x"93",x"CD",x"FD",x"1B",x"18",x"0B",
		x"32",x"29",x"80",x"32",x"00",x"85",x"3E",x"13",x"CD",x"FD",x"1B",x"D1",x"E1",x"C9",x"3A",x"29",
		x"80",x"FE",x"1B",x"F2",x"5A",x"15",x"3E",x"1B",x"18",x"13",x"FE",x"1E",x"28",x"06",x"38",x"04",
		x"3E",x"1B",x"18",x"09",x"3C",x"FE",x"1E",x"28",x"04",x"38",x"02",x"3E",x"1B",x"C9",x"3A",x"29",
		x"80",x"FE",x"1F",x"F2",x"7A",x"15",x"3E",x"1F",x"18",x"13",x"FE",x"22",x"28",x"06",x"38",x"04",
		x"3E",x"1F",x"18",x"09",x"3C",x"FE",x"22",x"28",x"04",x"38",x"02",x"3E",x"1F",x"C9",x"C5",x"D5",
		x"E5",x"DD",x"E5",x"DD",x"21",x"28",x"80",x"DD",x"7E",x"0B",x"FE",x"FF",x"CA",x"EE",x"16",x"DD",
		x"7E",x"1C",x"FE",x"02",x"CA",x"78",x"16",x"FE",x"01",x"CA",x"BC",x"15",x"DD",x"36",x"1D",x"28",
		x"DD",x"36",x"1E",x"00",x"DD",x"36",x"1F",x"00",x"DD",x"36",x"1C",x"01",x"3A",x"4B",x"80",x"FE",
		x"01",x"30",x"2A",x"3A",x"18",x"80",x"FE",x"00",x"20",x"07",x"3A",x"1A",x"80",x"FE",x"00",x"28",
		x"1C",x"DD",x"36",x"1D",x"00",x"DD",x"36",x"1E",x"00",x"DD",x"36",x"1F",x"00",x"DD",x"36",x"1C",
		x"02",x"21",x"00",x"00",x"22",x"42",x"80",x"22",x"31",x"80",x"C3",x"EE",x"16",x"DD",x"CB",x"00",
		x"DE",x"DD",x"7E",x"0B",x"FE",x"10",x"CA",x"3A",x"16",x"DA",x"3A",x"16",x"DD",x"36",x"1D",x"00",
		x"DD",x"36",x"1E",x"28",x"FE",x"20",x"CA",x"53",x"16",x"DA",x"53",x"16",x"DD",x"36",x"1E",x"04",
		x"DD",x"36",x"1C",x"02",x"DD",x"7E",x"19",x"E6",x"0A",x"28",x"0C",x"21",x"00",x"00",x"22",x"42",
		x"80",x"22",x"31",x"80",x"C3",x"6C",x"16",x"DD",x"7E",x"19",x"FE",x"00",x"28",x"06",x"CD",x"98",
		x"17",x"C3",x"6C",x"16",x"CD",x"73",x"17",x"C3",x"6C",x"16",x"DD",x"36",x"1D",x"00",x"DD",x"36",
		x"1E",x"04",x"DD",x"36",x"1F",x"02",x"01",x"FF",x"7F",x"CD",x"7A",x"17",x"DD",x"36",x"1C",x"02",
		x"C3",x"6C",x"16",x"3A",x"20",x"80",x"B7",x"C2",x"6C",x"16",x"DD",x"36",x"1E",x"04",x"DD",x"36",
		x"1F",x"02",x"01",x"00",x"1A",x"CD",x"7A",x"17",x"DD",x"36",x"1C",x"02",x"DD",x"7E",x"0B",x"FE",
		x"50",x"D2",x"78",x"16",x"3C",x"DD",x"77",x"0B",x"DD",x"7E",x"1D",x"FE",x"00",x"CA",x"8F",x"16",
		x"DD",x"36",x"0C",x"01",x"DD",x"36",x"0D",x"00",x"3D",x"DD",x"77",x"1D",x"C3",x"C9",x"16",x"DD",
		x"7E",x"1E",x"FE",x"00",x"CA",x"A6",x"16",x"DD",x"36",x"0C",x"01",x"DD",x"36",x"0D",x"01",x"3D",
		x"DD",x"77",x"1E",x"C3",x"C9",x"16",x"DD",x"7E",x"1F",x"FE",x"00",x"CA",x"BD",x"16",x"DD",x"36",
		x"0C",x"01",x"DD",x"36",x"0D",x"02",x"3D",x"DD",x"77",x"1F",x"C3",x"C9",x"16",x"DD",x"36",x"0C",
		x"00",x"DD",x"36",x"0D",x"00",x"DD",x"36",x"0B",x"FF",x"CD",x"B7",x"17",x"CD",x"FC",x"17",x"3A",
		x"20",x"80",x"FE",x"03",x"C2",x"EE",x"16",x"3E",x"12",x"CD",x"FD",x"1B",x"DD",x"36",x"0B",x"00",
		x"DD",x"36",x"1C",x"00",x"DD",x"7E",x"19",x"E6",x"0A",x"28",x"03",x"CD",x"73",x"17",x"DD",x"E1",
		x"E1",x"D1",x"C1",x"C9",x"3A",x"29",x"80",x"32",x"00",x"85",x"3A",x"2A",x"80",x"32",x"01",x"85",
		x"3A",x"2B",x"80",x"32",x"02",x"85",x"3A",x"2C",x"80",x"32",x"03",x"85",x"C9",x"3A",x"3B",x"80",
		x"CB",x"7F",x"28",x"0E",x"3A",x"3C",x"80",x"32",x"34",x"80",x"3A",x"3D",x"80",x"32",x"35",x"80",
		x"18",x"0A",x"CB",x"57",x"28",x"0C",x"3A",x"3E",x"80",x"32",x"35",x"80",x"CD",x"B7",x"17",x"CD",
		x"FC",x"17",x"C9",x"3A",x"3B",x"80",x"CB",x"77",x"28",x"08",x"3A",x"3D",x"80",x"32",x"34",x"80",
		x"18",x"0A",x"CB",x"4F",x"28",x"0C",x"3A",x"3D",x"80",x"32",x"35",x"80",x"CD",x"B7",x"17",x"CD",
		x"FC",x"17",x"C9",x"3A",x"3B",x"80",x"CB",x"6F",x"28",x"08",x"3A",x"3C",x"80",x"32",x"34",x"80",
		x"18",x"0A",x"CB",x"47",x"28",x"0C",x"3A",x"3C",x"80",x"32",x"35",x"80",x"CD",x"B7",x"17",x"CD",
		x"FC",x"17",x"C9",x"21",x"00",x"00",x"22",x"42",x"80",x"C9",x"E5",x"C5",x"3A",x"41",x"80",x"E6",
		x"0A",x"28",x"12",x"2A",x"42",x"80",x"09",x"CB",x"7C",x"28",x"03",x"21",x"FF",x"7F",x"22",x"42",
		x"80",x"DD",x"CB",x"00",x"C6",x"C1",x"E1",x"C9",x"E5",x"D5",x"21",x"00",x"00",x"3A",x"43",x"80",
		x"6F",x"CD",x"DD",x"17",x"65",x"DD",x"6E",x"1A",x"7C",x"B7",x"FE",x"08",x"30",x"03",x"21",x"00",
		x"00",x"22",x"42",x"80",x"D1",x"E1",x"C9",x"21",x"63",x"1E",x"DD",x"7E",x"0C",x"87",x"5F",x"16",
		x"00",x"19",x"5E",x"23",x"56",x"D5",x"FD",x"E1",x"DD",x"4E",x"0D",x"06",x"00",x"1E",x"07",x"16",
		x"00",x"79",x"B0",x"CA",x"DC",x"17",x"FD",x"19",x"0B",x"C3",x"D1",x"17",x"C9",x"D5",x"54",x"5D",
		x"B7",x"CB",x"15",x"CB",x"14",x"B7",x"CB",x"15",x"CB",x"14",x"19",x"B7",x"CB",x"1C",x"CB",x"1D",
		x"B7",x"CB",x"1C",x"CB",x"1D",x"B7",x"CB",x"1C",x"CB",x"1D",x"D1",x"C9",x"FD",x"7E",x"00",x"DD",
		x"77",x"01",x"FD",x"7E",x"01",x"DD",x"77",x"02",x"FD",x"7E",x"02",x"DD",x"77",x"12",x"FD",x"7E",
		x"03",x"DD",x"77",x"13",x"FD",x"7E",x"04",x"DD",x"77",x"14",x"FD",x"7E",x"05",x"DD",x"77",x"15",
		x"FD",x"7E",x"06",x"DD",x"77",x"16",x"C9",x"E5",x"D5",x"C5",x"DD",x"7E",x"19",x"CB",x"4F",x"CA",
		x"6C",x"18",x"DD",x"7E",x"01",x"B8",x"CA",x"6C",x"18",x"11",x"02",x"00",x"D2",x"42",x"18",x"11",
		x"FE",x"FF",x"D5",x"11",x"00",x"00",x"21",x"00",x"00",x"DD",x"6E",x"01",x"58",x"B7",x"ED",x"52",
		x"CD",x"C7",x"18",x"D1",x"7D",x"21",x"00",x"00",x"FE",x"01",x"28",x"06",x"38",x"04",x"19",x"3D",
		x"18",x"F6",x"11",x"00",x"00",x"DD",x"5E",x"04",x"19",x"DD",x"75",x"04",x"C1",x"D1",x"E1",x"C9",
		x"21",x"00",x"00",x"22",x"2F",x"80",x"3A",x"18",x"80",x"E6",x"03",x"FE",x"03",x"C2",x"89",x"18",
		x"2A",x"A2",x"1E",x"22",x"2F",x"80",x"C3",x"99",x"18",x"3A",x"1A",x"80",x"E6",x"03",x"FE",x"03",
		x"C2",x"99",x"18",x"2A",x"A6",x"1E",x"22",x"2F",x"80",x"C9",x"D5",x"E5",x"3A",x"3F",x"80",x"FE",
		x"00",x"C2",x"C4",x"18",x"2A",x"2F",x"80",x"DD",x"5E",x"05",x"DD",x"56",x"03",x"19",x"DD",x"75",
		x"05",x"DD",x"74",x"03",x"2A",x"31",x"80",x"DD",x"5E",x"06",x"DD",x"56",x"04",x"19",x"DD",x"75",
		x"06",x"DD",x"74",x"04",x"E1",x"D1",x"C9",x"D5",x"EB",x"B7",x"CB",x"7A",x"20",x"03",x"EB",x"18",
		x"06",x"21",x"00",x"00",x"B7",x"ED",x"52",x"D1",x"C9",x"D5",x"EB",x"21",x"00",x"00",x"B7",x"ED",
		x"52",x"D1",x"C9",x"E5",x"DD",x"E5",x"D5",x"21",x"00",x"00",x"22",x"5A",x"80",x"22",x"5C",x"80",
		x"DD",x"21",x"18",x"1C",x"2A",x"42",x"80",x"DD",x"56",x"01",x"DD",x"5E",x"00",x"B7",x"ED",x"52",
		x"CA",x"22",x"19",x"CB",x"7C",x"C2",x"22",x"19",x"DD",x"66",x"01",x"DD",x"6E",x"00",x"22",x"5C",
		x"80",x"DD",x"66",x"03",x"DD",x"6E",x"02",x"22",x"5A",x"80",x"11",x"04",x"00",x"DD",x"19",x"C3",
		x"F4",x"18",x"2A",x"42",x"80",x"ED",x"5B",x"5C",x"80",x"B7",x"ED",x"52",x"CA",x"4C",x"19",x"CB",
		x"7C",x"C2",x"4C",x"19",x"2A",x"5A",x"80",x"11",x"0A",x"00",x"19",x"22",x"5A",x"80",x"2A",x"5C",
		x"80",x"ED",x"5B",x"5A",x"80",x"19",x"22",x"5C",x"80",x"C3",x"22",x"19",x"D1",x"DD",x"E1",x"E1",
		x"C9",x"DD",x"E5",x"FD",x"E5",x"E5",x"D5",x"DD",x"21",x"6A",x"1C",x"3A",x"A1",x"81",x"87",x"11",
		x"00",x"00",x"5F",x"DD",x"19",x"DD",x"6E",x"00",x"DD",x"66",x"01",x"E5",x"DD",x"E1",x"FD",x"21",
		x"43",x"1E",x"3A",x"29",x"80",x"FE",x"19",x"20",x"06",x"FD",x"21",x"4D",x"1E",x"18",x"08",x"FE",
		x"1A",x"20",x"04",x"FD",x"21",x"57",x"1E",x"DD",x"7E",x"00",x"FE",x"FF",x"CA",x"C7",x"1A",x"21",
		x"00",x"00",x"11",x"00",x"00",x"DD",x"6E",x"00",x"FD",x"46",x"03",x"FD",x"4E",x"02",x"09",x"3A",
		x"2B",x"80",x"5F",x"B7",x"ED",x"52",x"CA",x"BF",x"1A",x"D2",x"BF",x"1A",x"CD",x"C7",x"18",x"22",
		x"5E",x"80",x"21",x"00",x"00",x"DD",x"6E",x"01",x"FD",x"46",x"05",x"FD",x"4E",x"04",x"09",x"B7",
		x"ED",x"52",x"CA",x"BF",x"1A",x"DA",x"BF",x"1A",x"22",x"60",x"80",x"21",x"00",x"00",x"DD",x"6E",
		x"02",x"FD",x"46",x"07",x"FD",x"4E",x"06",x"09",x"11",x"00",x"00",x"3A",x"2C",x"80",x"5F",x"B7",
		x"ED",x"52",x"CA",x"BF",x"1A",x"D2",x"BF",x"1A",x"CD",x"C7",x"18",x"22",x"62",x"80",x"21",x"00",
		x"00",x"DD",x"6E",x"03",x"FD",x"46",x"09",x"FD",x"4E",x"08",x"09",x"B7",x"ED",x"52",x"CA",x"BF",
		x"1A",x"DA",x"BF",x"1A",x"22",x"64",x"80",x"2A",x"5E",x"80",x"ED",x"5B",x"60",x"80",x"44",x"4D",
		x"B7",x"ED",x"52",x"38",x"0A",x"42",x"4B",x"21",x"00",x"00",x"22",x"5E",x"80",x"18",x"06",x"21",
		x"00",x"00",x"22",x"60",x"80",x"2A",x"62",x"80",x"ED",x"5B",x"64",x"80",x"B7",x"ED",x"52",x"38",
		x"08",x"21",x"00",x"00",x"22",x"62",x"80",x"18",x"0A",x"ED",x"5B",x"62",x"80",x"21",x"00",x"00",
		x"22",x"64",x"80",x"60",x"69",x"B7",x"ED",x"52",x"38",x"0B",x"21",x"00",x"00",x"22",x"5E",x"80",
		x"22",x"60",x"80",x"18",x"09",x"21",x"00",x"00",x"22",x"62",x"80",x"22",x"64",x"80",x"2A",x"5E",
		x"80",x"7C",x"B5",x"28",x"13",x"21",x"00",x"00",x"DD",x"6E",x"00",x"FD",x"56",x"03",x"FD",x"5E",
		x"02",x"19",x"7D",x"32",x"2B",x"80",x"18",x"5E",x"2A",x"60",x"80",x"7C",x"B5",x"28",x"13",x"21",
		x"00",x"00",x"DD",x"6E",x"01",x"FD",x"56",x"05",x"FD",x"5E",x"04",x"19",x"7D",x"32",x"2B",x"80",
		x"18",x"44",x"2A",x"62",x"80",x"7C",x"B5",x"28",x"13",x"21",x"00",x"00",x"DD",x"6E",x"02",x"FD",
		x"56",x"07",x"FD",x"5E",x"06",x"19",x"7D",x"32",x"2C",x"80",x"18",x"2A",x"21",x"00",x"00",x"DD",
		x"6E",x"03",x"FD",x"56",x"09",x"FD",x"5E",x"08",x"19",x"7D",x"32",x"2C",x"80",x"18",x"17",x"11",
		x"04",x"00",x"DD",x"19",x"C3",x"87",x"19",x"DD",x"7E",x"01",x"FE",x"FF",x"CA",x"D6",x"1A",x"DD",
		x"21",x"31",x"1E",x"C3",x"87",x"19",x"D1",x"E1",x"FD",x"E1",x"DD",x"E1",x"C9",x"C5",x"D5",x"11",
		x"00",x"00",x"3A",x"02",x"85",x"C6",x"04",x"47",x"3A",x"03",x"85",x"C6",x"00",x"4F",x"CD",x"DE",
		x"00",x"7E",x"CD",x"AF",x"1B",x"FE",x"00",x"28",x"02",x"CB",x"CB",x"3A",x"02",x"85",x"C6",x"0C",
		x"47",x"3A",x"03",x"85",x"C6",x"00",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",x"AF",x"1B",x"FE",x"00",
		x"28",x"02",x"CB",x"CB",x"3A",x"02",x"85",x"C6",x"04",x"47",x"3A",x"03",x"85",x"C6",x"0F",x"4F",
		x"CD",x"DE",x"00",x"7E",x"CD",x"AF",x"1B",x"FE",x"00",x"28",x"02",x"CB",x"DB",x"3A",x"02",x"85",
		x"C6",x"0C",x"47",x"3A",x"03",x"85",x"C6",x"0F",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",x"AF",x"1B",
		x"FE",x"00",x"28",x"02",x"CB",x"DB",x"3A",x"02",x"85",x"C6",x"02",x"47",x"3A",x"03",x"85",x"C6",
		x"04",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",x"D8",x"1B",x"FE",x"00",x"28",x"02",x"CB",x"C3",x"3A",
		x"02",x"85",x"C6",x"02",x"47",x"3A",x"03",x"85",x"C6",x"0C",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",
		x"D8",x"1B",x"FE",x"00",x"28",x"02",x"CB",x"C3",x"3A",x"02",x"85",x"C6",x"0D",x"47",x"3A",x"03",
		x"85",x"C6",x"04",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",x"D8",x"1B",x"FE",x"00",x"28",x"02",x"CB",
		x"C3",x"3A",x"02",x"85",x"C6",x"0D",x"47",x"3A",x"03",x"85",x"C6",x"0C",x"4F",x"CD",x"DE",x"00",
		x"7E",x"CD",x"D8",x"1B",x"FE",x"00",x"28",x"02",x"CB",x"C3",x"62",x"6B",x"D1",x"C1",x"C9",x"FE",
		x"60",x"38",x"22",x"FE",x"80",x"38",x"08",x"FE",x"A0",x"38",x"1A",x"FE",x"C0",x"30",x"16",x"E6",
		x"0F",x"FE",x"06",x"38",x"0C",x"FE",x"08",x"38",x"0C",x"FE",x"0C",x"38",x"04",x"FE",x"0E",x"38",
		x"04",x"3E",x"01",x"18",x"02",x"3E",x"00",x"C9",x"FE",x"60",x"38",x"1E",x"FE",x"80",x"38",x"08",
		x"FE",x"A0",x"38",x"16",x"FE",x"C0",x"30",x"12",x"E6",x"0F",x"FE",x"02",x"38",x"08",x"FE",x"04",
		x"38",x"08",x"FE",x"0E",x"30",x"04",x"3E",x"01",x"18",x"02",x"3E",x"00",x"C9",x"C5",x"FE",x"13",
		x"28",x"06",x"FE",x"93",x"28",x"02",x"18",x"08",x"47",x"3A",x"89",x"80",x"B8",x"28",x"07",x"78",
		x"32",x"89",x"80",x"CD",x"FC",x"00",x"C1",x"C9",x"96",x"00",x"32",x"00",x"C2",x"01",x"5A",x"00",
		x"8E",x"03",x"82",x"00",x"FA",x"05",x"AA",x"00",x"06",x"09",x"D2",x"00",x"B2",x"0C",x"FA",x"00",
		x"FE",x"10",x"22",x"01",x"EA",x"15",x"4A",x"01",x"76",x"1B",x"72",x"01",x"A2",x"21",x"9A",x"01",
		x"6E",x"28",x"C2",x"01",x"DA",x"2F",x"EA",x"01",x"E6",x"37",x"12",x"02",x"92",x"40",x"3A",x"02",
		x"DE",x"49",x"62",x"02",x"CA",x"53",x"8A",x"02",x"56",x"5E",x"B2",x"02",x"82",x"69",x"DA",x"02",
		x"4E",x"75",x"02",x"03",x"BA",x"81",x"2A",x"03",x"FF",x"FF",x"8C",x"1C",x"A1",x"1C",x"B2",x"1C",
		x"C7",x"1C",x"E9",x"1C",x"EA",x"1C",x"13",x"1D",x"2C",x"1D",x"3D",x"1D",x"52",x"1D",x"63",x"1D",
		x"94",x"1D",x"AD",x"1D",x"C6",x"1D",x"E7",x"1D",x"00",x"1E",x"FF",x"FF",x"7B",x"BD",x"31",x"46",
		x"33",x"5D",x"49",x"5E",x"63",x"9D",x"91",x"A6",x"1B",x"45",x"A9",x"BE",x"83",x"D5",x"C1",x"D6",
		x"FF",x"53",x"9D",x"31",x"46",x"33",x"45",x"51",x"9E",x"AB",x"BD",x"51",x"9E",x"53",x"9D",x"A9",
		x"BE",x"FF",x"6B",x"9D",x"31",x"46",x"0B",x"55",x"49",x"5E",x"9B",x"CD",x"61",x"76",x"93",x"A5",
		x"61",x"A6",x"33",x"A5",x"91",x"A6",x"FF",x"4B",x"5D",x"21",x"5E",x"93",x"A5",x"21",x"5E",x"23",
		x"5D",x"49",x"5E",x"93",x"CD",x"49",x"5E",x"23",x"55",x"91",x"A6",x"9B",x"CD",x"91",x"A6",x"4B",
		x"5D",x"91",x"CE",x"93",x"A5",x"91",x"CE",x"FF",x"00",x"FF",x"1B",x"45",x"31",x"46",x"63",x"8D",
		x"31",x"46",x"AB",x"D5",x"31",x"46",x"3B",x"6D",x"61",x"76",x"83",x"B5",x"61",x"76",x"1B",x"45",
		x"91",x"A6",x"63",x"8D",x"91",x"A6",x"AB",x"D5",x"91",x"A6",x"3B",x"6D",x"C1",x"D6",x"83",x"B5",
		x"C1",x"D6",x"FF",x"63",x"8D",x"31",x"46",x"33",x"6D",x"61",x"76",x"83",x"BD",x"61",x"76",x"33",
		x"6D",x"79",x"8E",x"83",x"BD",x"79",x"8E",x"63",x"8D",x"A9",x"BE",x"FF",x"23",x"55",x"31",x"46",
		x"9B",x"CD",x"31",x"46",x"23",x"55",x"A9",x"BE",x"9B",x"CD",x"A9",x"BE",x"FF",x"3B",x"6D",x"31",
		x"46",x"83",x"B5",x"31",x"46",x"63",x"8D",x"91",x"A6",x"1B",x"45",x"A9",x"BE",x"AB",x"D5",x"A9",
		x"BE",x"FF",x"3B",x"B5",x"31",x"46",x"33",x"45",x"31",x"9E",x"AB",x"BD",x"31",x"9E",x"63",x"8D",
		x"91",x"A6",x"FF",x"6B",x"85",x"19",x"2E",x"63",x"75",x"19",x"46",x"63",x"8D",x"31",x"46",x"4B",
		x"8D",x"49",x"5E",x"63",x"75",x"49",x"76",x"63",x"8D",x"61",x"76",x"6B",x"BD",x"79",x"8E",x"63",
		x"75",x"79",x"A6",x"63",x"8D",x"91",x"A6",x"1B",x"8D",x"A9",x"BE",x"63",x"75",x"B1",x"D6",x"63",
		x"8D",x"C1",x"D6",x"FF",x"0B",x"3D",x"49",x"5E",x"B3",x"E5",x"49",x"5E",x"23",x"55",x"79",x"8E",
		x"9B",x"CD",x"79",x"8E",x"3B",x"6D",x"A9",x"BE",x"83",x"B5",x"A9",x"BE",x"FF",x"3B",x"85",x"31",
		x"46",x"93",x"B5",x"31",x"46",x"33",x"45",x"31",x"BE",x"AB",x"BD",x"31",x"BE",x"33",x"5D",x"A9",
		x"BE",x"6B",x"BD",x"A9",x"BE",x"FF",x"33",x"85",x"19",x"2E",x"7B",x"8D",x"19",x"5E",x"23",x"5D",
		x"61",x"76",x"1B",x"2D",x"61",x"BE",x"C3",x"D5",x"31",x"8E",x"93",x"D5",x"79",x"8E",x"63",x"75",
		x"91",x"D6",x"63",x"BD",x"C1",x"D6",x"FF",x"B3",x"E5",x"31",x"46",x"0B",x"3D",x"49",x"5E",x"B3",
		x"E5",x"61",x"76",x"0B",x"3D",x"79",x"8E",x"B3",x"E5",x"91",x"A6",x"0B",x"3D",x"A9",x"BE",x"FF",
		x"3B",x"6D",x"19",x"2E",x"83",x"B5",x"19",x"2E",x"1B",x"2D",x"39",x"6E",x"C3",x"D5",x"39",x"6E",
		x"1B",x"2D",x"81",x"B6",x"C3",x"D5",x"81",x"B6",x"63",x"8D",x"49",x"5E",x"4B",x"5D",x"61",x"8E",
		x"93",x"A5",x"61",x"8E",x"63",x"8D",x"91",x"A6",x"3B",x"6D",x"C1",x"D6",x"83",x"B5",x"C1",x"D6",
		x"FF",x"04",x"FD",x"04",x"16",x"04",x"15",x"04",x"FE",x"DB",x"FD",x"04",x"FE",x"04",x"FD",x"D9",
		x"FE",x"FF",x"FF",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"19",x"00",x"FF",
		x"FF",x"01",x"00",x"00",x"00",x"FF",x"FF",x"1A",x"00",x"FF",x"FF",x"01",x"00",x"00",x"00",x"FF",
		x"FF",x"FF",x"FF",x"67",x"1E",x"6A",x"1E",x"18",x"00",x"FF",x"1A",x"00",x"20",x"04",x"FF",x"FF",
		x"00",x"19",x"00",x"28",x"04",x"FF",x"FF",x"00",x"18",x"00",x"04",x"04",x"FF",x"FF",x"00",x"18",
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"10",x"00",x"08",x"00",x"F0",x"FF",x"F8",x"FF",x"80",x"01",
		x"FF",x"FF",x"08",x"00",x"10",x"00",x"20",x"00",x"30",x"00",x"01",x"00",x"FF",x"FF",x"02",x"00",
		x"FE",x"FF",x"80",x"01",x"00",x"00",x"80",x"FE",x"00",x"00",x"D9",x"00",x"D8",x"00",x"D7",x"00",
		x"D6",x"00",x"33",x"00",x"34",x"00",x"35",x"00",x"D5",x"FF",x"C0",x"FF",x"00",x"FF",x"90",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CD",x"9F",x"02",x"3A",x"03",x"B0",x"C3",x"CB",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"27",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"5C",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"A4",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"1F",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"4C",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"60",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"32",x"03",x"B0",x"DD",x"36",x"00",x"30",x"C3",x"F8",x"05",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"72",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"8B",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"C3",x"98",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"11",x"08",x"00",x"C3",x"FC",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CD",x"D2",x"00",x"3A",x"03",x"B0",x"C3",x"F9",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C3",x"C7",x"18",x"C3",x"D9",x"18",x"00",x"3A",x"03",x"B0",x"CD",x"02",x"06",x"C3",x"AB",x"05",
		x"CD",x"05",x"22",x"3A",x"8D",x"80",x"FE",x"00",x"20",x"0A",x"3A",x"28",x"80",x"CB",x"57",x"20",
		x"03",x"CD",x"C0",x"20",x"3A",x"53",x"84",x"E6",x"03",x"FE",x"03",x"28",x"17",x"3A",x"A7",x"81",
		x"B7",x"FE",x"14",x"38",x"15",x"3E",x"00",x"32",x"A7",x"81",x"3E",x"03",x"32",x"53",x"84",x"3E",
		x"1B",x"CD",x"FC",x"00",x"CD",x"4B",x"23",x"CD",x"C9",x"00",x"3A",x"00",x"89",x"CB",x"47",x"28",
		x"06",x"CD",x"33",x"25",x"CD",x"C9",x"00",x"3A",x"60",x"84",x"FE",x"00",x"28",x"17",x"3D",x"32",
		x"60",x"84",x"FE",x"00",x"20",x"0F",x"21",x"00",x"00",x"22",x"08",x"85",x"22",x"0A",x"85",x"22",
		x"0C",x"85",x"22",x"0E",x"85",x"3A",x"02",x"89",x"FE",x"FF",x"28",x"16",x"3A",x"13",x"89",x"FE",
		x"00",x"28",x"3C",x"3D",x"32",x"13",x"89",x"FE",x"00",x"20",x"34",x"3A",x"0C",x"89",x"FE",x"02",
		x"20",x"0A",x"CD",x"36",x"60",x"3A",x"02",x"89",x"FE",x"FF",x"28",x"23",x"21",x"00",x"00",x"22",
		x"10",x"85",x"22",x"12",x"85",x"22",x"14",x"85",x"22",x"16",x"85",x"3A",x"0C",x"89",x"FE",x"03",
		x"20",x"08",x"3E",x"01",x"32",x"80",x"80",x"32",x"77",x"80",x"3E",x"00",x"32",x"0C",x"89",x"3A",
		x"8D",x"80",x"FE",x"00",x"CA",x"C3",x"00",x"3A",x"28",x"80",x"CB",x"57",x"C2",x"C3",x"00",x"C9",
		x"3A",x"28",x"80",x"CB",x"57",x"C2",x"75",x"21",x"DD",x"21",x"A2",x"81",x"FD",x"21",x"80",x"84",
		x"3A",x"A2",x"81",x"FE",x"00",x"CA",x"5D",x"21",x"FD",x"CB",x"00",x"76",x"C2",x"4B",x"21",x"3A",
		x"02",x"85",x"16",x"00",x"5F",x"21",x"08",x"00",x"19",x"54",x"5D",x"26",x"00",x"FD",x"6E",x"01",
		x"01",x"08",x"00",x"09",x"B7",x"ED",x"52",x"CD",x"F0",x"1F",x"11",x"0A",x"00",x"B7",x"ED",x"52",
		x"D2",x"4B",x"21",x"3A",x"03",x"85",x"16",x"00",x"5F",x"21",x"08",x"00",x"19",x"54",x"5D",x"26",
		x"00",x"FD",x"6E",x"02",x"01",x"08",x"00",x"09",x"B7",x"ED",x"52",x"CD",x"F0",x"1F",x"11",x"08",
		x"00",x"B7",x"ED",x"52",x"D2",x"4B",x"21",x"CD",x"76",x"21",x"3A",x"53",x"84",x"E6",x"03",x"FE",
		x"03",x"28",x"0A",x"3A",x"28",x"80",x"CB",x"7F",x"20",x"03",x"CD",x"06",x"29",x"CD",x"CF",x"22",
		x"3A",x"A2",x"81",x"FE",x"00",x"CA",x"5D",x"21",x"C3",x"75",x"21",x"FD",x"7E",x"00",x"E6",x"3F",
		x"FE",x"17",x"CA",x"75",x"21",x"11",x"05",x"00",x"FD",x"19",x"C3",x"D8",x"20",x"3A",x"70",x"80",
		x"FE",x"00",x"28",x"0A",x"3E",x"01",x"32",x"74",x"80",x"32",x"77",x"80",x"18",x"07",x"3E",x"01",
		x"32",x"78",x"80",x"18",x"00",x"C9",x"C5",x"DD",x"E5",x"FD",x"E5",x"FD",x"36",x"04",x"00",x"01",
		x"00",x"01",x"3E",x"19",x"FD",x"CB",x"00",x"7E",x"28",x"10",x"01",x"00",x"02",x"3A",x"AB",x"81",
		x"3C",x"32",x"AB",x"81",x"FD",x"36",x"04",x"01",x"3E",x"18",x"CD",x"FC",x"00",x"CD",x"E4",x"00",
		x"FD",x"46",x"01",x"FD",x"4E",x"02",x"CD",x"DE",x"00",x"E5",x"DD",x"E1",x"DD",x"36",x"00",x"86",
		x"DD",x"36",x"01",x"87",x"11",x"E0",x"FF",x"DD",x"19",x"DD",x"36",x"00",x"84",x"DD",x"36",x"01",
		x"85",x"FD",x"CB",x"00",x"F6",x"FD",x"36",x"03",x"01",x"3A",x"A2",x"81",x"FE",x"00",x"28",x"01",
		x"3D",x"32",x"A2",x"81",x"3A",x"A7",x"81",x"3C",x"FD",x"CB",x"00",x"7E",x"28",x"0C",x"3C",x"4F",
		x"FD",x"CB",x"00",x"BE",x"3E",x"00",x"32",x"A6",x"81",x"79",x"4F",x"3A",x"53",x"84",x"E6",x"03",
		x"FE",x"03",x"28",x"0B",x"3A",x"28",x"80",x"CB",x"7F",x"20",x"04",x"79",x"32",x"A7",x"81",x"FD",
		x"E1",x"DD",x"E1",x"C1",x"C9",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"DD",x"21",x"80",x"84",
		x"DD",x"7E",x"00",x"FE",x"FF",x"CA",x"C7",x"22",x"DD",x"CB",x"00",x"76",x"CA",x"BC",x"22",x"DD",
		x"7E",x"03",x"FE",x"00",x"CA",x"BC",x"22",x"DD",x"7E",x"03",x"3C",x"DD",x"77",x"03",x"FE",x"05",
		x"C2",x"57",x"22",x"DD",x"46",x"01",x"DD",x"4E",x"02",x"CD",x"DE",x"00",x"E5",x"FD",x"E1",x"FD",
		x"36",x"00",x"8A",x"FD",x"36",x"01",x"8B",x"11",x"E0",x"FF",x"FD",x"19",x"FD",x"36",x"00",x"88",
		x"FD",x"36",x"01",x"89",x"C3",x"BC",x"22",x"FE",x"09",x"C2",x"80",x"22",x"DD",x"46",x"01",x"DD",
		x"4E",x"02",x"CD",x"DE",x"00",x"E5",x"FD",x"E1",x"FD",x"36",x"00",x"8E",x"FD",x"36",x"01",x"8F",
		x"11",x"E0",x"FF",x"FD",x"19",x"FD",x"36",x"00",x"8C",x"FD",x"36",x"01",x"8D",x"C3",x"BC",x"22",
		x"FE",x"0D",x"DA",x"BC",x"22",x"DD",x"46",x"01",x"DD",x"4E",x"02",x"CD",x"DE",x"00",x"E5",x"FD",
		x"E1",x"FD",x"36",x"00",x"00",x"FD",x"36",x"01",x"00",x"11",x"E0",x"FF",x"FD",x"19",x"FD",x"36",
		x"00",x"00",x"FD",x"36",x"01",x"00",x"11",x"00",x"04",x"19",x"36",x"0A",x"23",x"36",x"0A",x"11",
		x"E0",x"FF",x"19",x"36",x"0A",x"2B",x"36",x"0A",x"DD",x"36",x"03",x"00",x"CD",x"2D",x"60",x"11",
		x"05",x"00",x"DD",x"19",x"C3",x"10",x"22",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",x"C5",
		x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"3A",x"A2",x"81",x"FE",x"00",x"CA",x"43",x"23",x"3A",x"A6",
		x"81",x"FE",x"01",x"CA",x"43",x"23",x"3E",x"01",x"32",x"A6",x"81",x"FD",x"7E",x"00",x"FE",x"FF",
		x"20",x"04",x"FD",x"21",x"80",x"84",x"FD",x"CB",x"00",x"76",x"28",x"07",x"11",x"05",x"00",x"FD",
		x"19",x"18",x"E8",x"FD",x"CB",x"00",x"FE",x"FD",x"46",x"01",x"FD",x"4E",x"02",x"CD",x"DE",x"00",
		x"E5",x"DD",x"E1",x"11",x"00",x"04",x"19",x"3A",x"A4",x"85",x"47",x"70",x"3A",x"A2",x"85",x"DD",
		x"77",x"00",x"23",x"DD",x"23",x"70",x"3A",x"A3",x"85",x"DD",x"77",x"00",x"11",x"DF",x"FF",x"19",
		x"DD",x"19",x"70",x"3A",x"A0",x"85",x"DD",x"77",x"00",x"23",x"DD",x"23",x"70",x"3A",x"A1",x"85",
		x"DD",x"77",x"00",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",x"3A",x"28",x"80",x"CB",x"57",
		x"C0",x"3A",x"8E",x"80",x"FE",x"00",x"C0",x"DD",x"21",x"53",x"84",x"3A",x"53",x"84",x"E6",x"03",
		x"FE",x"03",x"C2",x"46",x"24",x"DD",x"CB",x"00",x"56",x"20",x"2D",x"21",x"00",x"00",x"22",x"0C",
		x"85",x"22",x"0E",x"85",x"DD",x"CB",x"00",x"D6",x"DD",x"36",x"02",x"3D",x"DD",x"36",x"03",x"0E",
		x"DD",x"36",x"04",x"78",x"DD",x"36",x"05",x"78",x"DD",x"36",x"0C",x"01",x"DD",x"36",x"0D",x"00",
		x"3E",x"00",x"32",x"58",x"88",x"CD",x"A9",x"24",x"CD",x"47",x"24",x"FE",x"00",x"C2",x"01",x"24",
		x"DD",x"46",x"04",x"DD",x"4E",x"05",x"DD",x"36",x"01",x"00",x"FD",x"E5",x"FD",x"21",x"08",x"85",
		x"CD",x"F2",x"5F",x"FD",x"E1",x"FE",x"00",x"CA",x"DB",x"23",x"4F",x"E6",x"0C",x"28",x"09",x"2A",
		x"5D",x"84",x"CD",x"F3",x"1F",x"22",x"5D",x"84",x"3E",x"1C",x"CD",x"FC",x"00",x"79",x"E6",x"03",
		x"28",x"09",x"2A",x"5B",x"84",x"CD",x"F3",x"1F",x"22",x"5B",x"84",x"3A",x"53",x"84",x"E6",x"C0",
		x"FE",x"C0",x"20",x"1A",x"DD",x"CB",x"00",x"BE",x"DD",x"CB",x"00",x"B6",x"3A",x"5F",x"84",x"3C",
		x"FE",x"07",x"28",x"04",x"38",x"02",x"3E",x"01",x"32",x"5F",x"84",x"CD",x"A9",x"24",x"C3",x"38",
		x"24",x"3E",x"1A",x"CD",x"FC",x"00",x"3A",x"28",x"80",x"CB",x"FF",x"32",x"28",x"80",x"21",x"2C",
		x"01",x"22",x"36",x"80",x"21",x"00",x"00",x"22",x"53",x"84",x"22",x"55",x"84",x"CD",x"10",x"25",
		x"DD",x"66",x"0C",x"DD",x"36",x"0C",x"00",x"7C",x"21",x"00",x"00",x"FD",x"21",x"08",x"85",x"CD",
		x"F3",x"00",x"DD",x"36",x"0D",x"1E",x"18",x"03",x"CD",x"F3",x"2C",x"DD",x"21",x"54",x"84",x"FD",
		x"21",x"08",x"85",x"CD",x"24",x"2D",x"C9",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"3A",x"8D",
		x"80",x"FE",x"00",x"20",x"4A",x"3A",x"28",x"80",x"CB",x"57",x"20",x"43",x"11",x"00",x"00",x"3A",
		x"02",x"85",x"5F",x"21",x"08",x"00",x"19",x"EB",x"01",x"00",x"00",x"DD",x"4E",x"04",x"21",x"08",
		x"00",x"09",x"ED",x"52",x"CD",x"F0",x"1F",x"7D",x"FE",x"0A",x"D2",x"9F",x"24",x"11",x"00",x"00",
		x"3A",x"03",x"85",x"5F",x"21",x"0A",x"00",x"19",x"EB",x"01",x"00",x"00",x"DD",x"4E",x"05",x"21",
		x"08",x"00",x"09",x"ED",x"52",x"CD",x"F0",x"1F",x"7D",x"FE",x"0A",x"28",x"04",x"38",x"02",x"3E",
		x"00",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",
		x"FD",x"21",x"00",x"88",x"11",x"0A",x"00",x"FD",x"7E",x"00",x"E6",x"7F",x"FE",x"0E",x"28",x"04",
		x"FD",x"19",x"18",x"F3",x"21",x"48",x"0D",x"3A",x"5F",x"84",x"FE",x"00",x"28",x"0F",x"3D",x"21",
		x"9E",x"0D",x"11",x"12",x"00",x"FE",x"00",x"28",x"04",x"19",x"3D",x"18",x"F8",x"FD",x"75",x"01",
		x"FD",x"74",x"02",x"E5",x"DD",x"E1",x"06",x"07",x"FD",x"21",x"E2",x"8C",x"78",x"FE",x"00",x"28",
		x"17",x"DD",x"7E",x"00",x"FD",x"77",x"00",x"DD",x"7E",x"01",x"FD",x"77",x"01",x"DD",x"23",x"DD",
		x"23",x"FD",x"23",x"FD",x"23",x"05",x"18",x"E4",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",
		x"C5",x"FD",x"E5",x"3A",x"5F",x"84",x"3D",x"FD",x"21",x"7E",x"2F",x"FE",x"00",x"28",x"07",x"FD",
		x"23",x"FD",x"23",x"3D",x"18",x"F5",x"FD",x"46",x"01",x"FD",x"4E",x"00",x"CD",x"E4",x"00",x"FD",
		x"E1",x"C1",x"C9",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"DD",x"21",x"00",x"89",x"DD",x"CB",
		x"00",x"4E",x"20",x"06",x"CD",x"27",x"27",x"CD",x"00",x"28",x"DD",x"7E",x"11",x"FE",x"00",x"C2",
		x"95",x"26",x"DD",x"CB",x"00",x"7E",x"C2",x"E6",x"26",x"DD",x"CB",x"00",x"56",x"C2",x"9E",x"25",
		x"CD",x"C4",x"27",x"FE",x"00",x"C2",x"33",x"26",x"DD",x"36",x"03",x"0C",x"DD",x"36",x"0D",x"FF",
		x"DD",x"36",x"0E",x"03",x"DD",x"36",x"0F",x"00",x"DD",x"CB",x"00",x"D6",x"DD",x"36",x"07",x"00",
		x"DD",x"36",x"0A",x"00",x"DD",x"36",x"0B",x"00",x"21",x"AA",x"00",x"22",x"08",x"89",x"3A",x"2B",
		x"80",x"CB",x"47",x"28",x"06",x"21",x"56",x"FF",x"22",x"08",x"89",x"C3",x"1F",x"27",x"DD",x"46",
		x"04",x"DD",x"4E",x"05",x"DD",x"36",x"01",x"01",x"FD",x"E5",x"FD",x"21",x"10",x"85",x"CD",x"F2",
		x"5F",x"FD",x"E1",x"47",x"DD",x"4E",x"10",x"DD",x"36",x"10",x"00",x"E6",x"03",x"FE",x"00",x"28",
		x"01",x"0C",x"78",x"2A",x"0A",x"89",x"11",x"0A",x"00",x"19",x"22",x"0A",x"89",x"CB",x"57",x"CA",
		x"2B",x"26",x"ED",x"5B",x"0A",x"89",x"21",x"00",x"00",x"DD",x"71",x"10",x"22",x"0A",x"89",x"7B",
		x"FE",x"46",x"38",x"11",x"3E",x"1D",x"CD",x"FC",x"00",x"DD",x"36",x"0D",x"10",x"DD",x"36",x"0E",
		x"01",x"DD",x"36",x"0F",x"00",x"3A",x"0D",x"89",x"FE",x"FF",x"28",x"0C",x"FE",x"00",x"20",x"08",
		x"DD",x"36",x"0D",x"FF",x"DD",x"36",x"0E",x"03",x"78",x"E6",x"03",x"FE",x"00",x"28",x"24",x"3E",
		x"1D",x"CD",x"FC",x"00",x"2A",x"08",x"89",x"CD",x"F3",x"1F",x"22",x"08",x"89",x"DD",x"36",x"0D",
		x"10",x"DD",x"36",x"0E",x"01",x"DD",x"36",x"0F",x"00",x"18",x"08",x"DD",x"36",x"0D",x"FF",x"DD",
		x"36",x"0E",x"03",x"3A",x"10",x"89",x"FE",x"03",x"D2",x"C9",x"26",x"DD",x"46",x"04",x"DD",x"4E",
		x"05",x"CD",x"47",x"24",x"FE",x"00",x"CA",x"19",x"27",x"3A",x"0C",x"89",x"FE",x"02",x"20",x"05",
		x"3E",x"01",x"32",x"88",x"80",x"3A",x"0C",x"89",x"FE",x"03",x"3E",x"1E",x"20",x"0C",x"3E",x"01",
		x"CD",x"FC",x"00",x"3E",x"01",x"32",x"8E",x"80",x"3E",x"28",x"CD",x"FC",x"00",x"DD",x"36",x"11",
		x"10",x"DD",x"36",x"02",x"AD",x"DD",x"36",x"03",x"2B",x"3A",x"04",x"89",x"D6",x"08",x"32",x"04",
		x"89",x"3A",x"05",x"89",x"D6",x"08",x"32",x"05",x"89",x"21",x"00",x"00",x"22",x"08",x"89",x"22",
		x"0A",x"89",x"C3",x"1C",x"27",x"DD",x"35",x"11",x"DD",x"7E",x"11",x"FE",x"00",x"20",x"7D",x"3A",
		x"04",x"89",x"C6",x"08",x"32",x"04",x"89",x"3A",x"05",x"89",x"C6",x"08",x"32",x"05",x"89",x"DD",
		x"36",x"13",x"1E",x"3A",x"0C",x"89",x"3D",x"FD",x"21",x"10",x"85",x"21",x"01",x"00",x"CD",x"F3",
		x"00",x"CD",x"89",x"28",x"CD",x"FC",x"28",x"18",x"53",x"DD",x"CB",x"00",x"FE",x"DD",x"36",x"12",
		x"05",x"DD",x"36",x"0D",x"05",x"DD",x"36",x"0E",x"05",x"DD",x"36",x"0F",x"00",x"21",x"00",x"00",
		x"22",x"08",x"89",x"22",x"0A",x"89",x"DD",x"46",x"04",x"DD",x"4E",x"05",x"CD",x"47",x"24",x"FE",
		x"00",x"C2",x"49",x"26",x"CD",x"C4",x"27",x"FE",x"00",x"20",x"21",x"3A",x"12",x"89",x"FE",x"10",
		x"30",x"12",x"DD",x"34",x"12",x"3A",x"12",x"89",x"32",x"0D",x"89",x"32",x"0E",x"89",x"DD",x"36",
		x"0F",x"00",x"18",x"08",x"CD",x"A7",x"28",x"18",x"03",x"CD",x"C4",x"27",x"CD",x"3C",x"28",x"FD",
		x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"C9",x"E5",x"21",x"00",x"00",x"22",x"14",x"85",x"22",x"16",
		x"85",x"DD",x"CB",x"00",x"C6",x"DD",x"CB",x"00",x"CE",x"DD",x"36",x"03",x"1C",x"21",x"00",x"00",
		x"22",x"06",x"89",x"22",x"0A",x"89",x"21",x"80",x"FF",x"22",x"0A",x"89",x"DD",x"36",x"0D",x"20",
		x"DD",x"36",x"0E",x"01",x"DD",x"36",x"0F",x"00",x"DD",x"36",x"10",x"00",x"DD",x"36",x"11",x"00",
		x"DD",x"36",x"12",x"00",x"DD",x"36",x"13",x"00",x"CD",x"C9",x"00",x"3A",x"25",x"80",x"FE",x"AA",
		x"20",x"1F",x"3A",x"70",x"80",x"FE",x"00",x"28",x"18",x"3A",x"14",x"80",x"CB",x"7F",x"28",x"07",
		x"3A",x"24",x"80",x"CB",x"67",x"28",x"0A",x"DD",x"36",x"02",x"14",x"DD",x"36",x"0C",x"03",x"18",
		x"2E",x"3A",x"14",x"80",x"CB",x"7F",x"28",x"09",x"3A",x"B3",x"81",x"FE",x"3C",x"38",x"18",x"18",
		x"07",x"3A",x"B3",x"81",x"FE",x"28",x"38",x"0F",x"3E",x"00",x"32",x"B3",x"81",x"DD",x"36",x"02",
		x"10",x"DD",x"36",x"0C",x"02",x"18",x"08",x"DD",x"36",x"02",x"0C",x"DD",x"36",x"0C",x"01",x"CD",
		x"F0",x"3F",x"E1",x"C9",x"E5",x"3A",x"0D",x"89",x"FE",x"FF",x"28",x"08",x"FE",x"00",x"CA",x"FE",
		x"27",x"DD",x"35",x"0D",x"DD",x"34",x"0F",x"3A",x"0E",x"89",x"DD",x"BE",x"0F",x"28",x"03",x"D2",
		x"FC",x"27",x"3A",x"02",x"89",x"E6",x"03",x"FE",x"03",x"20",x"0A",x"DD",x"CB",x"02",x"86",x"DD",
		x"CB",x"02",x"8E",x"18",x"03",x"DD",x"34",x"02",x"DD",x"36",x"0F",x"00",x"3E",x"01",x"E1",x"C9",
		x"D5",x"E5",x"FD",x"E5",x"FD",x"21",x"00",x"88",x"11",x"0A",x"00",x"FD",x"7E",x"00",x"E6",x"7F",
		x"FE",x"0C",x"28",x"04",x"FD",x"19",x"18",x"F3",x"21",x"C4",x"0E",x"3A",x"0C",x"89",x"FE",x"00",
		x"28",x"0F",x"3D",x"21",x"D4",x"0E",x"11",x"12",x"00",x"FE",x"00",x"28",x"04",x"19",x"3D",x"18",
		x"F8",x"FD",x"75",x"01",x"FD",x"74",x"02",x"FD",x"E1",x"E1",x"D1",x"C9",x"D5",x"E5",x"3A",x"8D",
		x"80",x"FE",x"00",x"20",x"29",x"2A",x"0A",x"89",x"7C",x"B5",x"20",x"11",x"DD",x"66",x"04",x"DD",
		x"6E",x"06",x"ED",x"5B",x"08",x"89",x"19",x"DD",x"74",x"04",x"DD",x"75",x"06",x"DD",x"66",x"05",
		x"DD",x"6E",x"07",x"ED",x"5B",x"0A",x"89",x"19",x"DD",x"74",x"05",x"DD",x"75",x"07",x"3A",x"02",
		x"89",x"32",x"10",x"85",x"3A",x"03",x"89",x"32",x"11",x"85",x"3A",x"04",x"89",x"32",x"12",x"85",
		x"3A",x"05",x"89",x"32",x"13",x"85",x"E1",x"D1",x"C9",x"CD",x"C1",x"28",x"3A",x"0C",x"89",x"FE",
		x"01",x"20",x"0B",x"3A",x"AC",x"81",x"FE",x"04",x"30",x"04",x"3C",x"32",x"AC",x"81",x"3E",x"00",
		x"32",x"00",x"89",x"32",x"10",x"89",x"C9",x"E5",x"3E",x"00",x"32",x"00",x"89",x"32",x"10",x"89",
		x"21",x"00",x"00",x"22",x"02",x"89",x"22",x"06",x"89",x"22",x"08",x"89",x"22",x"0A",x"89",x"E1",
		x"C9",x"C5",x"FD",x"E5",x"3A",x"0C",x"89",x"3D",x"FD",x"21",x"8C",x"2F",x"FE",x"00",x"28",x"07",
		x"FD",x"23",x"FD",x"23",x"3D",x"18",x"F5",x"FD",x"46",x"01",x"FD",x"4E",x"00",x"CD",x"E4",x"00",
		x"FD",x"E1",x"C1",x"C9",x"C5",x"D5",x"E5",x"21",x"EA",x"2D",x"11",x"14",x"89",x"01",x"68",x"00",
		x"ED",x"B0",x"CD",x"CF",x"00",x"CA",x"2D",x"10",x"E1",x"D1",x"C1",x"C9",x"CD",x"10",x"29",x"CD",
		x"CF",x"00",x"CE",x"2D",x"02",x"C9",x"CD",x"50",x"29",x"CD",x"CF",x"00",x"D2",x"2D",x"0C",x"C9",
		x"D5",x"E5",x"FD",x"E5",x"FD",x"21",x"52",x"2E",x"3A",x"AC",x"81",x"11",x"08",x"00",x"FE",x"00",
		x"28",x"05",x"FD",x"19",x"3D",x"18",x"F7",x"FD",x"66",x"01",x"FD",x"6E",x"00",x"22",x"26",x"89",
		x"FD",x"66",x"03",x"FD",x"6E",x"02",x"22",x"28",x"89",x"FD",x"66",x"05",x"FD",x"6E",x"04",x"22",
		x"2E",x"89",x"FD",x"66",x"07",x"FD",x"6E",x"06",x"22",x"30",x"89",x"FD",x"E1",x"E1",x"D1",x"C9",
		x"D5",x"E5",x"FD",x"E5",x"21",x"24",x"24",x"22",x"36",x"89",x"22",x"3C",x"89",x"22",x"42",x"89",
		x"22",x"48",x"89",x"22",x"4E",x"89",x"22",x"54",x"89",x"22",x"5A",x"89",x"22",x"60",x"89",x"22",
		x"66",x"89",x"22",x"6C",x"89",x"22",x"72",x"89",x"22",x"78",x"89",x"FD",x"21",x"7A",x"2E",x"3A",
		x"A7",x"81",x"CB",x"3F",x"11",x"04",x"00",x"FE",x"00",x"28",x"0A",x"FD",x"19",x"3D",x"FE",x"00",
		x"28",x"03",x"FD",x"19",x"3D",x"FD",x"66",x"01",x"FD",x"6E",x"00",x"22",x"36",x"89",x"22",x"3C",
		x"89",x"FD",x"66",x"03",x"FD",x"6E",x"02",x"22",x"42",x"89",x"22",x"48",x"89",x"FE",x"00",x"CA",
		x"18",x"2A",x"FD",x"21",x"86",x"2E",x"3D",x"FE",x"00",x"28",x"11",x"FD",x"19",x"3D",x"FE",x"00",
		x"28",x"0A",x"FD",x"19",x"3D",x"FE",x"00",x"28",x"03",x"FD",x"19",x"3D",x"FD",x"66",x"01",x"FD",
		x"6E",x"00",x"22",x"4E",x"89",x"22",x"54",x"89",x"FD",x"66",x"03",x"FD",x"6E",x"02",x"22",x"5A",
		x"89",x"22",x"60",x"89",x"FE",x"00",x"CA",x"18",x"2A",x"FD",x"21",x"96",x"2E",x"3D",x"28",x"10",
		x"FD",x"19",x"3D",x"FE",x"00",x"28",x"09",x"FD",x"19",x"3D",x"FE",x"00",x"28",x"02",x"FD",x"19",
		x"FD",x"66",x"01",x"FD",x"6E",x"00",x"22",x"66",x"89",x"22",x"6C",x"89",x"FD",x"66",x"03",x"FD",
		x"6E",x"02",x"22",x"72",x"89",x"22",x"78",x"89",x"FD",x"E1",x"E1",x"D1",x"C9",x"DD",x"7E",x"10",
		x"FE",x"00",x"28",x"06",x"DD",x"35",x"10",x"C3",x"A9",x"2A",x"2A",x"5C",x"82",x"B7",x"CB",x"2C",
		x"CB",x"1D",x"DD",x"CB",x"09",x"7E",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"74",x"09",x"DD",x"75",
		x"08",x"2A",x"5C",x"82",x"DD",x"CB",x"0B",x"7E",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"74",x"0B",
		x"DD",x"75",x"0A",x"DD",x"46",x"04",x"DD",x"4E",x"05",x"CD",x"F2",x"5F",x"FE",x"00",x"CA",x"94",
		x"2A",x"DD",x"36",x"10",x"01",x"4F",x"E6",x"0C",x"FE",x"00",x"28",x"0F",x"DD",x"66",x"0B",x"DD",
		x"6E",x"0A",x"CD",x"F3",x"1F",x"DD",x"74",x"0B",x"DD",x"75",x"0A",x"79",x"E6",x"03",x"FE",x"00",
		x"28",x"0F",x"DD",x"66",x"09",x"DD",x"6E",x"08",x"CD",x"F3",x"1F",x"DD",x"74",x"09",x"DD",x"75",
		x"08",x"C3",x"A9",x"2A",x"21",x"6E",x"2F",x"CD",x"10",x"2B",x"FD",x"74",x"00",x"FD",x"75",x"01",
		x"CD",x"AA",x"2A",x"CD",x"F3",x"2C",x"CD",x"89",x"2B",x"C9",x"C5",x"D5",x"E5",x"21",x"A6",x"2E",
		x"DD",x"7E",x"01",x"FE",x"02",x"28",x"18",x"21",x"CE",x"2E",x"FE",x"03",x"28",x"11",x"21",x"F6",
		x"2E",x"FE",x"04",x"28",x"0A",x"21",x"1E",x"2F",x"FE",x"05",x"28",x"03",x"21",x"46",x"2F",x"DD",
		x"CB",x"09",x"7E",x"20",x"04",x"11",x"14",x"00",x"19",x"DD",x"34",x"11",x"DD",x"4E",x"11",x"7E",
		x"B9",x"28",x"02",x"30",x"27",x"23",x"54",x"5D",x"DD",x"34",x"12",x"DD",x"34",x"12",x"06",x"00",
		x"DD",x"4E",x"12",x"09",x"7E",x"FE",x"FF",x"20",x"07",x"DD",x"36",x"12",x"00",x"62",x"6B",x"7E",
		x"DD",x"77",x"02",x"23",x"7E",x"DD",x"77",x"03",x"DD",x"36",x"11",x"00",x"E1",x"D1",x"C1",x"C9",
		x"D5",x"11",x"00",x"00",x"DD",x"7E",x"08",x"DD",x"B6",x"09",x"20",x"07",x"DD",x"CB",x"0B",x"7E",
		x"C2",x"83",x"2B",x"23",x"23",x"DD",x"CB",x"09",x"7E",x"20",x"07",x"DD",x"CB",x"0B",x"7E",x"C2",
		x"83",x"2B",x"23",x"23",x"DD",x"7E",x"0A",x"DD",x"B6",x"0B",x"20",x"07",x"DD",x"CB",x"09",x"7E",
		x"CA",x"83",x"2B",x"23",x"23",x"DD",x"CB",x"09",x"7E",x"20",x"07",x"DD",x"CB",x"0B",x"7E",x"CA",
		x"83",x"2B",x"23",x"23",x"DD",x"7E",x"08",x"DD",x"B6",x"09",x"20",x"07",x"DD",x"CB",x"0B",x"7E",
		x"CA",x"83",x"2B",x"23",x"23",x"DD",x"CB",x"09",x"7E",x"28",x"06",x"DD",x"CB",x"0B",x"7E",x"20",
		x"12",x"23",x"23",x"DD",x"7E",x"0A",x"DD",x"B6",x"0B",x"20",x"06",x"DD",x"CB",x"09",x"7E",x"20",
		x"02",x"23",x"23",x"56",x"23",x"5E",x"EB",x"D1",x"C9",x"C5",x"DD",x"7E",x"04",x"FD",x"77",x"02",
		x"DD",x"7E",x"01",x"0E",x"04",x"CB",x"4F",x"28",x"02",x"0E",x"FC",x"DD",x"7E",x"05",x"81",x"FD",
		x"77",x"03",x"C1",x"C9",x"2A",x"60",x"82",x"DD",x"75",x"0C",x"DD",x"74",x"0D",x"DD",x"75",x"0E",
		x"DD",x"74",x"0F",x"DD",x"7E",x"01",x"FE",x"04",x"20",x"1C",x"DD",x"36",x"0C",x"00",x"DD",x"36",
		x"0D",x"00",x"2A",x"5C",x"82",x"DD",x"CB",x"09",x"7E",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"74",
		x"09",x"DD",x"75",x"08",x"18",x"19",x"3A",x"02",x"85",x"47",x"DD",x"7E",x"04",x"90",x"38",x"0F",
		x"DD",x"66",x"0D",x"DD",x"6E",x"0C",x"CD",x"F3",x"1F",x"DD",x"74",x"0D",x"DD",x"75",x"0C",x"DD",
		x"7E",x"01",x"FE",x"03",x"20",x"1C",x"DD",x"36",x"0E",x"00",x"DD",x"36",x"0F",x"00",x"2A",x"5C",
		x"82",x"DD",x"CB",x"0B",x"7E",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"74",x"0B",x"DD",x"75",x"0A",
		x"18",x"19",x"3A",x"03",x"85",x"47",x"DD",x"7E",x"05",x"90",x"38",x"0F",x"DD",x"66",x"0F",x"DD",
		x"6E",x"0E",x"CD",x"F3",x"1F",x"DD",x"74",x"0F",x"DD",x"75",x"0E",x"DD",x"46",x"04",x"DD",x"4E",
		x"05",x"CD",x"F2",x"5F",x"FE",x"00",x"CA",x"79",x"2C",x"DD",x"36",x"10",x"01",x"4F",x"E6",x"0C",
		x"FE",x"00",x"28",x"17",x"DD",x"66",x"0B",x"DD",x"6E",x"0A",x"CD",x"F3",x"1F",x"DD",x"74",x"0B",
		x"DD",x"75",x"0A",x"DD",x"36",x"0E",x"00",x"DD",x"36",x"0F",x"00",x"79",x"E6",x"03",x"FE",x"00",
		x"28",x"17",x"DD",x"66",x"09",x"DD",x"6E",x"08",x"CD",x"F3",x"1F",x"DD",x"74",x"09",x"DD",x"75",
		x"08",x"DD",x"36",x"0C",x"00",x"DD",x"36",x"0D",x"00",x"CD",x"92",x"2C",x"CD",x"F3",x"2C",x"21",
		x"6E",x"2F",x"CD",x"10",x"2B",x"FD",x"74",x"00",x"FD",x"75",x"01",x"CD",x"AA",x"2A",x"CD",x"89",
		x"2B",x"C9",x"C5",x"D5",x"E5",x"DD",x"7E",x"01",x"FE",x"04",x"28",x"26",x"DD",x"66",x"09",x"DD",
		x"6E",x"08",x"DD",x"56",x"0D",x"DD",x"5E",x"0C",x"19",x"44",x"4D",x"CD",x"F0",x"1F",x"ED",x"5B",
		x"5C",x"82",x"ED",x"52",x"7C",x"B5",x"28",x"04",x"CB",x"7C",x"28",x"06",x"DD",x"70",x"09",x"DD",
		x"71",x"08",x"DD",x"7E",x"01",x"FE",x"03",x"28",x"26",x"DD",x"66",x"0B",x"DD",x"6E",x"0A",x"DD",
		x"56",x"0F",x"DD",x"5E",x"0E",x"19",x"44",x"4D",x"CD",x"F0",x"1F",x"ED",x"5B",x"5C",x"82",x"ED",
		x"52",x"7C",x"B5",x"28",x"04",x"CB",x"7C",x"28",x"06",x"DD",x"70",x"0B",x"DD",x"71",x"0A",x"D1",
		x"E1",x"C1",x"C9",x"3A",x"8D",x"80",x"FE",x"00",x"C0",x"E5",x"D5",x"DD",x"66",x"04",x"DD",x"6E",
		x"06",x"DD",x"56",x"09",x"DD",x"5E",x"08",x"19",x"DD",x"74",x"04",x"DD",x"75",x"06",x"DD",x"66",
		x"05",x"DD",x"6E",x"07",x"DD",x"56",x"0B",x"DD",x"5E",x"0A",x"19",x"DD",x"74",x"05",x"DD",x"75",
		x"07",x"D1",x"E1",x"C9",x"DD",x"7E",x"01",x"FD",x"77",x"00",x"DD",x"7E",x"02",x"FD",x"77",x"01",
		x"DD",x"7E",x"03",x"FD",x"77",x"02",x"DD",x"7E",x"04",x"FD",x"77",x"03",x"C9",x"DD",x"46",x"04",
		x"DD",x"4E",x"05",x"CD",x"F2",x"5F",x"FE",x"00",x"CA",x"B4",x"2D",x"4F",x"16",x"00",x"DD",x"5E",
		x"04",x"3A",x"02",x"85",x"26",x"00",x"6F",x"B7",x"ED",x"52",x"3A",x"64",x"82",x"54",x"5D",x"FE",
		x"00",x"28",x"04",x"19",x"3D",x"18",x"F8",x"CB",x"7C",x"28",x"04",x"CB",x"49",x"20",x"08",x"CB",
		x"7C",x"20",x"07",x"CB",x"41",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"75",x"08",x"DD",x"74",x"09",
		x"16",x"00",x"DD",x"5E",x"05",x"3A",x"03",x"85",x"26",x"00",x"6F",x"B7",x"ED",x"52",x"3A",x"64",
		x"82",x"54",x"5D",x"FE",x"00",x"28",x"04",x"19",x"3D",x"18",x"F8",x"CB",x"7C",x"28",x"04",x"CB",
		x"59",x"20",x"08",x"CB",x"7C",x"20",x"07",x"CB",x"51",x"28",x"03",x"CD",x"F3",x"1F",x"DD",x"75",
		x"0A",x"DD",x"74",x"0B",x"CD",x"F3",x"2C",x"21",x"6E",x"2F",x"CD",x"10",x"2B",x"FD",x"74",x"00",
		x"FD",x"75",x"01",x"CD",x"AA",x"2A",x"CD",x"89",x"2B",x"C9",x"14",x"89",x"1C",x"89",x"24",x"89",
		x"2C",x"89",x"34",x"89",x"3A",x"89",x"40",x"89",x"46",x"89",x"4C",x"89",x"52",x"89",x"58",x"89",
		x"5E",x"89",x"64",x"89",x"6A",x"89",x"70",x"89",x"76",x"89",x"00",x"0E",x"C2",x"0E",x"C0",x"0E",
		x"FF",x"FF",x"01",x"0E",x"C3",x"0E",x"C1",x"0E",x"FF",x"FF",x"00",x"10",x"C6",x"0E",x"C4",x"0E",
		x"FF",x"FF",x"01",x"10",x"C7",x"0E",x"C5",x"0E",x"FF",x"FF",x"00",x"0D",x"E4",x"0E",x"FF",x"FF",
		x"01",x"0D",x"E4",x"0E",x"FF",x"FF",x"00",x"12",x"D8",x"0E",x"FF",x"FF",x"01",x"12",x"D8",x"0E",
		x"FF",x"FF",x"00",x"0C",x"00",x"0E",x"FF",x"FF",x"01",x"0C",x"00",x"0E",x"FF",x"FF",x"00",x"13",
		x"00",x"0E",x"FF",x"FF",x"01",x"13",x"00",x"0E",x"FF",x"FF",x"00",x"0B",x"00",x"0E",x"FF",x"FF",
		x"01",x"0B",x"00",x"0E",x"FF",x"FF",x"00",x"14",x"00",x"0E",x"FF",x"FF",x"01",x"14",x"00",x"0E",
		x"FF",x"FF",x"C6",x"0E",x"C4",x"0E",x"C7",x"0E",x"C5",x"0E",x"CA",x"0E",x"C8",x"0E",x"CB",x"0E",
		x"C9",x"0E",x"CE",x"0E",x"CC",x"0E",x"CF",x"0E",x"CD",x"0E",x"D2",x"0E",x"D0",x"0E",x"D3",x"0E",
		x"D1",x"0E",x"D6",x"0E",x"D4",x"0E",x"D7",x"0E",x"D5",x"0E",x"E4",x"0E",x"D8",x"0E",x"E5",x"0E",
		x"D9",x"0E",x"E6",x"0E",x"DA",x"0E",x"E8",x"0E",x"DC",x"0E",x"E9",x"0E",x"DD",x"0E",x"EA",x"0E",
		x"DE",x"0E",x"EB",x"0E",x"DF",x"0E",x"EC",x"0E",x"E0",x"0E",x"ED",x"0E",x"E1",x"0E",x"EE",x"0E",
		x"E2",x"0E",x"EF",x"0E",x"E3",x"0E",x"07",x"50",x"04",x"51",x"04",x"52",x"04",x"53",x"04",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"50",x"84",x"51",x"84",x"52",
		x"84",x"53",x"84",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"02",x"67",
		x"04",x"68",x"04",x"69",x"04",x"6A",x"04",x"6B",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"02",x"67",x"04",x"68",x"04",x"69",x"04",x"6A",x"04",x"6B",x"04",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"54",x"04",x"55",x"04",x"56",x"04",x"57",x"04",x"58",
		x"04",x"59",x"04",x"5A",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"5A",x"04",x"59",x"04",x"58",
		x"04",x"57",x"04",x"56",x"04",x"55",x"04",x"54",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"06",x"38",
		x"04",x"39",x"04",x"3A",x"04",x"3B",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"06",x"38",x"84",x"39",x"84",x"3A",x"84",x"3B",x"84",x"FF",x"FF",x"39",x"04",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"06",x"60",x"04",x"61",x"04",x"62",x"04",x"63",x"04",x"64",
		x"04",x"65",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"06",x"65",x"04",x"64",x"04",x"63",
		x"04",x"62",x"04",x"61",x"04",x"60",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",
		x"00",x"02",x"00",x"03",x"00",x"05",x"00",x"08",x"00",x"12",x"00",x"20",x"00",x"10",x"00",x"30",
		x"00",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C3",x"E4",x"28",x"C3",x"FC",x"28",x"C3",x"06",x"29",x"C3",x"05",x"22",x"C3",x"FF",x"FF",x"00",
		x"C3",x"1D",x"2A",x"C3",x"A4",x"2B",x"C3",x"3D",x"2D",x"C3",x"A9",x"24",x"00",x"00",x"00",x"00",
		x"3A",x"88",x"80",x"FE",x"03",x"CA",x"83",x"30",x"3A",x"8E",x"80",x"B7",x"C2",x"83",x"30",x"CD",
		x"8F",x"3C",x"3A",x"28",x"80",x"CB",x"7F",x"C2",x"3A",x"30",x"3A",x"8D",x"80",x"B7",x"C2",x"3A",
		x"30",x"CD",x"83",x"31",x"CD",x"1A",x"32",x"CD",x"5A",x"33",x"3E",x"01",x"CD",x"81",x"3D",x"C4",
		x"44",x"3D",x"3E",x"20",x"CD",x"81",x"3D",x"C4",x"C8",x"3C",x"DD",x"21",x"78",x"82",x"FD",x"21",
		x"18",x"85",x"11",x"19",x"00",x"06",x"09",x"0E",x"00",x"C5",x"D5",x"DD",x"7E",x"00",x"B7",x"CA",
		x"5E",x"30",x"1F",x"0C",x"D2",x"52",x"30",x"21",x"86",x"30",x"79",x"CD",x"EA",x"00",x"D1",x"C1",
		x"DD",x"19",x"D5",x"11",x"08",x"00",x"FD",x"19",x"D1",x"10",x"DE",x"CD",x"00",x"60",x"3A",x"8D",
		x"80",x"B7",x"CA",x"83",x"30",x"3A",x"28",x"80",x"CB",x"57",x"C2",x"83",x"30",x"3E",x"00",x"32",
		x"4B",x"82",x"C9",x"C3",x"C3",x"00",x"81",x"31",x"98",x"30",x"81",x"31",x"EF",x"30",x"81",x"31",
		x"81",x"31",x"35",x"31",x"81",x"31",x"81",x"31",x"DD",x"7E",x"01",x"21",x"CF",x"30",x"CD",x"EA",
		x"00",x"DD",x"7E",x"01",x"FE",x"0C",x"D2",x"CE",x"30",x"DD",x"7E",x"01",x"FE",x"01",x"CA",x"CE",
		x"30",x"DD",x"7E",x"01",x"FE",x"08",x"CA",x"CE",x"30",x"DD",x"7E",x"01",x"FE",x"07",x"CA",x"CE",
		x"30",x"3A",x"4A",x"82",x"B7",x"C2",x"CE",x"30",x"21",x"BB",x"3D",x"CD",x"07",x"36",x"C9",x"81",
		x"31",x"1C",x"32",x"73",x"32",x"81",x"31",x"10",x"33",x"81",x"31",x"81",x"31",x"1D",x"33",x"66",
		x"32",x"81",x"31",x"81",x"31",x"81",x"31",x"CE",x"39",x"1F",x"3A",x"C0",x"3A",x"81",x"31",x"00",
		x"DD",x"7E",x"01",x"21",x"15",x"31",x"CD",x"EA",x"00",x"DD",x"7E",x"01",x"FE",x"0C",x"D2",x"14",
		x"31",x"CD",x"CB",x"34",x"CD",x"32",x"3B",x"3A",x"4A",x"82",x"B7",x"C2",x"14",x"31",x"21",x"C3",
		x"3D",x"CD",x"07",x"36",x"C9",x"81",x"31",x"81",x"31",x"E2",x"33",x"63",x"34",x"81",x"31",x"81",
		x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"CE",x"39",x"1F",
		x"3A",x"C0",x"3A",x"81",x"31",x"00",x"DD",x"7E",x"01",x"21",x"61",x"31",x"CD",x"EA",x"00",x"DD",
		x"7E",x"01",x"FE",x"0C",x"30",x"1A",x"3A",x"4A",x"82",x"B7",x"C2",x"60",x"31",x"DD",x"7E",x"13",
		x"B7",x"CA",x"5A",x"31",x"DD",x"35",x"13",x"C3",x"60",x"31",x"21",x"C7",x"3D",x"CD",x"07",x"36",
		x"C9",x"81",x"31",x"6B",x"35",x"F2",x"35",x"F9",x"35",x"F9",x"35",x"F9",x"35",x"00",x"36",x"81",
		x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"81",x"31",x"CE",x"39",x"1F",x"3A",x"C0",x"3A",x"81",
		x"31",x"00",x"C9",x"21",x"D2",x"80",x"7E",x"23",x"BE",x"CA",x"19",x"32",x"2A",x"DA",x"80",x"2B",
		x"22",x"DA",x"80",x"7D",x"B4",x"C2",x"19",x"32",x"3A",x"D3",x"80",x"3C",x"32",x"D3",x"80",x"2A",
		x"D4",x"80",x"22",x"DA",x"80",x"DD",x"21",x"AA",x"82",x"06",x"07",x"CD",x"B7",x"38",x"B7",x"C2",
		x"19",x"32",x"21",x"CF",x"3D",x"CD",x"67",x"38",x"3A",x"2B",x"80",x"D6",x"78",x"38",x"09",x"DD",
		x"7E",x"04",x"FE",x"78",x"30",x"EC",x"18",x"07",x"DD",x"7E",x"04",x"FE",x"78",x"38",x"E3",x"DD",
		x"7E",x"04",x"C6",x"F8",x"DD",x"77",x"04",x"DD",x"7E",x"05",x"C6",x"F8",x"DD",x"77",x"05",x"DD",
		x"36",x"00",x"01",x"DD",x"36",x"01",x"01",x"DD",x"36",x"03",x"0F",x"DD",x"CB",x"03",x"EE",x"21",
		x"80",x"00",x"DD",x"75",x"08",x"DD",x"74",x"09",x"DD",x"36",x"0E",x"10",x"DD",x"36",x"0F",x"00",
		x"DD",x"36",x"14",x"01",x"2A",x"D6",x"80",x"DD",x"75",x"16",x"DD",x"74",x"17",x"3A",x"8D",x"80",
		x"B7",x"C2",x"19",x"32",x"3E",x"15",x"CD",x"FC",x"00",x"C9",x"00",x"C9",x"00",x"DD",x"35",x"14",
		x"C2",x"65",x"32",x"DD",x"36",x"14",x"06",x"21",x"73",x"3E",x"01",x"01",x"00",x"DD",x"7E",x"10",
		x"CD",x"F6",x"00",x"7E",x"FE",x"FF",x"CA",x"41",x"32",x"DD",x"77",x"02",x"DD",x"34",x"10",x"18",
		x"24",x"DD",x"36",x"02",x"04",x"DD",x"36",x"03",x"04",x"DD",x"36",x"10",x"00",x"DD",x"36",x"14",
		x"1E",x"DD",x"36",x"01",x"08",x"DD",x"7E",x"04",x"C6",x"08",x"DD",x"77",x"04",x"DD",x"7E",x"05",
		x"C6",x"08",x"DD",x"77",x"05",x"C9",x"DD",x"35",x"14",x"C2",x"6F",x"32",x"CD",x"AF",x"3B",x"CD",
		x"D6",x"32",x"C9",x"DD",x"6E",x"16",x"DD",x"66",x"17",x"7C",x"B5",x"CA",x"85",x"32",x"2B",x"DD",
		x"75",x"16",x"DD",x"74",x"17",x"CD",x"33",x"36",x"DD",x"7E",x"01",x"FE",x"02",x"C2",x"93",x"32",
		x"CD",x"09",x"60",x"CD",x"D6",x"32",x"CD",x"28",x"37",x"DD",x"7E",x"05",x"FE",x"D0",x"DA",x"D5",
		x"32",x"DD",x"36",x"01",x"07",x"DD",x"36",x"02",x"BC",x"DD",x"36",x"03",x"0F",x"DD",x"7E",x"04",
		x"C6",x"F8",x"DD",x"77",x"04",x"DD",x"7E",x"05",x"C6",x"F8",x"DD",x"77",x"05",x"DD",x"CB",x"03",
		x"EE",x"DD",x"36",x"10",x"00",x"DD",x"36",x"14",x"01",x"3A",x"8D",x"80",x"B7",x"C2",x"D5",x"32",
		x"3E",x"2D",x"CD",x"FC",x"00",x"C9",x"3A",x"4B",x"82",x"B7",x"C2",x"0F",x"33",x"3A",x"28",x"80",
		x"CB",x"7F",x"CA",x"0F",x"33",x"DD",x"E5",x"DD",x"E5",x"E1",x"11",x"E1",x"00",x"DD",x"19",x"DD",
		x"E5",x"D1",x"01",x"19",x"00",x"ED",x"B0",x"DD",x"E1",x"DD",x"36",x"01",x"0E",x"3E",x"22",x"DD",
		x"36",x"03",x"0B",x"DD",x"36",x"02",x"3F",x"FD",x"36",x"04",x"00",x"FD",x"36",x"05",x"00",x"C9",
		x"CD",x"03",x"60",x"CD",x"A9",x"36",x"CD",x"D6",x"32",x"CD",x"7A",x"37",x"C9",x"DD",x"35",x"14",
		x"C2",x"59",x"33",x"DD",x"36",x"14",x"06",x"21",x"73",x"3E",x"01",x"01",x"00",x"DD",x"7E",x"10",
		x"CD",x"F6",x"00",x"7E",x"FE",x"FF",x"CA",x"41",x"33",x"DD",x"77",x"02",x"DD",x"34",x"10",x"18",
		x"18",x"DD",x"36",x"00",x"20",x"DD",x"36",x"01",x"01",x"DD",x"7E",x"04",x"C6",x"08",x"DD",x"77",
		x"04",x"DD",x"7E",x"05",x"C6",x"08",x"DD",x"77",x"05",x"C9",x"21",x"C0",x"80",x"7E",x"23",x"BE",
		x"CA",x"E1",x"33",x"47",x"C5",x"DD",x"21",x"78",x"82",x"06",x"02",x"CD",x"B7",x"38",x"B7",x"C2",
		x"DE",x"33",x"DD",x"36",x"00",x"04",x"DD",x"36",x"01",x"02",x"DD",x"36",x"02",x"29",x"DD",x"36",
		x"03",x"84",x"DD",x"36",x"0D",x"01",x"DD",x"36",x"0E",x"00",x"DD",x"36",x"12",x"01",x"21",x"4F",
		x"3E",x"CD",x"70",x"38",x"3A",x"2B",x"80",x"D6",x"78",x"38",x"09",x"DD",x"7E",x"04",x"FE",x"78",
		x"30",x"EC",x"18",x"07",x"DD",x"7E",x"04",x"FE",x"78",x"38",x"E3",x"C1",x"C5",x"05",x"C2",x"C2",
		x"33",x"2A",x"4C",x"82",x"DD",x"5E",x"04",x"DD",x"56",x"05",x"B7",x"ED",x"52",x"CA",x"8E",x"33",
		x"18",x"09",x"DD",x"6E",x"04",x"DD",x"66",x"05",x"22",x"4C",x"82",x"21",x"C4",x"80",x"CD",x"87",
		x"38",x"3A",x"C1",x"80",x"3C",x"32",x"C1",x"80",x"3A",x"C8",x"80",x"DD",x"77",x"16",x"C1",x"10",
		x"83",x"C9",x"DD",x"7E",x"18",x"B7",x"C2",x"59",x"34",x"DD",x"36",x"18",x"01",x"CD",x"1D",x"3C",
		x"B7",x"C2",x"59",x"34",x"DD",x"35",x"12",x"C2",x"59",x"34",x"DD",x"36",x"12",x"03",x"2A",x"C4",
		x"80",x"DD",x"75",x"08",x"DD",x"74",x"09",x"DD",x"75",x"0A",x"DD",x"74",x"0B",x"DD",x"7E",x"11",
		x"DD",x"77",x"10",x"3A",x"C2",x"80",x"32",x"6C",x"84",x"32",x"6D",x"84",x"32",x"6E",x"84",x"32",
		x"6F",x"84",x"21",x"6C",x"84",x"CD",x"9E",x"38",x"CD",x"06",x"60",x"B7",x"C3",x"34",x"34",x"CD",
		x"DC",x"38",x"18",x"0E",x"CD",x"1C",x"39",x"DD",x"70",x"11",x"7A",x"BB",x"D2",x"42",x"34",x"DD",
		x"71",x"11",x"CD",x"FC",x"3B",x"CD",x"84",x"39",x"B7",x"CA",x"4F",x"34",x"CD",x"0D",x"37",x"CD",
		x"06",x"3B",x"DD",x"7E",x"0F",x"B7",x"C2",x"5F",x"34",x"CD",x"09",x"60",x"CD",x"7A",x"3B",x"CD",
		x"D6",x"32",x"C9",x"DD",x"35",x"12",x"C2",x"C7",x"34",x"DD",x"7E",x"13",x"DD",x"77",x"12",x"DD",
		x"6E",x"14",x"DD",x"66",x"15",x"7E",x"FE",x"FF",x"CA",x"87",x"34",x"DD",x"77",x"02",x"23",x"DD",
		x"75",x"14",x"DD",x"74",x"15",x"18",x"40",x"23",x"3E",x"04",x"B6",x"DD",x"77",x"03",x"23",x"7E",
		x"DD",x"77",x"02",x"DD",x"36",x"0D",x"06",x"DD",x"36",x"0E",x"00",x"DD",x"36",x"12",x"03",x"DD",
		x"36",x"13",x"00",x"DD",x"36",x"14",x"00",x"DD",x"36",x"15",x"00",x"DD",x"36",x"01",x"02",x"DD",
		x"7E",x"0F",x"B7",x"CA",x"C7",x"34",x"DD",x"7E",x"17",x"DD",x"77",x"11",x"DD",x"36",x"17",x"00",
		x"CD",x"CB",x"34",x"DD",x"36",x"0F",x"00",x"CD",x"D6",x"32",x"C9",x"DD",x"7E",x"10",x"DD",x"BE",
		x"11",x"CA",x"F0",x"34",x"21",x"F1",x"34",x"01",x"08",x"00",x"DD",x"7E",x"10",x"CD",x"F6",x"00",
		x"DD",x"7E",x"11",x"CD",x"EA",x"00",x"DD",x"7E",x"11",x"DD",x"77",x"10",x"DD",x"36",x"01",x"03",
		x"C9",x"81",x"31",x"11",x"35",x"16",x"35",x"1B",x"35",x"20",x"35",x"81",x"31",x"25",x"35",x"2A",
		x"35",x"2F",x"35",x"34",x"35",x"81",x"31",x"39",x"35",x"3E",x"35",x"43",x"35",x"48",x"35",x"81",
		x"31",x"21",x"78",x"3E",x"18",x"37",x"21",x"7F",x"3E",x"18",x"32",x"21",x"86",x"3E",x"18",x"2D",
		x"21",x"8D",x"3E",x"18",x"28",x"21",x"94",x"3E",x"18",x"23",x"21",x"9B",x"3E",x"18",x"1E",x"21",
		x"A2",x"3E",x"18",x"19",x"21",x"A9",x"3E",x"18",x"14",x"21",x"B0",x"3E",x"18",x"0F",x"21",x"B7",
		x"3E",x"18",x"0A",x"21",x"BE",x"3E",x"18",x"05",x"21",x"C5",x"3E",x"18",x"00",x"DD",x"7E",x"03",
		x"E6",x"0F",x"B6",x"DD",x"77",x"03",x"23",x"7E",x"DD",x"77",x"02",x"23",x"DD",x"75",x"14",x"DD",
		x"74",x"15",x"DD",x"36",x"12",x"06",x"DD",x"36",x"13",x"06",x"C9",x"3A",x"B0",x"81",x"21",x"68",
		x"82",x"01",x"01",x"00",x"CD",x"F6",x"00",x"7E",x"E6",x"0F",x"F5",x"C6",x"02",x"DD",x"77",x"01",
		x"F1",x"21",x"D2",x"3E",x"01",x"02",x"00",x"CD",x"F6",x"00",x"7E",x"DD",x"77",x"03",x"23",x"7E",
		x"DD",x"77",x"02",x"DD",x"E5",x"06",x"13",x"DD",x"36",x"06",x"00",x"DD",x"23",x"10",x"F8",x"DD",
		x"E1",x"DD",x"36",x"13",x"1E",x"3E",x"01",x"32",x"77",x"82",x"3A",x"B0",x"81",x"3C",x"32",x"B0",
		x"81",x"3A",x"B0",x"81",x"FE",x"08",x"DA",x"BE",x"35",x"3E",x"00",x"32",x"B0",x"81",x"DD",x"36",
		x"0A",x"0A",x"DD",x"7E",x"01",x"FE",x"04",x"C2",x"D3",x"35",x"2A",x"5C",x"82",x"DD",x"75",x"0A",
		x"DD",x"74",x"0B",x"DD",x"7E",x"01",x"FE",x"02",x"C2",x"F1",x"35",x"FD",x"36",x"00",x"69",x"FD",
		x"36",x"01",x"45",x"DD",x"7E",x"04",x"FD",x"77",x"02",x"DD",x"7E",x"05",x"C6",x"FC",x"FD",x"77",
		x"03",x"C9",x"CD",x"F0",x"2F",x"CD",x"D6",x"32",x"C9",x"CD",x"F3",x"2F",x"CD",x"D6",x"32",x"C9",
		x"CD",x"F6",x"2F",x"CD",x"D6",x"32",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3A",
		x"8D",x"80",x"B7",x"C2",x"32",x"36",x"3A",x"28",x"80",x"CB",x"7F",x"C2",x"32",x"36",x"CD",x"9E",
		x"38",x"CD",x"06",x"60",x"B7",x"CA",x"32",x"36",x"21",x"28",x"80",x"CB",x"D6",x"3E",x"01",x"32",
		x"4B",x"82",x"C9",x"DD",x"46",x"04",x"DD",x"4E",x"05",x"78",x"E6",x"07",x"C2",x"A8",x"36",x"CD",
		x"00",x"38",x"B7",x"CA",x"A8",x"36",x"DD",x"7E",x"11",x"3C",x"E6",x"01",x"DD",x"77",x"11",x"AF",
		x"B1",x"C2",x"A8",x"36",x"DD",x"7E",x"16",x"DD",x"B6",x"17",x"C2",x"A8",x"36",x"2A",x"D6",x"80",
		x"DD",x"75",x"16",x"DD",x"74",x"17",x"DD",x"36",x"01",x"04",x"DD",x"36",x"08",x"00",x"DD",x"36",
		x"09",x"00",x"21",x"80",x"00",x"DD",x"75",x"0A",x"DD",x"74",x"0B",x"DD",x"36",x"10",x"00",x"DD",
		x"7E",x"11",x"B7",x"C2",x"90",x"36",x"DD",x"7E",x"04",x"D6",x"08",x"DD",x"77",x"04",x"18",x"08",
		x"DD",x"7E",x"04",x"C6",x"08",x"DD",x"77",x"04",x"DD",x"36",x"14",x"01",x"3A",x"8D",x"80",x"B7",
		x"C2",x"A8",x"36",x"3E",x"16",x"CD",x"FC",x"00",x"C9",x"DD",x"7E",x"04",x"C6",x"08",x"47",x"DD",
		x"7E",x"05",x"C6",x"14",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",x"D6",x"5F",x"B7",x"CA",x"04",x"37",
		x"DD",x"36",x"0A",x"00",x"DD",x"36",x"0B",x"00",x"21",x"80",x"00",x"DD",x"75",x"08",x"DD",x"74",
		x"09",x"DD",x"36",x"0E",x"10",x"DD",x"36",x"0F",x"00",x"DD",x"36",x"10",x"00",x"DD",x"36",x"14",
		x"06",x"DD",x"36",x"15",x"00",x"DD",x"7E",x"05",x"E6",x"F8",x"C6",x"08",x"DD",x"77",x"05",x"DD",
		x"36",x"01",x"02",x"3A",x"8D",x"80",x"B7",x"C2",x"04",x"37",x"3E",x"17",x"CD",x"FC",x"00",x"3E",
		x"96",x"CD",x"FC",x"00",x"C9",x"11",x"F5",x"3E",x"CD",x"6B",x"39",x"B7",x"C9",x"21",x"57",x"3E",
		x"DD",x"7E",x"10",x"01",x"04",x"00",x"CD",x"F6",x"00",x"7E",x"DD",x"77",x"11",x"E5",x"CD",x"84",
		x"39",x"E1",x"23",x"B7",x"C2",x"19",x"37",x"C9",x"DD",x"7E",x"12",x"DD",x"BE",x"11",x"C2",x"4F",
		x"37",x"DD",x"35",x"14",x"C2",x"61",x"37",x"DD",x"36",x"14",x"06",x"CD",x"62",x"37",x"DD",x"34",
		x"10",x"DD",x"7E",x"10",x"FE",x"04",x"DA",x"61",x"37",x"DD",x"36",x"10",x"00",x"18",x"12",x"DD",
		x"7E",x"11",x"DD",x"77",x"12",x"DD",x"36",x"10",x"00",x"DD",x"36",x"14",x"06",x"DD",x"36",x"02",
		x"04",x"C9",x"DD",x"7E",x"11",x"B7",x"21",x"6F",x"3E",x"C2",x"6F",x"37",x"21",x"6B",x"3E",x"DD",
		x"5E",x"10",x"16",x"00",x"19",x"7E",x"DD",x"77",x"02",x"C9",x"DD",x"35",x"14",x"20",x"1A",x"DD",
		x"36",x"14",x"04",x"21",x"67",x"3E",x"DD",x"4E",x"10",x"06",x"00",x"09",x"7E",x"DD",x"77",x"02",
		x"DD",x"7E",x"10",x"3C",x"E6",x"03",x"DD",x"77",x"10",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"9F",x"3D",x"CD",x"30",x"38",x"CD",x"DE",x"00",x"7E",x"CD",x"D6",x"5F",x"B7",x"C2",x"26",
		x"38",x"21",x"97",x"3D",x"CD",x"30",x"38",x"CD",x"DE",x"00",x"7E",x"CD",x"D6",x"5F",x"B7",x"CA",
		x"2B",x"38",x"AF",x"C3",x"2F",x"38",x"0E",x"01",x"C3",x"2D",x"38",x"0E",x"00",x"3E",x"01",x"C9",
		x"DD",x"7E",x"11",x"E5",x"21",x"3A",x"38",x"C3",x"EA",x"00",x"42",x"38",x"47",x"38",x"4F",x"38",
		x"57",x"38",x"E1",x"CD",x"5B",x"38",x"C9",x"E1",x"CD",x"9B",x"38",x"CD",x"5B",x"38",x"C9",x"E1",
		x"CD",x"99",x"38",x"CD",x"5B",x"38",x"C9",x"E1",x"CD",x"97",x"38",x"DD",x"7E",x"04",x"86",x"47",
		x"23",x"DD",x"7E",x"05",x"86",x"4F",x"C9",x"01",x"08",x"00",x"3A",x"A1",x"81",x"CD",x"F6",x"00",
		x"CD",x"C9",x"00",x"3A",x"25",x"80",x"E6",x"03",x"87",x"16",x"00",x"5F",x"19",x"7E",x"DD",x"77",
		x"05",x"23",x"7E",x"DD",x"77",x"04",x"C9",x"5E",x"23",x"56",x"DD",x"73",x"08",x"DD",x"72",x"09",
		x"DD",x"73",x"0A",x"DD",x"72",x"0B",x"C9",x"23",x"23",x"23",x"23",x"23",x"23",x"C9",x"3A",x"2B",
		x"80",x"C6",x"08",x"47",x"3A",x"2C",x"80",x"C6",x"08",x"4F",x"DD",x"7E",x"04",x"C6",x"08",x"57",
		x"DD",x"7E",x"05",x"C6",x"08",x"5F",x"C9",x"11",x"19",x"00",x"AF",x"DD",x"B6",x"00",x"CA",x"CA",
		x"38",x"DD",x"19",x"10",x"F5",x"3E",x"01",x"C3",x"CC",x"38",x"3E",x"00",x"C9",x"DD",x"E5",x"06",
		x"19",x"DD",x"36",x"00",x"00",x"DD",x"23",x"10",x"F8",x"DD",x"E1",x"C9",x"CD",x"C9",x"00",x"3A",
		x"25",x"80",x"E6",x"03",x"21",x"EA",x"38",x"C3",x"EA",x"00",x"1B",x"39",x"F2",x"38",x"1B",x"39",
		x"08",x"39",x"DD",x"7E",x"11",x"FE",x"02",x"D2",x"01",x"39",x"DD",x"36",x"11",x"02",x"C3",x"1B",
		x"39",x"DD",x"36",x"11",x"00",x"C3",x"1B",x"39",x"DD",x"7E",x"11",x"FE",x"02",x"D2",x"17",x"39",
		x"DD",x"36",x"11",x"03",x"C3",x"1B",x"39",x"DD",x"36",x"11",x"01",x"C9",x"3A",x"2B",x"80",x"C6",
		x"08",x"6F",x"26",x"00",x"DD",x"7E",x"04",x"C6",x"08",x"5F",x"16",x"00",x"B7",x"ED",x"52",x"22",
		x"50",x"82",x"3A",x"2C",x"80",x"C6",x"08",x"6F",x"26",x"00",x"DD",x"7E",x"05",x"C6",x"08",x"5F",
		x"16",x"00",x"B7",x"ED",x"52",x"22",x"52",x"82",x"2A",x"50",x"82",x"7D",x"57",x"06",x"00",x"CB",
		x"7C",x"F2",x"59",x"39",x"ED",x"44",x"57",x"06",x"01",x"2A",x"52",x"82",x"7D",x"5F",x"0E",x"03",
		x"CB",x"7C",x"F2",x"6A",x"39",x"ED",x"44",x"5F",x"0E",x"02",x"C9",x"C5",x"E5",x"D5",x"E1",x"47",
		x"7E",x"23",x"FE",x"FF",x"CA",x"7F",x"39",x"B8",x"C2",x"70",x"39",x"AF",x"C3",x"81",x"39",x"3E",
		x"01",x"E1",x"C1",x"C9",x"21",x"AF",x"3D",x"CD",x"30",x"38",x"CD",x"DE",x"00",x"06",x"04",x"CD",
		x"A8",x"39",x"7E",x"C5",x"E5",x"CD",x"D6",x"5F",x"E1",x"C1",x"B7",x"C2",x"A5",x"39",x"10",x"EF",
		x"3E",x"00",x"C3",x"A7",x"39",x"3E",x"01",x"C9",x"E5",x"21",x"B0",x"39",x"78",x"C3",x"EA",x"00",
		x"CC",x"39",x"BA",x"39",x"BF",x"39",x"C7",x"39",x"CC",x"39",x"E1",x"23",x"C3",x"CD",x"39",x"E1",
		x"11",x"1F",x"00",x"19",x"C3",x"CD",x"39",x"E1",x"23",x"C3",x"CD",x"39",x"E1",x"C9",x"3A",x"49",
		x"82",x"FE",x"02",x"D2",x"DC",x"39",x"DD",x"35",x"14",x"C2",x"1E",x"3A",x"FD",x"36",x"04",x"00",
		x"FD",x"36",x"05",x"00",x"FD",x"36",x"06",x"00",x"FD",x"36",x"07",x"00",x"DD",x"7E",x"00",x"FE",
		x"01",x"C2",x"FE",x"39",x"3A",x"D3",x"80",x"3D",x"32",x"D3",x"80",x"C3",x"0D",x"3A",x"DD",x"7E",
		x"00",x"FE",x"20",x"CA",x"F4",x"39",x"3A",x"C1",x"80",x"3D",x"32",x"C1",x"80",x"CD",x"CD",x"38",
		x"3A",x"49",x"82",x"B7",x"CA",x"1E",x"3A",x"3A",x"49",x"82",x"3D",x"32",x"49",x"82",x"C9",x"DD",
		x"35",x"14",x"C2",x"81",x"3A",x"DD",x"7E",x"15",x"DD",x"77",x"14",x"21",x"DC",x"3E",x"16",x"00",
		x"DD",x"5E",x"10",x"19",x"7E",x"FE",x"FF",x"C2",x"7B",x"3A",x"DD",x"CB",x"03",x"AE",x"DD",x"7E",
		x"04",x"C6",x"08",x"DD",x"77",x"04",x"DD",x"7E",x"05",x"C6",x"08",x"DD",x"77",x"05",x"3A",x"47",
		x"82",x"21",x"03",x"00",x"CD",x"F3",x"00",x"CD",x"F1",x"3A",x"3A",x"47",x"82",x"FE",x"06",x"D2",
		x"69",x"3A",x"3A",x"47",x"82",x"3C",x"32",x"47",x"82",x"DD",x"36",x"14",x"1E",x"DD",x"36",x"01",
		x"0C",x"3A",x"49",x"82",x"3C",x"32",x"49",x"82",x"C3",x"81",x"3A",x"DD",x"77",x"02",x"DD",x"34",
		x"10",x"C9",x"21",x"CB",x"3D",x"CD",x"9E",x"38",x"CD",x"06",x"60",x"B7",x"CA",x"BF",x"3A",x"3E",
		x"2C",x"CD",x"FC",x"00",x"3A",x"B3",x"81",x"3C",x"32",x"B3",x"81",x"DD",x"36",x"10",x"00",x"DD",
		x"36",x"14",x"01",x"DD",x"36",x"15",x"04",x"DD",x"36",x"03",x"2D",x"DD",x"36",x"01",x"0D",x"DD",
		x"7E",x"04",x"C6",x"F8",x"DD",x"77",x"04",x"DD",x"7E",x"05",x"C6",x"F8",x"DD",x"77",x"05",x"C9",
		x"3A",x"28",x"80",x"CB",x"77",x"CA",x"CF",x"3A",x"DD",x"36",x"02",x"00",x"C3",x"D3",x"3A",x"DD",
		x"36",x"02",x"3F",x"3A",x"28",x"80",x"CB",x"7F",x"CA",x"E1",x"3A",x"CD",x"82",x"3A",x"C3",x"F0",
		x"3A",x"DD",x"E5",x"DD",x"E5",x"D1",x"E1",x"01",x"E1",x"00",x"09",x"01",x"19",x"00",x"ED",x"B0",
		x"C9",x"3A",x"47",x"82",x"01",x"02",x"00",x"21",x"01",x"3F",x"CD",x"F6",x"00",x"7E",x"4F",x"23",
		x"7E",x"47",x"CD",x"E4",x"00",x"C9",x"DD",x"35",x"16",x"C2",x"31",x"3B",x"3A",x"C8",x"80",x"DD",
		x"77",x"16",x"DD",x"7E",x"11",x"DD",x"77",x"17",x"CD",x"C9",x"00",x"3A",x"25",x"80",x"E6",x"03",
		x"DD",x"BE",x"10",x"28",x"F3",x"DD",x"BE",x"11",x"28",x"EE",x"DD",x"77",x"11",x"DD",x"36",x"0F",
		x"01",x"C9",x"3A",x"CC",x"80",x"3D",x"32",x"CC",x"80",x"C2",x"79",x"3B",x"3A",x"C6",x"80",x"32",
		x"CC",x"80",x"2A",x"C4",x"80",x"11",x"08",x"00",x"19",x"E5",x"11",x"00",x"02",x"B7",x"ED",x"52",
		x"E1",x"DA",x"55",x"3B",x"EB",x"22",x"C4",x"80",x"3A",x"4F",x"82",x"3D",x"32",x"4F",x"82",x"3A",
		x"C8",x"80",x"67",x"3A",x"C9",x"80",x"6F",x"7C",x"FE",x"18",x"D2",x"79",x"3B",x"11",x"20",x"00",
		x"19",x"7C",x"32",x"C8",x"80",x"7D",x"32",x"C9",x"80",x"C9",x"DD",x"35",x"0D",x"C2",x"AE",x"3B",
		x"DD",x"36",x"0D",x"06",x"21",x"CC",x"3E",x"DD",x"7E",x"11",x"FE",x"02",x"DA",x"92",x"3B",x"21",
		x"CF",x"3E",x"DD",x"7E",x"0E",x"01",x"01",x"00",x"CD",x"F6",x"00",x"7E",x"DD",x"77",x"02",x"DD",
		x"34",x"0E",x"DD",x"7E",x"0E",x"FE",x"03",x"DA",x"AE",x"3B",x"DD",x"36",x"0E",x"00",x"C9",x"DD",
		x"7E",x"04",x"C6",x"08",x"47",x"DD",x"7E",x"05",x"C6",x"14",x"4F",x"CD",x"DE",x"00",x"7E",x"CD",
		x"D6",x"5F",x"B7",x"C2",x"F3",x"3B",x"2A",x"D6",x"80",x"DD",x"75",x"16",x"DD",x"74",x"17",x"DD",
		x"36",x"08",x"00",x"DD",x"36",x"09",x"00",x"21",x"80",x"00",x"DD",x"75",x"0A",x"DD",x"74",x"0B",
		x"DD",x"36",x"10",x"00",x"DD",x"36",x"14",x"01",x"DD",x"36",x"01",x"04",x"3E",x"16",x"CD",x"FC",
		x"00",x"18",x"08",x"DD",x"36",x"14",x"06",x"DD",x"36",x"01",x"02",x"C9",x"DD",x"5E",x"10",x"16",
		x"00",x"21",x"11",x"3F",x"19",x"7E",x"DD",x"BE",x"11",x"C2",x"1C",x"3C",x"DD",x"7E",x"11",x"FE",
		x"02",x"D2",x"19",x"3C",x"DD",x"71",x"11",x"18",x"03",x"DD",x"70",x"11",x"C9",x"DD",x"7E",x"04",
		x"C6",x"08",x"E6",x"0F",x"11",x"88",x"3C",x"CD",x"6B",x"39",x"B7",x"20",x"54",x"DD",x"7E",x"05",
		x"C6",x"08",x"E6",x"0F",x"11",x"88",x"3C",x"CD",x"6B",x"39",x"B7",x"20",x"44",x"DD",x"7E",x"0C",
		x"B7",x"20",x"42",x"DD",x"36",x"0C",x"01",x"DD",x"7E",x"04",x"3C",x"E6",x"0F",x"FE",x"08",x"30",
		x"0D",x"3E",x"F0",x"DD",x"34",x"04",x"DD",x"A6",x"04",x"DD",x"77",x"04",x"18",x"04",x"3E",x"F8",
		x"18",x"F1",x"DD",x"7E",x"05",x"3C",x"E6",x"0F",x"FE",x"08",x"30",x"0D",x"3E",x"F0",x"DD",x"34",
		x"05",x"DD",x"A6",x"05",x"DD",x"77",x"05",x"18",x"04",x"3E",x"F8",x"18",x"F1",x"3E",x"00",x"18",
		x"06",x"DD",x"36",x"0C",x"00",x"3E",x"01",x"C9",x"0F",x"00",x"01",x"07",x"08",x"09",x"FF",x"3A",
		x"28",x"80",x"CB",x"7F",x"C2",x"C2",x"3C",x"DD",x"21",x"78",x"82",x"11",x"19",x"00",x"06",x"09",
		x"DD",x"7E",x"01",x"FE",x"0C",x"D2",x"C2",x"3C",x"DD",x"19",x"10",x"F4",x"3E",x"00",x"32",x"47",
		x"82",x"3A",x"4A",x"82",x"B7",x"CA",x"C7",x"3C",x"3A",x"4A",x"82",x"3D",x"32",x"4A",x"82",x"C3",
		x"C7",x"3C",x"3E",x"1E",x"32",x"4A",x"82",x"C9",x"2A",x"70",x"82",x"2B",x"22",x"70",x"82",x"7C",
		x"B5",x"C2",x"F3",x"3C",x"2A",x"5E",x"82",x"22",x"70",x"82",x"2A",x"5C",x"82",x"11",x"04",x"00",
		x"19",x"22",x"5C",x"82",x"01",x"40",x"04",x"B7",x"ED",x"42",x"DA",x"F3",x"3C",x"21",x"40",x"04",
		x"22",x"5C",x"82",x"2A",x"72",x"82",x"2B",x"22",x"72",x"82",x"7C",x"B5",x"C2",x"1C",x"3D",x"2A",
		x"62",x"82",x"22",x"72",x"82",x"2A",x"60",x"82",x"11",x"02",x"00",x"19",x"22",x"60",x"82",x"01",
		x"80",x"00",x"B7",x"ED",x"42",x"DA",x"1C",x"3D",x"ED",x"43",x"74",x"82",x"2A",x"74",x"82",x"2B",
		x"22",x"74",x"82",x"7C",x"B5",x"C2",x"43",x"3D",x"2A",x"66",x"82",x"22",x"74",x"82",x"3A",x"64",
		x"82",x"FE",x"0A",x"D2",x"3E",x"3D",x"C6",x"01",x"32",x"64",x"82",x"C3",x"43",x"3D",x"3E",x"0A",
		x"32",x"64",x"82",x"C9",x"2A",x"DC",x"80",x"2B",x"22",x"DC",x"80",x"7C",x"B5",x"C2",x"80",x"3D",
		x"2A",x"D8",x"80",x"22",x"DC",x"80",x"11",x"10",x"00",x"2A",x"D4",x"80",x"B7",x"ED",x"52",x"CA",
		x"65",x"3D",x"F2",x"68",x"3D",x"21",x"18",x"00",x"22",x"D4",x"80",x"2A",x"D6",x"80",x"11",x"10",
		x"00",x"B7",x"ED",x"52",x"CA",x"7A",x"3D",x"F2",x"7D",x"3D",x"21",x"01",x"00",x"22",x"D6",x"80",
		x"C9",x"21",x"78",x"82",x"11",x"19",x"00",x"06",x"09",x"BE",x"CA",x"93",x"3D",x"19",x"10",x"F9",
		x"AF",x"18",x"02",x"3E",x"01",x"B7",x"C9",x"0C",x"14",x"04",x"14",x"00",x"00",x"00",x"00",x"14",
		x"0C",x"FC",x"0C",x"00",x"00",x"00",x"00",x"10",x"14",x"00",x"14",x"10",x"FC",x"00",x"FC",x"1C",
		x"04",x"FC",x"04",x"0C",x"F4",x"0C",x"14",x"08",x"08",x"40",x"00",x"08",x"08",x"08",x"08",x"08",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0C",x"0C",x"0C",x"0C",x"48",
		x"48",x"30",x"A8",x"48",x"48",x"30",x"A8",x"30",x"60",x"30",x"A0",x"30",x"60",x"30",x"A0",x"48",
		x"30",x"60",x"A8",x"48",x"30",x"60",x"A8",x"48",x"48",x"48",x"C0",x"48",x"48",x"48",x"C0",x"48",
		x"48",x"48",x"A8",x"48",x"48",x"48",x"A8",x"30",x"30",x"30",x"C0",x"30",x"30",x"30",x"C0",x"60",
		x"48",x"60",x"A8",x"60",x"48",x"60",x"A8",x"30",x"30",x"30",x"C0",x"30",x"30",x"30",x"C0",x"30",
		x"48",x"30",x"90",x"30",x"48",x"30",x"90",x"30",x"48",x"30",x"A8",x"30",x"48",x"30",x"A8",x"48",
		x"60",x"48",x"A8",x"48",x"60",x"48",x"A8",x"48",x"30",x"48",x"C0",x"48",x"30",x"48",x"C0",x"30",
		x"60",x"30",x"A8",x"30",x"60",x"30",x"A8",x"18",x"60",x"78",x"A8",x"18",x"60",x"78",x"A8",x"48",
		x"30",x"30",x"C0",x"48",x"30",x"30",x"C0",x"18",x"60",x"18",x"A8",x"18",x"60",x"18",x"A8",x"18",
		x"D8",x"18",x"18",x"D8",x"18",x"D8",x"D8",x"00",x"02",x"03",x"01",x"01",x"03",x"02",x"00",x"02",
		x"01",x"00",x"03",x"03",x"00",x"01",x"02",x"04",x"05",x"04",x"05",x"06",x"07",x"08",x"07",x"09",
		x"0A",x"0B",x"0A",x"BC",x"BD",x"BE",x"BF",x"FF",x"00",x"30",x"2D",x"2F",x"FF",x"00",x"29",x"00",
		x"30",x"2D",x"2E",x"FF",x"00",x"2C",x"00",x"30",x"2D",x"2E",x"FF",x"00",x"2C",x"80",x"30",x"2D",
		x"2F",x"FF",x"80",x"29",x"80",x"30",x"2D",x"2E",x"FF",x"00",x"2C",x"80",x"30",x"2D",x"2E",x"FF",
		x"00",x"2C",x"80",x"2F",x"29",x"2A",x"FF",x"80",x"2B",x"00",x"2F",x"29",x"2A",x"FF",x"00",x"2B",
		x"00",x"2C",x"2D",x"2E",x"FF",x"00",x"2D",x"80",x"2F",x"29",x"2A",x"FF",x"80",x"2B",x"00",x"2F",
		x"29",x"2A",x"FF",x"00",x"2B",x"00",x"2C",x"2D",x"2E",x"FF",x"00",x"2D",x"29",x"2A",x"2B",x"2C",
		x"2D",x"2E",x"04",x"50",x"04",x"34",x"04",x"54",x"04",x"38",x"04",x"60",x"A0",x"A1",x"A2",x"A3",
		x"FF",x"00",x"01",x"02",x"03",x"04",x"05",x"80",x"81",x"82",x"83",x"90",x"91",x"92",x"93",x"FF",
		x"80",x"81",x"82",x"83",x"FF",x"60",x"61",x"62",x"63",x"66",x"67",x"68",x"69",x"6A",x"A0",x"A2",
		x"FF",x"00",x"01",x"00",x"02",x"00",x"03",x"00",x"05",x"00",x"08",x"00",x"12",x"00",x"20",x"00",
		x"00",x"01",x"00",x"03",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"FD",x"7E",x"03",x"C3",x"98",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"FD",x"7E",x"03",x"C3",x"D8",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"03",x"B0",x"3A",x"00",x"B0",x"E6",x"10",x"C2",x"39",x"05",x"2B",x"7C",x"B5",x"C3",x"2A",
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"21",x"CF",x"3D",x"C3",x"67",x"38",x"C3",x"81",x"31",x"C3",x"81",x"31",x"C3",x"81",x"31",x"00",
		x"CD",x"E4",x"42",x"06",x"00",x"3A",x"77",x"80",x"B7",x"CA",x"28",x"40",x"04",x"3A",x"74",x"80",
		x"B7",x"C2",x"28",x"40",x"04",x"3A",x"80",x"80",x"B7",x"C2",x"28",x"40",x"04",x"3A",x"9B",x"81",
		x"3D",x"32",x"9B",x"81",x"F2",x"28",x"40",x"04",x"78",x"21",x"2F",x"40",x"C3",x"EA",x"00",x"5C",
		x"40",x"AD",x"40",x"87",x"41",x"BA",x"41",x"75",x"42",x"E6",x"42",x"E6",x"42",x"CD",x"55",x"44",
		x"3E",x"00",x"32",x"4E",x"82",x"3E",x"00",x"32",x"4F",x"82",x"3E",x"00",x"32",x"49",x"82",x"3E",
		x"00",x"32",x"77",x"82",x"3E",x"01",x"32",x"03",x"80",x"C3",x"C0",x"00",x"CD",x"E8",x"42",x"CD",
		x"3D",x"43",x"3E",x"00",x"32",x"4B",x"82",x"3A",x"17",x"80",x"B7",x"CA",x"8C",x"40",x"3E",x"A0",
		x"CD",x"FC",x"00",x"AF",x"CD",x"D9",x"4B",x"CD",x"67",x"4B",x"3E",x"01",x"32",x"70",x"80",x"CD",
		x"FD",x"43",x"3E",x"00",x"32",x"70",x"80",x"CD",x"69",x"43",x"18",x"03",x"CD",x"CF",x"45",x"CD",
		x"95",x"44",x"CD",x"55",x"44",x"3E",x"00",x"32",x"81",x"80",x"3E",x"01",x"32",x"70",x"80",x"01",
		x"1E",x"00",x"CD",x"E1",x"00",x"3E",x"01",x"32",x"03",x"80",x"C3",x"C0",x"00",x"3E",x"00",x"32",
		x"28",x"80",x"32",x"77",x"80",x"32",x"74",x"80",x"32",x"88",x"80",x"00",x"CD",x"F8",x"5F",x"CD",
		x"30",x"60",x"3E",x"01",x"CD",x"FC",x"00",x"3E",x"25",x"CD",x"FC",x"00",x"3E",x"01",x"32",x"8D",
		x"80",x"01",x"F0",x"00",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"B7",x"C2",x"D9",x"40",
		x"C5",x"CD",x"33",x"60",x"CD",x"00",x"20",x"CD",x"10",x"30",x"C1",x"0B",x"78",x"B1",x"20",x"E4",
		x"21",x"48",x"0D",x"22",x"51",x"88",x"3E",x"00",x"32",x"8D",x"80",x"CD",x"20",x"4E",x"3E",x"00",
		x"32",x"AC",x"81",x"CD",x"67",x"4B",x"AF",x"CD",x"D9",x"4B",x"CD",x"F5",x"5F",x"CD",x"E0",x"2F",
		x"CD",x"E6",x"2F",x"CD",x"20",x"4E",x"21",x"A2",x"81",x"01",x"05",x"00",x"CD",x"CC",x"00",x"3E",
		x"00",x"32",x"AB",x"81",x"32",x"AC",x"81",x"32",x"B0",x"81",x"3A",x"A0",x"81",x"3C",x"32",x"A0",
		x"81",x"3A",x"A0",x"81",x"FE",x"41",x"DA",x"3E",x"41",x"3E",x"20",x"32",x"A0",x"81",x"3A",x"AF",
		x"81",x"FE",x"99",x"28",x"05",x"C6",x"01",x"27",x"18",x"02",x"3E",x"00",x"32",x"AF",x"81",x"3A",
		x"27",x"80",x"CD",x"40",x"44",x"3E",x"01",x"32",x"48",x"82",x"CD",x"CE",x"4E",x"CD",x"F4",x"4B",
		x"3E",x"18",x"32",x"A2",x"81",x"CD",x"0C",x"60",x"CD",x"E9",x"5F",x"CD",x"E8",x"42",x"CD",x"3D",
		x"43",x"CD",x"1F",x"44",x"C3",x"A0",x"4F",x"CD",x"E0",x"5F",x"3E",x"00",x"32",x"53",x"84",x"3E",
		x"01",x"32",x"54",x"84",x"C3",x"3D",x"40",x"3E",x"00",x"32",x"77",x"80",x"3E",x"00",x"32",x"80",
		x"80",x"3E",x"00",x"32",x"88",x"80",x"3E",x"00",x"32",x"8E",x"80",x"CD",x"20",x"4E",x"AF",x"CD",
		x"D9",x"4B",x"CD",x"F0",x"00",x"DD",x"21",x"4A",x"D2",x"CD",x"D2",x"00",x"3E",x"0D",x"CD",x"18",
		x"60",x"CD",x"FB",x"5F",x"CD",x"F8",x"5F",x"C3",x"F0",x"40",x"3E",x"00",x"32",x"77",x"80",x"3E",
		x"00",x"32",x"88",x"80",x"3E",x"00",x"32",x"95",x"80",x"3A",x"28",x"80",x"CB",x"97",x"32",x"28",
		x"80",x"3E",x"01",x"32",x"8D",x"80",x"06",x"7E",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",
		x"B7",x"C2",x"DD",x"41",x"C5",x"CD",x"00",x"20",x"CD",x"10",x"30",x"C1",x"78",x"FE",x"78",x"C2",
		x"F7",x"41",x"3E",x"01",x"CD",x"FC",x"00",x"10",x"DF",x"21",x"48",x"0D",x"22",x"51",x"88",x"3E",
		x"00",x"32",x"8D",x"80",x"3E",x"00",x"CD",x"D9",x"4B",x"CD",x"67",x"4B",x"3E",x"00",x"32",x"B0",
		x"81",x"CD",x"20",x"4E",x"CD",x"EF",x"5F",x"3A",x"27",x"80",x"CD",x"40",x"44",x"CD",x"87",x"45",
		x"3A",x"27",x"80",x"CD",x"2B",x"44",x"3A",x"AC",x"81",x"FE",x"00",x"28",x"05",x"CD",x"E3",x"2F",
		x"18",x"03",x"CD",x"E0",x"2F",x"CD",x"E6",x"2F",x"CD",x"0C",x"60",x"CD",x"EC",x"5F",x"3E",x"00",
		x"32",x"48",x"82",x"CD",x"CE",x"4E",x"CD",x"20",x"4E",x"CD",x"F4",x"4B",x"CD",x"E6",x"2F",x"CD",
		x"E9",x"5F",x"CD",x"E8",x"42",x"CD",x"1F",x"44",x"CD",x"C9",x"47",x"3A",x"9B",x"81",x"3C",x"32",
		x"9B",x"81",x"CD",x"3D",x"43",x"CD",x"E0",x"5F",x"3A",x"9B",x"81",x"3D",x"32",x"9B",x"81",x"CD",
		x"3D",x"43",x"C3",x"3D",x"40",x"3E",x"00",x"32",x"77",x"80",x"3E",x"00",x"32",x"88",x"80",x"3E",
		x"00",x"32",x"8D",x"80",x"3E",x"00",x"32",x"4B",x"82",x"3E",x"01",x"CD",x"FC",x"00",x"3E",x"26",
		x"CD",x"FC",x"00",x"3E",x"01",x"CD",x"D9",x"4B",x"3A",x"27",x"80",x"CD",x"40",x"44",x"CD",x"E3",
		x"5F",x"CD",x"20",x"4E",x"CD",x"67",x"4B",x"CD",x"00",x"48",x"3E",x"01",x"CD",x"FC",x"00",x"CD",
		x"20",x"4E",x"3A",x"8B",x"80",x"B7",x"C2",x"D3",x"42",x"3A",x"26",x"80",x"B7",x"CA",x"D3",x"42",
		x"3A",x"27",x"80",x"B7",x"C2",x"CC",x"42",x"3A",x"CD",x"81",x"18",x"03",x"3A",x"B4",x"81",x"B7",
		x"F2",x"11",x"42",x"CD",x"39",x"4B",x"3E",x"00",x"32",x"70",x"80",x"3E",x"01",x"32",x"03",x"80",
		x"C3",x"C6",x"00",x"C9",x"00",x"C9",x"00",x"C9",x"3A",x"70",x"80",x"B7",x"CA",x"14",x"43",x"3A",
		x"27",x"80",x"B7",x"CA",x"FE",x"42",x"CD",x"CF",x"00",x"91",x"CA",x"03",x"18",x"2A",x"3A",x"26",
		x"80",x"B7",x"20",x"08",x"CD",x"CF",x"00",x"89",x"CA",x"04",x"18",x"1C",x"CD",x"CF",x"00",x"83",
		x"CA",x"03",x"18",x"14",x"3A",x"26",x"80",x"B7",x"20",x"08",x"CD",x"CF",x"00",x"6D",x"CA",x"04",
		x"18",x"06",x"CD",x"CF",x"00",x"67",x"CA",x"03",x"3A",x"26",x"80",x"B7",x"20",x"08",x"CD",x"D8",
		x"00",x"7B",x"CA",x"02",x"18",x"06",x"CD",x"D8",x"00",x"75",x"CA",x"03",x"C9",x"CD",x"AC",x"44",
		x"DD",x"21",x"A7",x"CA",x"CD",x"D2",x"00",x"DD",x"21",x"C1",x"CA",x"CD",x"D5",x"00",x"DD",x"21",
		x"C7",x"CA",x"3A",x"AF",x"81",x"FE",x"10",x"DA",x"5E",x"43",x"DD",x"21",x"CF",x"CA",x"CD",x"D2",
		x"00",x"DD",x"21",x"D5",x"CA",x"CD",x"D2",x"00",x"C9",x"CD",x"E8",x"42",x"CD",x"3D",x"43",x"CD",
		x"E0",x"2F",x"CD",x"20",x"4E",x"3A",x"17",x"80",x"B7",x"CA",x"C8",x"43",x"3A",x"8B",x"80",x"B7",
		x"C2",x"8B",x"43",x"CD",x"DF",x"4C",x"3E",x"01",x"32",x"81",x"80",x"CD",x"0B",x"45",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"01",x"32",x"70",x"80",
		x"CD",x"20",x"4E",x"CD",x"2A",x"60",x"21",x"B4",x"81",x"01",x"32",x"00",x"CD",x"CC",x"00",x"CD",
		x"CC",x"43",x"AF",x"CD",x"40",x"44",x"3E",x"01",x"CD",x"40",x"44",x"3E",x"00",x"32",x"E5",x"81",
		x"3A",x"CD",x"81",x"32",x"75",x"80",x"18",x"03",x"CD",x"CC",x"43",x"C9",x"CD",x"20",x"4E",x"3E",
		x"00",x"32",x"48",x"82",x"CD",x"CE",x"4E",x"CD",x"F4",x"4B",x"CD",x"0C",x"60",x"CD",x"E9",x"5F",
		x"CD",x"C9",x"47",x"3A",x"17",x"80",x"B7",x"28",x"00",x"CD",x"E8",x"42",x"3A",x"9B",x"81",x"3D",
		x"32",x"9B",x"81",x"CD",x"1F",x"44",x"CD",x"E0",x"5F",x"CD",x"3D",x"43",x"C9",x"21",x"9B",x"81",
		x"01",x"19",x"00",x"CD",x"CC",x"00",x"3A",x"71",x"80",x"32",x"9B",x"81",x"3E",x"01",x"32",x"A0",
		x"81",x"3E",x"18",x"32",x"A2",x"81",x"3E",x"01",x"32",x"AF",x"81",x"CD",x"15",x"60",x"C9",x"CD",
		x"E7",x"00",x"CD",x"27",x"4E",x"3E",x"01",x"32",x"8C",x"80",x"C9",x"B7",x"C2",x"34",x"44",x"21",
		x"B4",x"81",x"18",x"03",x"21",x"CD",x"81",x"11",x"9B",x"81",x"01",x"19",x"00",x"ED",x"B0",x"C9",
		x"B7",x"C2",x"49",x"44",x"11",x"B4",x"81",x"18",x"03",x"11",x"CD",x"81",x"21",x"9B",x"81",x"01",
		x"19",x"00",x"ED",x"B0",x"C9",x"DD",x"21",x"28",x"80",x"DD",x"36",x"00",x"00",x"DD",x"36",x"01",
		x"18",x"DD",x"36",x"02",x"00",x"DD",x"36",x"03",x"78",x"DD",x"36",x"04",x"78",x"DD",x"36",x"05",
		x"00",x"DD",x"36",x"06",x"00",x"DD",x"36",x"09",x"80",x"DD",x"36",x"0B",x"FF",x"DD",x"36",x"0E",
		x"00",x"DD",x"36",x"0E",x"00",x"DD",x"36",x"12",x"FF",x"21",x"29",x"80",x"01",x"04",x"00",x"11",
		x"00",x"85",x"ED",x"B0",x"C9",x"3E",x"00",x"32",x"53",x"84",x"3E",x"01",x"32",x"54",x"84",x"21",
		x"E0",x"00",x"22",x"5B",x"84",x"21",x"E0",x"FE",x"22",x"5D",x"84",x"C9",x"3A",x"9B",x"81",x"B7",
		x"CA",x"D3",x"44",x"FE",x"01",x"CA",x"DA",x"44",x"FE",x"02",x"CA",x"E1",x"44",x"FE",x"03",x"CA",
		x"E8",x"44",x"FE",x"04",x"CA",x"EF",x"44",x"FE",x"05",x"CA",x"F6",x"44",x"FE",x"06",x"CA",x"FD",
		x"44",x"18",x"31",x"CD",x"CF",x"00",x"DB",x"CA",x"02",x"C9",x"CD",x"CF",x"00",x"DF",x"CA",x"02",
		x"C9",x"CD",x"CF",x"00",x"E3",x"CA",x"02",x"C9",x"CD",x"CF",x"00",x"E7",x"CA",x"02",x"C9",x"CD",
		x"CF",x"00",x"EB",x"CA",x"02",x"C9",x"CD",x"CF",x"00",x"EF",x"CA",x"02",x"C9",x"CD",x"CF",x"00",
		x"F3",x"CA",x"02",x"C9",x"CD",x"CF",x"00",x"F7",x"CA",x"02",x"C9",x"3E",x"02",x"32",x"8C",x"80",
		x"3A",x"8B",x"80",x"F5",x"3E",x"00",x"32",x"8B",x"80",x"F1",x"FE",x"02",x"CA",x"3E",x"45",x"FE",
		x"01",x"CA",x"68",x"45",x"3A",x"02",x"B0",x"E6",x"08",x"C2",x"36",x"45",x"3A",x"02",x"B0",x"E6",
		x"04",x"C2",x"68",x"45",x"18",x"D5",x"3A",x"17",x"80",x"FE",x"02",x"DA",x"0B",x"45",x"3E",x"01",
		x"32",x"26",x"80",x"3A",x"87",x"80",x"B7",x"CA",x"5D",x"45",x"3A",x"87",x"80",x"3D",x"32",x"87",
		x"80",x"CA",x"7D",x"45",x"3A",x"87",x"80",x"3D",x"32",x"87",x"80",x"18",x"29",x"3A",x"17",x"80",
		x"C6",x"98",x"27",x"32",x"17",x"80",x"18",x"1E",x"3E",x"00",x"32",x"26",x"80",x"3A",x"87",x"80",
		x"B7",x"CA",x"7D",x"45",x"3A",x"87",x"80",x"3D",x"32",x"87",x"80",x"18",x"09",x"3A",x"17",x"80",
		x"C6",x"99",x"27",x"32",x"17",x"80",x"C9",x"3A",x"26",x"80",x"B7",x"CA",x"CE",x"45",x"3A",x"75",
		x"80",x"B7",x"FA",x"CE",x"45",x"3A",x"27",x"80",x"3C",x"E6",x"01",x"32",x"27",x"80",x"3A",x"13",
		x"80",x"E6",x"40",x"C2",x"B9",x"45",x"3A",x"27",x"80",x"B7",x"CA",x"B4",x"45",x"3E",x"01",x"32",
		x"04",x"B0",x"18",x"05",x"3E",x"00",x"32",x"04",x"B0",x"3A",x"27",x"80",x"B7",x"C2",x"C8",x"45",
		x"3A",x"CD",x"81",x"32",x"75",x"80",x"18",x"06",x"3A",x"B4",x"81",x"32",x"75",x"80",x"C9",x"3E",
		x"00",x"32",x"88",x"80",x"3E",x"00",x"32",x"8D",x"80",x"3E",x"01",x"CD",x"FC",x"00",x"CD",x"20",
		x"4E",x"AF",x"CD",x"D9",x"4B",x"CD",x"E4",x"42",x"CD",x"67",x"4B",x"3A",x"AB",x"81",x"F5",x"CD",
		x"FD",x"43",x"F1",x"32",x"AB",x"81",x"CD",x"3D",x"43",x"3A",x"79",x"80",x"21",x"22",x"46",x"CD",
		x"EA",x"00",x"3A",x"79",x"80",x"3C",x"32",x"79",x"80",x"3A",x"79",x"80",x"FE",x"04",x"DA",x"16",
		x"46",x"3E",x"00",x"32",x"79",x"80",x"3E",x"00",x"32",x"78",x"80",x"3E",x"00",x"32",x"4B",x"82",
		x"18",x"AD",x"32",x"46",x"5A",x"46",x"50",x"47",x"C5",x"46",x"E6",x"42",x"E6",x"42",x"E6",x"42",
		x"E6",x"42",x"CD",x"CF",x"00",x"00",x"C0",x"0C",x"00",x"CD",x"D8",x"00",x"96",x"C1",x"0A",x"CD",
		x"CF",x"00",x"E6",x"C1",x"0A",x"CD",x"D8",x"00",x"FA",x"C1",x"0A",x"CD",x"9B",x"47",x"3E",x"0D",
		x"CD",x"18",x"60",x"01",x"2C",x"01",x"CD",x"E1",x"00",x"C9",x"CD",x"FD",x"43",x"CD",x"69",x"43",
		x"CD",x"95",x"44",x"CD",x"55",x"44",x"3E",x"00",x"32",x"7A",x"80",x"3E",x"00",x"32",x"7B",x"80",
		x"3A",x"E8",x"80",x"FE",x"00",x"20",x"05",x"2A",x"F8",x"CD",x"18",x"03",x"2A",x"FA",x"CD",x"22",
		x"7C",x"80",x"22",x"7E",x"80",x"01",x"1E",x"00",x"CD",x"E1",x"00",x"18",x"00",x"21",x"01",x"00",
		x"22",x"6E",x"80",x"CD",x"59",x"47",x"CD",x"00",x"10",x"3A",x"6E",x"80",x"B7",x"28",x"EE",x"CD",
		x"00",x"20",x"3A",x"6E",x"80",x"B7",x"28",x"E5",x"CD",x"00",x"30",x"3A",x"6E",x"80",x"B7",x"28",
		x"DC",x"CD",x"00",x"50",x"3A",x"78",x"80",x"B7",x"C2",x"C4",x"46",x"3A",x"6E",x"80",x"B7",x"CA",
		x"8D",x"46",x"18",x"F7",x"C9",x"3A",x"AB",x"81",x"FE",x"17",x"20",x"11",x"3E",x"3C",x"32",x"B3",
		x"81",x"21",x"E0",x"00",x"22",x"5B",x"84",x"21",x"E0",x"FE",x"22",x"5D",x"84",x"3E",x"00",x"32",
		x"AB",x"81",x"3E",x"02",x"32",x"A0",x"81",x"3E",x"18",x"32",x"A2",x"81",x"3E",x"02",x"32",x"AF",
		x"81",x"3A",x"71",x"80",x"32",x"9B",x"81",x"3A",x"E8",x"80",x"FE",x"00",x"20",x"0A",x"2A",x"FC",
		x"CD",x"3E",x"01",x"32",x"E8",x"80",x"18",x"08",x"2A",x"FE",x"CD",x"3E",x"00",x"32",x"E8",x"80",
		x"22",x"7C",x"80",x"22",x"7E",x"80",x"3E",x"01",x"32",x"48",x"82",x"3E",x"00",x"32",x"A7",x"81",
		x"18",x"00",x"CD",x"E0",x"2F",x"CD",x"CE",x"4E",x"CD",x"F4",x"4B",x"CD",x"0C",x"60",x"CD",x"E9",
		x"5F",x"3E",x"00",x"32",x"7A",x"80",x"3E",x"00",x"32",x"7B",x"80",x"CD",x"3D",x"43",x"CD",x"E8",
		x"42",x"CD",x"1F",x"44",x"CD",x"C9",x"47",x"CD",x"E0",x"5F",x"CD",x"55",x"44",x"C3",x"8D",x"46",
		x"3E",x"0D",x"CD",x"18",x"60",x"CD",x"21",x"60",x"C9",x"DD",x"21",x"7A",x"80",x"DD",x"7E",x"01",
		x"FE",x"00",x"C2",x"97",x"47",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"7E",x"DD",x"77",x"01",x"FE",
		x"FF",x"C2",x"8A",x"47",x"DD",x"36",x"00",x"00",x"DD",x"36",x"01",x"01",x"DD",x"7E",x"04",x"DD",
		x"77",x"02",x"DD",x"7E",x"05",x"DD",x"77",x"03",x"18",x"0C",x"23",x"7E",x"DD",x"77",x"00",x"23",
		x"DD",x"75",x"02",x"DD",x"74",x"03",x"C9",x"DD",x"35",x"01",x"C9",x"21",x"28",x"81",x"DD",x"21",
		x"87",x"94",x"06",x"0A",x"4E",x"DD",x"22",x"E6",x"80",x"7E",x"B9",x"38",x"07",x"28",x"05",x"DD",
		x"22",x"E6",x"80",x"4F",x"23",x"DD",x"23",x"DD",x"23",x"10",x"EE",x"2A",x"E6",x"80",x"36",x"0F",
		x"B7",x"11",x"20",x"00",x"ED",x"52",x"36",x"0F",x"C9",x"3E",x"21",x"CD",x"FC",x"00",x"21",x"3D",
		x"DE",x"01",x"06",x"00",x"3A",x"A0",x"81",x"CD",x"F6",x"00",x"7E",x"C6",x"22",x"CD",x"FC",x"00",
		x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"DD",x"21",x"00",x"81",x"06",x"0A",x"0E",x"00",x"FD",x"21",x"9C",x"81",x"FD",x"7E",x"03",x"DD",
		x"96",x"03",x"38",x"22",x"20",x"2D",x"FD",x"7E",x"02",x"DD",x"96",x"02",x"38",x"18",x"20",x"23",
		x"FD",x"7E",x"01",x"DD",x"96",x"01",x"38",x"0E",x"20",x"19",x"FD",x"7E",x"00",x"DD",x"96",x"00",
		x"38",x"04",x"28",x"02",x"18",x"0D",x"DD",x"23",x"DD",x"23",x"DD",x"23",x"DD",x"23",x"0C",x"10",
		x"CB",x"18",x"07",x"79",x"32",x"96",x"81",x"CD",x"4B",x"48",x"C9",x"CD",x"20",x"4E",x"21",x"00",
		x"85",x"01",x"60",x"00",x"CD",x"CC",x"00",x"CD",x"FC",x"48",x"CD",x"7C",x"49",x"CD",x"20",x"4B",
		x"3E",x"A6",x"CD",x"FC",x"00",x"3A",x"96",x"81",x"B7",x"C2",x"79",x"48",x"3E",x"29",x"CD",x"FC",
		x"00",x"3E",x"0D",x"CD",x"18",x"60",x"C3",x"83",x"48",x"3E",x"2A",x"CD",x"FC",x"00",x"3E",x"0D",
		x"CD",x"18",x"60",x"CD",x"9B",x"47",x"2A",x"E6",x"80",x"E5",x"DD",x"E1",x"DD",x"36",x"00",x"02",
		x"DD",x"36",x"E0",x"02",x"DD",x"21",x"87",x"96",x"DD",x"36",x"A0",x"02",x"DD",x"36",x"C0",x"02",
		x"DD",x"36",x"E0",x"02",x"DD",x"36",x"00",x"02",x"DD",x"36",x"20",x"02",x"DD",x"36",x"40",x"02",
		x"DD",x"36",x"60",x"02",x"DD",x"36",x"80",x"02",x"DD",x"21",x"1C",x"96",x"DD",x"36",x"80",x"01",
		x"DD",x"36",x"A0",x"01",x"DD",x"36",x"C0",x"01",x"DD",x"36",x"E0",x"01",x"DD",x"36",x"00",x"01",
		x"DD",x"36",x"20",x"01",x"3A",x"96",x"81",x"DD",x"21",x"07",x"94",x"FE",x"00",x"28",x"07",x"DD",
		x"23",x"DD",x"23",x"3D",x"18",x"F5",x"3E",x"20",x"11",x"20",x"00",x"FE",x"00",x"28",x"09",x"DD",
		x"36",x"00",x"0F",x"DD",x"19",x"3D",x"18",x"F3",x"CD",x"93",x"49",x"C9",x"3A",x"96",x"81",x"21",
		x"31",x"81",x"11",x"30",x"81",x"F5",x"47",x"3E",x"09",x"90",x"47",x"B7",x"28",x"06",x"1A",x"77",
		x"2B",x"1B",x"10",x"FA",x"3A",x"AF",x"81",x"77",x"F1",x"F5",x"47",x"3E",x"09",x"90",x"47",x"B7",
		x"28",x"41",x"21",x"20",x"81",x"11",x"24",x"81",x"0E",x"04",x"7E",x"12",x"23",x"13",x"0D",x"20",
		x"F9",x"C5",x"01",x"F8",x"FF",x"09",x"E5",x"EB",x"09",x"EB",x"E1",x"C1",x"10",x"EA",x"F1",x"F5",
		x"47",x"3E",x"09",x"90",x"47",x"21",x"84",x"81",x"11",x"8E",x"81",x"0E",x"03",x"7E",x"12",x"23",
		x"23",x"13",x"13",x"0D",x"20",x"F7",x"C5",x"01",x"F0",x"FF",x"09",x"E5",x"EB",x"09",x"EB",x"E1",
		x"C1",x"10",x"E8",x"F1",x"47",x"00",x"21",x"FC",x"80",x"11",x"04",x"00",x"04",x"19",x"10",x"FD",
		x"11",x"9C",x"81",x"06",x"04",x"1A",x"77",x"13",x"23",x"10",x"FA",x"C9",x"3A",x"96",x"81",x"3C",
		x"21",x"2A",x"81",x"11",x"0A",x"00",x"19",x"3D",x"20",x"FC",x"06",x"03",x"36",x"00",x"23",x"23",
		x"10",x"FA",x"C9",x"01",x"10",x"0E",x"ED",x"43",x"6E",x"80",x"3E",x"01",x"32",x"97",x"81",x"CD",
		x"41",x"4A",x"CD",x"CD",x"4A",x"CD",x"B4",x"4A",x"36",x"41",x"CD",x"CD",x"4A",x"3A",x"1B",x"80",
		x"CB",x"67",x"C2",x"05",x"4A",x"3A",x"19",x"80",x"CB",x"67",x"C2",x"DE",x"49",x"3A",x"20",x"80",
		x"FE",x"03",x"28",x"69",x"CD",x"83",x"4E",x"B7",x"C2",x"DD",x"49",x"ED",x"4B",x"6E",x"80",x"79",
		x"B0",x"20",x"DA",x"AF",x"CD",x"41",x"4A",x"01",x"B4",x"00",x"CD",x"E1",x"00",x"C9",x"3E",x"00",
		x"32",x"19",x"80",x"CD",x"B4",x"4A",x"7E",x"FE",x"00",x"20",x"04",x"36",x"41",x"18",x"11",x"FE",
		x"5A",x"20",x"04",x"36",x"2E",x"18",x"09",x"FE",x"2E",x"20",x"04",x"36",x"00",x"18",x"01",x"34",
		x"CD",x"CD",x"4A",x"18",x"BF",x"3E",x"00",x"32",x"1B",x"80",x"CD",x"B4",x"4A",x"7E",x"FE",x"00",
		x"20",x"04",x"36",x"2E",x"18",x"11",x"FE",x"41",x"20",x"04",x"36",x"00",x"18",x"09",x"FE",x"2E",
		x"20",x"04",x"36",x"5A",x"18",x"01",x"35",x"CD",x"CD",x"4A",x"C3",x"C4",x"49",x"3C",x"3C",x"32",
		x"20",x"80",x"3A",x"97",x"81",x"3C",x"FE",x"04",x"32",x"97",x"81",x"DA",x"A5",x"49",x"D2",x"D3",
		x"49",x"F5",x"11",x"00",x"00",x"21",x"82",x"4A",x"3A",x"96",x"81",x"87",x"5F",x"19",x"5E",x"23",
		x"56",x"EB",x"F1",x"11",x"96",x"4A",x"B7",x"28",x"03",x"11",x"A5",x"4A",x"06",x"05",x"0E",x"03",
		x"D5",x"E5",x"1A",x"FE",x"FF",x"28",x"01",x"77",x"FE",x"00",x"28",x"06",x"11",x"00",x"04",x"19",
		x"36",x"0F",x"E1",x"D1",x"23",x"13",x"0D",x"20",x"E7",x"D5",x"11",x"1D",x"00",x"19",x"D1",x"10",
		x"DD",x"C9",x"66",x"91",x"68",x"91",x"6A",x"91",x"6C",x"91",x"6E",x"91",x"70",x"91",x"72",x"91",
		x"74",x"91",x"76",x"91",x"78",x"91",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",
		x"FF",x"00",x"00",x"00",x"00",x"F2",x"F4",x"F7",x"F1",x"00",x"F6",x"F1",x"00",x"F6",x"F1",x"00",
		x"F6",x"F0",x"F3",x"F5",x"3A",x"96",x"81",x"21",x"32",x"81",x"11",x"0A",x"00",x"B7",x"28",x"04",
		x"19",x"3D",x"18",x"F9",x"3A",x"97",x"81",x"87",x"16",x"00",x"5F",x"19",x"C9",x"3A",x"96",x"81",
		x"21",x"32",x"81",x"11",x"0A",x"00",x"B7",x"28",x"05",x"19",x"3D",x"C3",x"D6",x"4A",x"E5",x"DD",
		x"E1",x"DD",x"7E",x"03",x"F5",x"DD",x"7E",x"05",x"F5",x"DD",x"7E",x"07",x"F5",x"DD",x"36",x"03",
		x"06",x"DD",x"36",x"05",x"06",x"DD",x"36",x"07",x"06",x"3A",x"97",x"81",x"FE",x"03",x"28",x"0C",
		x"FE",x"02",x"28",x"04",x"DD",x"36",x"03",x"03",x"DD",x"36",x"05",x"03",x"DD",x"36",x"07",x"03",
		x"CD",x"D2",x"00",x"F1",x"DD",x"77",x"07",x"F1",x"DD",x"77",x"05",x"F1",x"DD",x"77",x"03",x"C9",
		x"CD",x"CF",x"00",x"4A",x"C2",x"0D",x"CD",x"D8",x"00",x"96",x"C1",x"0A",x"CD",x"CF",x"00",x"E6",
		x"C1",x"0A",x"CD",x"D8",x"00",x"FA",x"C1",x"0A",x"C9",x"CD",x"67",x"4B",x"21",x"9B",x"81",x"01",
		x"19",x"00",x"CD",x"CC",x"00",x"21",x"B9",x"81",x"01",x"14",x"00",x"CD",x"CC",x"00",x"21",x"D2",
		x"81",x"01",x"14",x"00",x"CD",x"CC",x"00",x"3E",x"00",x"32",x"79",x"80",x"3E",x"00",x"32",x"04",
		x"B0",x"3E",x"00",x"32",x"27",x"80",x"C9",x"2A",x"5B",x"84",x"E5",x"2A",x"5D",x"84",x"E5",x"21",
		x"28",x"80",x"01",x"46",x"00",x"CD",x"CC",x"00",x"21",x"78",x"82",x"01",x"F4",x"01",x"CD",x"CC",
		x"00",x"21",x"D2",x"80",x"01",x"10",x"00",x"CD",x"CC",x"00",x"21",x"C0",x"80",x"01",x"12",x"00",
		x"CD",x"CC",x"00",x"21",x"00",x"89",x"01",x"14",x"00",x"CD",x"CC",x"00",x"E1",x"22",x"5D",x"84",
		x"E1",x"22",x"5B",x"84",x"C9",x"21",x"00",x"90",x"01",x"00",x"04",x"36",x"00",x"23",x"0B",x"78",
		x"B1",x"C2",x"AB",x"4B",x"21",x"00",x"98",x"01",x"00",x"04",x"36",x"00",x"23",x"0B",x"78",x"B1",
		x"C2",x"BA",x"4B",x"C9",x"F5",x"C5",x"E5",x"21",x"28",x"80",x"01",x"20",x"00",x"36",x"00",x"23",
		x"0B",x"78",x"B1",x"20",x"F8",x"E1",x"C1",x"F1",x"C9",x"C5",x"E5",x"B7",x"CA",x"E7",x"4B",x"21",
		x"08",x"85",x"06",x"58",x"C3",x"EC",x"4B",x"21",x"00",x"85",x"06",x"60",x"36",x"00",x"23",x"10",
		x"FB",x"E1",x"C1",x"C9",x"3E",x"01",x"32",x"8F",x"80",x"3A",x"A0",x"81",x"3D",x"01",x"06",x"00",
		x"21",x"38",x"DE",x"CD",x"F6",x"00",x"7E",x"32",x"A1",x"81",x"21",x"74",x"7C",x"CD",x"EA",x"00",
		x"3E",x"00",x"32",x"8F",x"80",x"21",x"3A",x"DE",x"01",x"06",x"00",x"3A",x"A0",x"81",x"3D",x"CD",
		x"F6",x"00",x"7E",x"E6",x"07",x"CD",x"18",x"60",x"C9",x"C5",x"D5",x"E5",x"57",x"3E",x"01",x"32",
		x"8F",x"80",x"1E",x"66",x"CD",x"D3",x"5F",x"06",x"0D",x"21",x"43",x"90",x"73",x"23",x"73",x"34",
		x"23",x"10",x"F9",x"21",x"A3",x"93",x"06",x"0D",x"73",x"23",x"73",x"34",x"23",x"10",x"F9",x"7A",
		x"21",x"43",x"94",x"06",x"1A",x"4F",x"77",x"23",x"10",x"FC",x"21",x"A3",x"97",x"06",x"1A",x"79",
		x"77",x"23",x"10",x"FC",x"11",x"80",x"87",x"21",x"A3",x"4C",x"01",x"3C",x"00",x"ED",x"B0",x"4F",
		x"CD",x"98",x"4C",x"DD",x"21",x"80",x"87",x"CD",x"D2",x"00",x"3E",x"1D",x"32",x"80",x"87",x"3E",
		x"6A",x"32",x"82",x"87",x"3E",x"6B",x"32",x"B8",x"87",x"79",x"CD",x"98",x"4C",x"DD",x"21",x"80",
		x"87",x"CD",x"D2",x"00",x"E1",x"D1",x"C1",x"C9",x"06",x"1C",x"21",x"83",x"87",x"77",x"23",x"23",
		x"10",x"FB",x"C9",x"02",x"02",x"68",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",
		x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",
		x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",
		x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"62",x"01",x"63",x"01",x"69",x"01",x"FF",x"FF",x"3E",
		x"0D",x"CD",x"18",x"60",x"CD",x"27",x"60",x"CD",x"24",x"60",x"CD",x"CF",x"00",x"00",x"D0",x"04",
		x"DD",x"21",x"14",x"D0",x"3A",x"17",x"80",x"FE",x"01",x"CA",x"00",x"4D",x"DD",x"21",x"40",x"D0",
		x"CD",x"D2",x"00",x"CD",x"F0",x"00",x"C3",x"63",x"4D",x"E6",x"07",x"21",x"11",x"4D",x"C3",x"EA",
		x"00",x"21",x"4D",x"24",x"4D",x"2D",x"4D",x"36",x"4D",x"3F",x"4D",x"48",x"4D",x"51",x"4D",x"5A",
		x"4D",x"C3",x"68",x"4D",x"CD",x"CF",x"00",x"AA",x"D0",x"02",x"C3",x"68",x"4D",x"CD",x"CF",x"00",
		x"AE",x"D0",x"02",x"C3",x"68",x"4D",x"CD",x"CF",x"00",x"B2",x"D0",x"02",x"C3",x"68",x"4D",x"CD",
		x"CF",x"00",x"B6",x"D0",x"02",x"C3",x"68",x"4D",x"CD",x"CF",x"00",x"BA",x"D0",x"04",x"C3",x"68",
		x"4D",x"CD",x"CF",x"00",x"C2",x"D0",x"04",x"C3",x"68",x"4D",x"CD",x"CF",x"00",x"CA",x"D0",x"06",
		x"C3",x"68",x"4D",x"3E",x"0D",x"CD",x"18",x"60",x"C9",x"3A",x"70",x"80",x"FE",x"00",x"28",x"08",
		x"3A",x"14",x"80",x"E6",x"18",x"0F",x"0F",x"0F",x"21",x"7E",x"4D",x"C3",x"EA",x"00",x"86",x"4D",
		x"90",x"4D",x"9B",x"4D",x"A6",x"4D",x"3A",x"A8",x"81",x"3C",x"32",x"A8",x"81",x"C3",x"B1",x"4D",
		x"3A",x"A8",x"81",x"C6",x"02",x"32",x"A8",x"81",x"C3",x"B1",x"4D",x"3A",x"A8",x"81",x"C6",x"04",
		x"32",x"A8",x"81",x"C3",x"B1",x"4D",x"3A",x"A8",x"81",x"C6",x"08",x"32",x"A8",x"81",x"C3",x"B1",
		x"4D",x"3A",x"A8",x"81",x"FE",x"20",x"DA",x"BE",x"4D",x"3E",x"1F",x"32",x"A8",x"81",x"C9",x"3A",
		x"70",x"80",x"FE",x"00",x"28",x"08",x"3A",x"14",x"80",x"E6",x"60",x"07",x"07",x"07",x"21",x"D4",
		x"4D",x"C3",x"EA",x"00",x"DC",x"4D",x"E6",x"4D",x"FC",x"4D",x"07",x"4E",x"3A",x"A9",x"81",x"3C",
		x"32",x"A9",x"81",x"C3",x"12",x"4E",x"3A",x"AA",x"81",x"3C",x"E6",x"01",x"32",x"AA",x"81",x"C2",
		x"12",x"4E",x"3A",x"A9",x"81",x"3C",x"32",x"A9",x"81",x"C3",x"12",x"4E",x"3A",x"A9",x"81",x"C6",
		x"02",x"32",x"A9",x"81",x"C3",x"12",x"4E",x"3A",x"A9",x"81",x"C6",x"04",x"32",x"A9",x"81",x"C3",
		x"12",x"4E",x"3A",x"A9",x"81",x"FE",x"20",x"DA",x"1F",x"4E",x"3E",x"13",x"32",x"A9",x"81",x"C9",
		x"01",x"1C",x"02",x"CD",x"ED",x"00",x"C9",x"21",x"39",x"DE",x"01",x"06",x"00",x"3A",x"A0",x"81",
		x"3D",x"CD",x"F6",x"00",x"23",x"7E",x"F5",x"2B",x"7E",x"21",x"00",x"D6",x"01",x"10",x"00",x"CD",
		x"F6",x"00",x"11",x"90",x"8C",x"ED",x"B0",x"F1",x"F5",x"21",x"00",x"D7",x"01",x"10",x"00",x"CD",
		x"F6",x"00",x"11",x"A0",x"8C",x"ED",x"B0",x"F1",x"21",x"80",x"D7",x"01",x"10",x"00",x"CD",x"F6",
		x"00",x"11",x"80",x"8C",x"ED",x"B0",x"21",x"3C",x"DE",x"01",x"06",x"00",x"3A",x"A0",x"81",x"3D",
		x"CD",x"F6",x"00",x"7E",x"21",x"80",x"D6",x"01",x"10",x"00",x"CD",x"F6",x"00",x"11",x"50",x"8C",
		x"ED",x"B0",x"C9",x"3A",x"17",x"80",x"B7",x"CA",x"B4",x"4E",x"3A",x"26",x"80",x"B7",x"CA",x"A4",
		x"4E",x"3A",x"27",x"80",x"B7",x"C2",x"9D",x"4E",x"3A",x"CD",x"81",x"18",x"03",x"3A",x"B4",x"81",
		x"B7",x"F2",x"B4",x"4E",x"3A",x"02",x"B0",x"E6",x"08",x"C2",x"BE",x"4E",x"3A",x"02",x"B0",x"E6",
		x"04",x"C2",x"B7",x"4E",x"3E",x"00",x"C9",x"3E",x"01",x"32",x"8B",x"80",x"18",x"0D",x"3A",x"17",
		x"80",x"FE",x"02",x"DA",x"B4",x"4E",x"3E",x"02",x"32",x"8B",x"80",x"3E",x"01",x"C9",x"00",x"21",
		x"D0",x"D8",x"3A",x"A0",x"81",x"3D",x"FE",x"20",x"DA",x"DD",x"4E",x"3E",x"1F",x"01",x"08",x"00",
		x"CD",x"F6",x"00",x"11",x"D2",x"80",x"ED",x"B0",x"11",x"01",x"00",x"ED",x"53",x"DA",x"80",x"2A",
		x"D8",x"80",x"22",x"DC",x"80",x"3A",x"48",x"82",x"FE",x"01",x"CA",x"02",x"4F",x"3A",x"A9",x"81",
		x"18",x"03",x"CD",x"BF",x"4D",x"21",x"B8",x"DB",x"01",x"14",x"00",x"CD",x"F6",x"00",x"11",x"5C",
		x"82",x"ED",x"B0",x"2A",x"5E",x"82",x"22",x"70",x"82",x"2A",x"62",x"82",x"22",x"72",x"82",x"2A",
		x"66",x"82",x"22",x"74",x"82",x"3A",x"48",x"82",x"FE",x"01",x"CA",x"32",x"4F",x"3A",x"A8",x"81",
		x"18",x"03",x"CD",x"69",x"4D",x"21",x"D8",x"D9",x"01",x"0C",x"00",x"CD",x"F6",x"00",x"11",x"C0",
		x"80",x"ED",x"B0",x"2A",x"C6",x"80",x"22",x"CC",x"80",x"2A",x"C8",x"80",x"22",x"CD",x"80",x"2A",
		x"CA",x"80",x"22",x"CF",x"80",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CD",x"C9",x"47",x"C3",x"77",x"41",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C3",x"29",x"4C",x"C3",x"3D",x"43",x"C3",x"D9",x"4B",x"C3",x"E6",x"42",x"C3",x"E6",x"42",x"00",
		x"CD",x"09",x"50",x"00",x"00",x"00",x"C3",x"C3",x"00",x"3A",x"70",x"80",x"B7",x"CA",x"30",x"50",
		x"CD",x"31",x"50",x"B7",x"CA",x"30",x"50",x"DD",x"21",x"21",x"CA",x"CD",x"D2",x"00",x"11",x"E2",
		x"80",x"21",x"9C",x"81",x"01",x"04",x"00",x"ED",x"B0",x"DD",x"21",x"55",x"CA",x"CD",x"D5",x"00",
		x"C9",x"DD",x"21",x"9F",x"81",x"21",x"E5",x"80",x"01",x"04",x"00",x"7E",x"DD",x"BE",x"00",x"DA",
		x"4D",x"50",x"C2",x"52",x"50",x"DD",x"2B",x"2B",x"10",x"F1",x"C3",x"52",x"50",x"3E",x"01",x"C3",
		x"53",x"50",x"AF",x"C9",x"0F",x"0F",x"0F",x"0F",x"C9",x"3A",x"00",x"B0",x"E6",x"40",x"CA",x"6B",
		x"50",x"3E",x"01",x"32",x"74",x"80",x"3E",x"01",x"32",x"77",x"80",x"C9",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"00",x"32",x"95",x"80",x"32",x"8D",x"80",x"32",x"88",x"80",x"3A",x"70",x"80",x"FE",x"00",
		x"20",x"15",x"DD",x"21",x"40",x"83",x"DD",x"36",x"02",x"AC",x"DD",x"36",x"03",x"2F",x"DD",x"36",
		x"04",x"70",x"DD",x"36",x"05",x"73",x"C9",x"3E",x"FF",x"32",x"94",x"80",x"3E",x"00",x"32",x"6C",
		x"84",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"28",x"03",x"00",x"18",x"F6",
		x"DD",x"21",x"6C",x"84",x"DD",x"7E",x"00",x"E6",x"07",x"FE",x"05",x"28",x"63",x"06",x"00",x"3E",
		x"14",x"FE",x"00",x"28",x"08",x"DD",x"70",x"00",x"DD",x"23",x"3D",x"18",x"F4",x"DD",x"21",x"6C",
		x"84",x"3E",x"8B",x"32",x"14",x"88",x"FD",x"21",x"00",x"88",x"FD",x"36",x"00",x"0B",x"21",x"48",
		x"0D",x"22",x"01",x"88",x"FD",x"36",x"03",x"02",x"FD",x"36",x"04",x"01",x"FD",x"36",x"05",x"01",
		x"FD",x"36",x"06",x"01",x"FD",x"36",x"07",x"02",x"FD",x"36",x"08",x"00",x"21",x"00",x"00",x"22",
		x"B4",x"8C",x"DD",x"CB",x"00",x"D6",x"DD",x"CB",x"00",x"8E",x"DD",x"CB",x"00",x"C6",x"DD",x"36",
		x"06",x"03",x"DD",x"36",x"08",x"EE",x"DD",x"36",x"0A",x"03",x"CD",x"43",x"52",x"C3",x"31",x"51",
		x"DD",x"7E",x"0B",x"FE",x"84",x"DA",x"D6",x"51",x"DD",x"CB",x"00",x"CE",x"DD",x"36",x"01",x"00",
		x"FD",x"21",x"00",x"85",x"3E",x"40",x"FE",x"00",x"28",x"09",x"FD",x"36",x"00",x"00",x"FD",x"23",
		x"3D",x"18",x"F3",x"C3",x"1E",x"52",x"DD",x"7E",x"0B",x"FE",x"48",x"DA",x"E1",x"51",x"C3",x"15",
		x"52",x"DD",x"7E",x"0B",x"FE",x"10",x"DA",x"F4",x"51",x"2A",x"75",x"84",x"11",x"0C",x"00",x"ED",
		x"52",x"22",x"75",x"84",x"2A",x"71",x"84",x"ED",x"5B",x"75",x"84",x"19",x"22",x"71",x"84",x"2A",
		x"73",x"84",x"ED",x"52",x"22",x"73",x"84",x"DD",x"7E",x"0C",x"FE",x"50",x"D2",x"15",x"52",x"DD",
		x"86",x"0A",x"DD",x"77",x"0C",x"CD",x"43",x"52",x"DD",x"34",x"0B",x"C3",x"31",x"51",x"3E",x"00",
		x"32",x"94",x"80",x"3E",x"89",x"32",x"00",x"88",x"3E",x"8B",x"32",x"14",x"88",x"3A",x"A0",x"81",
		x"FE",x"06",x"30",x"0E",x"3D",x"87",x"47",x"3E",x"0A",x"90",x"47",x"3A",x"B3",x"81",x"80",x"32",
		x"B3",x"81",x"C9",x"FD",x"E5",x"DD",x"36",x"02",x"0B",x"DD",x"7E",x"0B",x"FE",x"48",x"20",x"11",
		x"21",x"00",x"0D",x"22",x"01",x"88",x"3E",x"02",x"32",x"05",x"88",x"21",x"C0",x"00",x"22",x"B2",
		x"8C",x"DD",x"7E",x"0B",x"FE",x"48",x"38",x"10",x"CB",x"4F",x"28",x"0C",x"3A",x"B2",x"8C",x"FE",
		x"00",x"28",x"05",x"D6",x"10",x"32",x"B2",x"8C",x"DD",x"36",x"04",x"7A",x"DD",x"7E",x"0C",x"FE",
		x"10",x"DA",x"00",x"53",x"FE",x"20",x"DA",x"DA",x"52",x"FE",x"30",x"DA",x"B4",x"52",x"DD",x"36",
		x"01",x"40",x"DD",x"7E",x"06",x"D6",x"30",x"DD",x"77",x"03",x"FD",x"21",x"00",x"85",x"CD",x"25",
		x"53",x"DD",x"36",x"01",x"47",x"DD",x"7E",x"08",x"C6",x"30",x"DD",x"77",x"03",x"FD",x"21",x"38",
		x"85",x"CD",x"25",x"53",x"DD",x"36",x"01",x"41",x"DD",x"7E",x"06",x"D6",x"20",x"DD",x"77",x"03",
		x"FD",x"21",x"08",x"85",x"CD",x"25",x"53",x"DD",x"36",x"01",x"46",x"DD",x"7E",x"08",x"C6",x"20",
		x"DD",x"77",x"03",x"FD",x"21",x"30",x"85",x"CD",x"25",x"53",x"DD",x"36",x"01",x"42",x"DD",x"7E",
		x"06",x"D6",x"10",x"DD",x"77",x"03",x"FD",x"21",x"10",x"85",x"CD",x"25",x"53",x"DD",x"36",x"01",
		x"45",x"DD",x"7E",x"08",x"C6",x"10",x"DD",x"77",x"03",x"FD",x"21",x"28",x"85",x"CD",x"25",x"53",
		x"DD",x"36",x"01",x"43",x"DD",x"7E",x"06",x"DD",x"77",x"03",x"FD",x"21",x"18",x"85",x"CD",x"25",
		x"53",x"DD",x"36",x"01",x"44",x"DD",x"7E",x"08",x"DD",x"77",x"03",x"FD",x"21",x"20",x"85",x"CD",
		x"25",x"53",x"FD",x"E1",x"C9",x"DD",x"7E",x"01",x"FD",x"77",x"00",x"DD",x"7E",x"02",x"FD",x"77",
		x"01",x"DD",x"7E",x"03",x"FD",x"77",x"02",x"DD",x"7E",x"04",x"FD",x"77",x"03",x"C9",x"3E",x"FF",
		x"32",x"94",x"80",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"28",x"03",x"00",
		x"18",x"F6",x"DD",x"21",x"6C",x"84",x"DD",x"7E",x"00",x"E6",x"0F",x"FE",x"05",x"28",x"77",x"DD",
		x"36",x"00",x"05",x"DD",x"36",x"01",x"AC",x"DD",x"36",x"02",x"2B",x"3A",x"02",x"85",x"DD",x"77",
		x"03",x"3A",x"03",x"85",x"DD",x"77",x"04",x"21",x"00",x"00",x"22",x"71",x"84",x"22",x"77",x"84",
		x"21",x"FF",x"0F",x"22",x"BE",x"8C",x"3E",x"8B",x"32",x"14",x"88",x"DD",x"7E",x"03",x"21",x"80",
		x"01",x"FE",x"71",x"38",x"03",x"CD",x"F3",x"1F",x"22",x"73",x"84",x"DD",x"7E",x"04",x"21",x"80",
		x"01",x"FE",x"73",x"38",x"03",x"CD",x"F3",x"1F",x"22",x"75",x"84",x"11",x"71",x"00",x"21",x"00",
		x"00",x"DD",x"6E",x"03",x"ED",x"52",x"CD",x"F0",x"1F",x"4D",x"21",x"00",x"00",x"DD",x"6E",x"04",
		x"11",x"73",x"00",x"ED",x"52",x"CD",x"F0",x"1F",x"7D",x"B9",x"38",x"04",x"DD",x"CB",x"00",x"F6",
		x"CD",x"C2",x"54",x"C3",x"3E",x"53",x"DD",x"7E",x"0B",x"FE",x"10",x"30",x"09",x"CD",x"96",x"54",
		x"DD",x"34",x"0B",x"C3",x"3E",x"53",x"DD",x"7E",x"00",x"E6",x"30",x"FE",x"30",x"28",x"0F",x"CD",
		x"96",x"54",x"DD",x"34",x"0B",x"CD",x"24",x"54",x"CD",x"C2",x"54",x"C3",x"3E",x"53",x"DD",x"7E",
		x"0B",x"FE",x"FE",x"30",x"16",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"28",
		x"02",x"18",x"F7",x"CD",x"96",x"54",x"DD",x"34",x"0B",x"18",x"E3",x"3E",x"00",x"32",x"94",x"80",
		x"32",x"00",x"85",x"C9",x"DD",x"CB",x"00",x"76",x"C2",x"61",x"54",x"21",x"00",x"00",x"DD",x"6E",
		x"03",x"11",x"71",x"00",x"ED",x"52",x"CD",x"F0",x"1F",x"7D",x"FE",x"02",x"28",x"02",x"30",x"0E",
		x"DD",x"CB",x"00",x"E6",x"DD",x"CB",x"00",x"F6",x"DD",x"36",x"03",x"71",x"18",x"D6",x"DD",x"66",
		x"03",x"DD",x"6E",x"05",x"ED",x"5B",x"73",x"84",x"19",x"DD",x"74",x"03",x"DD",x"75",x"05",x"18",
		x"34",x"21",x"00",x"00",x"DD",x"6E",x"04",x"11",x"73",x"00",x"ED",x"52",x"CD",x"F0",x"1F",x"7D",
		x"FE",x"02",x"28",x"02",x"30",x"0E",x"DD",x"CB",x"00",x"EE",x"DD",x"CB",x"00",x"B6",x"DD",x"36",
		x"04",x"73",x"18",x"11",x"DD",x"66",x"04",x"DD",x"6E",x"06",x"ED",x"5B",x"75",x"84",x"19",x"DD",
		x"74",x"04",x"DD",x"75",x"06",x"C9",x"3A",x"77",x"84",x"E6",x"07",x"FE",x"00",x"20",x"22",x"DD",
		x"34",x"0C",x"DD",x"7E",x"0C",x"FE",x"07",x"38",x"05",x"3E",x"00",x"32",x"78",x"84",x"87",x"16",
		x"00",x"5F",x"FD",x"21",x"DB",x"54",x"FD",x"19",x"FD",x"66",x"01",x"FD",x"6E",x"00",x"22",x"BE",
		x"8C",x"C9",x"DD",x"7E",x"01",x"32",x"00",x"85",x"DD",x"7E",x"02",x"32",x"01",x"85",x"DD",x"7E",
		x"03",x"32",x"02",x"85",x"DD",x"7E",x"04",x"32",x"03",x"85",x"C9",x"FF",x"0F",x"AF",x"0A",x"5F",
		x"05",x"0F",x"00",x"0F",x"00",x"5F",x"05",x"AF",x"0A",x"C9",x"E5",x"DD",x"E5",x"C5",x"FD",x"E5",
		x"3E",x"00",x"32",x"A6",x"81",x"3A",x"A2",x"81",x"FE",x"00",x"CA",x"69",x"55",x"3A",x"A0",x"81",
		x"3D",x"26",x"00",x"6F",x"06",x"00",x"4F",x"29",x"29",x"09",x"09",x"01",x"38",x"DE",x"09",x"23",
		x"23",x"23",x"23",x"7E",x"26",x"00",x"6F",x"29",x"44",x"4D",x"29",x"29",x"09",x"01",x"80",x"D8",
		x"09",x"E5",x"FD",x"E1",x"FD",x"7E",x"05",x"32",x"A0",x"85",x"FD",x"7E",x"06",x"32",x"A1",x"85",
		x"FD",x"7E",x"07",x"32",x"A2",x"85",x"FD",x"7E",x"08",x"32",x"A3",x"85",x"FD",x"7E",x"09",x"32",
		x"A4",x"85",x"DD",x"21",x"80",x"84",x"DD",x"7E",x"00",x"FE",x"FF",x"CA",x"69",x"55",x"DD",x"CB",
		x"00",x"76",x"C2",x"61",x"55",x"DD",x"46",x"01",x"DD",x"4E",x"02",x"CD",x"DE",x"00",x"CD",x"70",
		x"55",x"01",x"05",x"00",x"DD",x"09",x"C3",x"46",x"55",x"FD",x"E1",x"C1",x"DD",x"E1",x"E1",x"C9",
		x"E5",x"D5",x"DD",x"E5",x"E5",x"DD",x"E1",x"11",x"00",x"04",x"DD",x"19",x"FD",x"46",x"04",x"FD",
		x"7E",x"02",x"77",x"DD",x"70",x"00",x"DD",x"23",x"23",x"FD",x"7E",x"03",x"77",x"DD",x"70",x"00",
		x"11",x"DF",x"FF",x"ED",x"5A",x"DD",x"19",x"FD",x"7E",x"00",x"77",x"DD",x"70",x"00",x"DD",x"23",
		x"23",x"FD",x"7E",x"01",x"77",x"DD",x"70",x"00",x"DD",x"E1",x"D1",x"E1",x"C9",x"C5",x"D5",x"DD",
		x"E5",x"FD",x"E5",x"DD",x"21",x"A3",x"81",x"FD",x"21",x"80",x"84",x"DD",x"46",x"00",x"0E",x"08",
		x"FD",x"7E",x"00",x"FE",x"FF",x"CA",x"E8",x"55",x"CB",x"40",x"28",x"04",x"FD",x"CB",x"00",x"F6",
		x"11",x"05",x"00",x"FD",x"19",x"0D",x"79",x"FE",x"00",x"28",x"05",x"CB",x"38",x"C3",x"C0",x"55",
		x"11",x"01",x"00",x"DD",x"19",x"C3",x"BB",x"55",x"FD",x"E1",x"DD",x"E1",x"D1",x"C1",x"C9",x"C5",
		x"D5",x"DD",x"E5",x"FD",x"E5",x"DD",x"21",x"A3",x"81",x"FD",x"21",x"80",x"84",x"06",x"00",x"0E",
		x"08",x"FD",x"7E",x"00",x"FE",x"FF",x"CA",x"2A",x"56",x"CB",x"38",x"FD",x"CB",x"00",x"76",x"28",
		x"02",x"CB",x"F8",x"11",x"05",x"00",x"FD",x"19",x"0D",x"79",x"FE",x"00",x"C2",x"01",x"56",x"DD",
		x"70",x"00",x"11",x"01",x"00",x"DD",x"19",x"C3",x"FD",x"55",x"FD",x"E1",x"DD",x"E1",x"D1",x"C1",
		x"C9",x"C5",x"D5",x"E5",x"FD",x"E5",x"21",x"00",x"70",x"DD",x"7E",x"01",x"FE",x"02",x"38",x"08",
		x"FD",x"23",x"FD",x"23",x"FD",x"23",x"FD",x"23",x"87",x"16",x"00",x"5F",x"19",x"FD",x"7E",x"02",
		x"56",x"82",x"47",x"FD",x"7E",x"03",x"23",x"56",x"82",x"4F",x"CD",x"DE",x"00",x"E5",x"FD",x"E1",
		x"11",x"00",x"00",x"DD",x"7E",x"01",x"FE",x"01",x"28",x"24",x"DD",x"CB",x"0B",x"7E",x"28",x"0C",
		x"FD",x"7E",x"FF",x"CD",x"FC",x"56",x"FE",x"00",x"28",x"02",x"CB",x"DB",x"DD",x"CB",x"0B",x"7E",
		x"20",x"0C",x"FD",x"7E",x"01",x"CD",x"FC",x"56",x"FE",x"00",x"28",x"02",x"CB",x"D3",x"DD",x"CB",
		x"09",x"7E",x"28",x"0C",x"FD",x"7E",x"20",x"CD",x"FC",x"56",x"FE",x"00",x"28",x"02",x"CB",x"CB",
		x"DD",x"CB",x"09",x"7E",x"20",x"0C",x"FD",x"7E",x"E0",x"CD",x"FC",x"56",x"FE",x"00",x"28",x"02",
		x"CB",x"C3",x"DD",x"7E",x"01",x"FE",x"01",x"C2",x"F5",x"56",x"FD",x"E1",x"FD",x"E5",x"FD",x"7E",
		x"02",x"C6",x"01",x"47",x"FD",x"7E",x"03",x"C6",x"08",x"4F",x"CD",x"DE",x"00",x"23",x"7E",x"CD",
		x"FC",x"56",x"FE",x"00",x"28",x"04",x"CB",x"D3",x"18",x"1B",x"FD",x"7E",x"02",x"C6",x"0E",x"47",
		x"FD",x"7E",x"03",x"C6",x"08",x"4F",x"CD",x"DE",x"00",x"23",x"7E",x"CD",x"FC",x"56",x"FE",x"00",
		x"CA",x"F5",x"56",x"CB",x"D3",x"7B",x"FD",x"E1",x"E1",x"D1",x"C1",x"C9",x"FE",x"60",x"38",x"0C",
		x"FE",x"80",x"38",x"0A",x"FE",x"A0",x"38",x"04",x"FE",x"C0",x"38",x"02",x"3E",x"00",x"C9",x"3A",
		x"AB",x"81",x"FE",x"14",x"DA",x"09",x"58",x"3E",x"2B",x"CD",x"FC",x"00",x"3E",x"00",x"32",x"82",
		x"89",x"32",x"83",x"89",x"32",x"84",x"89",x"3E",x"00",x"32",x"AC",x"81",x"CD",x"CF",x"00",x"0E",
		x"70",x"0F",x"3A",x"AB",x"81",x"FE",x"14",x"20",x"14",x"3E",x"0F",x"CD",x"18",x"60",x"CD",x"CF",
		x"00",x"D4",x"71",x"02",x"16",x"0A",x"3E",x"01",x"32",x"84",x"89",x"18",x"49",x"F5",x"3E",x"0F",
		x"CD",x"18",x"60",x"F1",x"FE",x"15",x"20",x"14",x"3E",x"0F",x"CD",x"18",x"60",x"CD",x"CF",x"00",
		x"D8",x"71",x"02",x"16",x"14",x"3E",x"02",x"32",x"84",x"89",x"18",x"2A",x"FE",x"16",x"20",x"14",
		x"3E",x"0F",x"CD",x"18",x"60",x"CD",x"CF",x"00",x"DC",x"71",x"02",x"16",x"1E",x"3E",x"03",x"32",
		x"84",x"89",x"18",x"12",x"3E",x"0E",x"CD",x"18",x"60",x"CD",x"CF",x"00",x"E0",x"71",x"02",x"16",
		x"32",x"3E",x"05",x"32",x"84",x"89",x"06",x"00",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",
		x"FE",x"00",x"20",x"F9",x"04",x"78",x"FE",x"78",x"20",x"EE",x"1E",x"00",x"3E",x"01",x"32",x"6E",
		x"80",x"3A",x"6E",x"80",x"FE",x"00",x"20",x"F9",x"7A",x"FE",x"00",x"28",x"28",x"1C",x"7B",x"E6",
		x"03",x"20",x"E9",x"01",x"00",x"10",x"CD",x"E4",x"00",x"3A",x"83",x"89",x"D6",x"0A",x"27",x"32",
		x"83",x"89",x"3A",x"84",x"89",x"DE",x"00",x"27",x"32",x"84",x"89",x"DD",x"21",x"44",x"72",x"CD",
		x"D5",x"00",x"15",x"18",x"C7",x"3E",x"00",x"32",x"F3",x"91",x"32",x"B3",x"91",x"32",x"93",x"91",
		x"06",x"00",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"20",x"F9",x"04",x"78",
		x"FE",x"3C",x"20",x"EE",x"3E",x"AB",x"CD",x"FC",x"00",x"3E",x"00",x"32",x"AB",x"81",x"32",x"00",
		x"89",x"32",x"01",x"89",x"C9",x"DD",x"21",x"28",x"80",x"DD",x"36",x"02",x"00",x"DD",x"36",x"03",
		x"00",x"DD",x"36",x"04",x"00",x"DD",x"36",x"05",x"00",x"DD",x"36",x"06",x"14",x"DD",x"36",x"07",
		x"15",x"FD",x"21",x"18",x"85",x"FD",x"36",x"00",x"14",x"FD",x"36",x"01",x"0C",x"FD",x"36",x"02",
		x"78",x"FD",x"36",x"03",x"78",x"FD",x"36",x"08",x"AE",x"FD",x"36",x"09",x"2B",x"FD",x"36",x"0A",
		x"60",x"FD",x"36",x"0B",x"60",x"FD",x"36",x"10",x"AF",x"FD",x"36",x"11",x"2B",x"FD",x"36",x"12",
		x"80",x"FD",x"36",x"13",x"60",x"FD",x"36",x"18",x"B0",x"FD",x"36",x"19",x"2B",x"FD",x"36",x"1A",
		x"60",x"FD",x"36",x"1B",x"80",x"FD",x"36",x"20",x"B1",x"FD",x"36",x"21",x"2B",x"FD",x"36",x"22",
		x"80",x"FD",x"36",x"23",x"80",x"3E",x"01",x"32",x"6E",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"28",
		x"03",x"00",x"18",x"F6",x"DD",x"34",x"02",x"3A",x"2A",x"80",x"FE",x"3C",x"38",x"07",x"DD",x"36",
		x"02",x"00",x"DD",x"34",x"03",x"DD",x"34",x"04",x"3A",x"2C",x"80",x"FE",x"04",x"38",x"07",x"CD",
		x"DB",x"59",x"DD",x"36",x"04",x"00",x"DD",x"34",x"05",x"3A",x"2D",x"80",x"FE",x"04",x"38",x"67",
		x"DD",x"36",x"05",x"00",x"3A",x"2E",x"80",x"FE",x"FF",x"28",x"06",x"CD",x"30",x"59",x"DD",x"35",
		x"06",x"3A",x"2F",x"80",x"FE",x"FF",x"28",x"06",x"CD",x"86",x"59",x"DD",x"35",x"07",x"3A",x"2B",
		x"80",x"FE",x"03",x"20",x"42",x"3A",x"2A",x"80",x"FE",x"10",x"20",x"0C",x"3E",x"00",x"32",x"40",
		x"85",x"3E",x"0A",x"32",x"41",x"85",x"18",x"2F",x"3A",x"2A",x"80",x"FE",x"0C",x"28",x"02",x"30",
		x"26",x"FE",x"00",x"20",x"1F",x"3A",x"17",x"80",x"FE",x"99",x"30",x"08",x"C6",x"01",x"27",x"32",
		x"17",x"80",x"18",x"09",x"3A",x"87",x"80",x"C6",x"01",x"27",x"32",x"87",x"80",x"CD",x"F0",x"00",
		x"DD",x"21",x"28",x"80",x"CD",x"F2",x"59",x"3A",x"2B",x"80",x"FE",x"0B",x"DA",x"85",x"58",x"C9",
		x"DD",x"E5",x"DD",x"21",x"B6",x"92",x"FD",x"21",x"B6",x"96",x"21",x"68",x"D2",x"01",x"00",x"00",
		x"79",x"FE",x"14",x"28",x"03",x"D2",x"83",x"59",x"DD",x"36",x"00",x"00",x"FD",x"36",x"00",x"0A",
		x"78",x"FE",x"00",x"20",x"1B",x"3A",x"2E",x"80",x"B9",x"28",x"02",x"30",x"13",x"7E",x"FE",x"FF",
		x"20",x"04",x"06",x"01",x"18",x"0A",x"7E",x"DD",x"77",x"00",x"23",x"7E",x"FD",x"77",x"00",x"23",
		x"79",x"FE",x"0E",x"38",x"04",x"DD",x"2B",x"FD",x"2B",x"11",x"E0",x"FF",x"DD",x"19",x"FD",x"19",
		x"0C",x"18",x"BD",x"DD",x"E1",x"C9",x"DD",x"E5",x"DD",x"21",x"37",x"91",x"FD",x"21",x"37",x"95",
		x"21",x"83",x"D2",x"01",x"00",x"00",x"79",x"FE",x"15",x"28",x"02",x"30",x"3B",x"DD",x"36",x"00",
		x"00",x"FD",x"36",x"00",x"0A",x"78",x"FE",x"00",x"20",x"1B",x"3A",x"2F",x"80",x"B9",x"28",x"02",
		x"30",x"13",x"7E",x"FE",x"FF",x"20",x"04",x"06",x"01",x"18",x"0A",x"7E",x"DD",x"77",x"00",x"23",
		x"7E",x"FD",x"77",x"00",x"23",x"79",x"FE",x"0D",x"38",x"04",x"DD",x"2B",x"FD",x"2B",x"11",x"20",
		x"00",x"DD",x"19",x"FD",x"19",x"0C",x"18",x"BE",x"DD",x"E1",x"C9",x"C5",x"3A",x"18",x"85",x"4F",
		x"E6",x"03",x"FE",x"03",x"20",x"05",x"79",x"E6",x"FC",x"18",x"02",x"0C",x"79",x"32",x"18",x"85",
		x"C1",x"C9",x"3E",x"AD",x"32",x"40",x"85",x"3E",x"3B",x"32",x"41",x"85",x"3E",x"8C",x"32",x"42",
		x"85",x"3E",x"D4",x"32",x"43",x"85",x"C9",x"C9",x"C5",x"D5",x"3A",x"AE",x"81",x"FE",x"FF",x"CA",
		x"E3",x"5A",x"3A",x"14",x"80",x"E6",x"07",x"FE",x"00",x"20",x"03",x"C3",x"E3",x"5A",x"FE",x"01",
		x"20",x"05",x"06",x"0A",x"C3",x"59",x"5A",x"FE",x"02",x"20",x"05",x"06",x"03",x"C3",x"59",x"5A",
		x"FE",x"03",x"20",x"05",x"06",x"05",x"C3",x"69",x"5A",x"FE",x"04",x"20",x"05",x"06",x"0A",x"C3",
		x"69",x"5A",x"FE",x"05",x"20",x"07",x"06",x"05",x"0E",x"0A",x"C3",x"7A",x"5A",x"FE",x"06",x"C2",
		x"9F",x"5A",x"06",x"0A",x"0E",x"1E",x"C3",x"7A",x"5A",x"16",x"00",x"3A",x"AD",x"81",x"B8",x"DA",
		x"D4",x"5A",x"14",x"90",x"32",x"AD",x"81",x"18",x"F2",x"3A",x"AD",x"81",x"B8",x"DA",x"E3",x"5A",
		x"16",x"01",x"3E",x"FF",x"32",x"AE",x"81",x"C3",x"D4",x"5A",x"16",x"00",x"3A",x"AE",x"81",x"FE",
		x"01",x"28",x"0D",x"3A",x"AD",x"81",x"B8",x"DA",x"E3",x"5A",x"14",x"3E",x"01",x"32",x"AE",x"81",
		x"3A",x"AD",x"81",x"B9",x"38",x"3E",x"14",x"3E",x"FF",x"32",x"AE",x"81",x"C3",x"D4",x"5A",x"16",
		x"00",x"3A",x"AE",x"81",x"FE",x"01",x"28",x"12",x"FE",x"02",x"28",x"1B",x"3A",x"AD",x"81",x"FE",
		x"05",x"DA",x"E3",x"5A",x"14",x"3E",x"01",x"32",x"AE",x"81",x"3A",x"AD",x"81",x"FE",x"0A",x"38",
		x"13",x"14",x"3E",x"02",x"32",x"AE",x"81",x"3A",x"AD",x"81",x"FE",x"1E",x"38",x"06",x"14",x"3E",
		x"FF",x"32",x"AE",x"81",x"7A",x"FE",x"00",x"28",x"0A",x"3A",x"9B",x"81",x"82",x"32",x"9B",x"81",
		x"CD",x"F3",x"4F",x"D1",x"C1",x"F1",x"C9",x"3A",x"04",x"B0",x"E6",x"03",x"FE",x"03",x"28",x"03",
		x"3C",x"18",x"02",x"3E",x"06",x"32",x"16",x"80",x"3A",x"04",x"B0",x"E6",x"0C",x"CB",x"3F",x"CB",
		x"3F",x"FE",x"01",x"20",x"0E",x"3E",x"FF",x"32",x"84",x"80",x"3E",x"00",x"32",x"85",x"80",x"3E",
		x"01",x"18",x"06",x"FE",x"00",x"20",x"02",x"3E",x"01",x"32",x"83",x"80",x"3A",x"04",x"B0",x"E6",
		x"30",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"FE",x"03",x"28",x"04",x"C6",x"03",x"18",
		x"02",x"3E",x"02",x"32",x"71",x"80",x"3A",x"04",x"B0",x"E6",x"40",x"28",x"02",x"3E",x"01",x"32",
		x"72",x"80",x"3A",x"04",x"B0",x"E6",x"80",x"28",x"02",x"3E",x"01",x"32",x"73",x"80",x"C9",x"DD",
		x"E5",x"DD",x"21",x"00",x"89",x"DD",x"CB",x"00",x"46",x"28",x"0F",x"CD",x"EC",x"2F",x"DD",x"7E",
		x"02",x"32",x"10",x"85",x"DD",x"7E",x"03",x"32",x"11",x"85",x"DD",x"E1",x"C9",x"F5",x"3A",x"8F",
		x"80",x"FE",x"00",x"28",x"52",x"7B",x"FE",x"00",x"28",x"4D",x"FE",x"FF",x"28",x"49",x"C5",x"E5",
		x"DD",x"E5",x"3A",x"A0",x"81",x"3D",x"26",x"00",x"6F",x"29",x"44",x"4D",x"29",x"09",x"DD",x"21",
		x"38",x"DE",x"44",x"4D",x"DD",x"09",x"DD",x"7E",x"02",x"DD",x"E1",x"E1",x"01",x"00",x"00",x"FE",
		x"04",x"38",x"06",x"06",x"10",x"3D",x"3D",x"3D",x"3D",x"FE",x"00",x"28",x"12",x"FE",x"01",x"20",
		x"04",x"0E",x"10",x"18",x"0A",x"FE",x"02",x"20",x"04",x"0E",x"40",x"18",x"02",x"0E",x"50",x"7A",
		x"B7",x"B0",x"57",x"7B",x"81",x"5F",x"C1",x"F1",x"C9",x"F5",x"C5",x"D5",x"E5",x"3A",x"94",x"80",
		x"FE",x"FF",x"CA",x"0B",x"5C",x"3A",x"91",x"80",x"3C",x"32",x"91",x"80",x"FE",x"03",x"DA",x"0B",
		x"5C",x"3E",x"00",x"32",x"91",x"80",x"21",x"0A",x"0F",x"11",x"B2",x"8C",x"01",x"0E",x"00",x"ED",
		x"B0",x"3A",x"92",x"80",x"3C",x"FE",x"07",x"38",x"02",x"3E",x"00",x"32",x"92",x"80",x"87",x"16",
		x"00",x"5F",x"21",x"B2",x"8C",x"19",x"36",x"FF",x"23",x"36",x"0F",x"E1",x"D1",x"C1",x"F1",x"C9",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C3",x"E7",x"5A",x"C3",x"6D",x"5B",x"C3",x"FC",x"56",x"C3",x"C9",x"5B",x"00",x"C3",x"07",x"5A",
		x"C3",x"00",x"51",x"C3",x"3E",x"53",x"C3",x"E9",x"54",x"C3",x"EA",x"54",x"C3",x"AD",x"55",x"C3",
		x"EF",x"55",x"C3",x"31",x"56",x"C3",x"0F",x"57",x"C3",x"09",x"50",x"C3",x"15",x"58",x"00",x"00",
		x"C3",x"02",x"61",x"C3",x"37",x"61",x"C3",x"74",x"61",x"C3",x"A6",x"61",x"C3",x"09",x"62",x"C3",
		x"81",x"62",x"C3",x"BE",x"62",x"C3",x"E5",x"62",x"C3",x"26",x"63",x"C3",x"9A",x"63",x"C3",x"BF",
		x"63",x"C3",x"79",x"64",x"C3",x"D8",x"64",x"C3",x"24",x"65",x"C3",x"69",x"65",x"C3",x"90",x"65",
		x"C3",x"FB",x"66",x"C3",x"18",x"67",x"C3",x"81",x"67",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C9",x"21",x"7A",x"82",x"11",x"18",x"85",x"06",x"09",x"C5",x"01",x"04",x"00",x"2B",x"2B",
		x"7E",x"FE",x"20",x"23",x"23",x"C2",x"29",x"61",x"2B",x"7E",x"FE",x"0C",x"23",x"D2",x"29",x"61",
		x"13",x"13",x"13",x"13",x"ED",x"B0",x"C3",x"2F",x"61",x"ED",x"B0",x"13",x"13",x"13",x"13",x"01",
		x"15",x"00",x"09",x"C1",x"10",x"D4",x"C9",x"3A",x"8D",x"80",x"B7",x"C2",x"73",x"61",x"DD",x"5E",
		x"0E",x"DD",x"56",x"0F",x"D5",x"01",x"80",x"01",x"21",x"10",x"00",x"EB",x"B7",x"ED",x"42",x"7D",
		x"B4",x"E1",x"C2",x"58",x"61",x"11",x"08",x"00",x"19",x"DD",x"75",x"0E",x"DD",x"74",x"0F",x"DD",
		x"5E",x"0A",x"DD",x"56",x"0B",x"19",x"DD",x"5E",x"07",x"DD",x"56",x"05",x"19",x"DD",x"75",x"07",
		x"DD",x"74",x"05",x"C9",x"78",x"92",x"57",x"79",x"93",x"5F",x"AF",x"B2",x"F2",x"8C",x"61",x"23",
		x"ED",x"44",x"57",x"7E",x"23",x"92",x"DA",x"A4",x"61",x"C3",x"91",x"61",x"7E",x"23",x"C3",x"84",
		x"61",x"AF",x"B3",x"F2",x"9A",x"61",x"23",x"ED",x"44",x"5F",x"7E",x"93",x"DA",x"A4",x"61",x"3E",
		x"01",x"C3",x"A5",x"61",x"AF",x"C9",x"3A",x"8D",x"80",x"B7",x"C2",x"08",x"62",x"DD",x"7E",x"11",
		x"FE",x"02",x"D2",x"C3",x"61",x"DD",x"5E",x"08",x"DD",x"56",x"09",x"DD",x"66",x"04",x"DD",x"6E",
		x"06",x"18",x"0F",x"DD",x"5E",x"0A",x"DD",x"56",x"0B",x"DD",x"66",x"05",x"DD",x"6E",x"07",x"3D",
		x"E6",x"01",x"B7",x"C2",x"D9",x"61",x"19",x"18",x"03",x"B7",x"ED",x"52",x"3E",x"01",x"DD",x"BE",
		x"11",x"DA",x"F7",x"61",x"7C",x"DD",x"BE",x"04",x"CA",x"EF",x"61",x"DD",x"36",x"18",x"00",x"DD",
		x"74",x"04",x"DD",x"75",x"06",x"18",x"11",x"7C",x"DD",x"BE",x"05",x"CA",x"02",x"62",x"DD",x"36",
		x"18",x"00",x"DD",x"74",x"05",x"DD",x"75",x"07",x"C9",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",
		x"DD",x"21",x"28",x"C8",x"3A",x"A0",x"81",x"3D",x"01",x"06",x"00",x"21",x"3B",x"DE",x"CD",x"F6",
		x"00",x"7E",x"87",x"16",x"00",x"5F",x"DD",x"19",x"DD",x"66",x"01",x"DD",x"6E",x"00",x"E5",x"DD",
		x"E1",x"FD",x"21",x"80",x"84",x"0E",x"00",x"79",x"FE",x"18",x"CA",x"75",x"62",x"FD",x"71",x"00",
		x"21",x"C8",x"C9",x"16",x"00",x"DD",x"7E",x"00",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",
		x"5F",x"19",x"7E",x"FD",x"77",x"01",x"21",x"C8",x"C9",x"16",x"00",x"DD",x"7E",x"00",x"E6",x"0F",
		x"5F",x"19",x"7E",x"FD",x"77",x"02",x"0C",x"DD",x"23",x"FD",x"23",x"FD",x"23",x"FD",x"23",x"FD",
		x"23",x"FD",x"23",x"18",x"C2",x"FD",x"36",x"00",x"FF",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",
		x"C9",x"C5",x"D5",x"E5",x"F5",x"3A",x"70",x"80",x"B7",x"20",x"16",x"3A",x"17",x"80",x"B7",x"C2",
		x"A1",x"62",x"3A",x"13",x"80",x"CB",x"7F",x"28",x"20",x"F1",x"F5",x"E6",x"7F",x"FE",x"20",x"20",
		x"18",x"21",x"01",x"87",x"01",x"01",x"00",x"3A",x"00",x"87",x"CD",x"F6",x"00",x"F1",x"77",x"3A",
		x"00",x"87",x"3C",x"32",x"00",x"87",x"C3",x"BA",x"62",x"F1",x"E1",x"D1",x"C1",x"C9",x"3A",x"00",
		x"87",x"B7",x"C8",x"21",x"01",x"87",x"7E",x"32",x"00",x"B8",x"3A",x"00",x"87",x"3D",x"32",x"00",
		x"87",x"C8",x"47",x"21",x"01",x"87",x"E5",x"DD",x"E1",x"DD",x"23",x"DD",x"7E",x"00",x"77",x"23",
		x"DD",x"23",x"10",x"F7",x"C9",x"3A",x"70",x"80",x"FE",x"00",x"28",x"08",x"3A",x"14",x"80",x"E6",
		x"18",x"0F",x"0F",x"0F",x"21",x"01",x"63",x"16",x"00",x"5F",x"19",x"7E",x"32",x"A8",x"81",x"18",
		x"04",x"00",x"01",x"03",x"07",x"3A",x"70",x"80",x"FE",x"00",x"28",x"08",x"3A",x"14",x"80",x"E6",
		x"60",x"07",x"07",x"07",x"21",x"21",x"63",x"16",x"00",x"5F",x"19",x"7E",x"32",x"A9",x"81",x"18",
		x"04",x"00",x"00",x"01",x"03",x"C9",x"C5",x"D5",x"E5",x"FE",x"11",x"D2",x"96",x"63",x"32",x"86",
		x"89",x"FE",x"10",x"CA",x"91",x"63",x"FE",x"08",x"D2",x"69",x"63",x"21",x"3A",x"DE",x"01",x"06",
		x"00",x"3A",x"A0",x"81",x"3D",x"CD",x"F6",x"00",x"7E",x"F5",x"21",x"00",x"D7",x"01",x"10",x"00",
		x"CD",x"F6",x"00",x"11",x"A0",x"8C",x"ED",x"B0",x"F1",x"21",x"80",x"D7",x"01",x"10",x"00",x"CD",
		x"F6",x"00",x"11",x"80",x"8C",x"ED",x"B0",x"18",x"28",x"D6",x"08",x"87",x"21",x"81",x"63",x"16",
		x"00",x"5F",x"19",x"5E",x"23",x"56",x"EB",x"11",x"70",x"8C",x"01",x"10",x"00",x"ED",x"B0",x"18",
		x"10",x"00",x"D8",x"10",x"D8",x"20",x"D8",x"30",x"D8",x"40",x"D8",x"50",x"D8",x"60",x"D8",x"70",
		x"D8",x"3E",x"01",x"32",x"85",x"89",x"E1",x"D1",x"C1",x"C9",x"3A",x"85",x"89",x"B7",x"C8",x"3A",
		x"86",x"89",x"FE",x"10",x"CA",x"B4",x"63",x"F5",x"21",x"70",x"8C",x"11",x"70",x"9C",x"01",x"40",
		x"00",x"ED",x"B0",x"F1",x"CB",x"E7",x"32",x"00",x"9E",x"3E",x"00",x"32",x"85",x"89",x"C9",x"F5",
		x"E5",x"DD",x"E5",x"D5",x"3A",x"9E",x"81",x"E6",x"0F",x"5F",x"F5",x"3A",x"AC",x"81",x"57",x"C5",
		x"B7",x"CB",x"38",x"CB",x"19",x"B7",x"CB",x"38",x"CB",x"19",x"B7",x"CB",x"38",x"CB",x"19",x"B7",
		x"CB",x"38",x"CB",x"19",x"B7",x"2A",x"B1",x"81",x"7D",x"81",x"27",x"6F",x"7C",x"88",x"27",x"67",
		x"22",x"B1",x"81",x"C1",x"21",x"9C",x"81",x"7E",x"81",x"27",x"77",x"23",x"7E",x"88",x"27",x"77",
		x"23",x"7E",x"CE",x"00",x"27",x"77",x"23",x"7E",x"CE",x"00",x"27",x"77",x"3A",x"AE",x"81",x"FE",
		x"FF",x"28",x"10",x"3A",x"9E",x"81",x"E6",x"0F",x"BB",x"28",x"08",x"5F",x"3A",x"AD",x"81",x"3C",
		x"32",x"AD",x"81",x"7A",x"FE",x"00",x"28",x"04",x"15",x"C3",x"CF",x"63",x"3A",x"27",x"80",x"B7",
		x"CA",x"3A",x"64",x"DD",x"21",x"61",x"CA",x"C3",x"3E",x"64",x"DD",x"21",x"4F",x"CA",x"3A",x"70",
		x"80",x"B7",x"CA",x"48",x"64",x"CD",x"D5",x"00",x"F1",x"3A",x"B2",x"81",x"FE",x"05",x"38",x"20",
		x"D6",x"05",x"27",x"FE",x"05",x"30",x"F9",x"32",x"B2",x"81",x"3A",x"88",x"80",x"FE",x"00",x"20",
		x"0F",x"3A",x"AC",x"81",x"FE",x"04",x"30",x"08",x"3A",x"00",x"89",x"CB",x"C7",x"32",x"00",x"89",
		x"CD",x"DD",x"5F",x"D1",x"DD",x"E1",x"E1",x"F1",x"C9",x"CD",x"24",x"65",x"CD",x"D8",x"64",x"3A",
		x"13",x"80",x"E6",x"03",x"FE",x"00",x"20",x"06",x"DD",x"21",x"2B",x"66",x"18",x"18",x"FE",x"01",
		x"20",x"06",x"DD",x"21",x"4B",x"66",x"18",x"0E",x"FE",x"02",x"20",x"06",x"DD",x"21",x"6B",x"66",
		x"18",x"04",x"DD",x"21",x"8B",x"66",x"CD",x"D2",x"00",x"DD",x"21",x"AB",x"66",x"CD",x"D2",x"00",
		x"3E",x"20",x"CD",x"FC",x"00",x"01",x"00",x"00",x"3E",x"01",x"32",x"6E",x"80",x"3E",x"02",x"32",
		x"8C",x"80",x"3A",x"6E",x"80",x"FE",x"00",x"20",x"F9",x"03",x"78",x"FE",x"02",x"20",x"E9",x"79",
		x"FE",x"58",x"20",x"E4",x"CD",x"69",x"65",x"C9",x"C3",x"00",x"6A",x"DD",x"E5",x"DD",x"21",x"00",
		x"85",x"06",x"A8",x"0E",x"06",x"26",x"21",x"79",x"FE",x"00",x"28",x"32",x"FE",x"04",x"20",x"02",
		x"06",x"B4",x"DD",x"70",x"00",x"DD",x"36",x"01",x"24",x"DD",x"74",x"02",x"DD",x"36",x"03",x"20",
		x"04",x"11",x"08",x"00",x"DD",x"19",x"DD",x"70",x"00",x"DD",x"36",x"01",x"24",x"DD",x"74",x"02",
		x"DD",x"36",x"03",x"40",x"DD",x"19",x"04",x"0D",x"3E",x"20",x"84",x"67",x"18",x"C9",x"DD",x"E1",
		x"E1",x"D1",x"C1",x"C9",x"C5",x"D5",x"E5",x"3A",x"64",x"88",x"F6",x"80",x"32",x"64",x"88",x"21",
		x"1A",x"0F",x"11",x"00",x"88",x"01",x"0A",x"00",x"ED",x"B0",x"21",x"FF",x"0F",x"22",x"42",x"8C",
		x"21",x"0F",x"00",x"22",x"44",x"8C",x"21",x"AF",x"00",x"22",x"46",x"8C",x"21",x"0F",x"08",x"22",
		x"48",x"8C",x"21",x"AD",x"0F",x"11",x"4A",x"8C",x"01",x"06",x"00",x"ED",x"B0",x"3A",x"00",x"88",
		x"E6",x"7F",x"32",x"00",x"88",x"E1",x"D1",x"C1",x"C9",x"C5",x"D5",x"E5",x"3A",x"00",x"88",x"F6",
		x"80",x"32",x"00",x"88",x"11",x"42",x"8C",x"21",x"42",x"D5",x"01",x"0E",x"00",x"ED",x"B0",x"3A",
		x"64",x"88",x"E6",x"7F",x"32",x"64",x"88",x"3E",x"00",x"CD",x"F6",x"4F",x"E1",x"D1",x"C1",x"C9",
		x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",x"DD",x"CB",x"00",x"76",x"CA",x"22",x"66",x"DD",
		x"7E",x"03",x"FE",x"00",x"C2",x"22",x"66",x"DD",x"7E",x"04",x"FE",x"00",x"CA",x"22",x"66",x"FE",
		x"01",x"20",x"45",x"DD",x"46",x"01",x"DD",x"4E",x"02",x"CD",x"DE",x"00",x"E5",x"FD",x"E1",x"3A",
		x"AC",x"81",x"26",x"00",x"6F",x"29",x"29",x"29",x"11",x"D3",x"66",x"19",x"7E",x"FD",x"77",x"E0",
		x"23",x"7E",x"FD",x"77",x"E1",x"23",x"7E",x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77",x"01",x"11",
		x"00",x"04",x"FD",x"19",x"23",x"7E",x"FD",x"77",x"E0",x"23",x"7E",x"FD",x"77",x"E1",x"23",x"7E",
		x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77",x"01",x"DD",x"34",x"04",x"DD",x"7E",x"04",x"FE",x"1F",
		x"38",x"20",x"DD",x"36",x"04",x"00",x"DD",x"46",x"01",x"DD",x"4E",x"02",x"CD",x"DE",x"00",x"E5",
		x"FD",x"E1",x"FD",x"36",x"00",x"00",x"FD",x"36",x"01",x"00",x"FD",x"36",x"E1",x"00",x"FD",x"36",
		x"E0",x"00",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",x"C9",x"13",x"09",x"31",x"05",x"43",
		x"00",x"4F",x"00",x"49",x"00",x"4E",x"00",x"02",x"FF",x"00",x"00",x"31",x"05",x"43",x"00",x"52",
		x"00",x"45",x"00",x"44",x"00",x"49",x"00",x"54",x"00",x"FF",x"FF",x"13",x"09",x"31",x"05",x"43",
		x"00",x"4F",x"00",x"49",x"00",x"4E",x"00",x"02",x"FF",x"00",x"00",x"32",x"05",x"43",x"00",x"52",
		x"00",x"45",x"00",x"44",x"00",x"49",x"00",x"54",x"00",x"FF",x"FF",x"13",x"09",x"31",x"05",x"43",
		x"00",x"4F",x"00",x"49",x"00",x"4E",x"00",x"02",x"FF",x"00",x"00",x"33",x"05",x"43",x"00",x"52",
		x"00",x"45",x"00",x"44",x"00",x"49",x"00",x"54",x"00",x"FF",x"FF",x"13",x"09",x"31",x"05",x"43",
		x"00",x"4F",x"00",x"49",x"00",x"4E",x"00",x"02",x"FF",x"00",x"00",x"36",x"05",x"43",x"00",x"52",
		x"00",x"45",x"00",x"44",x"00",x"49",x"00",x"54",x"00",x"FF",x"FF",x"1C",x"07",x"3A",x"05",x"3B",
		x"05",x"31",x"05",x"39",x"05",x"38",x"05",x"34",x"05",x"00",x"00",x"54",x"0F",x"45",x"0F",x"48",
		x"0F",x"4B",x"0F",x"41",x"0F",x"4E",x"0F",x"00",x"00",x"4C",x"05",x"54",x"05",x"44",x"05",x"2E",
		x"05",x"FF",x"FF",x"80",x"81",x"82",x"83",x"15",x"15",x"15",x"15",x"90",x"91",x"92",x"93",x"15",
		x"15",x"15",x"15",x"94",x"95",x"96",x"97",x"15",x"15",x"15",x"15",x"98",x"99",x"9A",x"9B",x"15",
		x"15",x"15",x"15",x"9C",x"9D",x"9E",x"9F",x"15",x"15",x"15",x"15",x"F5",x"E5",x"21",x"00",x"00",
		x"22",x"9F",x"80",x"22",x"A1",x"80",x"22",x"A3",x"80",x"3A",x"6D",x"67",x"32",x"00",x"85",x"3A",
		x"6E",x"67",x"32",x"01",x"85",x"E1",x"F1",x"C9",x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD",x"E5",
		x"DD",x"21",x"9F",x"80",x"DD",x"7E",x"00",x"FE",x"0E",x"38",x"36",x"FD",x"21",x"6D",x"67",x"ED",
		x"5B",x"A0",x"80",x"B7",x"FD",x"19",x"FD",x"7E",x"00",x"FE",x"FF",x"20",x"0C",x"FD",x"21",x"6D",
		x"67",x"DD",x"36",x"01",x"00",x"DD",x"36",x"02",x"00",x"FD",x"7E",x"00",x"32",x"00",x"85",x"FD",
		x"7E",x"01",x"32",x"01",x"85",x"DD",x"36",x"00",x"00",x"2A",x"A0",x"80",x"23",x"23",x"22",x"A0",
		x"80",x"DD",x"34",x"00",x"FD",x"E1",x"DD",x"E1",x"E1",x"D1",x"C1",x"F1",x"C9",x"31",x"00",x"32",
		x"00",x"31",x"00",x"32",x"80",x"31",x"00",x"33",x"00",x"31",x"00",x"33",x"00",x"FF",x"FF",x"FF",
		x"FF",x"DD",x"21",x"10",x"85",x"3A",x"02",x"89",x"FE",x"FF",x"28",x"3E",x"3E",x"FF",x"32",x"02",
		x"89",x"DD",x"36",x"00",x"18",x"DD",x"36",x"01",x"0B",x"DD",x"36",x"04",x"00",x"DD",x"36",x"05",
		x"00",x"DD",x"36",x"06",x"00",x"DD",x"36",x"07",x"00",x"3A",x"9B",x"81",x"3C",x"32",x"9B",x"81",
		x"FE",x"08",x"38",x"02",x"3E",x"07",x"4F",x"0D",x"06",x"10",x"79",x"FE",x"00",x"28",x"07",x"78",
		x"C6",x"10",x"47",x"0D",x"18",x"F4",x"78",x"32",x"03",x"89",x"3A",x"13",x"85",x"FE",x"F0",x"CA",
		x"FE",x"67",x"3A",x"12",x"85",x"FE",x"78",x"28",x"16",x"30",x"08",x"3C",x"FE",x"78",x"28",x"09",
		x"3C",x"18",x"06",x"3D",x"FE",x"78",x"28",x"01",x"3D",x"32",x"12",x"85",x"C3",x"7A",x"68",x"3A",
		x"13",x"85",x"3C",x"FE",x"F0",x"28",x"01",x"3C",x"32",x"13",x"85",x"C3",x"7A",x"68",x"3A",x"04",
		x"89",x"FE",x"01",x"28",x"24",x"3A",x"03",x"89",x"47",x"3A",x"12",x"85",x"B8",x"28",x"08",x"3D",
		x"B8",x"28",x"04",x"3D",x"B8",x"20",x"0C",x"47",x"3E",x"01",x"32",x"04",x"89",x"3E",x"30",x"32",
		x"05",x"89",x"78",x"32",x"12",x"85",x"C3",x"7A",x"68",x"3A",x"05",x"89",x"3D",x"32",x"05",x"89",
		x"FE",x"00",x"C2",x"7A",x"68",x"3E",x"1F",x"CD",x"FC",x"00",x"21",x"00",x"00",x"22",x"10",x"85",
		x"DD",x"46",x"02",x"DD",x"4E",x"03",x"CD",x"DE",x"00",x"E5",x"FD",x"E1",x"FD",x"36",x"00",x"0E",
		x"FD",x"36",x"01",x"0F",x"FD",x"36",x"E0",x"0C",x"FD",x"36",x"E1",x"0D",x"11",x"00",x"04",x"B7",
		x"FD",x"19",x"FD",x"36",x"00",x"00",x"FD",x"36",x"01",x"00",x"FD",x"36",x"E0",x"00",x"FD",x"36",
		x"E1",x"00",x"3E",x"00",x"32",x"02",x"89",x"32",x"88",x"80",x"C9",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"C5",x"D5",x"E5",x"CD",x"CF",x"00",x"10",x"6A",x"02",x"C3",x"DB",x"64",x"00",x"00",x"00",x"00",
		x"20",x"6A",x"60",x"6A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"04",x"22",x"14",x"20",x"14",x"26",x"14",x"24",x"14",x"2A",x"14",x"28",x"14",x"2E",x"14",
		x"2C",x"14",x"32",x"14",x"30",x"14",x"36",x"14",x"34",x"14",x"3A",x"14",x"38",x"14",x"3E",x"14",
		x"3C",x"14",x"42",x"14",x"40",x"14",x"46",x"14",x"44",x"14",x"4A",x"14",x"48",x"14",x"4E",x"14",
		x"4C",x"14",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0D",x"04",x"23",x"14",x"21",x"14",x"27",x"14",x"25",x"14",x"2B",x"14",x"29",x"14",x"2F",x"14",
		x"2D",x"14",x"33",x"14",x"31",x"14",x"37",x"14",x"35",x"14",x"3B",x"14",x"39",x"14",x"3F",x"14",
		x"3D",x"14",x"43",x"14",x"41",x"14",x"47",x"14",x"45",x"14",x"4B",x"14",x"49",x"14",x"4F",x"14",
		x"4D",x"14",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"18",x"08",x"06",x"10",x"1E",x"00",x"02",x"05",x"05",x"15",x"02",x"11",x"03",x"01",x"04",x"11",
		x"05",x"01",x"05",x"11",x"04",x"05",x"03",x"15",x"0A",x"05",x"04",x"15",x"04",x"05",x"05",x"15",
		x"06",x"05",x"03",x"01",x"42",x"09",x"01",x"08",x"01",x"00",x"45",x"06",x"02",x"16",x"3A",x"02",
		x"02",x"16",x"28",x"02",x"02",x"15",x"27",x"05",x"15",x"00",x"02",x"15",x"70",x"05",x"02",x"16",
		x"33",x"06",x"02",x"10",x"0E",x"0A",x"30",x"00",x"02",x"10",x"05",x"00",x"02",x"10",x"10",x"00",
		x"02",x"10",x"05",x"00",x"02",x"10",x"60",x"00",x"0A",x"01",x"0A",x"02",x"02",x"16",x"21",x"06",
		x"02",x"10",x"10",x"01",x"2D",x"0A",x"40",x"09",x"02",x"16",x"10",x"06",x"02",x"16",x"02",x"06",
		x"02",x"16",x"35",x"06",x"70",x"00",x"02",x"14",x"42",x"04",x"30",x"05",x"25",x"00",x"53",x"09",
		x"53",x"0A",x"0A",x"00",x"98",x"00",x"30",x"02",x"02",x"16",x"20",x"06",x"05",x"05",x"10",x"06",
		x"1C",x"05",x"02",x"15",x"24",x"08",x"02",x"10",x"05",x"00",x"02",x"10",x"10",x"00",x"02",x"10",
		x"05",x"00",x"02",x"10",x"10",x"00",x"02",x"10",x"05",x"00",x"02",x"10",x"10",x"00",x"05",x"01",
		x"02",x"11",x"20",x"01",x"02",x"11",x"40",x"01",x"42",x"08",x"27",x"02",x"02",x"16",x"35",x"06",
		x"30",x"08",x"60",x"01",x"02",x"10",x"20",x"04",x"10",x"06",x"10",x"05",x"18",x"04",x"02",x"16",
		x"30",x"06",x"02",x"15",x"30",x"05",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"06",x"05",
		x"1E",x"05",x"0E",x"02",x"02",x"10",x"1E",x"00",x"03",x"05",x"03",x"15",x"03",x"05",x"10",x"05",
		x"01",x"00",x"10",x"16",x"10",x"06",x"10",x"16",x"05",x"06",x"05",x"16",x"05",x"06",x"05",x"16",
		x"30",x"05",x"10",x"00",x"03",x"10",x"28",x"00",x"08",x"02",x"05",x"16",x"05",x"06",x"05",x"16",
		x"05",x"02",x"05",x"16",x"02",x"06",x"02",x"16",x"02",x"06",x"02",x"16",x"02",x"06",x"02",x"16",
		x"05",x"06",x"05",x"16",x"05",x"06",x"02",x"16",x"02",x"06",x"02",x"16",x"02",x"06",x"02",x"16",
		x"02",x"06",x"02",x"16",x"02",x"06",x"02",x"16",x"05",x"06",x"05",x"16",x"08",x"00",x"02",x"15",
		x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"15",x"02",x"05",
		x"80",x"05",x"50",x"00",x"45",x"02",x"40",x"00",x"02",x"10",x"53",x"00",x"05",x"15",x"05",x"05",
		x"02",x"15",x"05",x"06",x"02",x"16",x"02",x"06",x"03",x"16",x"03",x"06",x"03",x"16",x"03",x"06",
		x"03",x"16",x"03",x"06",x"03",x"16",x"03",x"06",x"03",x"16",x"18",x"06",x"32",x"08",x"01",x"00",
		x"02",x"10",x"2A",x"04",x"02",x"15",x"35",x"05",x"1C",x"00",x"05",x"16",x"05",x"06",x"05",x"16",
		x"05",x"02",x"03",x"12",x"10",x"00",x"03",x"02",x"02",x"05",x"02",x"05",x"02",x"05",x"18",x"01",
		x"50",x"00",x"02",x"10",x"13",x"00",x"02",x"15",x"05",x"00",x"3D",x"09",x"60",x"00",x"30",x"01",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3A",x"06",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",
		x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",x"02",x"05",x"02",x"15",
		x"02",x"05",x"02",x"15",x"02",x"05",x"40",x"01",x"30",x"00",x"40",x"02",x"02",x"10",x"10",x"04",
		x"18",x"05",x"02",x"15",x"20",x"01",x"10",x"02",x"02",x"10",x"20",x"04",x"02",x"10",x"05",x"05",
		x"05",x"15",x"05",x"05",x"05",x"15",x"10",x"05",x"20",x"02",x"20",x"08",x"02",x"10",x"20",x"04",
		x"02",x"10",x"10",x"01",x"20",x"00",x"02",x"10",x"02",x"00",x"02",x"10",x"05",x"00",x"02",x"10",
		x"02",x"00",x"02",x"10",x"05",x"00",x"02",x"10",x"02",x"00",x"02",x"10",x"05",x"00",x"02",x"10",
		x"02",x"00",x"02",x"10",x"05",x"00",x"15",x"0A",x"15",x"08",x"18",x"01",x"44",x"00",x"0C",x"01",
		x"28",x"02",x"22",x"0A",x"10",x"08",x"02",x"14",x"16",x"04",x"13",x"06",x"02",x"12",x"10",x"02",
		x"10",x"01",x"02",x"00",x"10",x"01",x"0E",x"00",x"02",x"14",x"02",x"06",x"02",x"16",x"02",x"06",
		x"02",x"16",x"02",x"06",x"02",x"16",x"12",x"06",x"40",x"00",x"44",x"01",x"10",x"00",x"02",x"10",
		x"40",x"04",x"02",x"16",x"0A",x"06",x"33",x"08",x"02",x"10",x"20",x"04",x"1E",x"05",x"02",x"10",
		x"05",x"06",x"05",x"16",x"05",x"06",x"05",x"16",x"05",x"06",x"05",x"16",x"05",x"06",x"05",x"16",
		x"05",x"06",x"05",x"16",x"05",x"06",x"05",x"16",x"10",x"06",x"08",x"00",x"05",x"15",x"05",x"05",
		x"05",x"15",x"05",x"05",x"05",x"15",x"05",x"05",x"10",x"08",x"10",x"0A",x"10",x"00",x"10",x"01",
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"2C",x"70",
		x"58",x"70",x"84",x"70",x"94",x"70",x"C0",x"70",x"D0",x"70",x"C0",x"70",x"F8",x"70",x"08",x"71",
		x"18",x"71",x"44",x"71",x"54",x"71",x"6C",x"71",x"7C",x"71",x"A8",x"71",x"09",x"06",x"12",x"0B",
		x"10",x"0B",x"12",x"1B",x"10",x"1B",x"12",x"1B",x"10",x"1B",x"12",x"1B",x"10",x"1B",x"12",x"1B",
		x"10",x"1B",x"12",x"1B",x"10",x"1B",x"12",x"1B",x"10",x"1B",x"12",x"1B",x"10",x"1B",x"12",x"1B",
		x"10",x"1B",x"1E",x"0B",x"1C",x"0B",x"FF",x"FF",x"0A",x"06",x"13",x"0B",x"11",x"0B",x"13",x"1B",
		x"11",x"1B",x"13",x"1B",x"11",x"1B",x"13",x"1B",x"11",x"1B",x"13",x"1B",x"11",x"1B",x"13",x"1B",
		x"11",x"1B",x"13",x"1B",x"11",x"1B",x"13",x"1B",x"11",x"1B",x"13",x"1B",x"11",x"1B",x"1F",x"0B",
		x"1D",x"0B",x"FF",x"FF",x"0B",x"06",x"16",x"1B",x"14",x"1B",x"10",x"FF",x"00",x"00",x"1E",x"1B",
		x"1C",x"1B",x"FF",x"FF",x"0C",x"06",x"17",x"1B",x"15",x"1B",x"00",x"00",x"59",x"00",x"4F",x"00",
		x"55",x"00",x"3D",x"00",x"56",x"00",x"45",x"00",x"00",x"00",x"47",x"00",x"4F",x"00",x"54",x"00",
		x"54",x"00",x"45",x"00",x"4E",x"00",x"00",x"00",x"00",x"00",x"1F",x"1B",x"1D",x"1B",x"FF",x"FF",
		x"0D",x"06",x"16",x"1B",x"14",x"1B",x"10",x"FF",x"00",x"00",x"1E",x"1B",x"1C",x"1B",x"FF",x"FF",
		x"0E",x"06",x"17",x"1B",x"15",x"1B",x"04",x"FF",x"00",x"00",x"46",x"00",x"49",x"00",x"52",x"00",
		x"45",x"00",x"00",x"00",x"42",x"00",x"4F",x"00",x"4D",x"00",x"42",x"00",x"53",x"00",x"2E",x"00",
		x"00",x"00",x"1F",x"1B",x"1D",x"1B",x"FF",x"FF",x"0F",x"06",x"16",x"1B",x"14",x"1B",x"10",x"FF",
		x"00",x"00",x"1E",x"1B",x"1C",x"1B",x"FF",x"FF",x"10",x"06",x"17",x"1B",x"15",x"1B",x"10",x"FF",
		x"00",x"00",x"1F",x"1B",x"1D",x"1B",x"FF",x"FF",x"11",x"06",x"16",x"1B",x"14",x"1B",x"00",x"00",
		x"53",x"05",x"50",x"05",x"45",x"05",x"43",x"05",x"49",x"05",x"41",x"05",x"4C",x"05",x"00",x"00",
		x"42",x"05",x"4F",x"05",x"4E",x"05",x"55",x"05",x"53",x"05",x"00",x"00",x"00",x"00",x"1E",x"1B",
		x"1C",x"1B",x"FF",x"FF",x"12",x"06",x"17",x"1B",x"15",x"1B",x"10",x"FF",x"00",x"00",x"1F",x"1B",
		x"1D",x"1B",x"FF",x"FF",x"13",x"06",x"16",x"1B",x"14",x"1B",x"0A",x"FF",x"00",x"00",x"3E",x"05",
		x"3C",x"05",x"04",x"FF",x"00",x"00",x"1E",x"1B",x"1C",x"1B",x"FF",x"FF",x"14",x"06",x"17",x"1B",
		x"15",x"1B",x"10",x"FF",x"00",x"00",x"1F",x"1B",x"1D",x"1B",x"FF",x"FF",x"15",x"06",x"16",x"0B",
		x"14",x"0B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",
		x"18",x"1B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",x"18",x"1B",x"1A",x"1B",
		x"18",x"1B",x"1A",x"0B",x"18",x"0B",x"FF",x"FF",x"16",x"06",x"17",x"0B",x"15",x"0B",x"1B",x"1B",
		x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"1B",
		x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"1B",x"19",x"1B",x"1B",x"0B",
		x"19",x"0B",x"FF",x"FF",x"E4",x"71",x"EC",x"71",x"FC",x"71",x"04",x"72",x"14",x"72",x"1C",x"72",
		x"2C",x"72",x"34",x"72",x"0E",x"09",x"32",x"0F",x"30",x"0F",x"FF",x"FF",x"13",x"0B",x"00",x"00",
		x"31",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",x"FF",x"FF",x"0E",x"09",x"32",x"0F",
		x"31",x"0F",x"FF",x"FF",x"13",x"0B",x"00",x"00",x"32",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",
		x"30",x"0F",x"FF",x"FF",x"0E",x"09",x"32",x"0F",x"32",x"0F",x"FF",x"FF",x"13",x"0B",x"00",x"00",
		x"33",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",x"FF",x"FF",x"0E",x"09",x"32",x"0F",
		x"33",x"0F",x"FF",x"FF",x"13",x"0B",x"00",x"00",x"35",x"0F",x"30",x"0F",x"30",x"0F",x"30",x"0F",
		x"30",x"0F",x"FF",x"FF",x"13",x"0B",x"82",x"89",x"0F",x"06",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0A",x"73",x"1C",x"73",x"28",x"73",x"38",x"73",x"44",x"73",x"08",x"11",x"60",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"0B",x"08",x"60",x"09",
		x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"14",x"0E",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"17",x"05",x"60",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"1A",x"12",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"6E",x"73",x"82",x"73",x"8E",x"73",
		x"9A",x"73",x"A6",x"73",x"B2",x"73",x"BE",x"73",x"CA",x"73",x"D6",x"73",x"E2",x"73",x"08",x"0C",
		x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",
		x"FF",x"FF",x"0C",x"08",x"64",x"09",x"0E",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"0D",x"08",
		x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0E",x"08",x"67",x"09",x"0E",x"FF",
		x"00",x"00",x"67",x"09",x"FF",x"FF",x"0F",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",
		x"FF",x"FF",x"10",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"11",x"08",
		x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"12",x"08",x"67",x"09",x"0E",x"FF",
		x"00",x"00",x"67",x"09",x"FF",x"FF",x"13",x"08",x"65",x"09",x"0E",x"FF",x"00",x"00",x"65",x"09",
		x"FF",x"FF",x"17",x"0C",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"63",x"09",x"61",x"09",x"FF",x"FF",x"08",x"74",x"16",x"74",x"2C",x"74",x"3C",x"74",x"42",x"74",
		x"48",x"74",x"4E",x"74",x"54",x"74",x"5A",x"74",x"08",x"0F",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"61",x"09",x"FF",x"FF",x"0B",x"02",x"6C",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"0E",x"14",x"68",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"0F",x"14",x"66",x"09",
		x"FF",x"FF",x"10",x"14",x"67",x"09",x"FF",x"FF",x"11",x"14",x"66",x"09",x"FF",x"FF",x"12",x"14",
		x"67",x"09",x"FF",x"FF",x"13",x"14",x"66",x"09",x"FF",x"FF",x"14",x"08",x"60",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"6B",x"09",x"FF",x"FF",x"90",x"74",x"9C",x"74",x"A8",x"74",x"B4",x"74",
		x"C0",x"74",x"CC",x"74",x"EC",x"74",x"0C",x"75",x"18",x"75",x"24",x"75",x"30",x"75",x"3C",x"75",
		x"06",x"0B",x"64",x"09",x"08",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"07",x"0B",x"66",x"09",
		x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"08",x"0B",x"67",x"09",x"08",x"FF",x"00",x"00",
		x"67",x"09",x"FF",x"FF",x"09",x"0B",x"66",x"09",x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",
		x"0A",x"0B",x"67",x"09",x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0B",x"06",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"6B",x"09",x"08",x"FF",x"00",x"00",x"6A",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"14",x"06",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"69",x"09",x"08",x"FF",x"00",x"00",x"68",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"15",x"0B",x"66",x"09",
		x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"16",x"0B",x"67",x"09",x"08",x"FF",x"00",x"00",
		x"67",x"09",x"FF",x"FF",x"17",x"0B",x"66",x"09",x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",
		x"18",x"0B",x"67",x"09",x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"19",x"0B",x"65",x"09",
		x"08",x"FF",x"00",x"00",x"65",x"09",x"FF",x"FF",x"50",x"75",x"74",x"75",x"90",x"75",x"B4",x"75",
		x"08",x"05",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"05",x"FF",x"00",x"00",x"60",x"09",
		x"62",x"09",x"63",x"09",x"61",x"09",x"05",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"0E",x"09",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",
		x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",
		x"14",x"05",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"05",x"FF",x"00",x"00",x"60",x"09",
		x"62",x"09",x"63",x"09",x"61",x"09",x"05",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"1A",x"09",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",
		x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",
		x"D8",x"75",x"E4",x"75",x"04",x"76",x"24",x"76",x"08",x"0E",x"60",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"0E",x"08",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"11",x"08",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"17",x"0E",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",
		x"34",x"76",x"50",x"76",x"08",x"06",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",
		x"0A",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",
		x"17",x"06",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"0A",x"FF",x"00",x"00",
		x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"72",x"76",x"8E",x"76",
		x"9A",x"76",x"08",x"09",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"04",x"FF",
		x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"14",x"0E",
		x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"17",x"05",x"60",x"09",x"62",x"09",
		x"63",x"09",x"61",x"09",x"0E",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",
		x"FF",x"FF",x"CC",x"76",x"F0",x"76",x"FC",x"76",x"08",x"77",x"14",x"77",x"20",x"77",x"2C",x"77",
		x"38",x"77",x"44",x"77",x"50",x"77",x"5C",x"77",x"68",x"77",x"74",x"77",x"08",x"08",x"68",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"69",x"09",x"FF",x"FF",
		x"09",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0A",x"08",x"67",x"09",
		x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0B",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",
		x"66",x"09",x"FF",x"FF",x"0C",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"0D",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0E",x"08",x"67",x"09",
		x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0F",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",
		x"66",x"09",x"FF",x"FF",x"10",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"11",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"12",x"08",x"67",x"09",
		x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"13",x"08",x"65",x"09",x"0E",x"FF",x"00",x"00",
		x"65",x"09",x"FF",x"FF",x"14",x"0E",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",
		x"A0",x"77",x"AA",x"77",x"B0",x"77",x"B6",x"77",x"C2",x"77",x"D4",x"77",x"DA",x"77",x"E0",x"77",
		x"EC",x"77",x"04",x"78",x"10",x"78",x"16",x"78",x"1C",x"78",x"3A",x"78",x"40",x"78",x"46",x"78",
		x"05",x"0E",x"68",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"06",x"0E",x"66",x"09",x"FF",x"FF",
		x"07",x"0E",x"67",x"09",x"FF",x"FF",x"08",x"0E",x"6A",x"09",x"62",x"09",x"63",x"09",x"61",x"09",
		x"FF",x"FF",x"0B",x"0B",x"60",x"09",x"62",x"09",x"63",x"09",x"6E",x"09",x"63",x"09",x"62",x"09",
		x"61",x"09",x"FF",x"FF",x"0C",x"0E",x"66",x"09",x"FF",x"FF",x"0D",x"0E",x"67",x"09",x"FF",x"FF",
		x"0E",x"0E",x"6A",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"11",x"0E",x"68",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"61",x"09",x"FF",x"FF",x"14",x"0E",x"6A",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",
		x"12",x"0E",x"66",x"09",x"FF",x"FF",x"13",x"0E",x"67",x"09",x"FF",x"FF",x"17",x"05",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"6E",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"18",x"0E",x"66",x"09",x"FF",x"FF",
		x"19",x"0E",x"67",x"09",x"FF",x"FF",x"1A",x"0E",x"6A",x"09",x"62",x"09",x"63",x"09",x"61",x"09",
		x"FF",x"FF",x"58",x"78",x"78",x"78",x"94",x"78",x"0B",x"02",x"6C",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"61",x"09",x"10",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"6D",x"09",x"FF",x"FF",x"11",x"06",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"61",x"09",x"0A",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"61",x"09",x"FF",x"FF",x"17",x"09",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",
		x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",
		x"D0",x"78",x"F2",x"78",x"FE",x"78",x"0A",x"79",x"16",x"79",x"22",x"79",x"2E",x"79",x"3A",x"79",
		x"46",x"79",x"52",x"79",x"5E",x"79",x"6A",x"79",x"76",x"79",x"82",x"79",x"8E",x"79",x"9A",x"79",
		x"08",x"08",x"68",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"61",x"09",x"03",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"69",x"09",
		x"FF",x"FF",x"09",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0A",x"08",
		x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0B",x"08",x"66",x"09",x"0E",x"FF",
		x"00",x"00",x"66",x"09",x"FF",x"FF",x"0C",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",
		x"FF",x"FF",x"0D",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0E",x"08",
		x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0F",x"08",x"66",x"09",x"0E",x"FF",
		x"00",x"00",x"66",x"09",x"FF",x"FF",x"10",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",
		x"FF",x"FF",x"11",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"12",x"08",
		x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"13",x"08",x"66",x"09",x"0E",x"FF",
		x"00",x"00",x"66",x"09",x"FF",x"FF",x"14",x"08",x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",
		x"FF",x"FF",x"15",x"08",x"66",x"09",x"0E",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"16",x"08",
		x"67",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"17",x"08",x"6A",x"09",x"62",x"09",
		x"63",x"09",x"61",x"09",x"03",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"6B",x"09",x"FF",x"FF",x"E8",x"79",x"00",x"7A",
		x"06",x"7A",x"0C",x"7A",x"18",x"7A",x"24",x"7A",x"30",x"7A",x"3C",x"7A",x"42",x"7A",x"48",x"7A",
		x"60",x"7A",x"6C",x"7A",x"78",x"7A",x"90",x"7A",x"96",x"7A",x"9C",x"7A",x"A8",x"7A",x"B4",x"7A",
		x"C0",x"7A",x"CC",x"7A",x"D2",x"7A",x"D8",x"7A",x"05",x"08",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"69",x"09",x"FF",x"FF",
		x"06",x"11",x"66",x"09",x"FF",x"FF",x"07",x"11",x"67",x"09",x"FF",x"FF",x"08",x"11",x"66",x"09",
		x"08",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"09",x"11",x"67",x"09",x"08",x"FF",x"00",x"00",
		x"66",x"09",x"FF",x"FF",x"0A",x"11",x"66",x"09",x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"0B",x"11",x"65",x"09",x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"0C",x"1A",x"67",x"09",
		x"FF",x"FF",x"0D",x"1A",x"66",x"09",x"FF",x"FF",x"0E",x"05",x"68",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"0E",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"0F",x"05",x"66",x"09",x"14",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"10",x"05",x"67",x"09",
		x"14",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"11",x"05",x"66",x"09",x"0E",x"FF",x"00",x"00",
		x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"6B",x"09",x"FF",x"FF",
		x"12",x"05",x"67",x"09",x"FF",x"FF",x"13",x"05",x"66",x"09",x"FF",x"FF",x"14",x"05",x"67",x"09",
		x"08",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"15",x"05",x"66",x"09",x"08",x"FF",x"00",x"00",
		x"66",x"09",x"FF",x"FF",x"16",x"05",x"67",x"09",x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"17",x"05",x"65",x"09",x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"18",x"0E",x"67",x"09",
		x"FF",x"FF",x"19",x"0E",x"66",x"09",x"FF",x"FF",x"1A",x"0E",x"6A",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",
		x"FC",x"7A",x"0C",x"7B",x"1C",x"7B",x"2C",x"7B",x"3C",x"7B",x"4C",x"7B",x"08",x"18",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"6D",x"09",x"FF",x"FF",x"0B",x"02",x"6C",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"0E",x"18",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"6D",x"09",x"FF",x"FF",x"11",x"02",x"6C",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"14",x"18",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"6D",x"09",x"FF",x"FF",x"17",x"02",x"6C",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"FF",x"FF",x"7C",x"7B",x"98",x"7B",
		x"A4",x"7B",x"B0",x"7B",x"C8",x"7B",x"D4",x"7B",x"E0",x"7B",x"EC",x"7B",x"F8",x"7B",x"04",x"7C",
		x"10",x"7C",x"1C",x"7C",x"28",x"7C",x"40",x"7C",x"4C",x"7C",x"58",x"7C",x"05",x"09",x"60",x"09",
		x"62",x"09",x"63",x"09",x"62",x"09",x"61",x"09",x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",
		x"63",x"09",x"62",x"09",x"61",x"09",x"FF",x"FF",x"09",x"05",x"64",x"09",x"14",x"FF",x"00",x"00",
		x"64",x"09",x"FF",x"FF",x"0A",x"05",x"66",x"09",x"14",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",
		x"0B",x"05",x"67",x"09",x"08",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",
		x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",x"0C",x"05",x"66",x"09",x"14",x"FF",x"00",x"00",
		x"66",x"09",x"FF",x"FF",x"0D",x"05",x"65",x"09",x"14",x"FF",x"00",x"00",x"65",x"09",x"FF",x"FF",
		x"0E",x"0B",x"64",x"09",x"08",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"0F",x"0B",x"66",x"09",
		x"08",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"10",x"0B",x"67",x"09",x"08",x"FF",x"00",x"00",
		x"67",x"09",x"FF",x"FF",x"11",x"0B",x"65",x"09",x"08",x"FF",x"00",x"00",x"65",x"09",x"FF",x"FF",
		x"12",x"05",x"64",x"09",x"14",x"FF",x"00",x"00",x"64",x"09",x"FF",x"FF",x"13",x"05",x"66",x"09",
		x"14",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"14",x"05",x"67",x"09",x"08",x"FF",x"00",x"00",
		x"60",x"09",x"62",x"09",x"63",x"09",x"61",x"09",x"08",x"FF",x"00",x"00",x"67",x"09",x"FF",x"FF",
		x"15",x"05",x"66",x"09",x"14",x"FF",x"00",x"00",x"66",x"09",x"FF",x"FF",x"16",x"05",x"65",x"09",
		x"14",x"FF",x"00",x"00",x"65",x"09",x"FF",x"FF",x"1A",x"09",x"60",x"09",x"62",x"09",x"63",x"09",
		x"62",x"09",x"61",x"09",x"04",x"FF",x"00",x"00",x"60",x"09",x"62",x"09",x"63",x"09",x"62",x"09",
		x"61",x"09",x"FF",x"FF",x"94",x"7C",x"9E",x"7C",x"A8",x"7C",x"B2",x"7C",x"BC",x"7C",x"C0",x"7C",
		x"CB",x"7C",x"D5",x"7C",x"DF",x"7C",x"EA",x"7C",x"F4",x"7C",x"FE",x"7C",x"09",x"7D",x"13",x"7D",
		x"1D",x"7D",x"28",x"7D",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"00",x"73",x"05",x"C9",x"CD",x"32",
		x"7D",x"CD",x"CF",x"00",x"5A",x"73",x"0A",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"F6",x"73",
		x"09",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"78",x"74",x"0C",x"C9",x"CD",x"32",x"7D",x"C9",
		x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"48",x"75",x"04",x"00",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",
		x"00",x"D0",x"75",x"04",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"30",x"76",x"02",x"C9",x"CD",
		x"32",x"7D",x"CD",x"CF",x"00",x"6C",x"76",x"03",x"00",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",
		x"B2",x"76",x"0D",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"80",x"77",x"10",x"C9",x"CD",x"32",
		x"7D",x"CD",x"CF",x"00",x"52",x"78",x"03",x"00",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"B0",
		x"78",x"10",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"BC",x"79",x"16",x"C9",x"CD",x"32",x"7D",
		x"CD",x"CF",x"00",x"F0",x"7A",x"06",x"00",x"C9",x"CD",x"32",x"7D",x"CD",x"CF",x"00",x"5C",x"7B",
		x"10",x"C9",x"3E",x"09",x"CD",x"F0",x"4F",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F2",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"60",x"C0",x"7C",x"C0",x"94",x"C0",x"AC",x"C0",x"C4",x"C0",x"DC",x"C0",x"F4",x"C0",x"0C",x"C1",
		x"24",x"C1",x"3C",x"C1",x"54",x"C1",x"6E",x"C1",x"03",x"08",x"46",x"0F",x"41",x"0F",x"4E",x"0F",
		x"54",x"0F",x"41",x"0F",x"53",x"0F",x"54",x"0F",x"49",x"0F",x"43",x"0F",x"00",x"00",x"53",x"0F",
		x"43",x"0F",x"4F",x"0F",x"52",x"0F",x"45",x"0F",x"3F",x"0F",x"FF",x"FF",x"05",x"08",x"52",x"05",
		x"45",x"05",x"43",x"05",x"4F",x"05",x"52",x"05",x"44",x"05",x"00",x"00",x"59",x"05",x"4F",x"05",
		x"55",x"05",x"52",x"05",x"00",x"00",x"4E",x"05",x"41",x"05",x"4D",x"05",x"45",x"05",x"FF",x"FF",
		x"04",x"0A",x"42",x"06",x"45",x"06",x"53",x"06",x"54",x"06",x"00",x"00",x"50",x"06",x"4C",x"06",
		x"41",x"06",x"59",x"06",x"45",x"06",x"52",x"06",x"53",x"06",x"FF",x"FF",x"07",x"04",x"31",x"05",
		x"53",x"05",x"54",x"05",x"0F",x"FF",x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",
		x"44",x"05",x"FF",x"FF",x"09",x"04",x"32",x"05",x"4E",x"05",x"44",x"05",x"0F",x"FF",x"00",x"00",
		x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",x"44",x"05",x"FF",x"FF",x"0B",x"04",x"33",x"05",
		x"52",x"05",x"44",x"05",x"0F",x"FF",x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",
		x"44",x"05",x"FF",x"FF",x"0D",x"04",x"34",x"05",x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",
		x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",x"44",x"05",x"FF",x"FF",x"0F",x"04",x"35",x"05",
		x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",
		x"44",x"05",x"FF",x"FF",x"11",x"04",x"36",x"05",x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",
		x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",x"44",x"05",x"FF",x"FF",x"13",x"04",x"37",x"05",
		x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",
		x"44",x"05",x"FF",x"FF",x"15",x"04",x"38",x"05",x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",
		x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",x"44",x"05",x"FF",x"FF",x"17",x"04",x"39",x"05",
		x"54",x"05",x"48",x"05",x"0F",x"FF",x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",
		x"44",x"05",x"FF",x"FF",x"19",x"03",x"31",x"05",x"30",x"05",x"54",x"05",x"48",x"05",x"0F",x"FF",
		x"00",x"00",x"52",x"05",x"4F",x"05",x"55",x"05",x"4E",x"05",x"44",x"05",x"FF",x"FF",x"1C",x"07",
		x"3A",x"05",x"3B",x"05",x"31",x"05",x"39",x"05",x"38",x"05",x"34",x"05",x"00",x"00",x"54",x"0F",
		x"45",x"0F",x"48",x"0F",x"4B",x"0F",x"41",x"0F",x"4E",x"0F",x"00",x"00",x"4C",x"05",x"54",x"05",
		x"44",x"05",x"2E",x"05",x"FF",x"FF",x"AA",x"C1",x"B0",x"C1",x"B6",x"C1",x"BC",x"C1",x"C2",x"C1",
		x"C8",x"C1",x"CE",x"C1",x"D4",x"C1",x"DA",x"C1",x"E0",x"C1",x"07",x"08",x"00",x"81",x"0F",x"08",
		x"09",x"08",x"04",x"81",x"05",x"08",x"0B",x"08",x"08",x"81",x"05",x"08",x"0D",x"08",x"0C",x"81",
		x"05",x"08",x"0F",x"08",x"10",x"81",x"05",x"08",x"11",x"08",x"14",x"81",x"05",x"08",x"13",x"08",
		x"18",x"81",x"05",x"08",x"15",x"08",x"1C",x"81",x"05",x"08",x"17",x"08",x"20",x"81",x"05",x"08",
		x"19",x"08",x"24",x"81",x"05",x"08",x"32",x"81",x"3C",x"81",x"46",x"81",x"50",x"81",x"5A",x"81",
		x"64",x"81",x"6E",x"81",x"78",x"81",x"82",x"81",x"8C",x"81",x"0E",x"C2",x"14",x"C2",x"1A",x"C2",
		x"20",x"C2",x"26",x"C2",x"2C",x"C2",x"32",x"C2",x"38",x"C2",x"3E",x"C2",x"44",x"C2",x"07",x"1B",
		x"28",x"81",x"05",x"02",x"09",x"1B",x"29",x"81",x"05",x"02",x"0B",x"1B",x"2A",x"81",x"05",x"02",
		x"0D",x"1B",x"2B",x"81",x"05",x"02",x"0F",x"1B",x"2C",x"81",x"05",x"02",x"11",x"1B",x"2D",x"81",
		x"05",x"02",x"13",x"1B",x"2E",x"81",x"05",x"02",x"15",x"1B",x"2F",x"81",x"05",x"02",x"17",x"1B",
		x"30",x"81",x"05",x"02",x"19",x"1B",x"31",x"81",x"05",x"02",x"18",x"C0",x"3C",x"C0",x"64",x"C2",
		x"7C",x"C2",x"94",x"C2",x"AC",x"C2",x"C4",x"C2",x"DC",x"C2",x"F4",x"C2",x"0C",x"C3",x"24",x"C3",
		x"3C",x"C3",x"6E",x"C1",x"07",x"04",x"31",x"02",x"53",x"02",x"54",x"02",x"0F",x"FF",x"00",x"00",
		x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",x"44",x"01",x"FF",x"FF",x"09",x"04",x"32",x"00",
		x"4E",x"00",x"44",x"00",x"0F",x"FF",x"00",x"00",x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",
		x"44",x"01",x"FF",x"FF",x"0B",x"04",x"33",x"00",x"52",x"00",x"44",x"00",x"0F",x"FF",x"00",x"00",
		x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",x"44",x"01",x"FF",x"FF",x"0D",x"04",x"34",x"00",
		x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",
		x"44",x"01",x"FF",x"FF",x"0F",x"04",x"35",x"00",x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",
		x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",x"44",x"01",x"FF",x"FF",x"11",x"04",x"36",x"00",
		x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",
		x"44",x"01",x"FF",x"FF",x"13",x"04",x"37",x"00",x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",
		x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",x"44",x"01",x"FF",x"FF",x"15",x"04",x"38",x"00",
		x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",
		x"44",x"01",x"FF",x"FF",x"17",x"04",x"39",x"00",x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",
		x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",x"01",x"44",x"01",x"FF",x"FF",x"19",x"03",x"31",x"00",
		x"30",x"00",x"54",x"00",x"48",x"00",x"0F",x"FF",x"00",x"00",x"52",x"01",x"4F",x"01",x"55",x"01",
		x"4E",x"01",x"44",x"01",x"FF",x"FF",x"00",x"00",x"00",x"20",x"21",x"0E",x"FC",x"C3",x"04",x"C4",
		x"DE",x"F1",x"00",x"20",x"00",x"40",x"7C",x"0E",x"44",x"C4",x"4C",x"C4",x"83",x"F1",x"00",x"40",
		x"00",x"60",x"21",x"0C",x"8C",x"C4",x"94",x"C4",x"DE",x"F3",x"00",x"60",x"00",x"80",x"57",x"0C",
		x"D4",x"C4",x"DC",x"C4",x"A8",x"F3",x"00",x"C0",x"00",x"E0",x"2F",x"0B",x"1C",x"C5",x"24",x"C5",
		x"E0",x"F4",x"FF",x"FF",x"00",x"80",x"00",x"84",x"20",x"C4",x"28",x"C4",x"00",x"84",x"00",x"88",
		x"68",x"C4",x"70",x"C4",x"00",x"88",x"00",x"8C",x"B0",x"C4",x"B8",x"C4",x"00",x"8C",x"00",x"90",
		x"F8",x"C4",x"00",x"C5",x"00",x"90",x"00",x"98",x"40",x"C5",x"48",x"C5",x"FF",x"FF",x"01",x"03",
		x"50",x"01",x"55",x"01",x"53",x"01",x"48",x"01",x"00",x"00",x"42",x"01",x"55",x"01",x"54",x"01",
		x"54",x"01",x"4F",x"01",x"4E",x"01",x"00",x"00",x"46",x"01",x"4F",x"01",x"52",x"01",x"00",x"00",
		x"00",x"00",x"43",x"08",x"48",x"08",x"45",x"08",x"43",x"08",x"4B",x"08",x"FF",x"FF",x"03",x"03",
		x"52",x"03",x"4F",x"03",x"4D",x"03",x"00",x"00",x"30",x"03",x"FF",x"FF",x"03",x"0A",x"4F",x"03",
		x"4B",x"03",x"FF",x"FF",x"03",x"0A",x"45",x"02",x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",
		x"FF",x"FF",x"03",x"11",x"52",x"03",x"41",x"03",x"4D",x"03",x"00",x"00",x"30",x"03",x"FF",x"FF",
		x"03",x"18",x"4F",x"03",x"4B",x"03",x"FF",x"FF",x"03",x"18",x"45",x"02",x"52",x"02",x"52",x"02",
		x"4F",x"02",x"52",x"02",x"FF",x"FF",x"04",x"03",x"52",x"03",x"4F",x"03",x"4D",x"03",x"00",x"00",
		x"31",x"03",x"FF",x"FF",x"04",x"0A",x"4F",x"03",x"4B",x"03",x"FF",x"FF",x"04",x"0A",x"45",x"02",
		x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",x"FF",x"FF",x"04",x"11",x"52",x"03",x"41",x"03",
		x"4D",x"03",x"00",x"00",x"31",x"03",x"FF",x"FF",x"04",x"18",x"4F",x"03",x"4B",x"03",x"FF",x"FF",
		x"04",x"18",x"45",x"02",x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",x"FF",x"FF",x"05",x"03",
		x"52",x"03",x"4F",x"03",x"4D",x"03",x"00",x"00",x"32",x"03",x"FF",x"FF",x"05",x"0A",x"4F",x"03",
		x"4B",x"03",x"FF",x"FF",x"05",x"0A",x"45",x"02",x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",
		x"FF",x"FF",x"05",x"11",x"52",x"03",x"41",x"03",x"4D",x"03",x"00",x"00",x"32",x"03",x"FF",x"FF",
		x"05",x"18",x"4F",x"03",x"4B",x"03",x"FF",x"FF",x"05",x"18",x"45",x"02",x"52",x"02",x"52",x"02",
		x"4F",x"02",x"52",x"02",x"FF",x"FF",x"06",x"03",x"52",x"03",x"4F",x"03",x"4D",x"03",x"00",x"00",
		x"33",x"03",x"FF",x"FF",x"06",x"0A",x"4F",x"03",x"4B",x"03",x"FF",x"FF",x"06",x"0A",x"45",x"02",
		x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",x"FF",x"FF",x"06",x"11",x"52",x"03",x"41",x"03",
		x"4D",x"03",x"00",x"00",x"33",x"03",x"FF",x"FF",x"06",x"18",x"4F",x"03",x"4B",x"03",x"FF",x"FF",
		x"06",x"18",x"45",x"02",x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",x"FF",x"FF",x"07",x"03",
		x"52",x"03",x"4F",x"03",x"4D",x"03",x"00",x"00",x"34",x"03",x"FF",x"FF",x"07",x"0A",x"4F",x"03",
		x"4B",x"03",x"FF",x"FF",x"07",x"0A",x"45",x"02",x"52",x"02",x"52",x"02",x"4F",x"02",x"52",x"02",
		x"FF",x"FF",x"07",x"11",x"52",x"03",x"41",x"03",x"4D",x"03",x"00",x"00",x"34",x"03",x"FF",x"FF",
		x"07",x"18",x"4F",x"03",x"4B",x"03",x"FF",x"FF",x"07",x"18",x"45",x"02",x"52",x"02",x"52",x"02",
		x"4F",x"02",x"52",x"02",x"FF",x"FF",x"08",x"03",x"43",x"01",x"4F",x"01",x"4C",x"01",x"4F",x"01",
		x"52",x"01",x"28",x"01",x"52",x"01",x"47",x"01",x"42",x"01",x"57",x"01",x"29",x"01",x"FF",x"FF",
		x"16",x"03",x"31",x"03",x"50",x"03",x"FF",x"FF",x"18",x"03",x"32",x"03",x"50",x"03",x"FF",x"FF",
		x"1A",x"03",x"43",x"03",x"4F",x"03",x"49",x"03",x"4E",x"03",x"FF",x"FF",x"1C",x"03",x"44",x"03",
		x"49",x"03",x"50",x"03",x"00",x"00",x"53",x"03",x"57",x"03",x"28",x"03",x"31",x"03",x"29",x"03",
		x"FF",x"FF",x"1E",x"03",x"44",x"03",x"49",x"03",x"50",x"03",x"00",x"00",x"53",x"03",x"57",x"03",
		x"28",x"03",x"32",x"03",x"29",x"03",x"FF",x"FF",x"BE",x"C3",x"EE",x"C3",x"36",x"C4",x"7E",x"C4",
		x"C6",x"C4",x"0E",x"C5",x"12",x"C4",x"5A",x"C4",x"A2",x"C4",x"EA",x"C4",x"32",x"C5",x"56",x"C5",
		x"80",x"C5",x"70",x"C5",x"78",x"C5",x"8C",x"C5",x"A2",x"C5",x"E4",x"C5",x"F8",x"C5",x"0C",x"C6",
		x"20",x"C6",x"34",x"C6",x"16",x"0E",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",
		x"30",x"02",x"30",x"02",x"30",x"02",x"FF",x"FF",x"18",x"0E",x"30",x"05",x"30",x"05",x"30",x"05",
		x"30",x"05",x"30",x"05",x"30",x"02",x"30",x"02",x"30",x"02",x"FF",x"FF",x"1A",x"0E",x"30",x"05",
		x"30",x"05",x"30",x"05",x"30",x"05",x"00",x"05",x"00",x"05",x"00",x"05",x"00",x"05",x"FF",x"FF",
		x"1C",x"0E",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",
		x"30",x"05",x"FF",x"FF",x"1E",x"0E",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",x"30",x"05",
		x"30",x"05",x"30",x"05",x"30",x"05",x"FF",x"FF",x"01",x"13",x"43",x"08",x"48",x"08",x"41",x"08",
		x"4E",x"08",x"47",x"08",x"45",x"08",x"00",x"00",x"44",x"08",x"49",x"08",x"53",x"08",x"50",x"08",
		x"FF",x"FF",x"00",x"00",x"0F",x"00",x"0D",x"00",x"0B",x"00",x"09",x"00",x"07",x"00",x"05",x"00",
		x"03",x"00",x"00",x"00",x"F0",x"00",x"D0",x"00",x"B0",x"00",x"90",x"00",x"70",x"00",x"50",x"00",
		x"30",x"00",x"00",x"00",x"00",x"0F",x"00",x"0D",x"00",x"0B",x"00",x"09",x"00",x"07",x"00",x"05",
		x"00",x"03",x"00",x"00",x"FF",x"0F",x"DD",x"0D",x"BB",x"0B",x"99",x"09",x"77",x"07",x"55",x"05",
		x"33",x"03",x"B2",x"C6",x"DE",x"C6",x"0A",x"C7",x"36",x"C7",x"62",x"C7",x"8E",x"C7",x"BA",x"C7",
		x"E6",x"C7",x"0A",x"03",x"03",x"FF",x"05",x"0C",x"00",x"00",x"03",x"FF",x"06",x"0C",x"00",x"00",
		x"03",x"FF",x"07",x"0C",x"00",x"00",x"03",x"FF",x"08",x"0C",x"00",x"00",x"03",x"FF",x"09",x"0C",
		x"00",x"00",x"03",x"FF",x"0A",x"0C",x"00",x"00",x"03",x"FF",x"0B",x"0C",x"FF",x"FF",x"0B",x"03",
		x"03",x"FF",x"05",x"0C",x"00",x"00",x"03",x"FF",x"06",x"0C",x"00",x"00",x"03",x"FF",x"07",x"0C",
		x"00",x"00",x"03",x"FF",x"08",x"0C",x"00",x"00",x"03",x"FF",x"09",x"0C",x"00",x"00",x"03",x"FF",
		x"0A",x"0C",x"00",x"00",x"03",x"FF",x"0B",x"0C",x"FF",x"FF",x"0D",x"03",x"03",x"FF",x"05",x"0D",
		x"00",x"00",x"03",x"FF",x"06",x"0D",x"00",x"00",x"03",x"FF",x"07",x"0D",x"00",x"00",x"03",x"FF",
		x"08",x"0D",x"00",x"00",x"03",x"FF",x"09",x"0D",x"00",x"00",x"03",x"FF",x"0A",x"0D",x"00",x"00",
		x"03",x"FF",x"0B",x"0D",x"FF",x"FF",x"0E",x"03",x"03",x"FF",x"05",x"0D",x"00",x"00",x"03",x"FF",
		x"06",x"0D",x"00",x"00",x"03",x"FF",x"07",x"0D",x"00",x"00",x"03",x"FF",x"08",x"0D",x"00",x"00",
		x"03",x"FF",x"09",x"0D",x"00",x"00",x"03",x"FF",x"0A",x"0D",x"00",x"00",x"03",x"FF",x"0B",x"0D",
		x"FF",x"FF",x"10",x"03",x"03",x"FF",x"05",x"0E",x"00",x"00",x"03",x"FF",x"06",x"0E",x"00",x"00",
		x"03",x"FF",x"07",x"0E",x"00",x"00",x"03",x"FF",x"08",x"0E",x"00",x"00",x"03",x"FF",x"09",x"0E",
		x"00",x"00",x"03",x"FF",x"0A",x"0E",x"00",x"00",x"03",x"FF",x"0B",x"0E",x"FF",x"FF",x"11",x"03",
		x"03",x"FF",x"05",x"0E",x"00",x"00",x"03",x"FF",x"06",x"0E",x"00",x"00",x"03",x"FF",x"07",x"0E",
		x"00",x"00",x"03",x"FF",x"08",x"0E",x"00",x"00",x"03",x"FF",x"09",x"0E",x"00",x"00",x"03",x"FF",
		x"0A",x"0E",x"00",x"00",x"03",x"FF",x"0B",x"0E",x"FF",x"FF",x"13",x"03",x"03",x"FF",x"05",x"0F",
		x"00",x"00",x"03",x"FF",x"06",x"0F",x"00",x"00",x"03",x"FF",x"07",x"0F",x"00",x"00",x"03",x"FF",
		x"08",x"0F",x"00",x"00",x"03",x"FF",x"09",x"0F",x"00",x"00",x"03",x"FF",x"0A",x"0F",x"00",x"00",
		x"03",x"FF",x"0B",x"0F",x"FF",x"FF",x"14",x"03",x"03",x"FF",x"05",x"0F",x"00",x"00",x"03",x"FF",
		x"06",x"0F",x"00",x"00",x"03",x"FF",x"07",x"0F",x"00",x"00",x"03",x"FF",x"08",x"0F",x"00",x"00",
		x"03",x"FF",x"09",x"0F",x"00",x"00",x"03",x"FF",x"0A",x"0F",x"00",x"00",x"03",x"FF",x"0B",x"0F",
		x"FF",x"FF",x"1C",x"0C",x"43",x"06",x"52",x"06",x"45",x"06",x"44",x"06",x"49",x"06",x"54",x"06",
		x"FF",x"FF",x"1C",x"12",x"17",x"80",x"05",x"02",x"48",x"C8",x"60",x"C8",x"78",x"C8",x"90",x"C8",
		x"A8",x"C8",x"C0",x"C8",x"D8",x"C8",x"F0",x"C8",x"08",x"C9",x"20",x"C9",x"38",x"C9",x"50",x"C9",
		x"68",x"C9",x"80",x"C9",x"98",x"C9",x"B0",x"C9",x"42",x"52",x"62",x"72",x"83",x"84",x"85",x"86",
		x"03",x"04",x"05",x"06",x"10",x"20",x"30",x"77",x"67",x"57",x"38",x"28",x"18",x"80",x"70",x"60",
		x"32",x"42",x"52",x"73",x"74",x"75",x"76",x"77",x"25",x"24",x"23",x"13",x"14",x"15",x"16",x"17",
		x"63",x"64",x"65",x"71",x"51",x"41",x"31",x"11",x"23",x"13",x"03",x"04",x"05",x"06",x"07",x"87",
		x"86",x"85",x"84",x"83",x"73",x"63",x"66",x"56",x"36",x"26",x"51",x"41",x"10",x"00",x"70",x"80",
		x"51",x"52",x"53",x"68",x"67",x"66",x"85",x"75",x"65",x"25",x"15",x"05",x"28",x"27",x"26",x"31",
		x"32",x"33",x"10",x"11",x"12",x"70",x"71",x"72",x"71",x"72",x"73",x"75",x"76",x"77",x"51",x"52",
		x"53",x"35",x"36",x"37",x"11",x"12",x"13",x"15",x"16",x"17",x"55",x"56",x"57",x"31",x"32",x"33",
		x"81",x"71",x"61",x"21",x"11",x"01",x"23",x"33",x"53",x"63",x"85",x"75",x"65",x"25",x"15",x"05",
		x"27",x"37",x"57",x"67",x"78",x"88",x"18",x"08",x"56",x"57",x"58",x"54",x"64",x"74",x"36",x"37",
		x"38",x"34",x"24",x"14",x"11",x"21",x"31",x"51",x"61",x"71",x"06",x"07",x"08",x"86",x"87",x"88",
		x"56",x"66",x"76",x"36",x"26",x"16",x"64",x"74",x"84",x"24",x"14",x"04",x"61",x"71",x"81",x"21",
		x"11",x"01",x"08",x"18",x"28",x"68",x"78",x"88",x"06",x"16",x"26",x"35",x"34",x"33",x"53",x"54",
		x"55",x"66",x"76",x"86",x"51",x"61",x"70",x"80",x"31",x"21",x"10",x"00",x"28",x"38",x"58",x"68",
		x"51",x"61",x"71",x"02",x"03",x"04",x"15",x"16",x"17",x"31",x"21",x"11",x"82",x"83",x"84",x"75",
		x"76",x"77",x"55",x"54",x"53",x"33",x"34",x"35",x"23",x"22",x"21",x"11",x"12",x"13",x"16",x"26",
		x"36",x"54",x"64",x"74",x"66",x"67",x"68",x"82",x"72",x"62",x"86",x"87",x"88",x"70",x"60",x"50",
		x"01",x"11",x"21",x"14",x"24",x"34",x"16",x"26",x"36",x"56",x"66",x"76",x"54",x"64",x"74",x"61",
		x"71",x"81",x"52",x"42",x"32",x"50",x"40",x"30",x"51",x"52",x"53",x"64",x"65",x"66",x"22",x"23",
		x"24",x"35",x"36",x"37",x"70",x"71",x"72",x"86",x"87",x"88",x"10",x"11",x"12",x"06",x"07",x"08",
		x"72",x"73",x"74",x"14",x"15",x"16",x"26",x"27",x"28",x"43",x"42",x"41",x"22",x"12",x"02",x"57",
		x"67",x"77",x"84",x"83",x"82",x"60",x"61",x"62",x"00",x"01",x"02",x"13",x"14",x"15",x"74",x"75",
		x"76",x"86",x"87",x"88",x"28",x"18",x"08",x"60",x"70",x"80",x"73",x"83",x"82",x"52",x"42",x"32",
		x"55",x"56",x"57",x"24",x"23",x"22",x"85",x"84",x"83",x"70",x"60",x"50",x"30",x"20",x"10",x"03",
		x"04",x"05",x"62",x"63",x"64",x"37",x"36",x"35",x"18",x"30",x"48",x"60",x"78",x"90",x"A8",x"C0",
		x"D8",x"00",x"03",x"53",x"00",x"49",x"00",x"44",x"00",x"45",x"00",x"2D",x"00",x"4F",x"00",x"4E",
		x"00",x"45",x"00",x"FF",x"FF",x"1E",x"16",x"48",x"00",x"49",x"00",x"2D",x"00",x"53",x"00",x"43",
		x"00",x"4F",x"00",x"52",x"00",x"45",x"00",x"FF",x"FF",x"00",x"15",x"53",x"00",x"49",x"00",x"44",
		x"00",x"45",x"00",x"2D",x"00",x"54",x"00",x"57",x"00",x"4F",x"00",x"FF",x"FF",x"00",x"03",x"53",
		x"0F",x"49",x"0F",x"44",x"0F",x"45",x"0F",x"2D",x"0F",x"4F",x"0F",x"4E",x"0F",x"45",x"0F",x"FF",
		x"FF",x"1E",x"16",x"48",x"0F",x"49",x"0F",x"2D",x"0F",x"53",x"0F",x"43",x"0F",x"4F",x"0F",x"52",
		x"0F",x"45",x"0F",x"FF",x"FF",x"00",x"15",x"53",x"0F",x"49",x"0F",x"44",x"0F",x"45",x"0F",x"2D",
		x"0F",x"54",x"0F",x"57",x"0F",x"30",x"0F",x"FF",x"FF",x"01",x"03",x"B5",x"81",x"05",x"08",x"01",
		x"03",x"9C",x"81",x"05",x"08",x"1F",x"16",x"E2",x"80",x"05",x"08",x"01",x"15",x"CE",x"81",x"05",
		x"08",x"01",x"15",x"9C",x"81",x"05",x"08",x"D1",x"C9",x"E5",x"C9",x"F9",x"C9",x"D1",x"C9",x"E5",
		x"C9",x"97",x"CA",x"9F",x"CA",x"49",x"CA",x"55",x"CA",x"5B",x"CA",x"49",x"CA",x"55",x"CA",x"97",
		x"CA",x"9F",x"CA",x"0D",x"CA",x"E5",x"C9",x"F9",x"C9",x"0D",x"CA",x"E5",x"C9",x"97",x"CA",x"9F",
		x"CA",x"D1",x"C9",x"E5",x"C9",x"35",x"CA",x"00",x"15",x"08",x"FF",x"24",x"00",x"FF",x"FF",x"01",
		x"15",x"08",x"FF",x"24",x"00",x"FF",x"FF",x"1E",x"10",x"52",x"01",x"4F",x"01",x"55",x"01",x"4E",
		x"01",x"44",x"01",x"FF",x"FF",x"1F",x"11",x"B9",x"81",x"03",x"02",x"1F",x"11",x"D2",x"81",x"03",
		x"02",x"1F",x"11",x"AF",x"81",x"03",x"02",x"1F",x"10",x"00",x"00",x"2D",x"03",x"FF",x"FF",x"1F",
		x"10",x"2D",x"03",x"FF",x"FF",x"1F",x"13",x"2D",x"03",x"FF",x"FF",x"FB",x"CA",x"03",x"CB",x"0B",
		x"CB",x"17",x"CB",x"23",x"CB",x"33",x"CB",x"43",x"CB",x"57",x"CB",x"6B",x"CB",x"83",x"CB",x"9B",
		x"CB",x"B7",x"CB",x"D3",x"CB",x"F3",x"CB",x"13",x"CC",x"33",x"CC",x"1E",x"02",x"0E",x"FF",x"24",
		x"00",x"FF",x"FF",x"1F",x"02",x"0E",x"FF",x"24",x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",
		x"00",x"0C",x"FF",x"24",x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0C",x"FF",x"24",
		x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0A",x"FF",x"24",
		x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0A",x"FF",x"24",
		x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",
		x"00",x"08",x"FF",x"24",x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"0F",x"00",x"0D",x"00",x"08",x"FF",x"24",x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",
		x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"06",x"FF",x"24",
		x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"0F",x"00",x"0D",x"00",x"06",x"FF",x"24",x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",
		x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",
		x"00",x"04",x"FF",x"24",x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"04",x"FF",x"24",
		x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",
		x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"02",x"FF",x"24",
		x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"02",x"FF",x"24",
		x"00",x"FF",x"FF",x"1E",x"02",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",
		x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",x"00",x"0E",x"00",x"0C",
		x"00",x"FF",x"FF",x"1F",x"02",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",x"00",x"0F",x"00",x"0D",
		x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"00",x"6D",x"00",x"6E",x"00",x"6F",
		x"18",x"08",x"06",x"10",x"1E",x"00",x"02",x"05",x"05",x"15",x"02",x"11",x"03",x"01",x"04",x"11",
		x"05",x"01",x"05",x"11",x"04",x"05",x"03",x"15",x"0A",x"05",x"04",x"15",x"04",x"05",x"05",x"15",
		x"06",x"05",x"03",x"01",x"42",x"09",x"01",x"08",x"01",x"00",x"06",x"10",x"03",x"00",x"0C",x"04",
		x"0C",x"06",x"0C",x"02",x"06",x"12",x"05",x"02",x"04",x"12",x"04",x"02",x"07",x"12",x"03",x"02",
		x"0C",x"12",x"05",x"02",x"0B",x"0A",x"0C",x"00",x"08",x"10",x"04",x"04",x"04",x"00",x"01",x"08",
		x"0F",x"09",x"03",x"01",x"11",x"00",x"03",x"10",x"01",x"12",x"02",x"16",x"37",x"06",x"06",x"16",
		x"06",x"06",x"05",x"16",x"02",x"02",x"33",x"00",x"03",x"10",x"05",x"11",x"01",x"01",x"08",x"11",
		x"04",x"01",x"09",x"11",x"01",x"19",x"21",x"09",x"0C",x"00",x"04",x"10",x"02",x"12",x"17",x"06",
		x"02",x"04",x"05",x"05",x"01",x"01",x"05",x"09",x"14",x"19",x"02",x"09",x"03",x"08",x"02",x"0A",
		x"01",x"02",x"07",x"00",x"04",x"10",x"08",x"00",x"06",x"10",x"04",x"18",x"0B",x"08",x"03",x"00",
		x"05",x"10",x"08",x"00",x"01",x"10",x"0B",x"18",x"0A",x"08",x"05",x"00",x"05",x"10",x"07",x"00",
		x"0A",x"18",x"08",x"08",x"07",x"00",x"04",x"10",x"06",x"00",x"03",x"08",x"0B",x"18",x"09",x"08",
		x"0C",x"00",x"20",x"00",x"0C",x"0A",x"0A",x"09",x"6B",x"00",x"12",x"02",x"05",x"12",x"0A",x"06",
		x"03",x"04",x"03",x"05",x"04",x"04",x"0C",x"06",x"04",x"16",x"09",x"12",x"04",x"10",x"1D",x"01",
		x"01",x"00",x"01",x"08",x"11",x"0A",x"01",x"08",x"21",x"00",x"02",x"01",x"03",x"11",x"01",x"10",
		x"02",x"12",x"06",x"02",x"06",x"12",x"0E",x"02",x"06",x"12",x"04",x"02",x"05",x"12",x"01",x"1A",
		x"0C",x"0A",x"57",x"00",x"05",x"10",x"03",x"00",x"38",x"04",x"15",x"05",x"1E",x"01",x"1B",x"09",
		x"05",x"08",x"0D",x"00",x"0C",x"01",x"08",x"11",x"05",x"01",x"06",x"11",x"04",x"01",x"07",x"11",
		x"04",x"01",x"07",x"11",x"06",x"01",x"03",x"09",x"05",x"00",x"05",x"02",x"0A",x"00",x"33",x"02",
		x"57",x"0A",x"05",x"02",x"02",x"12",x"05",x"16",x"3F",x"06",x"04",x"04",x"07",x"05",x"1A",x"01",
		x"A0",x"00",x"12",x"01",x"15",x"00",x"15",x"06",x"10",x"00",x"05",x"05",x"03",x"15",x"03",x"05",
		x"05",x"15",x"03",x"05",x"03",x"15",x"A0",x"05",x"03",x"10",x"5A",x"05",x"03",x"16",x"03",x"06",
		x"03",x"16",x"03",x"06",x"03",x"16",x"03",x"06",x"03",x"16",x"03",x"16",x"03",x"06",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"08",x"D0",x"6E",x"D0",x"84",x"D0",x"8C",x"D0",x"0F",x"0E",x"50",x"0F",x"55",x"0F",x"53",x"0F",
		x"48",x"0F",x"FF",x"FF",x"11",x"06",x"31",x"05",x"00",x"00",x"50",x"05",x"4C",x"05",x"41",x"05",
		x"59",x"05",x"45",x"05",x"52",x"05",x"00",x"00",x"42",x"05",x"55",x"05",x"54",x"05",x"54",x"05",
		x"4F",x"05",x"4E",x"05",x"00",x"00",x"4F",x"05",x"4E",x"05",x"4C",x"05",x"59",x"05",x"FF",x"FF",
		x"11",x"06",x"31",x"05",x"00",x"00",x"4F",x"05",x"52",x"05",x"00",x"00",x"32",x"05",x"00",x"00",
		x"50",x"05",x"4C",x"05",x"41",x"05",x"59",x"05",x"45",x"05",x"52",x"05",x"53",x"05",x"00",x"00",
		x"42",x"05",x"55",x"05",x"54",x"05",x"54",x"05",x"4F",x"05",x"4E",x"05",x"FF",x"FF",x"14",x"0B",
		x"50",x"05",x"52",x"05",x"45",x"05",x"53",x"05",x"45",x"05",x"4E",x"05",x"54",x"05",x"45",x"05",
		x"44",x"05",x"FF",x"FF",x"16",x"0F",x"42",x"05",x"59",x"05",x"FF",x"FF",x"18",x"0B",x"54",x"01",
		x"45",x"01",x"48",x"01",x"4B",x"01",x"41",x"01",x"4E",x"01",x"00",x"00",x"4C",x"05",x"54",x"05",
		x"44",x"05",x"2E",x"05",x"FF",x"FF",x"D6",x"D0",x"F0",x"D0",x"D6",x"D0",x"00",x"D1",x"D6",x"D0",
		x"10",x"D1",x"20",x"D1",x"2E",x"D1",x"20",x"D1",x"3E",x"D1",x"4E",x"D1",x"6A",x"D1",x"86",x"D1",
		x"A6",x"D1",x"4E",x"D1",x"6A",x"D1",x"96",x"D1",x"B6",x"D1",x"C6",x"D1",x"E2",x"D1",x"FE",x"D1",
		x"1A",x"D2",x"2A",x"D2",x"3A",x"D2",x"18",x"05",x"45",x"00",x"56",x"00",x"45",x"00",x"52",x"00",
		x"59",x"00",x"00",x"00",x"42",x"00",x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",x"FF",x"FF",
		x"18",x"12",x"35",x"05",x"04",x"FF",x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",
		x"18",x"11",x"31",x"05",x"05",x"FF",x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",
		x"18",x"12",x"33",x"05",x"04",x"FF",x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",
		x"18",x"08",x"42",x"00",x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",x"FF",x"FF",x"18",x"0F",
		x"35",x"05",x"04",x"FF",x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"18",x"0E",
		x"31",x"05",x"05",x"FF",x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"17",x"05",
		x"46",x"00",x"49",x"00",x"52",x"00",x"53",x"00",x"54",x"00",x"00",x"00",x"00",x"00",x"42",x"00",
		x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",x"FF",x"FF",x"19",x"05",x"53",x"00",x"45",x"00",
		x"43",x"00",x"4F",x"00",x"4E",x"00",x"44",x"00",x"00",x"00",x"42",x"00",x"4F",x"00",x"4E",x"00",
		x"55",x"00",x"53",x"00",x"FF",x"FF",x"17",x"13",x"35",x"05",x"04",x"FF",x"30",x"05",x"00",x"00",
		x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"17",x"12",x"31",x"05",x"05",x"FF",x"30",x"05",x"00",x"00",
		x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"19",x"12",x"31",x"05",x"05",x"FF",x"30",x"05",x"00",x"00",
		x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"19",x"12",x"33",x"05",x"05",x"FF",x"30",x"05",x"00",x"00",
		x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"16",x"05",x"46",x"00",x"49",x"00",x"52",x"00",x"53",x"00",
		x"54",x"00",x"00",x"00",x"00",x"00",x"42",x"00",x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",
		x"FF",x"FF",x"18",x"05",x"53",x"00",x"45",x"00",x"43",x"00",x"4F",x"00",x"4E",x"00",x"44",x"00",
		x"00",x"00",x"42",x"00",x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",x"FF",x"FF",x"1A",x"05",
		x"54",x"00",x"48",x"00",x"49",x"00",x"52",x"00",x"44",x"00",x"00",x"00",x"00",x"00",x"42",x"00",
		x"4F",x"00",x"4E",x"00",x"55",x"00",x"53",x"00",x"FF",x"FF",x"16",x"13",x"35",x"05",x"04",x"FF",
		x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"18",x"12",x"31",x"05",x"05",x"FF",
		x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"1A",x"12",x"33",x"05",x"05",x"FF",
		x"30",x"05",x"00",x"00",x"3E",x"05",x"3C",x"05",x"FF",x"FF",x"0A",x"09",x"59",x"0F",x"4F",x"0F",
		x"55",x"0F",x"00",x"00",x"41",x"0F",x"52",x"0F",x"45",x"0F",x"00",x"00",x"4C",x"0F",x"55",x"0F",
		x"43",x"0F",x"4B",x"0F",x"59",x"0F",x"FF",x"FF",x"59",x"05",x"4F",x"05",x"55",x"05",x"00",x"0A",
		x"43",x"05",x"41",x"05",x"4E",x"05",x"00",x"0A",x"45",x"05",x"4E",x"05",x"4A",x"05",x"4F",x"05",
		x"59",x"05",x"FF",x"59",x"05",x"41",x"05",x"4C",x"05",x"50",x"05",x"00",x"0A",x"45",x"05",x"52",
		x"05",x"4F",x"05",x"4D",x"05",x"00",x"0A",x"45",x"05",x"4E",x"05",x"4F",x"05",x"FF",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"FF",x"0F",x"CE",x"08",x"FF",x"0F",x"0F",x"00",x"A0",x"0F",x"FF",x"00",
		x"00",x"00",x"2A",x"00",x"50",x"00",x"A0",x"00",x"88",x"08",x"66",x"06",x"44",x"04",x"F0",x"00",
		x"00",x"00",x"0F",x"00",x"00",x"00",x"44",x"04",x"88",x"08",x"CC",x"0C",x"FF",x"0F",x"0F",x"00",
		x"00",x"00",x"0F",x"00",x"00",x"00",x"44",x"04",x"88",x"08",x"CC",x"0C",x"FF",x"0F",x"F0",x"0F",
		x"00",x"00",x"0F",x"00",x"00",x"00",x"55",x"05",x"88",x"08",x"BB",x"0B",x"DD",x"0D",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"0D",x"00",x"DD",x"00",x"AA",x"0A",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"0F",x"00",x"00",x"00",x"44",x"04",x"88",x"08",x"CC",x"0C",x"FF",x"0F",x"8F",x"00",
		x"00",x"00",x"88",x"00",x"FF",x"0F",x"FF",x"0F",x"F6",x"06",x"FF",x"0F",x"FF",x"00",x"00",x"0F",
		x"00",x"00",x"00",x"0F",x"6F",x"00",x"FF",x"00",x"F0",x"00",x"F0",x"0F",x"FF",x"0F",x"AF",x"0C",
		x"00",x"00",x"88",x"08",x"AA",x"08",x"CC",x"0C",x"80",x"00",x"A0",x"00",x"C0",x"00",x"0A",x"0F",
		x"00",x"00",x"88",x"08",x"88",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0A",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"0D",x"00",x"DD",x"00",x"AA",x"0A",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"44",x"04",x"66",x"06",x"88",x"08",x"AA",x"0A",x"FF",x"0F",x"CC",x"0C",x"47",x"0E",
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"07",x"00",x"17",x"00",x"27",x"00",x"37",x"00",x"47",x"00",x"57",x"00",x"67",x"00",
		x"00",x"00",x"77",x"00",x"77",x"01",x"77",x"02",x"77",x"03",x"77",x"04",x"77",x"05",x"77",x"06",
		x"00",x"00",x"3F",x"00",x"5F",x"00",x"7F",x"00",x"9F",x"00",x"BF",x"00",x"DF",x"00",x"FF",x"00",
		x"00",x"00",x"40",x"00",x"60",x"00",x"80",x"00",x"A0",x"00",x"C0",x"00",x"E0",x"00",x"F0",x"00",
		x"00",x"00",x"3F",x"00",x"5F",x"00",x"7F",x"00",x"9F",x"00",x"BF",x"00",x"DF",x"00",x"FF",x"00",
		x"00",x"00",x"55",x"00",x"77",x"00",x"99",x"00",x"BB",x"00",x"DD",x"00",x"FF",x"00",x"FF",x"04",
		x"00",x"00",x"00",x"08",x"00",x"0C",x"00",x"0F",x"80",x"0F",x"A0",x"0F",x"C0",x"0F",x"F0",x"0F",
		x"00",x"00",x"00",x"0F",x"C0",x"00",x"F0",x"00",x"F8",x"00",x"F0",x"00",x"FF",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"0F",x"5C",x"00",x"8F",x"00",x"FF",x"00",x"8F",x"00",x"FF",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"0F",x"0F",x"00",x"4F",x"04",x"8F",x"08",x"4F",x"04",x"CF",x"0C",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"00",x"08",x"00",x"0C",x"00",x"0F",x"00",x"00",x"00",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CC",x"0C",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CC",x"0C",x"FF",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CC",x"0C",x"FF",x"0F",
		x"00",x"00",x"58",x"0B",x"45",x"00",x"67",x"02",x"89",x"04",x"AB",x"06",x"CD",x"08",x"EF",x"0A",
		x"00",x"00",x"00",x"0C",x"00",x"0B",x"00",x"0A",x"00",x"09",x"00",x"08",x"00",x"07",x"00",x"06",
		x"00",x"00",x"00",x"0C",x"45",x"00",x"67",x"02",x"89",x"04",x"AB",x"06",x"CD",x"08",x"EF",x"0A",
		x"00",x"00",x"88",x"0C",x"50",x"00",x"A0",x"00",x"88",x"08",x"66",x"06",x"44",x"04",x"22",x"02",
		x"00",x"00",x"00",x"0C",x"00",x"0B",x"00",x"0A",x"00",x"09",x"00",x"08",x"88",x"08",x"AA",x"0A",
		x"00",x"00",x"44",x"04",x"44",x"04",x"00",x"00",x"30",x"03",x"50",x"05",x"70",x"07",x"05",x"07",
		x"00",x"00",x"44",x"04",x"44",x"04",x"00",x"00",x"33",x"00",x"55",x"00",x"77",x"00",x"05",x"07",
		x"00",x"00",x"44",x"04",x"44",x"04",x"00",x"00",x"33",x"03",x"55",x"05",x"77",x"07",x"05",x"07",
		x"00",x"00",x"05",x"00",x"50",x"00",x"80",x"00",x"28",x"00",x"4A",x"00",x"06",x"00",x"45",x"00",
		x"00",x"00",x"27",x"00",x"08",x"0C",x"40",x"00",x"CC",x"0C",x"0D",x"00",x"80",x"00",x"CC",x"00",
		x"00",x"00",x"0F",x"00",x"55",x"05",x"77",x"07",x"99",x"09",x"BB",x"0B",x"DD",x"0D",x"00",x"0F",
		x"00",x"00",x"88",x"0C",x"2A",x"00",x"AA",x"0A",x"88",x"08",x"66",x"06",x"44",x"04",x"22",x"02",
		x"00",x"00",x"60",x"0C",x"55",x"05",x"77",x"07",x"99",x"09",x"BB",x"0B",x"DD",x"0D",x"A0",x"00",
		x"00",x"00",x"00",x"07",x"37",x"00",x"77",x"00",x"10",x"01",x"30",x"03",x"50",x"05",x"57",x"06",
		x"00",x"00",x"00",x"07",x"37",x"00",x"77",x"00",x"11",x"00",x"33",x"00",x"55",x"00",x"57",x"06",
		x"00",x"00",x"00",x"07",x"37",x"00",x"77",x"00",x"11",x"01",x"33",x"03",x"55",x"05",x"57",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"55",x"00",x"77",x"00",x"99",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"44",x"04",x"66",x"06",x"88",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"55",x"00",x"66",x"00",x"77",x"00",x"88",x"00",x"88",x"00",x"88",x"00",x"88",x"00",
		x"00",x"00",x"44",x"04",x"55",x"05",x"66",x"06",x"77",x"07",x"77",x"07",x"77",x"07",x"77",x"07",
		x"CC",x"CD",x"CE",x"CF",x"15",x"94",x"95",x"96",x"97",x"0D",x"CC",x"CD",x"CE",x"CF",x"15",x"94",
		x"95",x"96",x"97",x"0D",x"CC",x"CD",x"CE",x"CF",x"15",x"94",x"95",x"96",x"97",x"0D",x"CC",x"CD",
		x"CE",x"CF",x"15",x"94",x"95",x"96",x"97",x"0D",x"CC",x"CD",x"CE",x"CF",x"15",x"94",x"95",x"96",
		x"97",x"0D",x"CC",x"CD",x"CE",x"CF",x"15",x"94",x"95",x"96",x"97",x"0D",x"D8",x"D9",x"DA",x"DB",
		x"15",x"90",x"91",x"92",x"93",x"0D",x"DC",x"DD",x"DE",x"DF",x"15",x"90",x"91",x"92",x"93",x"0D",
		x"04",x"00",x"00",x"01",x"C0",x"00",x"00",x"02",x"05",x"00",x"00",x"01",x"C0",x"00",x"00",x"02",
		x"06",x"00",x"C0",x"00",x"80",x"00",x"00",x"02",x"07",x"00",x"C0",x"00",x"80",x"00",x"00",x"01",
		x"07",x"00",x"80",x"00",x"60",x"00",x"00",x"02",x"04",x"00",x"80",x"00",x"40",x"00",x"00",x"01",
		x"05",x"00",x"60",x"00",x"60",x"00",x"00",x"01",x"06",x"00",x"60",x"00",x"40",x"00",x"00",x"01",
		x"07",x"00",x"60",x"00",x"40",x"00",x"00",x"01",x"07",x"00",x"20",x"00",x"40",x"00",x"00",x"01",
		x"04",x"00",x"80",x"00",x"30",x"00",x"00",x"01",x"05",x"00",x"80",x"00",x"30",x"00",x"00",x"01",
		x"06",x"00",x"60",x"00",x"30",x"00",x"00",x"01",x"07",x"00",x"60",x"00",x"30",x"00",x"00",x"01",
		x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"04",x"00",x"60",x"00",x"20",x"00",x"00",x"01",
		x"05",x"00",x"60",x"00",x"20",x"00",x"00",x"01",x"06",x"00",x"40",x"00",x"20",x"00",x"00",x"01",
		x"07",x"00",x"40",x"00",x"20",x"00",x"00",x"01",x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",
		x"04",x"00",x"40",x"00",x"20",x"00",x"00",x"01",x"05",x"00",x"40",x"00",x"20",x"00",x"00",x"01",
		x"06",x"00",x"40",x"00",x"20",x"00",x"00",x"01",x"07",x"00",x"40",x"00",x"20",x"00",x"00",x"01",
		x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"04",x"00",x"20",x"00",x"20",x"00",x"00",x"01",
		x"05",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"06",x"00",x"20",x"00",x"20",x"00",x"00",x"01",
		x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",
		x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",
		x"07",x"00",x"20",x"00",x"20",x"00",x"00",x"01",x"01",x"00",x"20",x"00",x"44",x"00",x"80",x"00",
		x"02",x"00",x"00",x"00",x"01",x"00",x"30",x"00",x"55",x"00",x"80",x"00",x"02",x"00",x"00",x"00",
		x"01",x"00",x"38",x"00",x"66",x"00",x"80",x"00",x"03",x"00",x"00",x"00",x"01",x"00",x"40",x"00",
		x"55",x"00",x"70",x"00",x"03",x"00",x"00",x"00",x"01",x"00",x"40",x"00",x"66",x"00",x"70",x"00",
		x"04",x"00",x"00",x"00",x"01",x"00",x"40",x"00",x"77",x"00",x"70",x"00",x"04",x"00",x"00",x"00",
		x"01",x"00",x"48",x"00",x"66",x"00",x"60",x"00",x"05",x"00",x"00",x"00",x"01",x"00",x"48",x"00",
		x"77",x"00",x"60",x"00",x"05",x"00",x"00",x"00",x"01",x"00",x"48",x"00",x"88",x"00",x"60",x"00",
		x"06",x"00",x"00",x"00",x"02",x"00",x"40",x"00",x"55",x"00",x"80",x"00",x"06",x"00",x"00",x"00",
		x"02",x"00",x"40",x"00",x"66",x"00",x"80",x"00",x"07",x"00",x"00",x"00",x"02",x"00",x"40",x"00",
		x"77",x"00",x"80",x"00",x"07",x"00",x"00",x"00",x"02",x"00",x"48",x"00",x"66",x"00",x"70",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"48",x"00",x"77",x"00",x"70",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"48",x"00",x"88",x"00",x"70",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"50",x"00",
		x"77",x"00",x"60",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"50",x"00",x"88",x"00",x"60",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"50",x"00",x"99",x"00",x"60",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"58",x"00",x"88",x"00",x"60",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"50",x"00",
		x"77",x"00",x"80",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"50",x"00",x"88",x"00",x"80",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"58",x"00",x"77",x"00",x"80",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"58",x"00",x"88",x"00",x"70",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"58",x"00",
		x"99",x"00",x"70",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"60",x"00",x"88",x"00",x"70",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"60",x"00",x"99",x"00",x"60",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"60",x"00",x"A2",x"00",x"60",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"68",x"00",
		x"99",x"00",x"60",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"68",x"00",x"A2",x"00",x"50",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"68",x"00",x"AA",x"00",x"50",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"70",x"00",x"A2",x"00",x"50",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"70",x"00",
		x"AA",x"00",x"48",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"70",x"00",x"B3",x"00",x"48",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"78",x"00",x"AA",x"00",x"48",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"78",x"00",x"B3",x"00",x"40",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"78",x"00",
		x"BB",x"00",x"40",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"80",x"00",x"B3",x"00",x"40",x"00",
		x"08",x"00",x"00",x"00",x"02",x"00",x"80",x"00",x"BB",x"00",x"38",x"00",x"08",x"00",x"00",x"00",
		x"02",x"00",x"80",x"00",x"C4",x"00",x"38",x"00",x"08",x"00",x"00",x"00",x"02",x"00",x"80",x"00",
		x"BB",x"00",x"38",x"00",x"08",x"00",x"00",x"00",x"80",x"00",x"00",x"01",x"01",x"00",x"00",x"02",
		x"01",x"00",x"00",x"04",x"B3",x"B3",x"B3",x"B4",x"B3",x"B3",x"B3",x"B4",x"91",x"00",x"C0",x"00",
		x"02",x"00",x"80",x"01",x"01",x"00",x"00",x"03",x"B1",x"B1",x"B1",x"B4",x"B1",x"B1",x"B1",x"B4",
		x"A2",x"00",x"C0",x"00",x"03",x"00",x"00",x"01",x"01",x"00",x"00",x"02",x"B2",x"B2",x"B2",x"B4",
		x"B2",x"B2",x"B2",x"B4",x"AE",x"00",x"80",x"00",x"04",x"00",x"C0",x"00",x"01",x"00",x"80",x"01",
		x"B0",x"B0",x"B0",x"B4",x"B0",x"B0",x"B0",x"B4",x"C0",x"00",x"80",x"00",x"05",x"00",x"C0",x"00",
		x"04",x"00",x"00",x"03",x"B4",x"B4",x"B4",x"B4",x"B4",x"B4",x"B4",x"B4",x"D1",x"00",x"80",x"00",
		x"06",x"00",x"C0",x"00",x"03",x"00",x"80",x"01",x"B2",x"B2",x"B1",x"B1",x"B2",x"B2",x"B3",x"B3",
		x"80",x"01",x"80",x"00",x"07",x"00",x"C0",x"00",x"03",x"00",x"80",x"01",x"B0",x"B1",x"B2",x"B3",
		x"B4",x"B3",x"B2",x"B1",x"EE",x"00",x"80",x"00",x"08",x"00",x"C0",x"00",x"03",x"00",x"80",x"01",
		x"B0",x"B0",x"B1",x"B1",x"B0",x"B0",x"B1",x"B1",x"00",x"01",x"80",x"00",x"09",x"00",x"C0",x"00",
		x"03",x"00",x"80",x"01",x"B3",x"B3",x"B4",x"B4",x"B3",x"B3",x"B4",x"B4",x"00",x"01",x"80",x"00",
		x"0A",x"00",x"C0",x"00",x"03",x"00",x"80",x"01",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",
		x"00",x"01",x"80",x"00",x"0B",x"00",x"C0",x"00",x"04",x"00",x"80",x"01",x"B4",x"B3",x"B4",x"B3",
		x"B0",x"B1",x"B0",x"B1",x"00",x"01",x"80",x"00",x"0C",x"00",x"C0",x"00",x"04",x"00",x"80",x"01",
		x"B1",x"B2",x"B1",x"B2",x"B1",x"B2",x"B1",x"B2",x"00",x"01",x"80",x"00",x"0D",x"00",x"C0",x"00",
		x"04",x"00",x"80",x"01",x"B3",x"B0",x"B3",x"B0",x"B3",x"B0",x"B3",x"B0",x"00",x"01",x"80",x"00",
		x"0E",x"00",x"C0",x"00",x"05",x"00",x"80",x"01",x"B4",x"B4",x"B4",x"B1",x"B4",x"B4",x"B4",x"B1",
		x"00",x"02",x"80",x"00",x"0F",x"00",x"C0",x"00",x"05",x"00",x"80",x"01",x"B0",x"B0",x"B0",x"B0",
		x"B0",x"B0",x"B0",x"B0",x"00",x"01",x"80",x"00",x"10",x"00",x"C0",x"00",x"05",x"00",x"80",x"01",
		x"B1",x"B1",x"B1",x"B1",x"B1",x"B1",x"B1",x"B1",x"80",x"01",x"80",x"00",x"11",x"00",x"C0",x"00",
		x"05",x"00",x"80",x"01",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",x"B2",x"80",x"01",x"80",x"00",
		x"12",x"00",x"C0",x"00",x"05",x"00",x"80",x"01",x"B3",x"B3",x"B3",x"B3",x"B3",x"B3",x"B3",x"B3",
		x"80",x"01",x"80",x"00",x"13",x"00",x"C0",x"00",x"06",x"00",x"80",x"01",x"B4",x"B4",x"B4",x"B4",
		x"B4",x"B4",x"B4",x"B4",x"80",x"01",x"80",x"00",x"14",x"00",x"C0",x"00",x"06",x"00",x"80",x"01",
		x"B0",x"B0",x"B4",x"B4",x"B2",x"B2",x"B4",x"B4",x"80",x"01",x"80",x"00",x"15",x"00",x"C0",x"00",
		x"06",x"00",x"80",x"01",x"B0",x"B0",x"B0",x"B0",x"B1",x"B1",x"B1",x"B1",x"80",x"01",x"80",x"00",
		x"16",x"00",x"C0",x"00",x"06",x"00",x"80",x"01",x"B1",x"B1",x"B1",x"B1",x"B2",x"B2",x"B2",x"B2",
		x"80",x"01",x"80",x"00",x"17",x"00",x"C0",x"00",x"06",x"00",x"80",x"01",x"B2",x"B2",x"B2",x"B2",
		x"B3",x"B3",x"B3",x"B3",x"80",x"01",x"80",x"00",x"18",x"00",x"C0",x"00",x"07",x"00",x"80",x"01",
		x"B3",x"B3",x"B3",x"B3",x"B4",x"B4",x"B4",x"B4",x"00",x"02",x"80",x"00",x"19",x"00",x"C0",x"00",
		x"07",x"00",x"80",x"01",x"B1",x"B3",x"B1",x"B3",x"B1",x"B3",x"B1",x"B3",x"00",x"02",x"80",x"00",
		x"1A",x"00",x"C0",x"00",x"07",x"00",x"80",x"01",x"B4",x"B4",x"B4",x"B4",x"B0",x"B0",x"B0",x"B0",
		x"00",x"02",x"80",x"00",x"1B",x"00",x"C0",x"00",x"07",x"00",x"80",x"01",x"B3",x"B3",x"B3",x"B3",
		x"B1",x"B1",x"B1",x"B1",x"00",x"02",x"80",x"00",x"1C",x"00",x"C0",x"00",x"08",x"00",x"80",x"01",
		x"B2",x"B2",x"B2",x"B2",x"B4",x"B4",x"B4",x"B4",x"00",x"02",x"80",x"00",x"1D",x"00",x"C0",x"00",
		x"08",x"00",x"80",x"01",x"B0",x"B0",x"B0",x"B0",x"B3",x"B3",x"B3",x"B3",x"00",x"02",x"80",x"00",
		x"1E",x"00",x"C0",x"00",x"09",x"00",x"80",x"01",x"B4",x"B3",x"B4",x"B2",x"B4",x"B1",x"B4",x"B0",
		x"00",x"02",x"80",x"00",x"1F",x"00",x"C0",x"00",x"09",x"00",x"80",x"01",x"B0",x"B1",x"B2",x"B3",
		x"B4",x"B0",x"B1",x"B2",x"00",x"02",x"80",x"00",x"20",x"00",x"C0",x"00",x"09",x"00",x"80",x"01",
		x"B3",x"B4",x"B0",x"B1",x"B2",x"B3",x"B4",x"B0",x"00",x"00",x"02",x"00",x"00",x"00",x"0B",x"01",
		x"00",x"0B",x"01",x"01",x"08",x"02",x"03",x"08",x"02",x"02",x"07",x"03",x"04",x"07",x"03",x"00",
		x"04",x"04",x"01",x"04",x"04",x"01",x"02",x"00",x"02",x"02",x"00",x"02",x"06",x"01",x"00",x"06",
		x"01",x"00",x"03",x"02",x"03",x"03",x"02",x"01",x"0A",x"03",x"04",x"0A",x"03",x"02",x"04",x"04",
		x"01",x"00",x"04",x"00",x"0C",x"00",x"02",x"0C",x"00",x"01",x"0E",x"01",x"00",x"0E",x"01",x"02",
		x"09",x"02",x"03",x"09",x"02",x"00",x"0F",x"03",x"04",x"0F",x"03",x"01",x"04",x"04",x"01",x"04",
		x"04",x"02",x"0D",x"00",x"02",x"0D",x"00",x"00",x"01",x"01",x"00",x"01",x"01",x"01",x"05",x"02",
		x"03",x"05",x"02",x"02",x"0B",x"03",x"04",x"0B",x"03",x"00",x"04",x"04",x"01",x"0D",x"04",x"01",
		x"0E",x"00",x"02",x"0E",x"00",x"02",x"06",x"01",x"00",x"06",x"01",x"00",x"07",x"02",x"03",x"07",
		x"02",x"01",x"09",x"03",x"04",x"09",x"03",x"02",x"04",x"04",x"01",x"0F",x"04",x"00",x"05",x"00",
		x"02",x"05",x"00",x"01",x"03",x"01",x"00",x"03",x"01",x"02",x"01",x"02",x"03",x"01",x"02",x"00",
		x"0C",x"03",x"04",x"0C",x"03",x"01",x"04",x"04",x"01",x"00",x"04",x"02",x"02",x"00",x"02",x"02",
		x"00",x"00",x"08",x"01",x"00",x"08",x"01",x"01",x"0F",x"02",x"03",x"0F",x"02",x"02",x"0D",x"03",
		x"04",x"0D",x"03",x"00",x"04",x"04",x"01",x"06",x"04",x"01",x"0A",x"00",x"02",x"0A",x"00",x"02",
		x"09",x"01",x"00",x"09",x"01",x"00",x"01",x"02",x"03",x"01",x"02",x"01",x"02",x"03",x"04",x"02",
		x"03",x"02",x"04",x"04",x"01",x"02",x"04",x"00",x"03",x"00",x"02",x"03",x"00",x"01",x"05",x"01",
		x"00",x"05",x"01",x"02",x"06",x"02",x"03",x"06",x"02",x"00",x"07",x"00",x"04",x"07",x"03",x"01",
		x"04",x"01",x"01",x"0E",x"04",x"02",x"08",x"02",x"02",x"08",x"00",x"00",x"09",x"03",x"00",x"09",
		x"01",x"01",x"0A",x"04",x"03",x"0A",x"02",x"02",x"0B",x"00",x"04",x"0B",x"03",x"00",x"04",x"01",
		x"01",x"0A",x"04",x"01",x"0C",x"02",x"02",x"0C",x"00",x"02",x"0D",x"03",x"00",x"0D",x"01",x"00",
		x"0E",x"04",x"03",x"0E",x"02",x"01",x"0F",x"00",x"04",x"0F",x"03",x"02",x"04",x"01",x"01",x"06",
		x"04",x"00",x"00",x"02",x"02",x"00",x"00",x"01",x"01",x"03",x"00",x"01",x"01",x"02",x"02",x"04",
		x"03",x"02",x"02",x"00",x"03",x"00",x"04",x"03",x"03",x"01",x"04",x"01",x"01",x"08",x"04",x"02",
		x"05",x"02",x"02",x"05",x"00",x"00",x"06",x"03",x"00",x"06",x"01",x"01",x"07",x"04",x"03",x"07",
		x"02",x"02",x"08",x"00",x"04",x"08",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"CB",x"01",x"E1",x"E1",x"E1",x"E1",x"08",x"80",x"02",x"E0",x"02",x"08",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"18",x"12",x"7D",x"7D",x"00",x"00",x"00",x"00",x"12",x"E2",x"72",x"2E",x"FE",
		x"00",x"6F",x"2F",x"31",x"0A",x"00",x"00",x"00",x"FC",x"4C",x"4E",x"A2",x"72",x"30",x"00",x"00",
		x"00",x"00",x"00",x"30",x"24",x"FA",x"FA",x"00",x"00",x"08",x"2C",x"46",x"E1",x"70",x"38",x"F8",
		x"00",x"DE",x"5E",x"62",x"34",x"00",x"00",x"00",x"F8",x"4C",x"42",x"B5",x"76",x"30",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0E",x"00",x"3C",x"00",x"00",x"00",x"00",x"10",x"30",x"30",x"62",
		x"6C",x"0D",x"13",x"67",x"33",x"39",x"0A",x"00",x"74",x"F0",x"F4",x"38",x"6E",x"38",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0E",x"00",x"3C",x"00",x"00",x"00",x"00",x"10",x"3C",x"36",x"66",
		x"6C",x"0D",x"13",x"67",x"33",x"39",x"0A",x"00",x"76",x"F6",x"B3",x"34",x"6E",x"1E",x"07",x"00",
		x"00",x"00",x"00",x"00",x"00",x"0C",x"00",x"3C",x"00",x"00",x"00",x"00",x"14",x"39",x"37",x"67",
		x"6C",x"0D",x"13",x"67",x"33",x"39",x"0A",x"00",x"7F",x"F8",x"F8",x"38",x"6C",x"37",x"0B",x"0E",
		x"00",x"0A",x"39",x"33",x"67",x"13",x"0D",x"6C",x"00",x"00",x"38",x"6E",x"38",x"F4",x"F0",x"74",
		x"20",x"1C",x"0C",x"00",x"00",x"00",x"00",x"00",x"62",x"30",x"30",x"10",x"00",x"00",x"00",x"00",
		x"00",x"0A",x"39",x"33",x"67",x"13",x"0D",x"6C",x"00",x"07",x"1E",x"6E",x"34",x"B3",x"F6",x"76",
		x"20",x"1C",x"0C",x"00",x"00",x"00",x"00",x"00",x"66",x"36",x"3C",x"10",x"00",x"00",x"00",x"00",
		x"00",x"0A",x"39",x"33",x"67",x"13",x"0D",x"6C",x"0E",x"0B",x"37",x"6C",x"38",x"FC",x"7C",x"78",
		x"20",x"1C",x"0C",x"00",x"00",x"00",x"00",x"00",x"22",x"36",x"3A",x"16",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"04",x"04",x"00",x"00",x"00",x"00",x"60",x"F0",x"90",x"90",
		x"04",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"90",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"08",x"1F",x"3F",x"3C",x"34",x"00",x"00",x"00",x"08",x"FC",x"FE",x"9E",x"96",
		x"34",x"3F",x"3F",x"18",x"0F",x"07",x"00",x"00",x"96",x"FE",x"FE",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"38",x"38",x"00",x"00",x"00",x"00",x"60",x"F0",x"00",x"00",
		x"38",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"0C",x"04",x"00",x"00",x"00",x"00",x"F0",x"F0",x"90",x"90",
		x"04",x"07",x"00",x"00",x"07",x"07",x"00",x"00",x"90",x"F2",x"06",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"10",x"90",x"90",x"90",
		x"04",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"90",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"08",x"1F",x"3F",x"3C",x"34",x"00",x"00",x"00",x"08",x"FC",x"FE",x"9E",x"96",
		x"34",x"3F",x"3F",x"18",x"0F",x"07",x"00",x"00",x"96",x"FE",x"FE",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"04",x"38",x"38",x"00",x"00",x"00",x"00",x"10",x"90",x"00",x"00",
		x"38",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"0C",x"04",x"00",x"00",x"00",x"00",x"F0",x"F0",x"90",x"90",
		x"04",x"07",x"00",x"00",x"07",x"07",x"00",x"00",x"90",x"F2",x"06",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"06",x"04",x"04",x"00",x"00",x"00",x"00",x"60",x"F0",x"90",x"90",
		x"04",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"90",x"B0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"08",x"1F",x"3F",x"3C",x"34",x"00",x"00",x"00",x"08",x"FC",x"FE",x"9E",x"96",
		x"34",x"3F",x"3B",x"18",x"0F",x"07",x"00",x"00",x"96",x"BE",x"2E",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"06",x"38",x"38",x"00",x"00",x"00",x"00",x"60",x"F0",x"00",x"00",
		x"38",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"B0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"0C",x"04",x"00",x"00",x"00",x"00",x"F0",x"F0",x"90",x"90",
		x"04",x"07",x"00",x"00",x"07",x"07",x"00",x"00",x"90",x"B2",x"06",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"06",x"1E",x"00",x"00",x"60",x"E0",x"C0",x"DA",x"DE",x"DE",
		x"06",x"1E",x"06",x"01",x"01",x"00",x"00",x"00",x"F8",x"DE",x"DE",x"DA",x"C0",x"E0",x"60",x"00",
		x"00",x"00",x"0C",x"0E",x"07",x"05",x"06",x"36",x"00",x"00",x"00",x"00",x"00",x"D9",x"DF",x"DE",
		x"0E",x"36",x"06",x"05",x"07",x"0E",x"0C",x"00",x"F8",x"DE",x"DF",x"D9",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"38",x"78",x"FC",x"6E",x"AE",x"AA",
		x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"B8",x"AA",x"AE",x"6E",x"FC",x"78",x"38",x"00",
		x"00",x"00",x"00",x"04",x"1E",x"06",x"00",x"0E",x"00",x"C2",x"C2",x"CE",x"DE",x"FC",x"D8",x"D0",
		x"0C",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"DA",x"DE",x"DE",x"CE",x"C4",x"E0",x"60",x"00",
		x"00",x"00",x"00",x"04",x"1E",x"06",x"00",x"0E",x"00",x"04",x"04",x"7C",x"FC",x"DA",x"5E",x"DE",
		x"0C",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"DE",x"FC",x"F8",x"78",x"00",x"00",x"00",x"00",
		x"00",x"01",x"01",x"04",x"1E",x"06",x"00",x"0E",x"00",x"82",x"C2",x"CE",x"DE",x"FC",x"58",x"D0",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DA",x"5E",x"1E",x"04",x"C0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"04",x"1E",x"06",x"00",x"0E",x"00",x"04",x"C4",x"DC",x"FC",x"DA",x"DE",x"DE",
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"F8",x"60",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"0C",x"00",x"60",x"E0",x"C4",x"CE",x"DE",x"DE",x"DA",
		x"0E",x"00",x"06",x"1E",x"04",x"00",x"00",x"00",x"D0",x"D8",x"FC",x"DE",x"CE",x"C2",x"C2",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"0C",x"00",x"00",x"00",x"00",x"78",x"F8",x"FC",x"DE",
		x"0E",x"00",x"06",x"1E",x"04",x"00",x"00",x"00",x"DE",x"DE",x"DA",x"FC",x"7C",x"04",x"04",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"00",x"00",x"C0",x"C0",x"04",x"1E",x"5E",x"DA",
		x"0E",x"00",x"06",x"1E",x"04",x"01",x"01",x"00",x"D0",x"D8",x"FC",x"DE",x"CE",x"C2",x"82",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"60",x"60",x"F8",x"FE",
		x"0E",x"00",x"06",x"1E",x"04",x"00",x"00",x"00",x"DE",x"DE",x"DE",x"FC",x"DC",x"C4",x"04",x"00",
		x"00",x"00",x"06",x"07",x"03",x"02",x"03",x"1B",x"00",x"00",x"00",x"00",x"80",x"ED",x"6F",x"6F",
		x"07",x"1B",x"03",x"02",x"03",x"07",x"06",x"00",x"7C",x"6F",x"6F",x"ED",x"80",x"00",x"00",x"00",
		x"00",x"00",x"03",x"03",x"01",x"01",x"01",x"03",x"00",x"00",x"00",x"80",x"C0",x"75",x"B7",x"B7",
		x"03",x"03",x"01",x"01",x"01",x"03",x"03",x"00",x"BC",x"B7",x"B7",x"75",x"C0",x"80",x"00",x"00",
		x"00",x"00",x"04",x"36",x"04",x"01",x"07",x"06",x"40",x"E0",x"F0",x"F9",x"7D",x"EF",x"4F",x"5E",
		x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"5C",x"DC",x"9C",x"CC",x"C6",x"E3",x"C0",x"00",
		x"00",x"00",x"01",x"03",x"03",x"03",x"05",x"1F",x"04",x"C6",x"CF",x"9F",x"BE",x"BC",x"B8",x"DC",
		x"06",x"0E",x"02",x"02",x"03",x"00",x"00",x"00",x"DE",x"DE",x"DE",x"D8",x"D8",x"F8",x"78",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"C0",x"E3",x"C6",x"CC",x"9C",x"DC",x"5C",
		x"06",x"07",x"01",x"04",x"36",x"04",x"00",x"00",x"5E",x"4F",x"EF",x"7D",x"F9",x"F0",x"E0",x"40",
		x"00",x"00",x"00",x"0D",x"02",x"02",x"0E",x"07",x"00",x"78",x"F8",x"D0",x"D8",x"DE",x"DE",x"DE",
		x"1E",x"05",x"03",x"03",x"03",x"01",x"00",x"00",x"DC",x"B8",x"BC",x"BE",x"9F",x"CF",x"C6",x"04",
		x"40",x"40",x"40",x"66",x"65",x"65",x"75",x"74",x"F4",x"70",x"C0",x"00",x"80",x"00",x"00",x"00",
		x"78",x"7C",x"7D",x"7E",x"1F",x"00",x"03",x"07",x"00",x"80",x"00",x"00",x"00",x"80",x"60",x"D0",
		x"03",x"25",x"24",x"34",x"35",x"3F",x"3F",x"3F",x"E0",x"D8",x"70",x"00",x"00",x"00",x"00",x"00",
		x"3F",x"3F",x"3E",x"1C",x"07",x"00",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"80",x"60",x"D0",
		x"03",x"01",x"00",x"02",x"00",x"00",x"00",x"00",x"80",x"C0",x"60",x"18",x"84",x"80",x"00",x"00",
		x"00",x"00",x"03",x"0C",x"07",x"00",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"80",x"20",x"D0",
		x"00",x"00",x"00",x"00",x"68",x"17",x"07",x"0F",x"00",x"00",x"00",x"00",x"00",x"80",x"FC",x"D7",
		x"07",x"1B",x"6F",x"40",x"20",x"20",x"10",x"00",x"38",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"04",x"08",x"08",x"10",x"03",x"07",x"0F",x"00",x"00",x"00",x"00",x"00",x"80",x"F8",x"D6",
		x"07",x"0B",x"07",x"00",x"10",x"08",x"04",x"00",x"38",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"00",x"00",x"10",x"03",x"07",x"0F",x"00",x"00",x"00",x"00",x"00",x"80",x"F0",x"D4",
		x"07",x"0B",x"07",x"08",x"08",x"0E",x"00",x"00",x"30",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"40",x"40",x"61",x"63",x"73",x"7B",x"7D",x"7D",x"00",x"82",x"70",x"00",x"00",x"00",x"00",x"00",
		x"59",x"7C",x"79",x"71",x"23",x"03",x"07",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"00",
		x"00",x"07",x"03",x"23",x"71",x"79",x"7C",x"59",x"00",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",
		x"7D",x"7D",x"7B",x"73",x"63",x"61",x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"70",x"82",x"00",
		x"00",x"00",x"00",x"00",x"01",x"05",x"06",x"1E",x"00",x"00",x"40",x"E0",x"E0",x"FA",x"DE",x"DE",
		x"0E",x"1E",x"06",x"05",x"01",x"00",x"00",x"00",x"F8",x"DE",x"DE",x"FA",x"E0",x"E0",x"40",x"00",
		x"00",x"00",x"07",x"07",x"01",x"01",x"01",x"06",x"00",x"00",x"80",x"8E",x"8E",x"DC",x"DC",x"D8",
		x"06",x"1E",x"0E",x"1C",x"00",x"03",x"03",x"00",x"D8",x"F8",x"DE",x"DE",x"CE",x"C2",x"C0",x"00",
		x"00",x"00",x"0C",x"0E",x"07",x"05",x"06",x"36",x"00",x"00",x"00",x"00",x"00",x"DA",x"DE",x"DE",
		x"0E",x"36",x"06",x"05",x"07",x"0E",x"0C",x"00",x"F8",x"DE",x"DE",x"DA",x"00",x"00",x"00",x"00",
		x"00",x"03",x"01",x"01",x"18",x"7D",x"7C",x"41",x"00",x"E0",x"80",x"38",x"A0",x"58",x"C0",x"30",
		x"01",x"12",x"1A",x"0D",x"01",x"00",x"01",x"00",x"30",x"A0",x"BC",x"5C",x"28",x"E0",x"C0",x"00",
		x"00",x"03",x"01",x"01",x"18",x"7D",x"7C",x"41",x"00",x"E0",x"80",x"3F",x"A0",x"59",x"C0",x"30",
		x"01",x"12",x"1A",x"0D",x"01",x"00",x"01",x"00",x"30",x"A0",x"BC",x"5C",x"2F",x"E0",x"C0",x"00",
		x"00",x"03",x"01",x"00",x"18",x"7E",x"7F",x"47",x"00",x"E0",x"F0",x"78",x"3C",x"3C",x"18",x"90",
		x"03",x"11",x"19",x"0C",x"00",x"00",x"01",x"00",x"D0",x"F8",x"FC",x"EC",x"E8",x"C0",x"C0",x"00",
		x"00",x"07",x"1B",x"22",x"2D",x"72",x"F9",x"82",x"00",x"CA",x"04",x"78",x"40",x"B0",x"80",x"60",
		x"02",x"25",x"35",x"1A",x"02",x"01",x"03",x"00",x"68",x"44",x"7C",x"BA",x"50",x"C0",x"80",x"00",
		x"80",x"E0",x"7C",x"5E",x"2C",x"3F",x"17",x"1B",x"04",x"06",x"06",x"0F",x"8F",x"76",x"24",x"8C",
		x"0B",x"0C",x"04",x"04",x"01",x"01",x"00",x"00",x"BC",x"6C",x"34",x"DA",x"EA",x"2C",x"08",x"00",
		x"80",x"E0",x"38",x"56",x"2D",x"2E",x"17",x"1F",x"00",x"02",x"06",x"0F",x"8F",x"66",x"44",x"CC",
		x"0B",x"0C",x"04",x"04",x"00",x"00",x"00",x"00",x"BC",x"6C",x"24",x"D2",x"6A",x"6C",x"C8",x"00",
		x"80",x"E0",x"38",x"77",x"2F",x"2C",x"17",x"1B",x"00",x"00",x"02",x"06",x"8F",x"66",x"84",x"8C",
		x"0B",x"0F",x"06",x"05",x"01",x"01",x"00",x"00",x"8C",x"7C",x"14",x"2A",x"2A",x"EC",x"E8",x"00",
		x"80",x"F0",x"28",x"72",x"2D",x"28",x"1B",x"13",x"00",x"00",x"00",x"02",x"C6",x"E6",x"04",x"8C",
		x"0B",x"0E",x"04",x"04",x"01",x"01",x"00",x"00",x"BC",x"6C",x"24",x"D2",x"8A",x"8C",x"C8",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"01",x"01",x"19",x"18",x"3A",x"3A",x"00",x"00",x"80",x"80",x"98",x"38",x"60",x"00",
		x"01",x"08",x"18",x"19",x"01",x"01",x"00",x"00",x"7C",x"1C",x"18",x"98",x"80",x"80",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"13",x"27",x"2F",x"2F",x"00",x"00",x"E0",x"10",x"88",x"C4",x"C4",x"E4",
		x"2F",x"2F",x"27",x"13",x"0F",x"07",x"00",x"00",x"E4",x"E4",x"C4",x"88",x"10",x"E0",x"00",x"00",
		x"CC",x"CC",x"C8",x"C8",x"C8",x"C8",x"C8",x"C0",x"C0",x"40",x"00",x"80",x"80",x"80",x"80",x"00",
		x"C4",x"CC",x"CC",x"4C",x"00",x"00",x"00",x"00",x"40",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",
		x"C0",x"CC",x"CC",x"CC",x"CC",x"C0",x"C0",x"CC",x"00",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"C0",
		x"CC",x"CC",x"CC",x"C0",x"C0",x"CC",x"CC",x"CC",x"C0",x"C0",x"C0",x"00",x"00",x"C0",x"C0",x"C0",
		x"C0",x"C0",x"CC",x"CC",x"CC",x"CC",x"C0",x"C0",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"80",x"00",
		x"CC",x"CC",x"CC",x"CC",x"C0",x"C0",x"CC",x"C0",x"00",x"40",x"C0",x"C0",x"00",x"00",x"C0",x"00",
		x"00",x"00",x"00",x"00",x"4C",x"CC",x"CC",x"C0",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",
		x"C0",x"C0",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"80",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"33",x"20",x"00",x"13",x"13",x"13",x"13",x"03",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"23",x"33",x"33",x"33",x"00",x"00",x"00",x"00",x"30",x"30",x"30",x"20",x"00",x"00",x"00",x"00",
		x"20",x"02",x"12",x"12",x"02",x"20",x"30",x"33",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"13",x"13",x"13",x"00",x"00",x"13",x"13",x"13",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"00",x"00",x"13",x"13",x"13",x"33",x"21",x"01",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"00",x"12",x"12",x"12",x"00",x"00",x"33",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"00",x"00",x"00",x"00",x"33",x"33",x"33",x"01",x"00",x"00",x"00",x"00",x"20",x"30",x"30",x"30",
		x"00",x"00",x"33",x"33",x"33",x"13",x"13",x"13",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
		x"00",x"00",x"0C",x"0E",x"07",x"05",x"06",x"36",x"00",x"00",x"00",x"00",x"00",x"D9",x"DF",x"DE",
		x"0E",x"36",x"06",x"05",x"07",x"0E",x"0C",x"00",x"F8",x"DE",x"DF",x"D9",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"A0",x"D9",x"5F",x"DE",
		x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"F8",x"DE",x"5F",x"D9",x"A0",x"F0",x"F0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"1C",x"0E",x"0F",x"1B",
		x"00",x"E0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"18",x"1B",x"0F",x"0E",x"1C",x"00",x"00",x"00",
		x"00",x"00",x"01",x"01",x"00",x"16",x"1E",x"1E",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"F0",x"E0",
		x"02",x"1E",x"1E",x"16",x"00",x"01",x"01",x"00",x"F0",x"E0",x"E0",x"F0",x"E0",x"C0",x"80",x"00",
		x"00",x"00",x"03",x"03",x"03",x"02",x"03",x"13",x"00",x"00",x"40",x"E0",x"F8",x"FC",x"5E",x"5E",
		x"07",x"13",x"03",x"02",x"03",x"03",x"03",x"00",x"7E",x"5E",x"5E",x"FC",x"F8",x"E0",x"40",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"0F",x"00",x"3C",x"3E",x"4F",x"03",x"00",x"00",x"80",x"E0",x"30",x"18",x"88",x"CC",
		x"00",x"1C",x"1E",x"0E",x"06",x"00",x"00",x"00",x"C4",x"E4",x"74",x"74",x"30",x"30",x"40",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"20",x"11",x"09",x"03",x"08",x"1C",x"1E",x"00",x"00",x"80",x"80",x"3C",x"60",x"62",x"80",
		x"0B",x"09",x"01",x"00",x"00",x"00",x"00",x"21",x"90",x"98",x"62",x"20",x"9C",x"80",x"00",x"80",
		x"00",x"00",x"00",x"01",x"43",x"28",x"1C",x"1E",x"00",x"00",x"00",x"80",x"BC",x"30",x"40",x"81",
		x"03",x"01",x"01",x"10",x"20",x"40",x"00",x"00",x"90",x"D8",x"40",x"24",x"9C",x"80",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"08",x"1C",x"1E",x"00",x"00",x"00",x"00",x"BC",x"28",x"40",x"80",
		x"E3",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"D1",x"98",x"40",x"28",x"9C",x"00",x"00",x"00",
		x"00",x"00",x"80",x"01",x"03",x"08",x"1C",x"1E",x"00",x"00",x"00",x"80",x"BC",x"24",x"40",x"C0",
		x"03",x"09",x"09",x"28",x"40",x"00",x"00",x"00",x"90",x"99",x"00",x"30",x"9C",x"80",x"00",x"00",
		x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"20",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"02",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"20",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",
		x"01",x"09",x"0C",x"06",x"00",x"00",x"00",x"00",x"C0",x"C0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"02",x"09",x"0D",x"05",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"20",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"0E",x"05",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"00",x"00",
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"02",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"00",
		x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"20",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"0F",x"00",x"3C",x"3E",x"4F",x"01",x"00",x"00",x"80",x"E0",x"30",x"18",x"88",x"4C",
		x"01",x"1C",x"1E",x"0E",x"06",x"00",x"00",x"00",x"C4",x"64",x"74",x"74",x"30",x"30",x"40",x"00",
		x"00",x"00",x"0F",x"00",x"3C",x"3E",x"4F",x"05",x"00",x"00",x"80",x"E0",x"30",x"18",x"88",x"CC",
		x"03",x"1D",x"1E",x"0E",x"06",x"00",x"00",x"00",x"C4",x"64",x"74",x"74",x"30",x"30",x"40",x"00",
		x"00",x"00",x"0F",x"00",x"3C",x"3E",x"4C",x"07",x"00",x"00",x"80",x"E0",x"30",x"18",x"88",x"CC",
		x"07",x"1B",x"1D",x"0E",x"06",x"00",x"00",x"00",x"84",x"A4",x"F4",x"74",x"30",x"30",x"40",x"00",
		x"00",x"00",x"0F",x"00",x"3C",x"3D",x"4F",x"0F",x"00",x"00",x"80",x"E0",x"30",x"98",x"C8",x"EC",
		x"07",x"17",x"1B",x"0C",x"06",x"00",x"00",x"00",x"E4",x"C4",x"F4",x"F4",x"30",x"30",x"40",x"00",
		x"00",x"00",x"06",x"04",x"18",x"1C",x"0E",x"06",x"00",x"20",x"F0",x"F0",x"E0",x"00",x"20",x"30",
		x"26",x"34",x"18",x"1C",x"0E",x"06",x"00",x"00",x"F0",x"E0",x"C0",x"20",x"20",x"10",x"E0",x"C0",
		x"00",x"00",x"06",x"08",x"18",x"1C",x"0E",x"06",x"00",x"20",x"E0",x"D0",x"E0",x"00",x"20",x"30",
		x"34",x"38",x"1C",x"1E",x"0E",x"06",x"00",x"00",x"F0",x"E0",x"C0",x"20",x"30",x"30",x"E0",x"C0",
		x"00",x"00",x"02",x"00",x"1C",x"1C",x"0E",x"26",x"00",x"20",x"F0",x"F0",x"E0",x"00",x"20",x"20",
		x"32",x"38",x"1C",x"1E",x"0E",x"06",x"00",x"00",x"D0",x"E0",x"C0",x"20",x"30",x"30",x"E0",x"C0",
		x"00",x"00",x"02",x"04",x"1C",x"1C",x"0E",x"06",x"00",x"20",x"F0",x"F0",x"E0",x"00",x"20",x"30",
		x"22",x"34",x"1C",x"1C",x"0E",x"06",x"00",x"00",x"F0",x"E0",x"C0",x"20",x"20",x"10",x"E0",x"C0",
		x"00",x"00",x"06",x"06",x"1E",x"1C",x"0C",x"26",x"00",x"20",x"E0",x"D0",x"E0",x"00",x"20",x"30",
		x"36",x"3E",x"1C",x"1C",x"0E",x"06",x"00",x"00",x"F0",x"E0",x"C0",x"20",x"30",x"30",x"E0",x"C0",
		x"00",x"00",x"06",x"0E",x"0C",x"1C",x"2E",x"26",x"00",x"20",x"F0",x"F0",x"E0",x"00",x"20",x"20",
		x"36",x"3C",x"1C",x"1C",x"0E",x"06",x"00",x"00",x"D0",x"E0",x"C0",x"20",x"30",x"30",x"E0",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0C",x"14",x"0F",x"4F",x"07",x"00",x"00",x"80",x"D0",x"28",x"90",x"C8",x"EC",
		x"03",x"1D",x"0E",x"1E",x"0E",x"04",x"00",x"00",x"C4",x"A4",x"70",x"68",x"10",x"00",x"40",x"00",
		x"00",x"00",x"0E",x"1E",x"2C",x"32",x"0F",x"62",x"00",x"00",x"80",x"E8",x"34",x"18",x"68",x"F4",
		x"60",x"1C",x"16",x"0E",x"1F",x"0F",x"02",x"00",x"F4",x"64",x"14",x"74",x"38",x"30",x"40",x"00",
		x"00",x"03",x"07",x"07",x"3B",x"3C",x"7F",x"73",x"00",x"00",x"80",x"A0",x"B0",x"00",x"98",x"BC",
		x"78",x"6C",x"1F",x"0B",x"07",x"07",x"03",x"00",x"BC",x"D8",x"64",x"F4",x"F0",x"F0",x"C0",x"00",
		x"00",x"00",x"0D",x"01",x"3C",x"3E",x"7F",x"7B",x"00",x"C0",x"E0",x"E0",x"D0",x"18",x"86",x"DE",
		x"78",x"74",x"0E",x"0E",x"05",x"01",x"00",x"00",x"CE",x"E6",x"30",x"F4",x"F0",x"F0",x"C0",x"00",
		x"00",x"00",x"0F",x"10",x"3C",x"3E",x"4F",x"0F",x"00",x"00",x"E0",x"70",x"30",x"08",x"88",x"CC",
		x"1F",x"16",x"18",x"2E",x"16",x"00",x"00",x"00",x"C4",x"E4",x"74",x"3C",x"78",x"70",x"00",x"00",
		x"00",x"00",x"07",x"0E",x"38",x"3C",x"4F",x"07",x"00",x"00",x"80",x"D0",x"18",x"0C",x"80",x"CC",
		x"07",x"1F",x"1F",x"1E",x"0E",x"04",x"00",x"00",x"CC",x"FC",x"F8",x"78",x"30",x"20",x"40",x"00",
		x"00",x"01",x"07",x"0E",x"30",x"3E",x"4F",x"03",x"00",x"00",x"80",x"E0",x"70",x"F8",x"78",x"74",
		x"1C",x"1E",x"1F",x"1F",x"0E",x"00",x"00",x"00",x"86",x"EC",x"6C",x"58",x"10",x"20",x"40",x"00",
		x"00",x"00",x"05",x"0E",x"1E",x"04",x"4F",x"03",x"00",x"00",x"B0",x"78",x"7C",x"3C",x"98",x"C4",
		x"1E",x"3F",x"1F",x"2F",x"17",x"0E",x"00",x"00",x"C4",x"E6",x"EC",x"D8",x"10",x"00",x"40",x"00",
		x"00",x"00",x"05",x"0C",x"18",x"16",x"0F",x"07",x"00",x"40",x"B0",x"B8",x"1C",x"0C",x"84",x"CC",
		x"1F",x"1F",x"1F",x"0F",x"07",x"00",x"00",x"00",x"C4",x"E4",x"E8",x"D8",x"30",x"00",x"40",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"00",x"07",x"04",x"00",x"00",x"00",x"00",x"00",x"40",x"C0",x"40",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"05",x"05",x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"05",x"05",x"00",x"00",x"00",x"00",x"00",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"05",x"05",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"05",x"05",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"00",x"07",x"04",x"00",x"C0",x"40",x"C0",x"00",x"40",x"C0",x"40",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"05",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"40",x"C0",x"00",x"00",x"00",x"00",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"00",x"07",x"04",x"00",x"C0",x"40",x"C0",x"00",x"40",x"C0",x"40",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"05",x"05",x"00",x"00",x"07",x"04",x"00",x"40",x"40",x"C0",x"00",x"40",x"C0",x"40",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"07",x"05",x"05",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"40",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"07",x"05",x"05",x"00",x"C0",x"40",x"C0",x"00",x"40",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"07",x"04",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"C0",
		x"00",x"07",x"04",x"07",x"00",x"05",x"05",x"07",x"00",x"C0",x"40",x"C0",x"00",x"C0",x"40",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"07",x"05",x"05",x"00",x"01",x"00",x"01",x"00",x"40",x"40",x"C0",x"00",x"40",x"80",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"07",x"05",x"05",x"00",x"01",x"00",x"01",x"00",x"C0",x"40",x"40",x"00",x"40",x"80",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"00",x"07",x"00",x"01",x"00",x"01",x"00",x"C0",x"80",x"80",x"00",x"40",x"80",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"05",x"05",x"07",x"00",x"01",x"00",x"01",x"00",x"C0",x"40",x"40",x"00",x"40",x"80",x"40",
		x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"10",x"11",x"11",x"01",x"01",
		x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"0F",x"08",x"08",x"25",x"11",x"C9",x"20",x"03",x"3B",
		x"00",x"00",x"00",x"08",x"88",x"88",x"80",x"80",x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"80",
		x"10",x"10",x"A4",x"88",x"93",x"04",x"C0",x"DC",x"00",x"00",x"00",x"38",x"00",x"00",x"00",x"F0",
		x"0F",x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"3B",x"03",x"20",x"C9",x"11",x"25",x"08",x"08",
		x"01",x"02",x"04",x"08",x"00",x"00",x"00",x"00",x"01",x"01",x"11",x"11",x"10",x"00",x"00",x"00",
		x"DC",x"C0",x"04",x"93",x"88",x"A4",x"10",x"10",x"F0",x"00",x"00",x"00",x"38",x"00",x"00",x"00",
		x"80",x"80",x"88",x"88",x"08",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"00",x"00",x"00",x"00",
		x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",x"00",x"01",x"21",x"21",x"20",x"01",x"01",x"11",
		x"00",x"00",x"1C",x"01",x"00",x"00",x"00",x"73",x"90",x"48",x"20",x"80",x"40",x"00",x"00",x"80",
		x"00",x"80",x"80",x"84",x"04",x"04",x"80",x"88",x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",
		x"89",x"12",x"04",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"1C",x"80",x"00",x"00",x"00",x"EE",
		x"77",x"00",x"00",x"00",x"01",x"38",x"00",x"00",x"00",x"00",x"00",x"40",x"80",x"20",x"48",x"91",
		x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",x"11",x"01",x"20",x"20",x"21",x"01",x"01",x"00",
		x"01",x"00",x"00",x"02",x"01",x"04",x"12",x"09",x"CE",x"00",x"00",x"00",x"80",x"38",x"00",x"00",
		x"88",x"80",x"80",x"04",x"84",x"84",x"80",x"00",x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"02",x"01",x"81",x"81",x"01",x"00",x"21",x"21",x"00",x"00",
		x"60",x"00",x"0C",x"00",x"00",x"00",x"00",x"EC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"84",x"84",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"40",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"30",x"00",x"00",x"00",x"00",x"37",
		x"EC",x"00",x"00",x"00",x"00",x"0C",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"02",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"21",x"21",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"37",x"00",x"00",x"00",x"00",x"30",x"00",x"06",
		x"00",x"00",x"84",x"84",x"00",x"80",x"81",x"81",x"80",x"40",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"00",x"00",x"81",x"81",x"01",x"00",x"00",x"00",x"00",x"00",
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
		x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
		x"00",x"00",x"00",x"00",x"00",x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"9B",x"FB",x"7A",x"1B",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"30",x"70",x"E0",x"C0",x"A0",x"60",x"E0",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"7A",x"FB",x"9B",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E0",x"60",x"A0",x"C0",x"E0",x"70",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"19",x"31",x"38",x"3D",x"1D",x"0D",x"0D",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"C0",x"C0",x"E0",x"A0",x"60",x"60",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0D",x"1D",x"3D",x"38",x"31",x"19",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"60",x"60",x"A0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"0C",x"8C",x"D8",x"F0",x"70",x"70",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"70",x"70",x"F0",x"D8",x"8C",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"18",x"1E",x"0F",x"07",x"03",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"06",x"0E",x"1C",x"38",x"70",x"70",x"70",x"B8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"1E",x"18",x"10",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"70",x"70",x"70",x"38",x"1C",x"0E",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"03",x"02",x"02",x"06",x"04",x"04",x"04",x"08",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"08",x"00",x"00",x"00",x"00",x"00",x"20",x"30",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"3F",x"1F",x"4F",x"07",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"83",x"F0",x"FE",x"FF",x"FF",x"FF",x"7F",x"7F",
		x"80",x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"70",x"70",x"70",x"F8",x"FE",x"FF",x"FF",x"FF",
		x"83",x"83",x"87",x"C7",x"43",x"60",x"38",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"02",x"02",x"02",x"03",x"07",x"87",x"E3",x"F8",x"7F",x"0F",x"01",x"1C",x"1F",x"1F",x"7F",x"7F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"80",x"80",x"00",x"C0",x"C0",x"C0",x"80",x"80",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"0F",x"0F",x"0F",x"87",x"87",x"87",x"C3",x"C3",x"FC",x"FC",x"FC",x"FC",x"FE",x"FE",x"FE",x"FE",
		x"C3",x"E3",x"E3",x"E1",x"E1",x"E1",x"F1",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"08",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"FF",
		x"F1",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"78",x"0B",x"C3",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"83",x"87",x"8E",x"9E",x"9A",x"9B",x"99",x"9C",x"FB",x"FA",x"F8",x"F8",x"78",x"38",x"3F",x"9F",
		x"9C",x"9E",x"98",x"9E",x"9F",x"80",x"98",x"9C",x"8F",x"45",x"01",x"00",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"0F",x"0F",x"1F",x"0F",x"C1",x"F8",x"F0",x"F0",x"E0",x"E0",x"E0",x"C0",x"C0",
		x"C0",x"80",x"00",x"30",x"4C",x"46",x"43",x"40",x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"80",x"81",x"00",x"C0",x"C0",x"80",x"00",x"00",
		x"9E",x"9E",x"9C",x"9C",x"98",x"98",x"90",x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",
		x"42",x"82",x"06",x"06",x"07",x"0F",x"0F",x"18",x"00",x"00",x"00",x"00",x"00",x"08",x"8E",x"07",
		x"00",x"00",x"00",x"40",x"80",x"80",x"80",x"00",x"03",x"00",x"00",x"00",x"01",x"03",x"17",x"17",
		x"3E",x"20",x"00",x"30",x"7E",x"7E",x"7C",x"00",x"00",x"0F",x"00",x"00",x"00",x"08",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3C",x"FC",x"FC",x"0C",x"0E",x"0E",x"8E",x"8E",x"1F",x"0F",x"0F",x"07",x"07",x"07",x"03",x"03",
		x"8F",x"8F",x"8F",x"0F",x"0F",x"0F",x"0F",x"0F",x"01",x"01",x"01",x"00",x"80",x"80",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"60",x"78",x"0F",x"00",x"00",x"C0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"04",x"0E",x"0E",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"C0",x"C0",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",
		x"0F",x"1F",x"1F",x"3F",x"3F",x"1F",x"1F",x"1F",x"F0",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"7F",x"38",x"1C",x"38",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"39",x"7B",x"4F",x"46",x"44",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"1F",x"3F",x"64",x"44",x"64",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"4F",x"4F",x"49",x"49",x"63",x"3E",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"78",x"7C",x"0E",x"07",x"0E",x"7C",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"7F",x"41",x"41",x"41",x"7F",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"02",x"04",x"09",x"12",x"24",x"49",x"92",x"FF",x"00",x"FF",x"00",x"7F",x"80",x"3F",x"40",
		x"A4",x"A9",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"00",x"FF",x"00",x"FE",x"01",x"FC",x"02",x"80",x"40",x"20",x"90",x"48",x"24",x"92",x"49",
		x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"95",x"55",x"55",x"55",x"55",x"55",x"55",
		x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"A9",x"A4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",
		x"92",x"49",x"24",x"12",x"09",x"04",x"02",x"01",x"40",x"3F",x"80",x"7F",x"00",x"FF",x"00",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"55",x"55",x"55",x"55",x"55",x"55",x"95",x"25",
		x"02",x"FC",x"01",x"FE",x"00",x"FF",x"00",x"FF",x"49",x"92",x"24",x"48",x"90",x"20",x"40",x"80",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"30",x"30",x"3F",x"3F",x"00",x"00",
		x"33",x"33",x"30",x"30",x"3F",x"3F",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"00",x"00",x"3F",x"3F",x"30",x"30",x"33",x"33",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"00",x"00",x"3F",x"3F",x"30",x"30",x"33",x"33",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",x"33",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",
		x"CC",x"CC",x"0C",x"0C",x"FC",x"FC",x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"CC",x"CC",x"0C",x"0C",x"FC",x"FC",x"00",x"00",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FC",x"FC",x"0C",x"0C",x"CC",x"CC",
		x"00",x"00",x"FC",x"FC",x"0C",x"0C",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9C",x"80",x"80",x"F0",x"F0",x"F1",x"F7",x"87",x"03",x"03",x"00",
		x"80",x"80",x"81",x"87",x"9F",x"9F",x"9F",x"9F",x"0C",x"3E",x"FE",x"F8",x"FA",x"FB",x"FB",x"FB",
		x"04",x"3C",x"FC",x"FC",x"F8",x"E0",x"80",x"00",x"80",x"F0",x"C1",x"07",x"1E",x"3C",x"78",x"11",
		x"06",x"0E",x"06",x"00",x"00",x"F8",x"E0",x"C1",x"03",x"00",x"0F",x"00",x"00",x"00",x"F8",x"F8",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FB",x"FB",x"F8",x"F8",x"E0",x"C0",x"80",x"01",
		x"9C",x"98",x"80",x"80",x"80",x"80",x"80",x"81",x"03",x"07",x"0F",x"1E",x"3E",x"78",x"FB",x"FB",
		x"83",x"07",x"0F",x"1F",x"3F",x"7F",x"1F",x"C6",x"F0",x"F0",x"E1",x"C3",x"83",x"07",x"0E",x"0F",
		x"F0",x"FC",x"E0",x"00",x"00",x"00",x"81",x"03",x"1F",x"3E",x"3E",x"06",x"3C",x"FC",x"F8",x"F8",
		x"00",x"00",x"80",x"98",x"3F",x"7A",x"F6",x"F6",x"A8",x"28",x"28",x"28",x"68",x"68",x"4C",x"4C",
		x"EC",x"4C",x"08",x"00",x"00",x"00",x"00",x"60",x"CC",x"CC",x"CC",x"CC",x"0C",x"04",x"00",x"00",
		x"3C",x"1F",x"4F",x"27",x"23",x"31",x"38",x"3C",x"3F",x"0F",x"C3",x"F0",x"FC",x"FE",x"F8",x"40",
		x"3C",x"3E",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"00",x"0E",x"0F",x"07",x"43",x"41",x"60",x"70",
		x"E3",x"E3",x"C3",x"C3",x"87",x"87",x"07",x"07",x"80",x"8E",x"8E",x"8E",x"8E",x"8F",x"0F",x"0F",
		x"00",x"08",x"0E",x"0F",x"1F",x"1F",x"1E",x"1E",x"0F",x"00",x"00",x"00",x"00",x"08",x"0E",x"0F",
		x"07",x"07",x"03",x"03",x"01",x"01",x"01",x"00",x"78",x"7C",x"7C",x"3E",x"1F",x"1F",x"00",x"FF",
		x"70",x"70",x"F0",x"30",x"08",x"08",x"08",x"B8",x"FF",x"7F",x"7F",x"7F",x"3F",x"3F",x"1F",x"1F",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"8F",x"83",x"81",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"80",x"80",x"80",x"98",x"9E",x"9F",x"9F",x"7F",x"3F",x"0F",x"03",x"00",x"00",x"C0",x"F0",
		x"01",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F",x"0F",
		x"FE",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",x"07",x"07",x"03",x"81",x"C1",x"E0",x"F0",x"F8",x"FC",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FC",x"FF",x"FF",x"FF",x"FE",x"FC",x"FD",x"F9",
		x"80",x"80",x"80",x"80",x"9F",x"9F",x"9F",x"9F",x"7B",x"00",x"00",x"00",x"F7",x"F7",x"F7",x"F0",
		x"00",x"80",x"80",x"04",x"00",x"00",x"C0",x"F8",x"7E",x"1F",x"07",x"02",x"00",x"00",x"03",x"01",
		x"FF",x"3F",x"00",x"00",x"FC",x"FC",x"C0",x"00",x"80",x"F8",x"1F",x"00",x"9F",x"00",x"07",x"06",
		x"07",x"87",x"87",x"C7",x"C3",x"C3",x"E3",x"E2",x"D0",x"D1",x"D1",x"D1",x"D1",x"81",x"81",x"00",
		x"E0",x"F0",x"F0",x"F8",x"F8",x"78",x"7C",x"3C",x"60",x"70",x"33",x"33",x"33",x"33",x"33",x"33",
		x"03",x"00",x"C0",x"E0",x"C0",x"C0",x"C3",x"47",x"00",x"00",x"10",x"1E",x"10",x"03",x"01",x"00",
		x"06",x"06",x"10",x"00",x"07",x"00",x"00",x"00",x"10",x"3C",x"7E",x"7C",x"18",x"C1",x"01",x"00",
		x"E0",x"80",x"00",x"04",x"62",x"32",x"88",x"E4",x"B2",x"B2",x"96",x"96",x"D4",x"55",x"55",x"54",
		x"7A",x"1C",x"C2",x"00",x"FF",x"02",x"00",x"09",x"55",x"55",x"38",x"17",x"C0",x"21",x"98",x"48",
		x"60",x"EF",x"DE",x"BC",x"F9",x"73",x"E6",x"CC",x"00",x"00",x"20",x"78",x"E0",x"81",x"1F",x"F8",
		x"9B",x"40",x"80",x"C6",x"00",x"C7",x"47",x"11",x"80",x"03",x"7F",x"07",x"00",x"FC",x"FE",x"FF",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"8F",x"8F",x"87",x"83",x"81",x"80",x"80",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",
		x"E0",x"F0",x"F0",x"F8",x"F8",x"F8",x"FC",x"FC",x"07",x"07",x"07",x"07",x"03",x"03",x"03",x"03",
		x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"00",x"80",x"80",x"80",
		x"80",x"80",x"80",x"80",x"80",x"90",x"98",x"9C",x"3F",x"1F",x"0F",x"0F",x"07",x"03",x"01",x"00",
		x"9E",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F8",
		x"FF",x"7F",x"3F",x"1F",x"0F",x"0F",x"07",x"03",x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"70",x"70",x"70",x"60",x"00",x"90",x"30",x"70",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"70",x"70",x"70",x"30",x"B0",x"90",x"D0",x"C0",
		x"0F",x"0F",x"1F",x"1F",x"1F",x"03",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"00",x"C0",
		x"01",x"13",x"07",x"07",x"01",x"00",x"00",x"30",x"FF",x"FE",x"F8",x"F0",x"F8",x"3C",x"02",x"00",
		x"7F",x"7F",x"7F",x"7F",x"3F",x"3F",x"3F",x"3F",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"0F",x"C0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
		x"3E",x"3E",x"7E",x"7E",x"7C",x"7C",x"1C",x"04",x"00",x"00",x"07",x"07",x"07",x"0F",x"0F",x"1F",
		x"00",x"78",x"D8",x"C8",x"C0",x"E0",x"F0",x"F6",x"1F",x"1F",x"00",x"3F",x"5E",x"0C",x"08",x"00",
		x"0F",x"38",x"60",x"43",x"C7",x"8F",x"9F",x"9F",x"FF",x"00",x"00",x"00",x"00",x"80",x"80",x"80",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"C0",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F8",
		x"FF",x"00",x"00",x"07",x"03",x"03",x"03",x"03",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7F",x"7F",x"7F",x"3F",x"3F",x"3F",x"3F",
		x"00",x"80",x"80",x"80",x"C0",x"C0",x"E0",x"E0",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"0F",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"F0",x"F0",x"C0",x"C0",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"40",x"60",x"70",x"70",x"70",x"70",x"70",x"70",
		x"FF",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"01",x"03",x"03",x"03",x"03",x"01",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"70",x"70",x"10",x"C0",x"E0",x"F0",x"F0",x"C0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"60",x"70",x"70",x"70",x"70",x"70",
		x"00",x"00",x"00",x"04",x"06",x"07",x"07",x"07",x"7F",x"3F",x"0E",x"04",x"00",x"80",x"C4",x"EC",
		x"07",x"07",x"07",x"01",x"00",x"0F",x"0F",x"0F",x"F8",x"F8",x"F8",x"F8",x"70",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"0D",x"00",x"00",x"78",x"E4",x"92",x"86",x"09",x"10",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"60",x"F0",x"96",x"8B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"14",x"28",x"28",x"24",x"02",x"03",x"05",x"06",x"90",x"01",x"40",x"88",x"88",x"45",x"37",x"87",
		x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"38",x"01",x"03",x"00",x"00",x"00",x"00",
		x"91",x"05",x"0A",x"26",x"98",x"80",x"08",x"18",x"08",x"A0",x"60",x"00",x"00",x"00",x"00",x"00",
		x"A0",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"02",x"42",x"23",x"1F",x"0C",x"06",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"10",x"30",x"E0",x"BF",x"06",x"0C",x"18",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"06",x"0C",x"19",x"3F",x"02",x"02",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"03",x"8F",x"DC",x"78",x"34",x"22",x"01",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"42",x"00",x"40",x"00",
		x"00",x"00",x"09",x"00",x"00",x"02",x"00",x"24",x"00",x"04",x"00",x"00",x"20",x"02",x"00",x"88",
		x"00",x"00",x"00",x"40",x"00",x"00",x"02",x"90",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",
		x"00",x"00",x"10",x"82",x"00",x"00",x"50",x"00",x"00",x"20",x"00",x"00",x"88",x"00",x"00",x"02",
		x"00",x"10",x"00",x"01",x"00",x"10",x"02",x"00",x"02",x"00",x"10",x"00",x"40",x"01",x"00",x"00",
		x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"08",x"00",x"40",x"08",x"00",x"01",x"00",
		x"04",x"01",x"40",x"00",x"00",x"08",x"00",x"00",x"10",x"00",x"00",x"08",x"00",x"40",x"00",x"00",
		x"10",x"00",x"04",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1E",x"0F",x"13",x"13",x"6E",x"00",x"00",x"30",x"1B",x"89",x"C1",x"B1",x"8F",
		x"7E",x"62",x"62",x"32",x"1C",x"00",x"00",x"00",x"87",x"31",x"3D",x"CB",x"4B",x"30",x"00",x"00",
		x"00",x"00",x"00",x"3C",x"1E",x"26",x"26",x"DC",x"00",x"0C",x"36",x"4B",x"8F",x"CC",x"B0",x"84",
		x"FC",x"C4",x"C4",x"64",x"38",x"00",x"00",x"00",x"84",x"16",x"2B",x"CD",x"4C",x"2C",x"08",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"02",x"00",x"00",x"00",x"00",x"08",x"28",x"29",x"D9",
		x"12",x"72",x"6C",x"78",x"7C",x"3E",x"1C",x"00",x"AF",x"AB",x"EB",x"6F",x"7F",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"10",x"1E",x"02",x"00",x"00",x"00",x"00",x"0A",x"2A",x"29",x"D9",
		x"12",x"72",x"6C",x"78",x"7C",x"3E",x"1C",x"00",x"A9",x"AC",x"AB",x"69",x"79",x"39",x"07",x"00",
		x"00",x"00",x"00",x"00",x"00",x"12",x"1E",x"02",x"00",x"00",x"00",x"03",x"0F",x"2B",x"29",x"DD",
		x"12",x"72",x"6C",x"78",x"7C",x"3E",x"1C",x"00",x"AF",x"AC",x"EF",x"69",x"79",x"09",x"0D",x"0E",
		x"00",x"1C",x"3E",x"7C",x"78",x"6C",x"72",x"12",x"00",x"00",x"00",x"7F",x"6F",x"EB",x"AB",x"AF",
		x"1E",x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"D9",x"29",x"28",x"08",x"00",x"00",x"00",x"00",
		x"00",x"1C",x"3E",x"7C",x"78",x"6C",x"72",x"12",x"00",x"07",x"39",x"79",x"69",x"AB",x"AC",x"A9",
		x"1E",x"02",x"12",x"00",x"00",x"00",x"00",x"00",x"D9",x"29",x"2A",x"0A",x"00",x"00",x"00",x"00",
		x"00",x"1C",x"3E",x"7C",x"78",x"6C",x"72",x"12",x"0E",x"0D",x"09",x"79",x"69",x"EF",x"AC",x"AF",
		x"1E",x"02",x"12",x"00",x"00",x"00",x"00",x"00",x"DD",x"29",x"29",x"0D",x"03",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"04",x"04",x"00",x"00",x"00",x"00",x"60",x"F0",x"90",x"90",
		x"04",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"90",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"18",x"30",x"24",x"04",x"00",x"00",x"F0",x"F0",x"00",x"00",x"90",x"90",
		x"04",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"90",x"F8",x"F8",x"F0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"F0",x"0E",x"0E",
		x"00",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"0E",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"1B",x"3F",x"3C",x"34",x"00",x"00",x"F0",x"F8",x"6C",x"FE",x"9E",x"96",
		x"34",x"3F",x"3F",x"1F",x"08",x"00",x"00",x"00",x"96",x"FE",x"FE",x"FC",x"08",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"10",x"90",x"90",x"90",
		x"04",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"90",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"18",x"30",x"24",x"04",x"00",x"00",x"F0",x"F0",x"00",x"00",x"90",x"90",
		x"04",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"90",x"F8",x"F8",x"F0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"90",x"0E",x"0E",
		x"00",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"0E",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"1C",x"3C",x"3C",x"34",x"00",x"00",x"F0",x"F8",x"1C",x"9E",x"9E",x"96",
		x"34",x"3F",x"3F",x"1F",x"08",x"00",x"00",x"00",x"96",x"FE",x"FE",x"FC",x"08",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"06",x"04",x"04",x"00",x"00",x"00",x"00",x"60",x"F0",x"90",x"90",
		x"04",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"90",x"B0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"18",x"30",x"24",x"04",x"00",x"00",x"F0",x"F0",x"00",x"00",x"90",x"90",
		x"04",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"90",x"B8",x"F8",x"F0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"F0",x"0E",x"0E",
		x"00",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"0E",x"B0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"1A",x"3E",x"3C",x"34",x"00",x"00",x"F0",x"F8",x"6C",x"FE",x"9E",x"96",
		x"34",x"3F",x"3F",x"1F",x"08",x"00",x"00",x"00",x"96",x"BE",x"FE",x"FC",x"08",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"70",x"7A",x"C7",x"C7",x"00",x"00",x"1C",x"1C",x"3C",x"24",x"20",x"20",
		x"FF",x"C7",x"C7",x"7A",x"70",x"E0",x"00",x"00",x"24",x"20",x"20",x"24",x"3C",x"1C",x"18",x"00",
		x"00",x"00",x"00",x"E1",x"70",x"7E",x"C7",x"C7",x"00",x"18",x"FC",x"FC",x"F8",x"24",x"20",x"20",
		x"FF",x"C7",x"C7",x"7E",x"70",x"E0",x"00",x"00",x"24",x"20",x"20",x"24",x"FC",x"F8",x"38",x"08",
		x"00",x"00",x"00",x"1C",x"0E",x"0F",x"18",x"38",x"00",x"00",x"00",x"06",x"02",x"D0",x"D0",x"D4",
		x"3E",x"38",x"18",x"0F",x"0E",x"1C",x"00",x"00",x"D6",x"D4",x"D0",x"D0",x"02",x"06",x"00",x"00",
		x"00",x"00",x"00",x"24",x"46",x"E7",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"2C",
		x"FF",x"7D",x"78",x"E0",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"30",x"38",x"1C",x"0C",x"00",
		x"00",x"00",x"00",x"24",x"46",x"E7",x"FF",x"FF",x"00",x"00",x"00",x"00",x"20",x"20",x"A0",x"20",
		x"FF",x"7D",x"78",x"E0",x"00",x"00",x"00",x"00",x"20",x"00",x"04",x"84",x"7C",x"3C",x"18",x"00",
		x"00",x"00",x"00",x"24",x"46",x"E7",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"20",x"A0",x"20",
		x"FF",x"7D",x"79",x"E0",x"00",x"00",x"00",x"00",x"20",x"A0",x"E0",x"F8",x"3C",x"08",x"00",x"00",
		x"00",x"00",x"00",x"24",x"46",x"E7",x"FF",x"FF",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",
		x"FF",x"7D",x"79",x"F0",x"00",x"00",x"00",x"00",x"00",x"04",x"9C",x"FC",x"7C",x"18",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"78",x"7D",x"FF",x"00",x"0C",x"1C",x"38",x"30",x"20",x"20",x"24",
		x"FF",x"FF",x"E7",x"46",x"24",x"00",x"00",x"00",x"2C",x"24",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"78",x"7D",x"FF",x"00",x"18",x"3C",x"7C",x"84",x"04",x"00",x"20",
		x"FF",x"FF",x"E7",x"46",x"24",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"79",x"7D",x"FF",x"00",x"00",x"08",x"3C",x"F8",x"E0",x"A0",x"20",
		x"FF",x"FF",x"E7",x"46",x"24",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"79",x"7D",x"FF",x"00",x"00",x"18",x"7C",x"9C",x"9C",x"04",x"00",
		x"FF",x"FF",x"E7",x"46",x"24",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"70",x"38",x"3F",x"63",x"E3",x"00",x"06",x"1E",x"3C",x"7E",x"12",x"90",x"90",
		x"FF",x"E3",x"63",x"3F",x"38",x"70",x"00",x"00",x"92",x"90",x"90",x"12",x"7C",x"3E",x"0E",x"00",
		x"00",x"60",x"78",x"FC",x"FE",x"7F",x"F1",x"F1",x"00",x"00",x"00",x"00",x"00",x"88",x"C8",x"C8",
		x"FF",x"F1",x"F1",x"7F",x"FE",x"FC",x"78",x"00",x"C8",x"C8",x"C8",x"88",x"00",x"00",x"00",x"00",
		x"00",x"00",x"3D",x"47",x"C7",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"90",x"10",x"B0",x"A0",
		x"7F",x"3F",x"3A",x"70",x"01",x"00",x"00",x"00",x"A2",x"22",x"62",x"32",x"38",x"1C",x"3E",x"1C",
		x"00",x"00",x"00",x"00",x"E0",x"78",x"46",x"C6",x"00",x"00",x"00",x"00",x"00",x"40",x"64",x"22",
		x"FF",x"E3",x"E3",x"FF",x"7E",x"3D",x"38",x"70",x"20",x"20",x"20",x"26",x"26",x"06",x"86",x"3C",
		x"00",x"00",x"00",x"01",x"00",x"72",x"3F",x"3F",x"1C",x"3E",x"1C",x"38",x"32",x"62",x"22",x"A2",
		x"7F",x"FF",x"FF",x"C7",x"47",x"3D",x"00",x"00",x"A0",x"B0",x"10",x"90",x"00",x"00",x"00",x"00",
		x"70",x"38",x"3D",x"7E",x"FF",x"E3",x"E3",x"FE",x"3C",x"86",x"06",x"2E",x"26",x"20",x"20",x"20",
		x"C7",x"46",x"78",x"E0",x"00",x"00",x"00",x"00",x"22",x"64",x"40",x"00",x"00",x"00",x"00",x"00",
		x"40",x"46",x"47",x"67",x"67",x"66",x"76",x"74",x"F3",x"0C",x"30",x"C0",x"C0",x"40",x"40",x"40",
		x"78",x"7C",x"7C",x"7C",x"19",x"07",x"04",x"04",x"40",x"00",x"00",x"00",x"00",x"80",x"A0",x"30",
		x"03",x"22",x"25",x"36",x"36",x"38",x"3C",x"3C",x"E0",x"18",x"8E",x"70",x"40",x"40",x"40",x"40",
		x"3C",x"3C",x"3C",x"1E",x"01",x"07",x"04",x"04",x"40",x"00",x"00",x"00",x"00",x"80",x"A0",x"30",
		x"03",x"16",x"1F",x"1B",x"1C",x"1E",x"1E",x"1F",x"80",x"40",x"A0",x"E8",x"9C",x"C0",x"40",x"40",
		x"1F",x"1F",x"1C",x"1C",x"01",x"07",x"04",x"04",x"40",x"00",x"00",x"00",x"00",x"80",x"E0",x"30",
		x"10",x"30",x"20",x"60",x"7F",x"1F",x"04",x"04",x"00",x"00",x"00",x"00",x"80",x"C0",x"FC",x"10",
		x"0C",x"17",x"30",x"60",x"20",x"30",x"10",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"06",x"0C",x"18",x"18",x"1F",x"0F",x"04",x"04",x"00",x"00",x"00",x"00",x"80",x"C0",x"F8",x"10",
		x"0C",x"0F",x"18",x"18",x"18",x"0C",x"06",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"16",x"18",x"18",x"1F",x"0F",x"04",x"04",x"00",x"00",x"00",x"00",x"80",x"C0",x"F0",x"10",
		x"0C",x"0F",x"18",x"18",x"18",x"1E",x"07",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"80",x"00",
		x"40",x"47",x"67",x"64",x"74",x"7C",x"7E",x"7E",x"00",x"00",x"88",x"E0",x"40",x"40",x"40",x"40",
		x"1E",x"07",x"05",x"16",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"00",x"00",
		x"00",x"00",x"04",x"24",x"16",x"05",x"07",x"1E",x"00",x"00",x"20",x"40",x"80",x"00",x"00",x"00",
		x"7E",x"7E",x"7C",x"74",x"64",x"67",x"47",x"40",x"40",x"40",x"40",x"40",x"E0",x"88",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"70",x"7E",x"C7",x"C7",x"00",x"00",x"0C",x"1C",x"1C",x"04",x"20",x"20",
		x"FF",x"C7",x"C7",x"7E",x"70",x"E0",x"00",x"00",x"24",x"20",x"20",x"04",x"1C",x"1C",x"08",x"00",
		x"00",x"00",x"00",x"70",x"38",x"3C",x"7E",x"FF",x"00",x"1C",x"3C",x"70",x"70",x"20",x"20",x"24",
		x"C7",x"C7",x"FF",x"44",x"78",x"F0",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E1",x"70",x"7E",x"C3",x"C3",x"00",x"18",x"FC",x"FC",x"F8",x"24",x"20",x"20",
		x"FB",x"C3",x"C3",x"7E",x"70",x"E0",x"00",x"00",x"24",x"20",x"20",x"24",x"FC",x"F8",x"38",x"08",
		x"00",x"03",x"01",x"01",x"01",x"03",x"02",x"3C",x"00",x"E0",x"F0",x"F8",x"BC",x"24",x"20",x"F0",
		x"7C",x"7E",x"7E",x"3F",x"1F",x"0F",x"02",x"00",x"F0",x"60",x"64",x"3C",x"08",x"60",x"00",x"00",
		x"00",x"03",x"01",x"01",x"01",x"03",x"02",x"3C",x"00",x"E0",x"F1",x"FF",x"BC",x"24",x"21",x"F0",
		x"7C",x"7E",x"7E",x"3F",x"1F",x"0F",x"02",x"00",x"F0",x"60",x"64",x"3C",x"08",x"61",x"00",x"00",
		x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"38",x"00",x"E0",x"F0",x"78",x"3C",x"24",x"00",x"10",
		x"7C",x"7E",x"7E",x"3F",x"1F",x"0F",x"02",x"00",x"10",x"00",x"04",x"0C",x"08",x"00",x"00",x"00",
		x"00",x"07",x"03",x"1B",x"27",x"76",x"64",x"79",x"00",x"CA",x"E4",x"F8",x"78",x"48",x"40",x"E0",
		x"F9",x"FC",x"FC",x"7E",x"3E",x"1E",x"04",x"00",x"E0",x"C0",x"C8",x"78",x"1C",x"C4",x"0A",x"00",
		x"00",x"90",x"08",x"27",x"30",x"20",x"08",x"1C",x"00",x"02",x"04",x"0A",x"44",x"62",x"00",x"39",
		x"0C",x"0B",x"03",x"06",x"00",x"00",x"00",x"00",x"79",x"89",x"09",x"02",x"02",x"C0",x"D0",x"00",
		x"00",x"B0",x"44",x"67",x"10",x"10",x"18",x"18",x"00",x"00",x"02",x"04",x"C2",x"54",x"00",x"39",
		x"04",x"07",x"07",x"06",x"01",x"01",x"00",x"00",x"79",x"89",x"09",x"02",x"82",x"80",x"10",x"00",
		x"00",x"B0",x"4C",x"46",x"11",x"30",x"18",x"14",x"00",x"00",x"00",x"02",x"C4",x"32",x"00",x"39",
		x"04",x"0C",x"05",x"06",x"00",x"00",x"00",x"00",x"49",x"89",x"09",x"C2",x"C2",x"00",x"30",x"00",
		x"00",x"A0",x"4C",x"41",x"31",x"30",x"14",x"0C",x"00",x"00",x"00",x"00",x"82",x"70",x"00",x"39",
		x"0C",x"0D",x"03",x"02",x"00",x"00",x"00",x"00",x"79",x"89",x"09",x"02",x"62",x"60",x"10",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"03",x"0F",x"07",x"00",x"39",x"3A",x"00",x"00",x"80",x"80",x"80",x"00",x"1C",x"7C",
		x"3B",x"30",x"00",x"01",x"01",x"01",x"00",x"00",x"7C",x"1C",x"00",x"E0",x"F0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"08",x"18",x"20",x"23",x"22",x"00",x"00",x"E0",x"10",x"28",x"24",x"F4",x"74",
		x"20",x"23",x"22",x"10",x"08",x"07",x"00",x"00",x"74",x"F4",x"64",x"28",x"10",x"E0",x"00",x"00",
		x"00",x"00",x"04",x"04",x"04",x"04",x"04",x"0C",x"00",x"80",x"C0",x"40",x"40",x"40",x"40",x"C0",
		x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"00",x"00",x"00",x"00",x"0C",x"0C",x"00",x"C0",x"00",x"00",x"00",x"00",x"C0",x"C0",x"00",
		x"00",x"00",x"00",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"00",x"00",x"00",
		x"0C",x"0C",x"00",x"00",x"00",x"00",x"0C",x"0C",x"C0",x"C0",x"00",x"00",x"00",x"00",x"40",x"C0",
		x"00",x"00",x"00",x"00",x"0C",x"0C",x"00",x"0C",x"C0",x"80",x"00",x"00",x"C0",x"C0",x"00",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"13",x"33",x"20",x"20",x"20",x"20",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"13",x"31",x"21",x"21",x"31",x"13",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"20",x"20",x"33",x"33",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"20",x"20",x"20",x"00",x"12",x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"21",x"21",x"21",x"33",x"33",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"33",x"33",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E1",x"70",x"7E",x"C7",x"C7",x"00",x"18",x"FC",x"FC",x"F8",x"24",x"20",x"20",
		x"FF",x"C7",x"C7",x"7E",x"70",x"E0",x"00",x"00",x"24",x"20",x"20",x"24",x"FC",x"F8",x"38",x"08",
		x"00",x"00",x"00",x"1C",x"0E",x"1F",x"3E",x"3E",x"00",x"18",x"0C",x"0C",x"5E",x"26",x"20",x"20",
		x"3F",x"3E",x"3E",x"1F",x"0E",x"1C",x"00",x"00",x"A4",x"20",x"20",x"26",x"5E",x"0C",x"0C",x"18",
		x"00",x"18",x"3F",x"3F",x"1F",x"3F",x"1F",x"3F",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"88",x"88",
		x"3F",x"1F",x"3F",x"3F",x"1F",x"3F",x"3F",x"18",x"F8",x"88",x"88",x"F0",x"E0",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"00",x"06",x"07",x"0E",x"1F",x"1F",x"0F",x"1E",
		x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"0F",x"1F",x"1F",x"0E",x"1F",x"0F",x"07",x"02",
		x"00",x"00",x"00",x"70",x"38",x"3D",x"63",x"E3",x"00",x"04",x"1C",x"1C",x"04",x"00",x"A0",x"A0",
		x"FF",x"E3",x"63",x"3D",x"38",x"70",x"00",x"00",x"A0",x"A0",x"A0",x"00",x"04",x"1C",x"3C",x"18",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"00",x"30",x"7C",x"00",x"C0",x"F0",x"F8",x"3C",x"1C",x"0E",x"0E",
		x"7F",x"7F",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"06",x"06",x"84",x"84",x"C0",x"C0",x"80",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"11",x"09",x"03",x"00",x"00",x"00",x"00",x"80",x"80",x"F8",x"FC",x"E0",x"FE",x"BE",
		x"14",x"16",x"1E",x"0F",x"07",x"01",x"01",x"01",x"BE",x"BE",x"FE",x"C0",x"60",x"78",x"80",x"80",
		x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"F0",x"DC",x"BF",
		x"1C",x"1E",x"1E",x"0F",x"07",x"01",x"01",x"00",x"BE",x"FE",x"DC",x"C4",x"60",x"78",x"80",x"00",
		x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"FC",x"E8",x"DC",x"BE",
		x"1C",x"1E",x"1E",x"0F",x"07",x"00",x"00",x"00",x"FF",x"BE",x"DC",x"C8",x"60",x"38",x"00",x"00",
		x"00",x"00",x"01",x"41",x"23",x"10",x"00",x"00",x"00",x"00",x"80",x"F8",x"FC",x"E4",x"DC",x"FE",
		x"1C",x"16",x"16",x"07",x"07",x"01",x"00",x"00",x"BE",x"BF",x"9C",x"D0",x"60",x"78",x"00",x"00",
		x"00",x"00",x"06",x"0E",x"1F",x"1F",x"3F",x"3F",x"00",x"00",x"10",x"18",x"DC",x"FC",x"FE",x"FE",
		x"3F",x"3F",x"1F",x"1F",x"0F",x"07",x"00",x"00",x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"00",x"00",
		x"00",x"01",x"04",x"0E",x"1E",x"1E",x"3F",x"3F",x"00",x"C0",x"10",x"18",x"1C",x"1C",x"DE",x"FE",
		x"3F",x"3F",x"1F",x"1F",x"0F",x"07",x"01",x"00",x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"C0",x"00",
		x"00",x"01",x"07",x"0F",x"1C",x"1E",x"3E",x"3E",x"00",x"C0",x"F0",x"F8",x"1C",x"1C",x"1E",x"1E",
		x"3F",x"3F",x"1F",x"1F",x"0F",x"07",x"01",x"00",x"DE",x"FE",x"FC",x"FC",x"F8",x"F0",x"C0",x"00",
		x"00",x"01",x"07",x"0F",x"1F",x"1F",x"3C",x"3E",x"00",x"C0",x"F0",x"F8",x"FC",x"FC",x"1E",x"1E",
		x"3E",x"3E",x"1F",x"1F",x"0F",x"07",x"01",x"00",x"1E",x"1E",x"DC",x"FC",x"F8",x"F0",x"C0",x"00",
		x"00",x"01",x"07",x"0F",x"1F",x"1F",x"3F",x"3F",x"00",x"C0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",
		x"3C",x"3E",x"1E",x"1E",x"0F",x"07",x"01",x"00",x"1E",x"1E",x"1C",x"1C",x"D8",x"F0",x"C0",x"00",
		x"00",x"01",x"07",x"0F",x"1F",x"1F",x"3F",x"3F",x"00",x"C0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",
		x"3F",x"3F",x"1C",x"1E",x"0E",x"06",x"01",x"00",x"FE",x"FE",x"1C",x"1C",x"18",x"10",x"C0",x"00",
		x"00",x"00",x"07",x"0F",x"1F",x"1F",x"3F",x"3F",x"00",x"00",x"D0",x"F8",x"FC",x"FC",x"FE",x"FE",
		x"3F",x"3F",x"1F",x"1F",x"0C",x"06",x"00",x"00",x"FE",x"FE",x"FC",x"FC",x"18",x"10",x"00",x"00",
		x"00",x"00",x"06",x"0E",x"1F",x"1F",x"3F",x"3F",x"00",x"00",x"10",x"18",x"DC",x"FC",x"FE",x"FE",
		x"3F",x"3F",x"1F",x"1F",x"0F",x"07",x"00",x"00",x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"00",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"00",x"30",x"7D",x"00",x"C0",x"F0",x"F8",x"3C",x"1C",x"0E",x"8E",
		x"7E",x"7F",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"86",x"06",x"84",x"84",x"C0",x"C0",x"80",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"00",x"31",x"78",x"00",x"C0",x"F0",x"F8",x"3C",x"1C",x"0E",x"8E",
		x"7C",x"7E",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"46",x"06",x"84",x"84",x"C0",x"C0",x"80",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"00",x"33",x"7C",x"00",x"C0",x"F0",x"F8",x"3C",x"1C",x"8E",x"4E",
		x"7C",x"7C",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"46",x"46",x"84",x"84",x"C0",x"C0",x"80",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"02",x"30",x"78",x"00",x"C0",x"F0",x"F8",x"3C",x"9C",x"4E",x"2E",
		x"78",x"78",x"3C",x"3F",x"1F",x"0F",x"03",x"00",x"06",x"26",x"04",x"84",x"C0",x"C0",x"80",x"00",
		x"00",x"01",x"03",x"01",x"01",x"01",x"31",x"39",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",
		x"39",x"3B",x"1F",x"1F",x"0B",x"03",x"01",x"00",x"00",x"00",x"00",x"C0",x"D0",x"F0",x"E0",x"C0",
		x"00",x"01",x"03",x"01",x"01",x"01",x"31",x"39",x"C0",x"C0",x"D0",x"F0",x"E0",x"00",x"00",x"00",
		x"3B",x"3F",x"1F",x"1B",x"0B",x"03",x"01",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"01",x"03",x"01",x"01",x"01",x"31",x"39",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"10",
		x"3D",x"3F",x"1B",x"1B",x"0B",x"03",x"01",x"00",x"30",x"20",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"01",x"03",x"01",x"01",x"01",x"31",x"39",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",
		x"3D",x"3B",x"1B",x"1B",x"0B",x"07",x"01",x"00",x"00",x"00",x"00",x"C0",x"D0",x"F0",x"E0",x"C0",
		x"00",x"01",x"03",x"03",x"03",x"01",x"31",x"39",x"C0",x"C0",x"D0",x"F0",x"E0",x"00",x"00",x"00",
		x"39",x"39",x"1B",x"1B",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"01",x"03",x"0B",x"01",x"01",x"31",x"39",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"10",
		x"39",x"3B",x"1B",x"1F",x"0F",x"03",x"01",x"00",x"30",x"20",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"03",x"07",x"04",x"00",x"31",x"32",x"7C",x"00",x"C0",x"C0",x"E0",x"30",x"9C",x"4E",x"2E",
		x"7C",x"7E",x"0F",x"0F",x"07",x"07",x"03",x"00",x"26",x"46",x"8C",x"80",x"E0",x"E0",x"80",x"00",
		x"00",x"03",x"01",x"01",x"12",x"0C",x"70",x"3C",x"00",x"C0",x"F0",x"F0",x"38",x"7C",x"9E",x"0E",
		x"3F",x"7F",x"3B",x"31",x"01",x"01",x"03",x"00",x"06",x"96",x"E4",x"80",x"C0",x"C0",x"80",x"00",
		x"00",x"00",x"08",x"08",x"04",x"23",x"10",x"0C",x"00",x"C0",x"70",x"78",x"3C",x"1C",x"26",x"42",
		x"07",x"1F",x"3F",x"3C",x"18",x"08",x"00",x"00",x"42",x"22",x"9C",x"84",x"40",x"40",x"80",x"00",
		x"00",x"03",x"0E",x"02",x"01",x"30",x"08",x"04",x"00",x"00",x"10",x"18",x"3C",x"DC",x"08",x"10",
		x"07",x"0F",x"3F",x"3F",x"1E",x"0E",x"03",x"00",x"10",x"08",x"44",x"24",x"10",x"10",x"00",x"00",
		x"00",x"03",x"0F",x"00",x"00",x"06",x"39",x"60",x"00",x"C0",x"00",x"88",x"4C",x"3C",x"0C",x"88",
		x"70",x"79",x"3F",x"1F",x"0F",x"0F",x"03",x"00",x"80",x"04",x"B4",x"CC",x"80",x"80",x"C0",x"00",
		x"00",x"03",x"00",x"00",x"18",x"03",x"34",x"7C",x"00",x"C0",x"E0",x"E0",x"20",x"90",x"4E",x"2E",
		x"7C",x"6E",x"07",x"03",x"03",x"03",x"03",x"00",x"22",x"50",x"90",x"A0",x"E0",x"E0",x"80",x"00",
		x"00",x"00",x"00",x"10",x"0C",x"01",x"30",x"7C",x"00",x"C0",x"F0",x"98",x"8C",x"04",x"86",x"8E",
		x"7F",x"47",x"03",x"01",x"01",x"03",x"03",x"00",x"70",x"00",x"90",x"A0",x"E0",x"D0",x"80",x"00",
		x"00",x"03",x"03",x"00",x"00",x"38",x"30",x"7C",x"00",x"C0",x"C0",x"80",x"80",x"40",x"26",x"1E",
		x"73",x"61",x"00",x"00",x"01",x"07",x"03",x"00",x"02",x"08",x"90",x"A0",x"E0",x"E0",x"80",x"00",
		x"00",x"03",x"03",x"00",x"00",x"00",x"70",x"7F",x"00",x"C0",x"C0",x"C0",x"20",x"10",x"0E",x"0E",
		x"70",x"70",x"30",x"18",x"0F",x"07",x"03",x"00",x"86",x"4E",x"54",x"A0",x"C0",x"C0",x"80",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"00",x"03",x"07",x"04",x"00",x"00",x"00",x"00",x"20",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"00",x"00",x"00",x"A0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"02",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"02",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"03",x"07",x"04",x"E0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"03",x"07",x"04",x"E0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"03",x"07",x"04",x"A0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"05",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"05",x"E0",x"E0",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"05",x"00",x"01",x"00",x"01",x"A0",x"E0",x"E0",x"C0",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"05",x"00",x"01",x"00",x"01",x"E0",x"E0",x"E0",x"40",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"03",x"03",x"07",x"00",x"01",x"00",x"01",x"E0",x"C0",x"C0",x"80",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"02",x"07",x"07",x"07",x"00",x"01",x"00",x"01",x"E0",x"E0",x"E0",x"40",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"10",x"11",x"11",x"01",x"01",
		x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"0F",x"08",x"08",x"25",x"11",x"C9",x"20",x"03",x"3B",
		x"00",x"00",x"00",x"08",x"88",x"88",x"80",x"80",x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"80",
		x"10",x"10",x"A4",x"88",x"93",x"04",x"C0",x"DC",x"00",x"00",x"00",x"38",x"00",x"00",x"00",x"F0",
		x"0F",x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"3B",x"03",x"20",x"C9",x"11",x"25",x"08",x"08",
		x"01",x"02",x"04",x"08",x"00",x"00",x"00",x"00",x"01",x"01",x"11",x"11",x"10",x"00",x"00",x"00",
		x"DC",x"C0",x"04",x"93",x"88",x"A4",x"10",x"10",x"F0",x"00",x"00",x"00",x"38",x"00",x"00",x"00",
		x"80",x"80",x"88",x"88",x"08",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"00",x"00",x"00",x"00",
		x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",x"00",x"01",x"21",x"21",x"20",x"01",x"01",x"11",
		x"00",x"00",x"1C",x"01",x"00",x"00",x"00",x"73",x"90",x"48",x"20",x"80",x"40",x"00",x"00",x"80",
		x"00",x"80",x"80",x"84",x"04",x"04",x"80",x"88",x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",
		x"89",x"12",x"04",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"1C",x"80",x"00",x"00",x"00",x"EE",
		x"77",x"00",x"00",x"00",x"01",x"38",x"00",x"00",x"00",x"00",x"00",x"40",x"80",x"20",x"48",x"91",
		x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",x"11",x"01",x"20",x"20",x"21",x"01",x"01",x"00",
		x"01",x"00",x"00",x"02",x"01",x"04",x"12",x"09",x"CE",x"00",x"00",x"00",x"80",x"38",x"00",x"00",
		x"88",x"80",x"80",x"04",x"84",x"84",x"80",x"00",x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"02",x"01",x"81",x"81",x"01",x"00",x"21",x"21",x"00",x"00",
		x"60",x"00",x"0C",x"00",x"00",x"00",x"00",x"EC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"84",x"84",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"40",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"30",x"00",x"00",x"00",x"00",x"37",
		x"EC",x"00",x"00",x"00",x"00",x"0C",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"02",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"21",x"21",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"37",x"00",x"00",x"00",x"00",x"30",x"00",x"06",
		x"00",x"00",x"84",x"84",x"00",x"80",x"81",x"81",x"80",x"40",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"00",x"00",x"81",x"81",x"01",x"00",x"00",x"00",x"00",x"00",
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
		x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
		x"00",x"00",x"00",x"00",x"00",x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"7C",x"7E",x"64",x"04",x"05",x"60",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0E",x"7E",x"E3",x"63",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"04",x"64",x"7E",x"7B",x"30",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"63",x"E3",x"7E",x"0E",x"07",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4E",x"47",x"02",x"62",x"72",x"30",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0E",x"7E",x"E3",x"E3",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"72",x"62",x"42",x"07",x"4E",x"60",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E3",x"E3",x"7E",x"0E",x"07",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"71",x"73",x"27",x"1F",x"B9",x"B9",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"B9",x"B9",x"1F",x"27",x"73",x"71",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"20",x"71",x"E3",x"C7",x"9F",x"B9",x"B9",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"B9",x"B9",x"9F",x"C7",x"E3",x"71",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FB",x"FA",x"F2",x"F6",x"F4",x"F4",x"E4",x"E8",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"E8",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"3F",x"1F",x"4F",x"07",x"03",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"83",x"F0",x"FE",x"FF",x"FF",x"FF",x"7F",x"7F",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9E",x"9E",x"9E",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",
		x"9C",x"9C",x"88",x"C0",x"40",x"60",x"38",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
		x"02",x"02",x"02",x"03",x"07",x"07",x"03",x"00",x"7F",x"0F",x"01",x"1C",x"1F",x"1F",x"7F",x"7F",
		x"0F",x"0F",x"0F",x"0F",x"1F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"9C",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"86",x"80",x"00",x"C0",x"C0",x"C0",x"80",x"80",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"07",x"07",x"07",x"87",x"87",x"87",x"C3",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C3",x"E3",x"E3",x"E1",x"E1",x"E1",x"F1",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"80",x"80",x"00",x"80",x"F0",x"FE",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"C3",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"FF",
		x"F1",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"78",x"08",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",
		x"9C",x"98",x"90",x"80",x"80",x"80",x"80",x"80",x"03",x"02",x"00",x"00",x"08",x"08",x"1F",x"1F",
		x"80",x"80",x"80",x"80",x"83",x"80",x"89",x"8C",x"0F",x"45",x"01",x"40",x"40",x"50",x"FC",x"78",
		x"03",x"07",x"07",x"0F",x"0F",x"1F",x"0F",x"E1",x"F8",x"F0",x"F0",x"E0",x"E0",x"E0",x"C0",x"C0",
		x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"04",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"BC",x"B8",x"0C",x"EE",x"E8",x"E4",x"E5",x"F7",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"F7",x"FF",x"FF",x"FE",x"FE",x"FC",x"FD",x"F9",
		x"0C",x"1C",x"38",x"98",x"C8",x"60",x"30",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E0",x"80",x"00",x"40",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"17",x"17",
		x"3E",x"20",x"00",x"30",x"7E",x"7E",x"7C",x"00",x"00",x"30",x"00",x"00",x"00",x"08",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3F",x"7F",x"7F",x"0F",x"0F",x"0F",x"8F",x"8F",x"E0",x"F0",x"F0",x"F8",x"F8",x"F8",x"FC",x"FC",
		x"8F",x"8F",x"8F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"04",x"0E",x"0E",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"7F",x"38",x"1C",x"38",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"39",x"7B",x"4F",x"46",x"44",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"1F",x"3F",x"64",x"44",x"64",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"4F",x"4F",x"49",x"49",x"63",x"3E",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"78",x"7C",x"0E",x"07",x"0E",x"7C",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"7F",x"41",x"41",x"41",x"7F",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"03",x"07",x"0E",x"1C",x"38",x"71",x"E3",x"FF",x"FF",x"00",x"00",x"7F",x"FF",x"C0",x"80",
		x"C7",x"CE",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"00",x"00",x"FE",x"FF",x"03",x"01",x"80",x"C0",x"E0",x"70",x"38",x"1C",x"8E",x"C7",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E3",x"73",x"33",x"33",x"33",x"33",x"33",x"33",
		x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CE",x"C7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"E3",x"71",x"38",x"1C",x"0E",x"07",x"03",x"01",x"80",x"C0",x"FF",x"7F",x"00",x"00",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"33",x"33",x"33",x"33",x"33",x"33",x"73",x"E3",
		x"01",x"03",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"C7",x"8E",x"1C",x"38",x"70",x"E0",x"C0",x"80",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",
		x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"F0",x"F0",x"F1",x"F7",x"F7",x"F3",x"FB",x"F8",
		x"9F",x"9F",x"9E",x"98",x"80",x"80",x"80",x"80",x"F0",x"C0",x"00",x"00",x"02",x"0B",x"3B",x"7B",
		x"04",x"3C",x"FC",x"FC",x"F8",x"E0",x"80",x"00",x"80",x"F0",x"C1",x"07",x"1E",x"3C",x"78",x"11",
		x"06",x"0E",x"06",x"00",x"00",x"F8",x"E0",x"C1",x"03",x"38",x"70",x"00",x"00",x"00",x"F8",x"F8",
		x"81",x"83",x"8F",x"9F",x"9F",x"9F",x"9F",x"9F",x"FB",x"FB",x"F8",x"F8",x"F8",x"FC",x"FF",x"FE",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9E",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"03",x"03",
		x"83",x"07",x"0F",x"1F",x"3F",x"7F",x"1F",x"06",x"F0",x"F0",x"E1",x"C3",x"83",x"07",x"0E",x"0F",
		x"00",x"04",x"00",x"00",x"00",x"00",x"81",x"03",x"1F",x"3E",x"3E",x"06",x"3C",x"FC",x"F8",x"F8",
		x"00",x"00",x"80",x"98",x"3F",x"7A",x"F6",x"F6",x"A8",x"28",x"28",x"28",x"68",x"68",x"4C",x"4C",
		x"EC",x"4C",x"08",x"00",x"00",x"00",x"00",x"60",x"CC",x"CC",x"CC",x"CC",x"0C",x"04",x"00",x"00",
		x"4F",x"67",x"73",x"39",x"3C",x"3E",x"3F",x"3F",x"C0",x"F0",x"FC",x"FF",x"7F",x"3F",x"18",x"80",
		x"1F",x"1F",x"2F",x"27",x"27",x"F3",x"31",x"39",x"C0",x"0E",x"0F",x"07",x"43",x"41",x"60",x"70",
		x"E3",x"E3",x"C3",x"C3",x"87",x"87",x"07",x"07",x"80",x"8E",x"8E",x"8E",x"8E",x"8F",x"0F",x"0F",
		x"00",x"08",x"0E",x"0F",x"1F",x"1F",x"1E",x"1E",x"0F",x"00",x"00",x"00",x"00",x"08",x"0E",x"0F",
		x"38",x"38",x"1C",x"1C",x"1E",x"1E",x"1E",x"1F",x"78",x"7C",x"7C",x"3E",x"1F",x"1F",x"00",x"07",
		x"7F",x"7F",x"FF",x"3F",x"0F",x"0F",x"0F",x"BF",x"07",x"83",x"81",x"81",x"C0",x"C0",x"E0",x"E0",
		x"9E",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"01",x"00",x"C0",x"E0",x"F8",x"FC",x"FF",x"FF",
		x"9F",x"9F",x"9F",x"9F",x"87",x"81",x"80",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",
		x"FF",x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"83",x"F0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FF",x"FF",
		x"C1",x"E0",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"8F",x"C7",x"E3",
		x"80",x"80",x"9C",x"9F",x"9F",x"9F",x"9F",x"9F",x"03",x"00",x"00",x"80",x"F0",x"FC",x"FD",x"F9",
		x"9F",x"9F",x"9F",x"9F",x"80",x"80",x"80",x"80",x"FB",x"F8",x"F0",x"F0",x"07",x"07",x"07",x"30",
		x"F0",x"40",x"00",x"04",x"00",x"00",x"C0",x"F8",x"71",x"1C",x"06",x"02",x"00",x"00",x"03",x"01",
		x"FF",x"3F",x"00",x"00",x"FC",x"FC",x"C0",x"00",x"80",x"F8",x"1F",x"00",x"1F",x"00",x"07",x"06",
		x"FF",x"7F",x"7F",x"3F",x"3F",x"3F",x"1F",x"1E",x"10",x"11",x"91",x"91",x"91",x"81",x"81",x"00",
		x"1E",x"8E",x"8E",x"C6",x"C6",x"E6",x"F2",x"F2",x"60",x"70",x"33",x"33",x"33",x"33",x"33",x"33",
		x"00",x"00",x"C0",x"E0",x"C0",x"C0",x"C3",x"47",x"F0",x"70",x"F0",x"1E",x"10",x"03",x"01",x"00",
		x"06",x"06",x"00",x"1C",x"07",x"00",x"00",x"00",x"10",x"3C",x"7E",x"7C",x"18",x"01",x"11",x"00",
		x"00",x"00",x"00",x"04",x"62",x"32",x"88",x"E4",x"B2",x"B2",x"96",x"96",x"D4",x"55",x"55",x"54",
		x"7A",x"1C",x"C2",x"00",x"FF",x"02",x"30",x"01",x"55",x"55",x"38",x"17",x"C0",x"21",x"98",x"48",
		x"60",x"EF",x"DE",x"BC",x"F9",x"73",x"E6",x"CC",x"00",x"00",x"20",x"78",x"E0",x"81",x"1F",x"F8",
		x"9B",x"40",x"80",x"C1",x"07",x"C3",x"58",x"1E",x"80",x"03",x"7F",x"07",x"F0",x"FC",x"0E",x"00",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"00",x"00",x"80",x"C0",x"C0",x"E0",x"F0",x"F0",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"F8",x"FC",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",
		x"1F",x"0F",x"0F",x"07",x"07",x"07",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"01",x"01",x"01",x"00",x"00",x"00",x"80",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",
		x"9F",x"9F",x"9F",x"9F",x"9F",x"8F",x"87",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"81",x"80",x"80",x"80",x"80",x"80",x"98",x"9C",x"FF",x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"03",
		x"C0",x"E0",x"E0",x"F0",x"F0",x"F8",x"F8",x"FC",x"3F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",
		x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"07",x"03",x"03",x"81",x"C1",x"C1",x"E0",
		x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"70",x"70",x"70",x"60",x"00",x"10",x"30",x"70",
		x"F8",x"F8",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"70",x"70",x"70",x"30",x"30",x"10",x"10",x"00",
		x"0F",x"0F",x"1F",x"1F",x"1F",x"03",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"00",x"C0",
		x"01",x"13",x"07",x"07",x"01",x"00",x"00",x"30",x"80",x"80",x"80",x"80",x"00",x"00",x"01",x"00",
		x"FC",x"FC",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"08",x"0C",x"0E",x"00",x"00",
		x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
		x"3E",x"3E",x"7E",x"7E",x"7C",x"7C",x"1C",x"04",x"00",x"00",x"07",x"07",x"07",x"0F",x"0F",x"1F",
		x"00",x"78",x"D8",x"C8",x"C0",x"E0",x"F0",x"F0",x"1F",x"1F",x"00",x"3F",x"5E",x"0C",x"28",x"E0",
		x"0F",x"38",x"60",x"40",x"C0",x"80",x"80",x"80",x"FF",x"00",x"00",x"FF",x"FF",x"7F",x"7F",x"7F",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"3F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"07",x"07",x"03",x"03",x"01",x"01",x"01",x"00",
		x"90",x"90",x"98",x"98",x"9C",x"9C",x"9E",x"9E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"7F",x"7F",x"7F",x"3F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"00",x"00",x"80",x"80",x"80",x"80",x"80",x"FF",x"00",x"00",x"0F",x"0F",x"07",x"03",x"01",
		x"80",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"40",x"60",x"70",x"70",x"70",x"70",x"70",x"70",
		x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"01",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"70",x"70",x"10",x"00",x"00",x"00",x"08",x"02",
		x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"60",x"70",x"70",x"70",x"70",x"70",
		x"00",x"00",x"00",x"04",x"06",x"07",x"07",x"07",x"7E",x"3E",x"0E",x"04",x"00",x"80",x"C4",x"EC",
		x"07",x"07",x"07",x"01",x"00",x"0F",x"0F",x"0F",x"F8",x"F8",x"F8",x"F8",x"70",x"F0",x"F0",x"F0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"60",x"30",x"1C",x"0E",x"07",x"00",x"00",x"20",x"20",x"10",x"10",x"18",x"0C",
		x"03",x"03",x"01",x"00",x"00",x"0F",x"03",x"00",x"8E",x"CF",x"E7",x"F7",x"7F",x"3F",x"FF",x"FF",
		x"00",x"00",x"01",x"02",x"02",x"04",x"0C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"38",x"78",x"F9",x"FF",x"FF",x"FF",x"FF",x"FE",x"00",x"0F",x"FC",x"F0",x"C0",x"80",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"1E",x"3F",x"1F",x"3F",x"7F",x"FF",x"FF",x"C7",x"07",
		x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"04",x"0C",x"08",x"08",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"7F",x"77",x"80",x"E0",x"F8",x"FC",x"00",x"00",x"00",x"80",
		x"33",x"31",x"30",x"10",x"10",x"10",x"00",x"00",x"C0",x"C0",x"E0",x"60",x"30",x"18",x"08",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"42",x"00",x"40",x"00",
		x"00",x"00",x"09",x"00",x"00",x"02",x"00",x"24",x"00",x"04",x"00",x"00",x"20",x"02",x"00",x"88",
		x"00",x"00",x"00",x"40",x"00",x"00",x"02",x"90",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",
		x"00",x"00",x"10",x"82",x"00",x"00",x"50",x"00",x"00",x"20",x"00",x"00",x"88",x"00",x"00",x"02",
		x"00",x"10",x"00",x"01",x"00",x"10",x"02",x"00",x"02",x"00",x"10",x"00",x"40",x"01",x"00",x"00",
		x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"08",x"00",x"40",x"08",x"00",x"01",x"00",
		x"04",x"01",x"40",x"00",x"00",x"08",x"00",x"00",x"10",x"00",x"00",x"08",x"00",x"40",x"00",x"00",
		x"10",x"00",x"04",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"10",x"00",x"00",x"00",x"00",
		x"04",x"00",x"11",x"00",x"08",x"00",x"00",x"40",x"01",x"10",x"00",x"00",x"24",x"00",x"00",x"82",
		x"00",x"00",x"00",x"00",x"00",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",
		x"00",x"10",x"01",x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"12",x"00",x"00",
		x"00",x"08",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"40",x"00",x"00",x"04",x"20",x"00",x"00",
		x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",x"01",x"00",x"00",
		x"00",x"81",x"00",x"10",x"00",x"00",x"80",x"00",x"10",x"00",x"00",x"00",x"90",x"00",x"00",x"10",
		x"01",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"3C",x"62",x"62",x"73",x"00",x"00",x"00",x"60",x"72",x"7E",x"7E",x"7E",
		x"7F",x"73",x"73",x"3F",x"1E",x"00",x"00",x"00",x"78",x"CE",x"EE",x"F2",x"72",x"30",x"00",x"00",
		x"00",x"00",x"00",x"00",x"78",x"C4",x"C4",x"E6",x"00",x"00",x"08",x"34",x"76",x"77",x"7E",x"78",
		x"FE",x"E6",x"E6",x"7E",x"3C",x"00",x"00",x"00",x"78",x"E8",x"F4",x"F2",x"73",x"3E",x"0C",x"00",
		x"00",x"00",x"00",x"00",x"00",x"12",x"23",x"3F",x"00",x"00",x"00",x"00",x"10",x"30",x"32",x"22",
		x"63",x"63",x"73",x"7F",x"7F",x"3F",x"1E",x"00",x"72",x"76",x"36",x"F6",x"F6",x"38",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"02",x"23",x"3F",x"00",x"00",x"00",x"00",x"14",x"34",x"36",x"26",
		x"63",x"63",x"73",x"7F",x"7F",x"3F",x"1E",x"00",x"76",x"72",x"74",x"F6",x"F6",x"3E",x"06",x"00",
		x"00",x"00",x"00",x"00",x"00",x"02",x"23",x"3F",x"00",x"00",x"00",x"00",x"12",x"36",x"36",x"26",
		x"63",x"63",x"73",x"7F",x"7F",x"3F",x"1E",x"00",x"76",x"70",x"30",x"F6",x"F6",x"3E",x"0E",x"0C",
		x"00",x"1E",x"3F",x"7F",x"7F",x"73",x"63",x"63",x"00",x"00",x"38",x"F6",x"F6",x"36",x"76",x"72",
		x"23",x"3F",x"12",x"00",x"00",x"00",x"00",x"00",x"22",x"32",x"30",x"10",x"00",x"00",x"00",x"00",
		x"00",x"1E",x"3F",x"7F",x"7F",x"73",x"63",x"63",x"00",x"06",x"3E",x"F6",x"F6",x"74",x"72",x"76",
		x"23",x"3F",x"02",x"00",x"00",x"00",x"00",x"00",x"26",x"36",x"34",x"14",x"00",x"00",x"00",x"00",
		x"00",x"1E",x"3F",x"7F",x"7F",x"73",x"63",x"63",x"0C",x"0E",x"3E",x"F6",x"F6",x"30",x"70",x"76",
		x"23",x"3F",x"02",x"00",x"00",x"00",x"00",x"00",x"26",x"36",x"36",x"12",x"00",x"00",x"00",x"00",
		x"00",x"07",x"0F",x"1C",x"3B",x"37",x"34",x"34",x"00",x"F0",x"F8",x"1C",x"6E",x"F6",x"96",x"96",
		x"34",x"37",x"3F",x"1C",x"0F",x"07",x"00",x"00",x"96",x"F6",x"FE",x"1C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"1C",x"34",x"00",x"00",x"00",x"00",x"F0",x"F8",x"9C",x"96",
		x"34",x"37",x"37",x"18",x"0F",x"07",x"00",x"00",x"96",x"F6",x"F6",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"3F",x"3F",x"00",x"00",x"00",x"00",x"60",x"F0",x"F0",x"F0",
		x"3F",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"07",x"04",x"04",x"00",x"00",x"00",x"00",x"F0",x"F8",x"98",x"90",
		x"04",x"27",x"30",x"18",x"0F",x"07",x"00",x"00",x"90",x"F0",x"00",x"00",x"F0",x"F0",x"00",x"00",
		x"00",x"07",x"0F",x"1C",x"3C",x"34",x"34",x"34",x"00",x"F0",x"F8",x"1C",x"1E",x"96",x"96",x"96",
		x"34",x"37",x"3F",x"1C",x"0F",x"07",x"00",x"00",x"96",x"F6",x"FE",x"1C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"1C",x"34",x"00",x"00",x"00",x"00",x"F0",x"F8",x"9C",x"96",
		x"34",x"37",x"37",x"18",x"0F",x"07",x"00",x"00",x"96",x"F6",x"F6",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"04",x"3F",x"3F",x"00",x"00",x"00",x"00",x"10",x"90",x"F0",x"F0",
		x"3F",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"07",x"04",x"04",x"00",x"00",x"00",x"00",x"F0",x"F8",x"98",x"90",
		x"04",x"27",x"30",x"18",x"0F",x"07",x"00",x"00",x"90",x"F0",x"00",x"00",x"F0",x"F0",x"00",x"00",
		x"00",x"07",x"0F",x"1C",x"3A",x"36",x"34",x"34",x"00",x"F0",x"F8",x"1C",x"6E",x"F6",x"96",x"96",
		x"34",x"37",x"3B",x"1C",x"0F",x"07",x"00",x"00",x"96",x"B6",x"2E",x"1C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"0F",x"1C",x"34",x"00",x"00",x"00",x"00",x"F0",x"F8",x"9C",x"96",
		x"34",x"37",x"33",x"18",x"0F",x"07",x"00",x"00",x"96",x"B6",x"26",x"0C",x"F8",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"02",x"06",x"3F",x"3F",x"00",x"00",x"00",x"00",x"60",x"F0",x"F0",x"F0",
		x"3F",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"F0",x"B0",x"20",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"07",x"07",x"04",x"04",x"00",x"00",x"00",x"00",x"F0",x"F8",x"98",x"90",
		x"04",x"27",x"30",x"18",x"0F",x"07",x"00",x"00",x"90",x"B0",x"00",x"00",x"F0",x"F0",x"00",x"00",
		x"00",x"00",x"00",x"E0",x"71",x"79",x"F8",x"E0",x"00",x"00",x"00",x"80",x"C0",x"F8",x"FC",x"7C",
		x"F8",x"E0",x"F8",x"79",x"71",x"E0",x"00",x"00",x"F8",x"7C",x"FC",x"F8",x"C0",x"80",x"00",x"00",
		x"00",x"00",x"00",x"E2",x"77",x"79",x"F8",x"C8",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"7C",
		x"F0",x"C8",x"F8",x"79",x"77",x"E2",x"00",x"00",x"F8",x"7C",x"FC",x"F8",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1C",x"0E",x"0F",x"1F",x"3E",x"00",x"00",x"20",x"60",x"EC",x"7C",x"3C",x"18",
		x"3F",x"3E",x"1F",x"0F",x"0E",x"1C",x"00",x"00",x"38",x"18",x"3C",x"7C",x"EC",x"60",x"20",x"00",
		x"00",x"00",x"00",x"38",x"60",x"F8",x"FE",x"F0",x"00",x"00",x"C0",x"CC",x"5C",x"FC",x"78",x"F0",
		x"F2",x"7C",x"79",x"E1",x"00",x"00",x"00",x"00",x"F8",x"FC",x"FC",x"C8",x"C0",x"80",x"00",x"00",
		x"00",x"00",x"00",x"38",x"60",x"F8",x"FE",x"F0",x"00",x"00",x"00",x"18",x"78",x"F8",x"7C",x"FC",
		x"F2",x"7C",x"79",x"E0",x"00",x"00",x"00",x"00",x"FC",x"EC",x"E0",x"60",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"38",x"60",x"F8",x"FE",x"F0",x"00",x"00",x"40",x"CC",x"5C",x"FC",x"78",x"F0",
		x"F2",x"7C",x"78",x"E0",x"00",x"00",x"00",x"00",x"F8",x"7C",x"18",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"38",x"60",x"F8",x"FE",x"F0",x"00",x"00",x"00",x"D8",x"78",x"F8",x"7C",x"EC",
		x"F2",x"7C",x"78",x"F0",x"00",x"00",x"00",x"00",x"E4",x"E0",x"60",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F1",x"79",x"7C",x"F2",x"00",x"00",x"80",x"C0",x"C8",x"FC",x"FC",x"F8",
		x"F0",x"FE",x"F8",x"60",x"38",x"00",x"00",x"00",x"F0",x"78",x"FC",x"5C",x"CC",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"79",x"7C",x"F2",x"00",x"00",x"00",x"00",x"60",x"E0",x"EC",x"FC",
		x"F0",x"FE",x"F8",x"60",x"38",x"00",x"00",x"00",x"FC",x"7C",x"F8",x"78",x"18",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"78",x"7C",x"F2",x"00",x"00",x"00",x"C0",x"00",x"18",x"7C",x"F8",
		x"F0",x"FE",x"F8",x"60",x"38",x"00",x"00",x"00",x"F0",x"78",x"FC",x"5C",x"CC",x"40",x"00",x"00",
		x"00",x"00",x"00",x"00",x"F0",x"78",x"7C",x"F2",x"00",x"00",x"00",x"00",x"60",x"60",x"E0",x"E4",
		x"F0",x"FE",x"F8",x"60",x"38",x"00",x"00",x"00",x"EC",x"7C",x"FC",x"78",x"D8",x"00",x"00",x"00",
		x"00",x"00",x"00",x"71",x"3B",x"3C",x"7C",x"E4",x"00",x"00",x"00",x"00",x"80",x"FC",x"7E",x"3E",
		x"F8",x"E4",x"7C",x"3C",x"3B",x"71",x"00",x"00",x"7C",x"3E",x"7E",x"FC",x"80",x"00",x"00",x"00",
		x"00",x"00",x"00",x"38",x"1D",x"1E",x"3E",x"7C",x"00",x"00",x"00",x"80",x"C0",x"7C",x"3E",x"1E",
		x"7C",x"7C",x"3E",x"1E",x"1D",x"38",x"00",x"00",x"3C",x"1E",x"3E",x"7C",x"C0",x"80",x"00",x"00",
		x"00",x"00",x"38",x"48",x"FB",x"FE",x"F8",x"F8",x"40",x"E0",x"C0",x"48",x"7C",x"7E",x"7E",x"7E",
		x"7E",x"3C",x"39",x"71",x"00",x"00",x"00",x"00",x"7C",x"FC",x"9C",x"C0",x"C0",x"00",x"00",x"00",
		x"00",x"00",x"01",x"03",x"E3",x"7A",x"79",x"E0",x"00",x"00",x"0C",x"9E",x"BE",x"FC",x"F8",x"FC",
		x"F8",x"F0",x"FC",x"FC",x"7D",x"3C",x"38",x"70",x"FC",x"FC",x"FC",x"F8",x"C8",x"E0",x"60",x"00",
		x"00",x"00",x"00",x"00",x"01",x"71",x"3C",x"3E",x"00",x"00",x"00",x"C0",x"C0",x"9C",x"FC",x"7C",
		x"79",x"F8",x"FE",x"FB",x"48",x"38",x"00",x"00",x"7E",x"7E",x"7E",x"7C",x"48",x"C0",x"E0",x"40",
		x"70",x"38",x"3C",x"73",x"FC",x"FC",x"F0",x"F8",x"00",x"60",x"E0",x"C0",x"F8",x"FC",x"FC",x"FC",
		x"E0",x"79",x"7A",x"E3",x"03",x"01",x"00",x"00",x"FC",x"F8",x"FC",x"BE",x"9E",x"0C",x"00",x"00",
		x"43",x"47",x"41",x"64",x"66",x"67",x"67",x"77",x"0F",x"FC",x"F0",x"40",x"00",x"80",x"80",x"80",
		x"77",x"63",x"63",x"42",x"06",x"07",x"04",x"04",x"80",x"80",x"00",x"00",x"00",x"00",x"C0",x"20",
		x"04",x"27",x"27",x"37",x"37",x"3F",x"3F",x"3F",x"00",x"E0",x"FE",x"F0",x"80",x"80",x"80",x"80",
		x"3F",x"3B",x"33",x"00",x"06",x"07",x"04",x"04",x"80",x"80",x"00",x"00",x"00",x"00",x"C0",x"20",
		x"00",x"17",x"19",x"1C",x"1F",x"1F",x"1F",x"1F",x"00",x"80",x"C0",x"70",x"58",x"00",x"80",x"80",
		x"1F",x"1F",x"1F",x"12",x"06",x"07",x"04",x"04",x"80",x"80",x"00",x"00",x"00",x"00",x"C0",x"20",
		x"10",x"20",x"20",x"40",x"60",x"18",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2F",
		x"04",x"0F",x"7F",x"40",x"20",x"20",x"10",x"00",x"FC",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"06",x"08",x"10",x"10",x"18",x"08",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2E",
		x"04",x"0F",x"1F",x"10",x"10",x"08",x"06",x"00",x"F8",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
		x"07",x"18",x"10",x"10",x"18",x"08",x"0C",x"0C",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"2C",
		x"04",x"0F",x"1F",x"10",x"10",x"18",x"07",x"00",x"F0",x"C0",x"80",x"00",x"00",x"00",x"80",x"00",
		x"40",x"47",x"60",x"67",x"77",x"77",x"63",x"43",x"00",x"FE",x"F8",x"60",x"80",x"80",x"80",x"80",
		x"67",x"7B",x"7A",x"67",x"07",x"04",x"04",x"00",x"80",x"00",x"00",x"00",x"80",x"C0",x"20",x"00",
		x"00",x"04",x"04",x"07",x"67",x"7A",x"7B",x"67",x"00",x"20",x"C0",x"80",x"00",x"00",x"00",x"80",
		x"43",x"63",x"77",x"77",x"67",x"60",x"47",x"40",x"80",x"80",x"80",x"80",x"60",x"F8",x"FE",x"00",
		x"00",x"00",x"00",x"E0",x"71",x"79",x"F8",x"E0",x"00",x"00",x"40",x"E0",x"80",x"98",x"FC",x"7C",
		x"F0",x"E0",x"F8",x"79",x"71",x"E0",x"00",x"00",x"F8",x"7C",x"FC",x"98",x"80",x"E0",x"40",x"00",
		x"00",x"00",x"01",x"71",x"39",x"3D",x"7F",x"F8",x"00",x"00",x"80",x"80",x"8C",x"FC",x"FC",x"F8",
		x"F8",x"E0",x"F0",x"60",x"78",x"F0",x"00",x"00",x"78",x"F8",x"7C",x"DC",x"CC",x"C0",x"C0",x"00",
		x"00",x"00",x"00",x"E2",x"77",x"79",x"F8",x"C8",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"7C",
		x"F0",x"C8",x"F8",x"79",x"77",x"E2",x"00",x"00",x"F8",x"7C",x"FC",x"F8",x"00",x"00",x"00",x"00",
		x"00",x"00",x"0E",x"1E",x"3E",x"7C",x"7D",x"7B",x"00",x"00",x"00",x"00",x"40",x"C0",x"C0",x"80",
		x"7B",x"7D",x"7D",x"3E",x"1E",x"0F",x"03",x"00",x"80",x"C0",x"C0",x"E0",x"F0",x"90",x"E0",x"00",
		x"00",x"00",x"0E",x"1E",x"3E",x"7C",x"7D",x"7B",x"00",x"00",x"00",x"00",x"43",x"C1",x"C1",x"80",
		x"7B",x"7D",x"7D",x"3E",x"1E",x"0F",x"03",x"00",x"80",x"C1",x"C1",x"E3",x"F7",x"91",x"E0",x"00",
		x"00",x"00",x"0E",x"1F",x"3F",x"7F",x"7F",x"7F",x"00",x"00",x"00",x"80",x"C0",x"C0",x"E0",x"E0",
		x"7F",x"7F",x"7F",x"3F",x"1F",x"0F",x"03",x"00",x"E0",x"E0",x"E0",x"F0",x"F0",x"F0",x"E0",x"00",
		x"00",x"00",x"1C",x"3C",x"58",x"09",x"9B",x"F7",x"00",x"00",x"00",x"00",x"84",x"82",x"88",x"04",
		x"F7",x"FB",x"FB",x"7D",x"3D",x"1F",x"07",x"00",x"0A",x"94",x"84",x"C2",x"EC",x"24",x"CA",x"00",
		x"C0",x"C0",x"30",x"30",x"37",x"2E",x"0E",x"1D",x"00",x"02",x"04",x"0A",x"04",x"82",x"C6",x"CE",
		x"0D",x"0B",x"02",x"05",x"02",x"00",x"00",x"00",x"8E",x"7E",x"FE",x"3C",x"1C",x"1C",x"38",x"00",
		x"C0",x"80",x"70",x"68",x"1E",x"1D",x"1B",x"1B",x"00",x"00",x"02",x"04",x"02",x"84",x"A6",x"8E",
		x"07",x"07",x"06",x"05",x"02",x"00",x"00",x"00",x"0E",x"7E",x"FE",x"3C",x"1C",x"1C",x"38",x"00",
		x"40",x"C0",x"60",x"58",x"1C",x"3B",x"1B",x"17",x"00",x"00",x"00",x"02",x"04",x"82",x"66",x"4E",
		x"06",x"0D",x"04",x"04",x"02",x"00",x"00",x"00",x"BE",x"7E",x"FE",x"1C",x"1C",x"1C",x"18",x"00",
		x"C0",x"C0",x"50",x"5C",x"3A",x"37",x"16",x"0E",x"00",x"00",x"00",x"00",x"02",x"00",x"E6",x"CE",
		x"0D",x"0D",x"02",x"01",x"02",x"00",x"00",x"00",x"8E",x"7E",x"FE",x"3C",x"1C",x"1C",x"38",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"3B",x"00",x"00",x"40",x"70",x"78",x"78",x"7C",x"7C",
		x"3A",x"38",x"18",x"1E",x"0E",x"02",x"00",x"00",x"7C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"07",x"0F",x"1F",x"3F",x"3F",x"3E",x"00",x"00",x"E0",x"F0",x"D8",x"DC",x"8C",x"0C",
		x"3F",x"3F",x"3E",x"1F",x"0F",x"07",x"00",x"00",x"8C",x"8C",x"1C",x"D8",x"F0",x"E0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"E2",x"77",x"79",x"F8",x"C8",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"7C",
		x"F0",x"C8",x"F8",x"79",x"77",x"E2",x"00",x"00",x"F8",x"7C",x"FC",x"F8",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1D",x"0F",x"1F",x"3F",x"3F",x"00",x"00",x"C0",x"C0",x"80",x"F8",x"FC",x"7C",
		x"3F",x"3F",x"3F",x"1F",x"0F",x"1D",x"00",x"00",x"78",x"7C",x"FC",x"F8",x"80",x"C0",x"C0",x"00",
		x"00",x"00",x"00",x"01",x"00",x"41",x"63",x"43",x"00",x"00",x"00",x"C0",x"FC",x"FE",x"F4",x"E0",
		x"03",x"63",x"43",x"41",x"00",x"01",x"00",x"00",x"E0",x"E0",x"F4",x"FE",x"FC",x"C0",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"0F",x"00",x"00",x"00",x"40",x"E0",x"E0",x"F0",x"E0",
		x"03",x"0F",x"0F",x"07",x"01",x"00",x"00",x"00",x"F0",x"E0",x"E0",x"F0",x"E0",x"40",x"00",x"00",
		x"00",x"00",x"00",x"70",x"3B",x"3E",x"7C",x"EC",x"00",x"00",x"00",x"80",x"D8",x"FC",x"7E",x"3E",
		x"F8",x"EC",x"7C",x"3E",x"3B",x"70",x"00",x"00",x"7E",x"3E",x"7E",x"FC",x"D8",x"80",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"1F",x"3F",x"3F",x"7F",x"7F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"7F",x"7F",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"04",x"0F",x"1F",x"17",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"41",
		x"17",x"17",x"1F",x"0F",x"07",x"09",x"11",x"01",x"51",x"59",x"22",x"3C",x"BC",x"B8",x"80",x"80",
		x"00",x"00",x"00",x"00",x"04",x"27",x"17",x"17",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"41",
		x"1F",x"1F",x"1F",x"1F",x"27",x"01",x"01",x"00",x"51",x"59",x"22",x"3C",x"BC",x"B8",x"80",x"00",
		x"00",x"00",x"00",x"00",x"04",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"41",
		x"7F",x"1F",x"1F",x"0F",x"07",x"00",x"00",x"00",x"51",x"59",x"22",x"3C",x"BC",x"38",x"00",x"00",
		x"00",x"00",x"00",x"40",x"24",x"1F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"1C",x"22",x"41",
		x"1F",x"17",x"17",x"27",x"07",x"01",x"00",x"00",x"51",x"59",x"62",x"3C",x"BC",x"B8",x"00",x"00",
		x"00",x"00",x"02",x"02",x"03",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"E0",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",
		x"00",x"00",x"03",x"02",x"02",x"02",x"03",x"00",x"00",x"00",x"E0",x"20",x"20",x"20",x"E0",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"02",x"02",x"02",x"00",x"00",x"00",x"00",x"E0",x"20",x"20",x"20",
		x"03",x"08",x"0C",x"06",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"20",
		x"02",x"0A",x"0F",x"06",x"00",x"00",x"00",x"00",x"20",x"20",x"E0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"0A",x"0E",x"06",x"03",x"00",x"00",x"00",x"E0",x"20",x"20",x"20",x"E0",x"00",x"00",x"00",
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"0F",x"06",x"02",x"02",x"01",x"00",x"00",x"00",x"E0",x"20",x"20",x"20",x"C0",x"00",
		x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"03",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"20",x"00",x"00",
		x"00",x"00",x"02",x"02",x"03",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"E0",x"00",x"00",x"00",
		x"00",x"08",x"0C",x"06",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",
		x"00",x"00",x"00",x"1F",x"3F",x"3F",x"7F",x"7F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"7C",x"7E",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"1F",x"3F",x"3F",x"7F",x"7E",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"78",x"7C",x"3E",x"3F",x"1F",x"0F",x"03",x"00",x"78",x"F8",x"F8",x"F8",x"F8",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"1F",x"3F",x"3F",x"7F",x"78",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"70",
		x"78",x"78",x"3C",x"3F",x"1F",x"0F",x"03",x"00",x"78",x"78",x"78",x"F8",x"F8",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"1F",x"3F",x"3F",x"7C",x"70",x"00",x"00",x"00",x"00",x"C0",x"E0",x"70",x"30",
		x"70",x"70",x"38",x"3C",x"1F",x"0F",x"03",x"00",x"38",x"38",x"78",x"78",x"F8",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"0A",x"1E",x"1E",x"3A",x"3A",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",
		x"3A",x"3A",x"1E",x"1E",x"0A",x"02",x"00",x"00",x"C0",x"C0",x"C0",x"E0",x"F0",x"F0",x"E0",x"C0",
		x"00",x"00",x"00",x"0E",x"1E",x"1A",x"3A",x"3A",x"00",x"20",x"30",x"30",x"20",x"C0",x"C0",x"C0",
		x"3A",x"3E",x"1E",x"1A",x"0A",x"02",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"00",x"04",x"0E",x"1A",x"1A",x"3A",x"3A",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",
		x"3E",x"3E",x"1A",x"1A",x"0A",x"02",x"00",x"00",x"F0",x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"00",x"04",x"0A",x"1A",x"1A",x"3A",x"3E",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",
		x"3E",x"3A",x"1A",x"1A",x"0A",x"06",x"00",x"00",x"C0",x"C0",x"C0",x"E0",x"F0",x"F0",x"E0",x"C0",
		x"00",x"00",x"00",x"08",x"18",x"1A",x"3E",x"3E",x"00",x"20",x"30",x"30",x"20",x"C0",x"C0",x"C0",
		x"3A",x"3A",x"1A",x"1A",x"0E",x"06",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"00",x"00",x"00",x"1A",x"1E",x"3E",x"3A",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",
		x"3A",x"3A",x"1A",x"1E",x"0E",x"02",x"00",x"00",x"F0",x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"04",x"07",x"0F",x"0F",x"7E",x"78",x"00",x"00",x"20",x"00",x"C0",x"EC",x"70",x"10",
		x"78",x"7C",x"3E",x"07",x"07",x"07",x"03",x"00",x"18",x"38",x"7C",x"F0",x"C0",x"C0",x"C0",x"00",
		x"00",x"02",x"01",x"01",x"21",x"33",x"7F",x"1F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"90",x"08",
		x"1E",x"3F",x"37",x"23",x"01",x"01",x"03",x"00",x"08",x"08",x"98",x"F8",x"F0",x"F0",x"C0",x"00",
		x"00",x"00",x"00",x"10",x"38",x"3C",x"1F",x"0F",x"00",x"80",x"40",x"40",x"C0",x"F8",x"E4",x"82",
		x"0F",x"0F",x"1F",x"38",x"10",x"00",x"00",x"00",x"82",x"C4",x"E0",x"F8",x"78",x"70",x"C0",x"00",
		x"00",x"00",x"00",x"1C",x"3E",x"3F",x"0F",x"07",x"00",x"00",x"10",x"10",x"20",x"24",x"F8",x"E0",
		x"07",x"07",x"0F",x"3E",x"1C",x"0C",x"02",x"00",x"E0",x"F0",x"F8",x"38",x"18",x"10",x"00",x"00",
		x"00",x"00",x"00",x"0F",x"1F",x"3F",x"79",x"70",x"00",x"40",x"80",x"08",x"88",x"C0",x"F0",x"F0",
		x"60",x"70",x"39",x"1F",x"0F",x"0F",x"03",x"00",x"F8",x"F8",x"F8",x"88",x"00",x"00",x"80",x"00",
		x"00",x"02",x"01",x"03",x"27",x"3F",x"78",x"78",x"00",x"00",x"00",x"00",x"C0",x"E0",x"70",x"30",
		x"78",x"7C",x"2E",x"07",x"07",x"07",x"03",x"00",x"3C",x"22",x"64",x"C0",x"C0",x"C0",x"C0",x"00",
		x"00",x"01",x"01",x"03",x"33",x"3E",x"7F",x"7F",x"00",x"00",x"00",x"60",x"10",x"08",x"08",x"00",
		x"7F",x"67",x"23",x"21",x"13",x"0F",x"03",x"00",x"8E",x"F8",x"E0",x"C0",x"C0",x"E0",x"C0",x"00",
		x"00",x"02",x"02",x"03",x"07",x"07",x"7F",x"7F",x"00",x"00",x"30",x"08",x"04",x"84",x"C0",x"E0",
		x"63",x"41",x"20",x"30",x"19",x"0F",x"03",x"00",x"FC",x"F2",x"E0",x"C0",x"C0",x"C0",x"C0",x"00",
		x"00",x"02",x"02",x"03",x"07",x"0F",x"0F",x"7F",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",
		x"60",x"60",x"20",x"10",x"08",x"07",x"03",x"00",x"F8",x"78",x"64",x"C0",x"80",x"80",x"C0",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"00",x"03",x"07",x"04",x"00",x"00",x"00",x"00",x"20",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"00",x"00",x"00",x"A0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"02",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"02",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"03",x"07",x"04",x"E0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"00",x"03",x"07",x"04",x"E0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"05",x"00",x"03",x"07",x"04",x"A0",x"E0",x"E0",x"C0",x"20",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"05",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"40",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"05",x"E0",x"E0",x"E0",x"C0",x"A0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",
		x"03",x"07",x"07",x"07",x"03",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"05",x"00",x"01",x"00",x"01",x"A0",x"E0",x"E0",x"C0",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"03",x"07",x"07",x"05",x"00",x"01",x"00",x"01",x"E0",x"E0",x"E0",x"40",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"03",x"03",x"07",x"00",x"01",x"00",x"01",x"E0",x"C0",x"C0",x"80",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"02",x"07",x"07",x"07",x"00",x"01",x"00",x"01",x"E0",x"E0",x"E0",x"40",x"A0",x"40",x"A0",x"40",
		x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"10",x"11",x"11",x"01",x"01",
		x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"0F",x"08",x"08",x"25",x"11",x"C9",x"20",x"03",x"3B",
		x"00",x"00",x"00",x"08",x"88",x"88",x"80",x"80",x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"80",
		x"10",x"10",x"A4",x"88",x"93",x"04",x"C0",x"DC",x"00",x"00",x"00",x"38",x"00",x"00",x"00",x"F0",
		x"0F",x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"3B",x"03",x"20",x"C9",x"11",x"25",x"08",x"08",
		x"01",x"02",x"04",x"08",x"00",x"00",x"00",x"00",x"01",x"01",x"11",x"11",x"10",x"00",x"00",x"00",
		x"DC",x"C0",x"04",x"93",x"88",x"A4",x"10",x"10",x"F0",x"00",x"00",x"00",x"38",x"00",x"00",x"00",
		x"80",x"80",x"88",x"88",x"08",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"00",x"00",x"00",x"00",
		x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",x"00",x"01",x"21",x"21",x"20",x"01",x"01",x"11",
		x"00",x"00",x"1C",x"01",x"00",x"00",x"00",x"73",x"90",x"48",x"20",x"80",x"40",x"00",x"00",x"80",
		x"00",x"80",x"80",x"84",x"04",x"04",x"80",x"88",x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",
		x"89",x"12",x"04",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"1C",x"80",x"00",x"00",x"00",x"EE",
		x"77",x"00",x"00",x"00",x"01",x"38",x"00",x"00",x"00",x"00",x"00",x"40",x"80",x"20",x"48",x"91",
		x"00",x"00",x"04",x"08",x"10",x"20",x"00",x"00",x"11",x"01",x"20",x"20",x"21",x"01",x"01",x"00",
		x"01",x"00",x"00",x"02",x"01",x"04",x"12",x"09",x"CE",x"00",x"00",x"00",x"80",x"38",x"00",x"00",
		x"88",x"80",x"80",x"04",x"84",x"84",x"80",x"00",x"00",x"00",x"20",x"10",x"08",x"04",x"00",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"02",x"01",x"81",x"81",x"01",x"00",x"21",x"21",x"00",x"00",
		x"60",x"00",x"0C",x"00",x"00",x"00",x"00",x"EC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"84",x"84",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"40",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"30",x"00",x"00",x"00",x"00",x"37",
		x"EC",x"00",x"00",x"00",x"00",x"0C",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"02",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"21",x"21",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"37",x"00",x"00",x"00",x"00",x"30",x"00",x"06",
		x"00",x"00",x"84",x"84",x"00",x"80",x"81",x"81",x"80",x"40",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"40",x"20",x"10",x"00",x"00",x"00",x"00",x"81",x"81",x"01",x"00",x"00",x"00",x"00",x"00",
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"04",x"08",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
		x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
		x"00",x"00",x"00",x"00",x"00",x"80",x"81",x"81",x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"1F",x"3F",x"3E",x"1F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"40",x"E7",x"CE",x"9E",x"1F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"3F",x"1F",x"01",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0F",x"1F",x"9E",x"CE",x"E7",x"40",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3F",x"1F",x"0E",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"40",x"47",x"EE",x"9E",x"1F",x"0B",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"1F",x"3F",x"18",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0B",x"1F",x"9E",x"EE",x"47",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"F0",x"78",x"38",x"08",x"04",x"0E",x"0A",x"00",x"00",x"01",x"03",x"06",x"04",x"47",x"57",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"01",x"8F",x"1F",x"6F",x"CF",x"8D",x"87",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0E",x"04",x"08",x"38",x"78",x"F0",x"F0",x"A0",x"47",x"04",x"06",x"03",x"01",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"8D",x"CF",x"6F",x"1F",x"8F",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"0E",x"00",x"00",x"00",x"00",x"C0",x"00",x"80",x"00",
		x"0C",x"0C",x"0C",x"08",x"08",x"04",x"0E",x"0A",x"00",x"00",x"00",x"06",x"07",x"07",x"43",x"51",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"09",x"1F",x"3F",x"EF",x"CF",x"8D",x"87",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"0E",x"04",x"08",x"08",x"0C",x"0C",x"0C",x"0E",x"43",x"07",x"07",x"06",x"00",x"00",x"00",x"00",
		x"07",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",
		x"8D",x"CF",x"EF",x"3F",x"1F",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F8",x"F9",x"F1",x"F1",x"F3",x"F3",x"E3",x"E7",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"E7",x"EF",x"EF",x"EF",x"EF",x"EF",x"E7",x"F7",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"FC",x"C0",x"C0",x"C0",x"C0",x"00",x"40",x"00",x"00",
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F7",x"F7",x"F3",x"F8",x"FE",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"4F",x"27",x"33",x"18",x"07",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",
		x"FC",x"FC",x"FC",x"FC",x"38",x"88",x"E0",x"F8",x"00",x"00",x"00",x"1C",x"1F",x"1F",x"7F",x"7F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",
		x"1F",x"1F",x"1F",x"1F",x"1F",x"07",x"01",x"1C",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
		x"06",x"00",x"00",x"00",x"3C",x"3F",x"7F",x"7F",x"70",x"30",x"10",x"10",x"00",x"80",x"F0",x"F0",
		x"0F",x"0F",x"0F",x"07",x"07",x"07",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"03",x"03",x"03",x"01",x"01",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"7F",x"7F",x"7F",x"3F",x"87",x"F0",x"FE",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"10",x"C0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"F8",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",
		x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"03",x"C3",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",
		x"5F",x"5F",x"5E",x"5E",x"5A",x"5B",x"59",x"5C",x"F8",x"F9",x"FB",x"FB",x"7B",x"38",x"3F",x"9F",
		x"5C",x"5E",x"58",x"5E",x"5F",x"40",x"58",x"5C",x"8F",x"45",x"01",x"00",x"00",x"00",x"00",x"00",
		x"FC",x"F8",x"F8",x"F0",x"F0",x"60",x"00",x"E0",x"07",x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"3E",
		x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"04",x"20",x"80",x"40",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"80",x"80",x"00",x"E0",x"E0",x"E4",x"E5",x"F7",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F7",x"FF",x"FF",x"FE",x"FE",x"FC",x"FC",x"F8",
		x"0E",x"1E",x"3E",x"9E",x"CF",x"6F",x"3F",x"B8",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",
		x"E0",x"80",x"1E",x"3F",x"7F",x"7F",x"7F",x"FF",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",
		x"C1",x"C0",x"00",x"C0",x"81",x"81",x"83",x"00",x"00",x"3F",x"00",x"00",x"00",x"F0",x"F0",x"30",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3F",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"0F",x"1F",x"1F",x"3F",x"3F",x"1F",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"7F",x"7F",x"38",x"1C",x"38",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"39",x"7B",x"4F",x"46",x"44",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"41",x"49",x"49",x"49",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"1F",x"3F",x"64",x"44",x"64",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"4F",x"4F",x"49",x"49",x"63",x"3E",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"78",x"7C",x"0E",x"07",x"0E",x"7C",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"3E",x"7F",x"41",x"41",x"41",x"7F",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7E",x"FC",x"FF",x"FF",x"FF",x"FF",x"80",x"00",x"00",x"00",
		x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"01",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"7E",x"3F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FC",x"7E",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"80",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"1F",
		x"00",x"00",x"00",x"01",x"FF",x"FF",x"FF",x"FF",x"3F",x"7E",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F7",x"F7",x"F6",x"F0",x"F0",x"F0",x"F8",x"F9",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FC",x"FE",x"FE",x"F8",x"F8",x"F8",x"F8",x"F8",
		x"F8",x"C0",x"00",x"00",x"04",x"1C",x"7C",x"FE",x"03",x"08",x"3E",x"F8",x"E1",x"43",x"07",x"0E",
		x"78",x"10",x"00",x"00",x"00",x"04",x"1F",x"3E",x"00",x"38",x"7F",x"00",x"00",x"00",x"00",x"07",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F8",x"F8",x"FB",x"FB",x"F9",x"FC",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FE",x"FE",x"F8",x"F8",x"F8",
		x"7C",x"F8",x"F0",x"E0",x"C0",x"00",x"00",x"C1",x"0F",x"0F",x"1E",x"3C",x"7C",x"F8",x"F0",x"F0",
		x"F1",x"FC",x"E0",x"00",x"00",x"3F",x"7E",x"FC",x"E0",x"41",x"01",x"01",x"03",x"03",x"07",x"07",
		x"00",x"00",x"00",x"60",x"C0",x"85",x"09",x"09",x"54",x"54",x"54",x"14",x"94",x"94",x"B2",x"B2",
		x"13",x"33",x"07",x"01",x"00",x"00",x"00",x"90",x"32",x"32",x"32",x"32",x"32",x"02",x"00",x"00",
		x"7F",x"7F",x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"C0",
		x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"3F",x"3F",x"C1",x"01",x"70",x"78",x"3C",x"3E",x"1F",x"0F",
		x"1C",x"1C",x"3C",x"3C",x"78",x"78",x"38",x"88",x"40",x"70",x"70",x"70",x"70",x"70",x"F0",x"F0",
		x"E0",x"F0",x"F0",x"F0",x"E0",x"E0",x"E1",x"E1",x"30",x"00",x"00",x"80",x"E0",x"F0",x"F0",x"F0",
		x"3F",x"3F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"07",x"03",x"03",x"41",x"60",x"60",x"00",x"FF",
		x"7F",x"7F",x"FF",x"3F",x"0F",x"0F",x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"FC",x"F8",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"F8",x"FB",x"F3",x"F7",x"F0",x"F0",x"F0",x"F7",
		x"F0",x"C0",x"80",x"18",x"7F",x"FF",x"3F",x"07",x"7F",x"1F",x"07",x"02",x"00",x"C1",x"E0",x"F6",
		x"00",x"C0",x"FE",x"FC",x"00",x"00",x"3C",x"FC",x"77",x"07",x"60",x"3F",x"80",x"0F",x"08",x"01",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"CC",x"CE",x"CE",x"CE",x"CE",x"86",x"80",x"00",
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"80",x"8C",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",
		x"03",x"00",x"00",x"00",x"38",x"38",x"30",x"38",x"F3",x"77",x"F0",x"1E",x"10",x"00",x"00",x"20",
		x"19",x"01",x"11",x"1C",x"07",x"00",x"00",x"C0",x"60",x"40",x"80",x"03",x"07",x"C6",x"10",x"00",
		x"E0",x"80",x"00",x"3A",x"9C",x"CC",x"76",x"1A",x"4D",x"4D",x"69",x"69",x"2B",x"AA",x"AA",x"AB",
		x"84",x"E2",x"3C",x"FF",x"00",x"85",x"33",x"08",x"AA",x"AA",x"47",x"08",x"07",x"D0",x"64",x"B4",
		x"98",x"10",x"21",x"43",x"06",x"8C",x"19",x"33",x"00",x"00",x"C0",x"84",x"1F",x"7E",x"E0",x"07",
		x"64",x"87",x"40",x"07",x"C7",x"07",x"1F",x"1F",x"7F",x"FC",x"00",x"00",x"F1",x"FC",x"FE",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"01",x"00",x"88",x"0E",x"0F",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"0F",x"8F",x"8F",x"CF",x"CF",
		x"F0",x"F0",x"E0",x"E0",x"E0",x"00",x"00",x"80",x"1F",x"1F",x"1F",x"1F",x"3F",x"3F",x"1F",x"C0",
		x"E1",x"E3",x"C7",x"87",x"81",x"80",x"C0",x"C0",x"FF",x"FE",x"F8",x"F3",x"F9",x"3C",x"03",x"00",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"E7",x"F3",x"F9",x"FC",x"FE",x"F0",x"F0",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",
		x"C0",x"C1",x"81",x"81",x"83",x"03",x"03",x"03",x"00",x"E0",x"F8",x"F8",x"F8",x"F0",x"F0",x"E0",
		x"01",x"84",x"07",x"07",x"07",x"01",x"00",x"06",x"E0",x"60",x"00",x"C0",x"81",x"80",x"21",x"E1",
		x"00",x"07",x"18",x"33",x"27",x"4F",x"5F",x"5F",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"C7",x"C3",x"01",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"08",x"0C",x"0E",x"0F",x"0F",
		x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"01",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F",x"CF",x"E7",x"F3",x"F8",x"C2",
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"0E",x"0F",x"0F",x"0F",x"0F",
		x"C0",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"78",x"7F",x"3F",x"0E",x"04",x"00",x"03",x"03",x"03",
		x"18",x"08",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"07",x"07",x"07",x"07",x"0F",x"0E",x"08",x"0F",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"01",x"03",x"01",x"02",x"00",x"00",x"00",x"78",x"FC",x"FE",x"FF",x"FF",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"F6",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"1A",
		x"0F",x"1F",x"1F",x"1F",x"3F",x"1D",x"03",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"73",x"07",x"06",x"00",x"00",x"00",x"00",x"00",
		x"EF",x"FB",x"FD",x"FC",x"FC",x"FC",x"F0",x"E0",x"F0",x"50",x"B0",x"E0",x"00",x"00",x"00",x"00",
		x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"40",x"F8",x"F0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"06",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"F0",x"FC",x"70",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"10",x"00",x"00",x"00",x"00",
		x"04",x"00",x"11",x"00",x"08",x"00",x"00",x"40",x"01",x"10",x"00",x"00",x"24",x"00",x"00",x"82",
		x"00",x"00",x"00",x"00",x"00",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",
		x"00",x"10",x"01",x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"12",x"00",x"00",
		x"00",x"08",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"40",x"00",x"00",x"04",x"20",x"00",x"00",
		x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"20",x"00",x"01",x"00",x"00",
		x"00",x"81",x"00",x"10",x"00",x"00",x"80",x"00",x"10",x"00",x"00",x"00",x"90",x"00",x"00",x"10",
		x"01",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
	);

begin
	process (ROM_A)
	begin
		if (ROM_nCS='1') or (ROM_nOE='1') then
			ROM_D <= (others => 'Z');
		else
			ROM_D <= my_rom(conv_integer(ROM_A)) after 10 ns;
		end if;
	end process;
end architecture behavioral;
