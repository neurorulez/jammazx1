-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "72063040F244AB3AED2A5FF11FE0600B082324221A22644EFFFFFFFFFF249BD1";
    attribute INIT_01 of inst : label is "80C462225C8623C298426E31C478276E227FF65FFF786CC4C119464433FA4A19";
    attribute INIT_02 of inst : label is "E8443A26F0FAF8918DF0122827CE8C1610FC240B0E518412169541C343070301";
    attribute INIT_03 of inst : label is "301A20FD1886210C0FA8008061723FFFE018C84F73E1C416441A1DCC1B441D10";
    attribute INIT_04 of inst : label is "06DC95AD6B4BB9343030EF98C082A055DF20CD9C3704090803D007E6E10C1837";
    attribute INIT_05 of inst : label is "BB667AF83BC4CA329B14253AC668D1E922F78C726003598E06231180C0CBEF63";
    attribute INIT_06 of inst : label is "4248F199CC69967039188C4603011C8D9DD9085C6F03A0A3C83B781381102602";
    attribute INIT_07 of inst : label is "000000000000003EBB3CD2203067603602965BBE8466A4591870311576382092";
    attribute INIT_08 of inst : label is "3100000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "7BFF178D9635A001CEDA97BB37FE09FF05CC1935584C0DB4F3F219964CBB2660";
    attribute INIT_0A of inst : label is "0CEF9B0ED0D1D91A3635BDD02C8DEC01870C71C31C30C39DF6F9B7B2E093D960";
    attribute INIT_0B of inst : label is "D0377AEC20D6CB35B1A3637607EC24D5D81A37C46BB080DD55FC51BA823180D3";
    attribute INIT_0C of inst : label is "46305A966C229078CC4B0042EBAE80B88AEB800002060C193264FBF80401BED6";
    attribute INIT_0D of inst : label is "6238B2D6E5D27DD7FE7EC91637480110988C004C3012CC46082644910515458C";
    attribute INIT_0E of inst : label is "8061D030C884470AC467084EBD88D089118EB1709FCFBF963FE4EF810FBF9894";
    attribute INIT_0F of inst : label is "9C1CC18530984C260C434D25C324C9820E230E20288494C02A521430C230C284";
    attribute INIT_10 of inst : label is "FF3FF3FF34AFF5DD3FF2ECEEB77DEBF800008880808800008088808384830018";
    attribute INIT_11 of inst : label is "F3A7D7CFBEFBEF3ECBAF7DF36F3FFFED2BFD77F9F79FF9FF9FF9E5CBAE7F3EF3";
    attribute INIT_12 of inst : label is "74AFF577ADFFFE7DF7DE7DE6DE7FFFDB79EFBE7972AB987D8B1B360DB7748C87";
    attribute INIT_13 of inst : label is "4A4FDB6549F27F9BEEF51BFFBEFFEFFFFFFFFFFFFFFFFFF5DF5D77D75DF5D77D";
    attribute INIT_14 of inst : label is "DDEF6D236D72EF522DAE5DC521DB97F2496C9A143E6CCFC6CC7C49136308D11A";
    attribute INIT_15 of inst : label is "A5707D91268B192E8D486DEECC13C692E69A4BA903BC091B6B9764DDAE2916E5";
    attribute INIT_16 of inst : label is "290536DB2A41DF15DF6A90FE0652C020521D210ED104F8000001F4FCAA9F250B";
    attribute INIT_17 of inst : label is "C0C90C0623138C23183363094C460C64300D6309B23415ED9D0313C8743F7948";
    attribute INIT_18 of inst : label is "CE074D638E084870678CD81CD1870461C75399CCBABB66038E539C1AC6C1C1C0";
    attribute INIT_19 of inst : label is "3168420E2C5A4E6E30CE98168EF7A1070E9F8838E084C673988C464F25A30461";
    attribute INIT_1A of inst : label is "833210661C87A7573079E0C366264BBD222444C3F0908908908908B6A7906840";
    attribute INIT_1B of inst : label is "9A0E3B8E3324642914C3F9D3E32D73CBF3BD716A3E883E0A002502EA0DBEB580";
    attribute INIT_1C of inst : label is "50799CF62AA00B3283E4C82300E61D021CC0ECC6188881EBD8D756C98816C626";
    attribute INIT_1D of inst : label is "C42E6E0402175C8FB605333FCC5743E4C605D17BE2F7C5EF0BDE17BC2FC17AB4";
    attribute INIT_1E of inst : label is "9318D4B6C74B8646C6324023384C46180B18CC462EECF5EFFCCA6085033B11BE";
    attribute INIT_1F of inst : label is "43720C6449028920C6449011242B249849A0608D206891C111240481A2444901";
    attribute INIT_20 of inst : label is "716A81B83140FFD49510E98DEEC30C0C63192C71AA190A39952D062233433678";
    attribute INIT_21 of inst : label is "4F11A1E0401B1018FAC597068D991240907F19B634518DB9EB11B63405B6216E";
    attribute INIT_22 of inst : label is "D36233B6193F541AD703F818F35839CE73858A9FFFFFE7FFFF83CFE95EAC29B0";
    attribute INIT_23 of inst : label is "4D0BB1884C20F988C576316C1F254102CED8F9725DC1CDE7BD276C94B92EE0E6";
    attribute INIT_24 of inst : label is "AFF0BDF90BDE85EF42F7A17BF0BDF85D8C41F268C5768D850BEF47F68F8F883E";
    attribute INIT_25 of inst : label is "49ADECD820A8CD8B118962312C4626110A085B6B34D9B6DB6C643174006D0B6E";
    attribute INIT_26 of inst : label is "C88206440CA4BD083484A864908C3861B6C61C59435E6CDC2DED888B2540DA5E";
    attribute INIT_27 of inst : label is "95C7FC8C9A622062F70CC0D8626334DFB6C890E818C9626636B16228DAF74240";
    attribute INIT_28 of inst : label is "D2DA365E65EE8C599A624B6488BDC7617997BA35EEE653DEDC4897BBE894B200";
    attribute INIT_29 of inst : label is "E8571304C3038E0CC41C19CA61C0AF74C9D0B0A8732DCBD09269644911EE6746";
    attribute INIT_2A of inst : label is "C4C61C6A3C762CEDB0A95B6E46D82719898C38782A735EE46D8CC038C457BA64";
    attribute INIT_2B of inst : label is "B4C19E60ECF6DB170C1F5A2CF67E8421FD6F2D8B4DCDD8A8C28DAB6C9ADE2B78";
    attribute INIT_2C of inst : label is "3FC3361390950C9840BDC410329334A489C31F6220B6E69A71B63C0CB110B90D";
    attribute INIT_2D of inst : label is "A2E4E2CAE4EE8B5D6D16B1D2F23FD38A5643682ED0F487F21FDA2E34A106C2EE";
    attribute INIT_2E of inst : label is "A9FEECC450866920DE1263D031806F32217062131E83D021A69A437898C07816";
    attribute INIT_2F of inst : label is "000000000000001FF555567859DB2F08BEA3E403E819B4961C542A1221119A19";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000001044000000000000";
    attribute INIT_31 of inst : label is "8000000000000A20AAAA82AAA0882AAAAA82A82000080080AA00000000000080";
    attribute INIT_32 of inst : label is "8302E87C984C03E60C574C5A1F2430C09E0085012FE519158F3221FFC5B2D04B";
    attribute INIT_33 of inst : label is "1F9A266D211EC809445322ECF7F5B8A48BCFBD5017AC93224E400AA802AA83CF";
    attribute INIT_34 of inst : label is "E0E49FCAEDEBCAEAFBDAD935D5BAAEA1C5104307F818016600785ECC8999AF91";
    attribute INIT_35 of inst : label is "094C08A0B04B3F4CC4C6B94F9087FCCA0740B3C4CDBC588280EA194729FFD4E0";
    attribute INIT_36 of inst : label is "06BFFC2EF6628E5F865E1CF3E19A6495A19FBC05070A48E6D3C8000002CE5200";
    attribute INIT_37 of inst : label is "09FE23F000FF004FFB4F4732853D1C94566FFFE76A8A9713375C5F15DBB8EBFF";
    attribute INIT_38 of inst : label is "94056347FE9F3F977BB060CB48108244440E0A49863651887110910069EDCFE0";
    attribute INIT_39 of inst : label is "540055001540055001540000003EC6843CEDFE88F9A7CC7F602F188C83B64480";
    attribute INIT_3A of inst : label is "10880C4604224311A5B966C3B870000040401540055001540015400540015041";
    attribute INIT_3B of inst : label is "BE0C82D01434084298B433EB235B09B3484D9A426CD0FCA349813D94F348C638";
    attribute INIT_3C of inst : label is "3D806C033EC66E07B98119F333ECE510A03C9B087C9B09FB42711B13C2423E98";
    attribute INIT_3D of inst : label is "8BE89FAB75843E07029EAAF8DEFE5955600E34C4A70429443E6296F03999BD37";
    attribute INIT_3E of inst : label is "7DF75F7FEC91FE7B37FF79BFD58FCFFFBE3693749BF336A7FFCBB7F366937F57";
    attribute INIT_3F of inst : label is "7FFB56E7EBA4FD756E7EBA5FAEFF9F7DF7DFFB76CA5CDFBCFBEFBDFEC9943CBE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "9B29586135843A7B81B31E99B934E7534D35BE01A373766E1600000000A4F2DA";
    attribute INIT_01 of inst : label is "DDC2F5FFAED736EADD68F27AE6DC34F6F315502571100A880D8DE3761A7B630D";
    attribute INIT_02 of inst : label is "80FFE03F01DF80FF7F043DFC780FFF1BEF00D7E73FBF67F9F35CF5FF2A6E572B";
    attribute INIT_03 of inst : label is "FC4DE207084210845DFC1C67DEFE7800F3EFFCFDDF10047FFE3DCF5E3C07F01F";
    attribute INIT_04 of inst : label is "AD695ADEB5BCBD2EE746CFDB9827E3FFB83FBFE23EFE06FC3EF87C07DF8304BE";
    attribute INIT_05 of inst : label is "700D0057DD485D8FBDBB5F6797FDFBFCF7739C68D6BF4D9CEE77BBD5CA4F4767";
    attribute INIT_06 of inst : label is "B0E475D9EC53CCE57BB85EAE57AFEADDEEEB1C5EEDA659F695DDEDCFDCDB95AF";
    attribute INIT_07 of inst : label is "AAAABBFFFFEAEFFEDD1B27D57B3CEA9ED64353A6CFE7BABBFAE572FFBAF3153B";
    attribute INIT_08 of inst : label is "AFAAAAEFFFFFABAAAABBFFFFEAEAAAAEFFFFFABAAAABBFFFFEAEAAAAEFFFFFAB";
    attribute INIT_09 of inst : label is "98F8C930C1E31C94D0F3D73330E94754A5993249320DF932E6BBFBD25EF5F39A";
    attribute INIT_0A of inst : label is "FFB55DFF246BAF1A1D32DFF556CDC297AFAEB3CF3CF2CFAF0904E8339F4C19DF";
    attribute INIT_0B of inst : label is "064CAFF7FCDAADF2F9A9533BFEF7F8DDEFF9375265DFF6D3789B0983B165F3DD";
    attribute INIT_0C of inst : label is "73B6989C480240DAF92B68AB4D34AAD3574D1DDDDFAB162D5AE1E5E818083A7B";
    attribute INIT_0D of inst : label is "844DA76F4A9B199B0D8C49DA6B175F3AB85E739C709A5E6E1C266A7292EAE4EC";
    attribute INIT_0E of inst : label is "914AD070E8662DD8CDE3A956BB3C59F9B8C4EDD291FE323C16368CBDFE32304A";
    attribute INIT_0F of inst : label is "39B861927E3F1F8FDDEB6D84E9B3E8D25662766A6C6236634CD91C30C6E546E2";
    attribute INIT_10 of inst : label is "00020020291082088100000048800006EEEFF6EEE666E66677FF7FFB8E833FFD";
    attribute INIT_11 of inst : label is "6BFF882000082082080082080080000840208104100104104105080400200208";
    attribute INIT_12 of inst : label is "A91082028000000000410410010000000010414201001CAF5EEFA1BE79DE6E06";
    attribute INIT_13 of inst : label is "24C2932509A48804000000000000000000000000800020000820020800820020";
    attribute INIT_14 of inst : label is "BE83833C3DE5DE3BC7BCBBE33E8F2EEBFDBEF7F9C768C3BE63D664FB6B47F0FE";
    attribute INIT_15 of inst : label is "DBDED6FBB87D2EE6F5EFE3C0CC8D779F695E7CBDFC7939E1EF2EFF87BD19E3CB";
    attribute INIT_16 of inst : label is "DFBBF0335FFC9DB7BA21DFDB5458BD0A3BE919FE69A637FFFFFB419DFFE76FDE";
    attribute INIT_17 of inst : label is "EA795CAE57BBCC7E3DE16F89EB3FD9DAE3FB4ED7F766AF55A8921F96BCD5D2F9";
    attribute INIT_18 of inst : label is "E42A494F1C7D0D6577BE90A97537BD4DEAEF3DE8D1674F550F6F3E6E959783D5";
    attribute INIT_19 of inst : label is "AAFF35D4F2B9FEF5E79CD2A4D4A735AB54CB2CF1C7D0DF593D5C274596EA7D4D";
    attribute INIT_1A of inst : label is "D59F5AB636D76D7D0EE95DEB4E124DE9E5FEBFDEA44A3EA3EA3EA3FC72DEFFFF";
    attribute INIT_1B of inst : label is "935D316F5AE44007FC49928413FBF0FEC0F7C1FE7F8FC1008BDF07DF87FDCDFF";
    attribute INIT_1C of inst : label is "B9FEFBFED5F57667BC2D9DE7BA1659A7CC3ECCFF397CD2C1B39213BF2FBF94A4";
    attribute INIT_1D of inst : label is "739996F2796BAA71A751B1858FBFCF5BE7CFF3F787EF0FDE1FBC3F787E03F77B";
    attribute INIT_1E of inst : label is "850EC4E3424E8E47EF364BBBBD5C2E384FBC5E2F3806810B2620F7533C4CC859";
    attribute INIT_1F of inst : label is "CDF24763D9287B24763D928F6493ECA84FA4BC9D24A7B3C90F2C84929EC3CB22";
    attribute INIT_20 of inst : label is "E3DFC7F7EFC6DF7C7BF83F9F7ED31C3EF7893D96B379D971B3BA7433320000E4";
    attribute INIT_21 of inst : label is "5BB5B5D734F4ED3773B713AA7B3B734A3380E1FDDBBF87E03EF1FDDB9EFDC7BB";
    attribute INIT_22 of inst : label is "F3DFEDEE76F6FC77FDF007F76EF80000001F9F0000000000001B0FF9F2E7B9D5";
    attribute INIT_23 of inst : label is "BE1FE1F0FBC3D6F0FBFC3EF87ADE478FB7B9F7EDFBC77BE0FBDBDCFBF6FDE3BD";
    attribute INIT_24 of inst : label is "C091FBC01FBC0FDE07EF03F781FBC0FF0F87ADF0FBFC8F0E1FDE07FC8F0F70F5";
    attribute INIT_25 of inst : label is "DB2F48DA6DB86DBCB72F96F5F2DCBE3F1B7849F20040000001D7E0B02E3F3FFB";
    attribute INIT_26 of inst : label is "C5B6E62DCC76133D24C5987419F63BE837A4A8A2A46428E900491F9B6CC0484C";
    attribute INIT_27 of inst : label is "2A7EF9DE924664246709E5BD15152497348CDEEF0D19677326B9636CC4663ACC";
    attribute INIT_28 of inst : label is "825B00495DCCAE4B9246D94D98198F6AA5773290CEB425365CD993339DC10AB5";
    attribute INIT_29 of inst : label is "EC2B371CC71B1E6DC23CDBC473CC8665FDD9B9B8CAED95D482502DDB30CE3766";
    attribute INIT_2A of inst : label is "97E6B941B9BC25C925984E2D3D934E532FCD72326E210CE3D9ADC339C2433AFE";
    attribute INIT_2B of inst : label is "340218608BB0DAAB490AE7BBE6598FE6D13A451D15B9D5B8D27B09C5B2748BD2";
    attribute INIT_2C of inst : label is "00EB97BB1AB30E8CCD19CDB731D316AE85A67E67E493E491272499686B30998D";
    attribute INIT_2D of inst : label is "E7DBDF87DBDF1FF7BF3FF0F3EF1FF07E7BF1F9FBF3D7E39F877E7C7BE7E38FBA";
    attribute INIT_2E of inst : label is "C8C5AFB7E9FC7B6D89F0659A7FDD1637313AF3332CD1BB6FE49068B3F2E8F73F";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFEABFF55557F1F6F73EFF7F6AD7E5B1DC6E935CCC6616E3F0E75F";
    attribute INIT_30 of inst : label is "FFFFFFFFFFFFFFF7FF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1407FFFFFFFFFFF";
    attribute INIT_31 of inst : label is "55555555555575D555F57FF5FF77D555557D5FDFFFF7FF7F57FFFFFFFFFFFFFF";
    attribute INIT_32 of inst : label is "73E7F9EB7CFBCF5BCFBFCFBE7ADE73CF9E73CF9F3D8DB34E4466BE0D3E72D9ED";
    attribute INIT_33 of inst : label is "F6CBD3F99FCEA0D47FF38F666E65E76485BB3D777306DA3446E80822A80003CF";
    attribute INIT_34 of inst : label is "DADD8DCADCAECEDBF3539F2D9C60E4EEA046C6436EFD619F5047D0CF859F29CC";
    attribute INIT_35 of inst : label is "CFFAD5FF4DC7ADCA67E631645F51F0A666B9C63DD19DD568EF67CB6F043B00DA";
    attribute INIT_36 of inst : label is "ABF6BEAED3F65E5723D45293C8F2C633B4DB13A8A27E63ECADBBFDFFCFFBEF7F";
    attribute INIT_37 of inst : label is "62499B85A774AB12F11A46470469193814CFFACC69888C8845DFDE8019A775E2";
    attribute INIT_38 of inst : label is "7B9EF1E003E0E389492F368EDBCE76EAA4163B4F8E57A4CD7370BF3C6D033557";
    attribute INIT_39 of inst : label is "BEAFAFABEBEAFAFABEBEAFFFFFECD7D69890017D03201806FCC607FB7EEE7BCF";
    attribute INIT_3A of inst : label is "F1FCF8FE7C7F7E3FAC9B66F3CF8FFFFFAAEBEAEAFABABEAEAFABABEAEAFABABE";
    attribute INIT_3B of inst : label is "00000000000000000000028B1B568D586C6AC363561B59730CD17596A727DB5B";
    attribute INIT_3C of inst : label is "DDD98ECC7F314379ACE89DD22767EF8DF570D9AD28D9ACB71F59B29000000000";
    attribute INIT_3D of inst : label is "0000332AD733993D94C8EBB289BEF67F13F5A6E32BBEBDE68D137D9BD41CE3CE";
    attribute INIT_3E of inst : label is "04100104052210414D002A4000A0180010080009240080802200002481B68000";
    attribute INIT_3F of inst : label is "936157A5B222B6C17A5B6016C880410400410508040020820800820A10080040";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "3B69DB66193645E459022FBB9FF55BE77CB7AD89F3A634C6FF000000000BCDD8";
    attribute INIT_01 of inst : label is "66F379A71E97626BB940B299CE4DB796AA700C50A4488C010D29EB74D2FA436C";
    attribute INIT_02 of inst : label is "78921E13D1AF681ED2F02FDC5FC30E1DB1FC636F35EEA0E2249DA4F7289DBE4F";
    attribute INIT_03 of inst : label is "981320F814E7394A1AF000853BAE5FFFB37F4CF2EBE1341D403E9FDC3F40ED0A";
    attribute INIT_04 of inst : label is "5FBA2042C6354DF41DD513DB22A283DDEF0772FC0D3801A029F053E1B40A140D";
    attribute INIT_05 of inst : label is "FCDD603F6F74FB61FDF683FB61AF5E9EAFB9A9EBE5618DBB7C9ADDAFB75BD36B";
    attribute INIT_06 of inst : label is "0C9D32666DEDF7DBEFDE6F3C9EFDB986DF79184E778FBE6FFC6F734B749FE4FA";
    attribute INIT_07 of inst : label is "5555555555555F84EBEB7BF246E5B92C643B2196DFBA4A14D1CBE7DFD6960727";
    attribute INIT_08 of inst : label is "3555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_09 of inst : label is "6FFFDB10D5AE176DCEF5411157FD45FFA199DE9EAA3C2B1763FA5F3ADCB7DE39";
    attribute INIT_0A of inst : label is "DCEEFB068F85C9C2BB8495D584A1EA5056C92D92C96C96CCFA754B5E2ADDAF05";
    attribute INIT_0B of inst : label is "85CA7B6C22177B1CB42BB876076C3616D85A86D709B88C1CFDF55427ABA48A13";
    attribute INIT_0C of inst : label is "CF432151D624D21ADBB739FE4186A7924461919912EBD5AB5EBD75F4E2903E16";
    attribute INIT_0D of inst : label is "2CDD17334A937F9FFFFE190A605F949BDE79AFACEEFF6FBCDD67465D204537D0";
    attribute INIT_0E of inst : label is "9B2E0DBFED543CED14BBAD4EBB4F52F7929D0E13EFE757537FF4D5D7E7575DA3";
    attribute INIT_0F of inst : label is "FAFBD7CDE5F2F97CA96F4DADEBB6EDDA207930FDA852D4F28FD399FAEBCA6ED6";
    attribute INIT_10 of inst : label is "AEFAEFEEB4AA458D7E5F7F54F72FBD204444D04CCCCCC4454CCC55F4D2EFBFD2";
    attribute INIT_11 of inst : label is "EBA9EBAEBAFBEF3EFFECBAEBBEBCF3CF2E91E3F9B7BF7BF7BF79A576CE3EB2EF";
    attribute INIT_12 of inst : label is "648A41A27CBE9E7DF7DF79F77D69E79FF9F7DF593DC3191CFDFB63E8AB3EC48F";
    attribute INIT_13 of inst : label is "E0578FEBA9924EFBFFBAABFFFEFFFEBBEBAEFADDF7D77DFFFFDFFFF7BEF9EFBE";
    attribute INIT_14 of inst : label is "E7EF87534C70F375298E1E6753D387F9369A6D0E22449FFE567EEC566A5FF7FE";
    attribute INIT_15 of inst : label is "8081FEEB44637D9C48D44E47DC9F87AAE21EAB1A82CE9A9A638787098FDA94E1";
    attribute INIT_16 of inst : label is "BFF3EC7F5D4FE2889A2BA8FF4406DDCDB5183A84B534FC510545F5D440355A75";
    attribute INIT_17 of inst : label is "B3E7FB3DBE4DAEECF245B11B7A01D05084072684CF4546EED57831040FABA1DB";
    attribute INIT_18 of inst : label is "62F1770E1099291599BE4BC5524990D26AEE2A6180548334136E2CAA11571727";
    attribute INIT_19 of inst : label is "283820326A0E7E7F47E8C2488DFE31D3A07E2EE10996DE7BDE6F3F6FBAA4B0D2";
    attribute INIT_1A of inst : label is "C5FB12BE5E97CBDB2D762FE0F7DA5BD16BFF7FAFD239A99A9989988A2FCCFEC0";
    attribute INIT_1B of inst : label is "D75B5097B6C0A1003D47F5D4F0F7A335335A70FA5087FE1F02FF043C8BFDDF80";
    attribute INIT_1C of inst : label is "786D5F4677D7F7EB427FE8D913D5FFA37B73C34377EA99CDE4962639ED52C623";
    attribute INIT_1D of inst : label is "77958165BACA2E0EFF4D1BBFCB768AE7658DA3AD475A8EB59D6B3AD475E3AFDE";
    attribute INIT_1E of inst : label is "DDBD0B8E6AA88A4E625B43B44DEF367779096FBCDEE6306FFEAB77B4C5919F55";
    attribute INIT_1F of inst : label is "7BDB5F8FDFAFFBF1F8FDF8FF7EB3AFECC9227EC9227FBD493F7E1489FEFFDFA6";
    attribute INIT_20 of inst : label is "71348659D043E4A4F6E0DE16976BB9A6312B2DA4031B3FA7FEE615265E11E27C";
    attribute INIT_21 of inst : label is "68DE31F26617D894F43837A7DB57276BD0FF987E666E8BF9FDD07E661D7F275D";
    attribute INIT_22 of inst : label is "73FB17FE697BFC6CA6D3FE7CBD28FFFFFF991F9FFFFFE7FFFF8FC2309E5E11EB";
    attribute INIT_23 of inst : label is "779B596CAFB2B94CB76B2DE65735860B5FF96E5797C6AEC757EFFC572BCBE357";
    attribute INIT_24 of inst : label is "FFF1D6BD9D6ACEB5E75AF3AD59D6ACDACB6573BCB76B0BC59DB5E11B07C79CAE";
    attribute INIT_25 of inst : label is "D94405423FF77C2C9FBDB3D7B27EF5D6EA36DD25AC6A800824162E940E5F0E44";
    attribute INIT_26 of inst : label is "1EFB50F7A5FEF66C82969FF650FE218CD610C48A1807C084D880AB6DBFB5E56F";
    attribute INIT_27 of inst : label is "406BFFC4CE7FCEFC4DA047C8CCCDAC6FD0DE9F87BB5204C89026204DA05FDF7A";
    attribute INIT_28 of inst : label is "5B4A6369D6BF64DFD63A3E97F217E02AA75AFDC89BFFA57C577F22FFD526086C";
    attribute INIT_29 of inst : label is "86017E7C2E78BFE39B7FC7FE17FC45FCDF0F8BF38EB7556F418427EFAC9BBC30";
    attribute INIT_2A of inst : label is "DEBB156E4F0B6F9DA3D2B876EBA1C509BD762A62F4F489BE9A039F0B9A226E6F";
    attribute INIT_2B of inst : label is "B8ACFA6C2EC358C160BEEEEF5DFF3789FAE0340BD6273FD367DAD70D95C29108";
    attribute INIT_2C of inst : label is "3FEBB9FCDBD3FEDD6B1377DE97F8649573E19D0AD9BA739F2802154B7FAEDD24";
    attribute INIT_2D of inst : label is "27A6F14FA6F292995F2531B15A2463F415F2F9D5F2E3E5EF9BBE7A2EC6A4CB4E";
    attribute INIT_2E of inst : label is "D008369D44372F37FB8E5DFA3489D7B7A37A3252EFD5E63CB58F46BFDFE0FC25";
    attribute INIT_2F of inst : label is "8AAA8AAA8000A978D2D2D7F96BFF15E9D367FC33D448F9DB7D4FEDFEDD6FC7AD";
    attribute INIT_30 of inst : label is "FFF5FDFFFFF7FFFD7F7FFFFDFFFF7FF7FFFF7FFFF7FDFFFFDBBBA0000AAA8AAA";
    attribute INIT_31 of inst : label is "D5555555555547564A2DBFD7556FED6CD4FA846DE9A0929F015BFD6A7427D05F";
    attribute INIT_32 of inst : label is "92C6D15CECAF8AE50B768B785734508784328D8A2FFDF520ABEA413FA6F752FB";
    attribute INIT_33 of inst : label is "5FDFDF159F09F487A06EB80EF4F90A5ED3F7C68E5F85DB63C67A0208A0A081C7";
    attribute INIT_34 of inst : label is "C0C7DE84DCE4C4F97BD959ADCAEA465CC4FEF6FFF649D7127DE16F8EF71977D5";
    attribute INIT_35 of inst : label is "C57A5BAFFD793EFCE64CBF4FC0F4FDE307B28B3F3C92684F500837F43B7F80D0";
    attribute INIT_36 of inst : label is "AD5FFFD17F1FE83FAE6E6733EBCFE6DA71DFF7726525AE1EABF77A2FC2F5DAAF";
    attribute INIT_37 of inst : label is "F23F3BFC72FEAF87FF9E2654FE789907B2F7FFE1B9E6CE46F1DEDFCD699154EE";
    attribute INIT_38 of inst : label is "F61DB247FD3FAC7E2EED2477FD7F7ABB14CCBA598A3A6EEDF7EFDE4D2982AF95";
    attribute INIT_39 of inst : label is "040450450515405011055400017F6BC6BC66D3FCFDBEECFF4CBF1EC59DBE278B";
    attribute INIT_3A of inst : label is "F4FAF2797D3EFC9E6DB927431054000055051505405110050450051515445111";
    attribute INIT_3B of inst : label is "EB6C3C9244D33B444750D3D59D0098EEC4E77727333AFBE768D7BEB4EF67EF3F";
    attribute INIT_3C of inst : label is "DF863C317F696B7DC898C8FBB7FCF51AA5FE99A97ED9ADFF7B9B0F53D4F1D10F";
    attribute INIT_3D of inst : label is "E10867C4883F7F07B9DB143EFB6DE36F58FCF4780D1C9CE6CE8AF2DBF65D97CF";
    attribute INIT_3E of inst : label is "75D7DD75D5930A3135E2FBB6968BCFD79E25BF7DFB4F9B4AF3CE9F7A4E9B7E7F";
    attribute INIT_3F of inst : label is "320DB89C26D784DB89C26D709B6F9F7DD7DF79366756FF3EFBAFBEF248EE187D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "258BCD164953EAAEB840C0FDDE889961A38C1B55B88CB9970000000000B54CFD";
    attribute INIT_01 of inst : label is "B55AAF957774AAFA7B30B0AB115E8FF7D980065000007D46FCE7B9E3CFFC91E6";
    attribute INIT_02 of inst : label is "970505E62E45978D4E2BB4CB683980FA84034D14CA213CE48A3A6933F98AF5FA";
    attribute INIT_03 of inst : label is "33A11D00EF3BCE73A45BE319409DA000CC8D0389500FFB8B01E8A931E8BCE2F2";
    attribute INIT_04 of inst : label is "79D23184339DDF528CD954FD66D8188010E70D81C039F82B8A9714180576EF40";
    attribute INIT_05 of inst : label is "D457F2057AAFD5ED2DAB9A47F3162C3F9DFBC78E9FA38FD7EBF57ABD7FB1D7F5";
    attribute INIT_06 of inst : label is "98A57AAEFEA8AEAF55AB55EBF54C2266F3D6A1212A64D774E67A5E4AEC8FC0F9";
    attribute INIT_07 of inst : label is "FFFFEEAAAAFFFBE67E7F74476C01B3B7707BA3D7E8F0EFB49CAF5DC6FDA7832B";
    attribute INIT_08 of inst : label is "80FFFFBAAAABFFFFFFEEAAAAFFFFFFFBAAAABFFFFFFEEAAAAFFFFFFFBAAAABFF";
    attribute INIT_09 of inst : label is "0C3EC8576B9BEBECE92D4445983DD41FE933DC92AEBEA65A48394AFDA137F033";
    attribute INIT_0A of inst : label is "D6AEBCA163860E46BA88CE548623EFD059679E5D779E5D74482E59E0E864D0E5";
    attribute INIT_0B of inst : label is "7BC88B7212375C80C46BA8B913720636E40B8ED511CA583DD3F75456DAF5D831";
    attribute INIT_0C of inst : label is "08CB87C6A90CE6FACE4D3AF43043AD0CC410F131BAE1C983260CB4F77A344E97";
    attribute INIT_0D of inst : label is "289339343A6CBC480081661898DC858F2B57BD815E8D97EAF299934CD45BF213";
    attribute INIT_0E of inst : label is "2D1E375412F1ABF52AD8674A86E7851B4E7BA1E7706389EB5F8BE27EE389ED19";
    attribute INIT_0F of inst : label is "86A2B4390782C1E0A43D1E68184C1238B198B10D437AA15BDE85AD8434FB357A";
    attribute INIT_10 of inst : label is "000200001364BE01268000009B40080666677E6EE664EEEE77FFF77B36687FCE";
    attribute INIT_11 of inst : label is "57DE0C00000000800020820800000006DD2B00840040040040049B247C300200";
    attribute INIT_12 of inst : label is "9364BE01C0002104104000000000000104104136E958128B76FC81F6DADB532F";
    attribute INIT_13 of inst : label is "B33887F3A6649205E80004104104104104104100020000800020000800020000";
    attribute INIT_14 of inst : label is "4D7C92D0CA48A7E5194914EED13245F64B25BD42289328F4337F760ED397EEFD";
    attribute INIT_15 of inst : label is "9AA9849AC7E2D4814AB41CFF23B2AB68932DA152829C968652453CF94BD68C91";
    attribute INIT_16 of inst : label is "D6DECC3F9D3ED5D7D7FF687FC1A6DCDDAD02DE81FC7101515005FE5515350041";
    attribute INIT_17 of inst : label is "5A0A55EBF5680357AF5E02B477A3D23B1BE73DF0CD4AE9781229E06F89044797";
    attribute INIT_18 of inst : label is "F110E33CD33363C9ABE72443B72BDDCEFDE8E2F2C540946457E8E136312672F5";
    attribute INIT_19 of inst : label is "FEB1FC33DFAC27994FC32EC367F4497AF1A2EECD3132F0E7ABD5A0905F6E7DCE";
    attribute INIT_1A of inst : label is "35808EB409714BE4FDCA5D13EABDA0225DDBAB37DE3B27B27B27B25B18F4F6BF";
    attribute INIT_1B of inst : label is "2CC58041E8ED4B53BB17ABEF0F407CDC0C844D118A6B00E07602FA52753FD97E";
    attribute INIT_1C of inst : label is "0610803500028B5CC2B8555A3942A669C5613A012AC2293C7671D1E4E540339F";
    attribute INIT_1D of inst : label is "3190637138C02348D8DC44403621F000BB387C7238E471C8E391C7238EDC7102";
    attribute INIT_1E of inst : label is "7CE33E39396728B8A501B9955795A0AF429597EAD9BE083FD1F68D70E4C4C705";
    attribute INIT_1F of inst : label is "102DD09AB6EF565D09AB2EEADB900B67319A4E6CDE5565B8EADBB37955BAB2EE";
    attribute INIT_20 of inst : label is "0C1A39B1C1B800470217317B6E00D7EA5234CDA423CC151E2BEAD3C938B44B76";
    attribute INIT_21 of inst : label is "D7E24DF77ECD5EA61E87A06D72CAF4B9ED8007A4D0217526228FA4D060A4182A";
    attribute INIT_22 of inst : label is "1E490529C00483C0714C0104485700000060706000001A31CF60300711E03F40";
    attribute INIT_23 of inst : label is "0A70E6C3608C00C3621CD82980083C7194A69004023C6938A00A538802011E34";
    attribute INIT_24 of inst : label is "9E0E391A639131C898E44C722639138736180053621C77326208980079393300";
    attribute INIT_25 of inst : label is "92F9B62E9D1A94E4CED4B9DA933B52AA50DA820A5BEC5925B6F29919FDA9C562";
    attribute INIT_26 of inst : label is "2D147168E2E986429E395A094671C495A9F3E6EBB883E6E6DE9257E808FC2D97";
    attribute INIT_27 of inst : label is "58683C4A25F4EA0C19E68455CDCC5BE183E22D3B831D16EAF1371667E819FC9E";
    attribute INIT_28 of inst : label is "7CA0FB92B333B0822DF8C7E13B066C988ACCCED833F37C642613A0CFD136DC9C";
    attribute INIT_29 of inst : label is "3BE1A54C65599565572ACAA632A6C19E3275191B559AC477DBE5B382343349D2";
    attribute INIT_2A of inst : label is "6A50473DE70B4032591BD382BB65C9CCD4A08E8E469D833BB64553195760CF19";
    attribute INIT_2B of inst : label is "0E74399D36CEA7C1E683ED571AFD2AAC1F4D9066B3262D1A0576EAF12E9BAEEE";
    attribute INIT_2C of inst : label is "C09A7A854F2B41229B0669A38BA8B1E9DBB0CC956904097D8C492362CA7F2D77";
    attribute INIT_2D of inst : label is "9CC000B4C01C61C4A9C38E7E84C00C1DCA0D4E729C141A106453CDD0789A31A1";
    attribute INIT_2E of inst : label is "EE2BE06B3CA38E8C4315AC669D1CD1858A0610CD6334749C0B7D168E0E1314C3";
    attribute INIT_2F of inst : label is "AAAAAAAA8AAA280FFA857BFE3294E82524EBEB9415C0DD59EEAD4E84EAB40685";
    attribute INIT_30 of inst : label is "FFDFFD7FFFE7FFFDFFFFFFF9FFFF5FF7FFFE7FFFDFFFFFFF9AFAAAAA2AAAAAAA";
    attribute INIT_31 of inst : label is "0000000000001F778758555F67D7C8A68878D8F7E9749F5F567CFE096617B39F";
    attribute INIT_32 of inst : label is "3D9C3E001760B0033621F60B80098C31E19C3865C1EBAEB0A95D4147FED80594";
    attribute INIT_33 of inst : label is "BF3ED03857D125DDA87ED81103FFBEEB602FBCDF4851E5B9571F55F555D5FE79";
    attribute INIT_34 of inst : label is "969121BEA56EBEAB913F845D5687EAB0458595A5F5D4F415352512402484C84C";
    attribute INIT_35 of inst : label is "FC7B7A7FEC123ED02282AA1140F47D30C0AC0119752395EB51100AF8970FA886";
    attribute INIT_36 of inst : label is "ED408BAAF0357136E113338FB814B1A3C83F86306665B6106833E7DFF00A0F7F";
    attribute INIT_37 of inst : label is "B2A1BBEB561FE588F48E2836FA38A097BD387FE74DE14CC84ED1D342F0AF54D7";
    attribute INIT_38 of inst : label is "0060CD380280FAF75CDF5634D5EF5099B3CB98E569E07A67BAF423CD839207FC";
    attribute INIT_39 of inst : label is "EAE5BBB97EEE5EBED7BFF455547E2F2181C20932069934CF7F9062411C89D038";
    attribute INIT_3A of inst : label is "6F37B79BDFCFAFE7F36E920D10455551FFBD7EFE5ABFD6BFB5EEED7BBB5FEAD6";
    attribute INIT_3B of inst : label is "E3CDA92B34D148849F86C7EF9E57F6C437B621BDB98E1ECBE3F21C412BB57C9F";
    attribute INIT_3C of inst : label is "DD4EAA75877938D8D7B9C671186262DC5C9E3FE33E3FE33FA8FC4FC5C915BD92";
    attribute INIT_3D of inst : label is "00207FEB9DDFC1A6582FBBFDC395632BDBB0F31BDCCB93BBCF9165C6C206264A";
    attribute INIT_3E of inst : label is "04000004026C97C0E90024D400402A0000DB24D9255080000012010DB324B911";
    attribute INIT_3F of inst : label is "4424A0702050040E0702070081404000000004DBA560200008008001B74AC040";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "BB51BE734C55D9388356B8C2016342849BA92C0087228C5150FFFFFFFF839100";
    attribute INIT_01 of inst : label is "42A150A0488F4390D0EC3E34EE33BC21728002102EAB3E283B8FE3AE1F024F0E";
    attribute INIT_02 of inst : label is "0720C1D80F080730200BC00B803264E04A038893C4045B0549220AA6511C0E97";
    attribute INIT_03 of inst : label is "C3ACDD06E358D6B5B083E77A860188008E2A4B40050E03F059D92A2DD83B00E5";
    attribute INIT_04 of inst : label is "001E95AD6B4B12E00070DD2340DFDC5D80D80001E4C1FE53D4A7A81C8A70E364";
    attribute INIT_05 of inst : label is "93A8134003D03A4A7674D4E00C68C1C0A0026831C81062381C0A1503A5E9041A";
    attribute INIT_06 of inst : label is "02254BFA91C509D0E0542A1D2E8501C9081D7BFC3D1EA69ED80320B10B10070A";
    attribute INIT_07 of inst : label is "000001545540480581358A0AE8E2245A1F1096403D2E942009C0E85002BE498B";
    attribute INIT_08 of inst : label is "4800000551550100000154554040000055155010000015455404000005515501";
    attribute INIT_09 of inst : label is "32211797D577FB2305F8B7DE6A20051104CEC07C08004DA4302A8F4F7E208E44";
    attribute INIT_0A of inst : label is "A6A4A709592EAF9E503ADED276CF0D6DAB2EB2CFACBAEB3B93D9129090916858";
    attribute INIT_0B of inst : label is "3FA74A5CC4F2172AD1E503AE625CC4F4B98A3C49757108F05A8125DBFADBA9FC";
    attribute INIT_0C of inst : label is "D7B07E65738EC65197FD177B5D5596D7AB555133121F3E68D9E3C56F6AFE38D1";
    attribute INIT_0D of inst : label is "EAB87BC641BA82F020A02F56C77AC3BDD4384A6DE057EA1D09BF64508C0FA5EF";
    attribute INIT_0E of inst : label is "B059E0AAC6171EBAF40B38DE19959EA098EE2651C474F8FA10673E2534F8FA6D";
    attribute INIT_0F of inst : label is "1898F3B33A9C4EA71C767104CD63C6AA8F62AF29AE905720A1DD9076FA04FE14";
    attribute INIT_10 of inst : label is "EF7EF7EF36EFFD9FFE7FFD7DB73FBDE9111089991999999988000004A0874037";
    attribute INIT_11 of inst : label is "08C21BDFFFFFDFFDFBDFFFFBEF7DF7CFBFFFE6FFE7FF7FE7FF7DF7FEFEFF7EF7";
    attribute INIT_12 of inst : label is "F6EFEDB73FFE9FFFFFFFFBFFDEFBEF9F7FFFFF6DDFFF3D3CA9112B03872D0DAC";
    attribute INIT_13 of inst : label is "426057F73DDB7FFBFFFA5BFFBEFFEFFEFBFFBEDFFDF7FF7FF7FFFDFFFF7FFFDF";
    attribute INIT_14 of inst : label is "8182ABA00524403A00A48803A181228400492E140CC8D8D4EC40885105281903";
    attribute INIT_15 of inst : label is "32700383204998178CC87012DE0B8DD0EA37403D0080DD0121220000A4FD0048";
    attribute INIT_16 of inst : label is "E919256046108C99CE019040261C0AE9F204110E21F70011555102E000281061";
    attribute INIT_17 of inst : label is "8D41BA5C4EA5AFF175A7B3ED7C26AEE735497F0926BD7FC69E5BD1C8661BBB6D";
    attribute INIT_18 of inst : label is "94D6895F058CCFA3FE39935B49E6763D9BDF6C99B53B57B964DF6EA98C8F8F5B";
    attribute INIT_19 of inst : label is "50C05A4FF43038543EAD995FC28B62040D031AF058C81FD0542A16315293F63D";
    attribute INIT_1A of inst : label is "8E5239CBDCC923BE18A5F3C5150FE8DDB6E4CC9A32A11E11E11E10E630EC1C00";
    attribute INIT_1B of inst : label is "9A30759E12409FFD0629FB9EFC000C008C018EAF91F040F5744DF900F15062C0";
    attribute INIT_1C of inst : label is "96E4294BF7FD5EFFBCBCAB935514793E3892D52EF138FBC3888AE4A92A7E8C62";
    attribute INIT_1D of inst : label is "D50ECC44E2269C45262DCD54391437085CB50C00180030006000C001802C0229";
    attribute INIT_1E of inst : label is "EBDEFA66FB3682E2D6DB65533EEA16F02B5BEA5D2334D5282C496A64A1331230";
    attribute INIT_1F of inst : label is "609B2E7469948D32E7469951A64964DF7B3AFCB9F0E8D265D1A667C3A344699D";
    attribute INIT_20 of inst : label is "AF81B806063FD21B20470860034BFA0D6BFDE8B074AF7AA8F48C44EAC9FE4BC8";
    attribute INIT_21 of inst : label is "6C75E30AC59050701D93133289B70244FE0066290984F146201E2909E828DA00";
    attribute INIT_22 of inst : label is "2E86C94782527F810C2C00E32097000000726F6000001800007F3996627E4E55";
    attribute INIT_23 of inst : label is "84EA0F271B1DC2279141E4B3B844B874251E448921F8189802128F024490FC0C";
    attribute INIT_24 of inst : label is "0C1E0004E000700038001C000E000750793B84279141787CEC803CC974744770";
    attribute INIT_25 of inst : label is "C98149D9E3E17B2E713DEE27B9C4F5542BA04DECCBACDB6C9355306A218AF891";
    attribute INIT_26 of inst : label is "FAEB97D62F94782BA8F685639F85B8E511859AFBFD2CAA1B31C928051F05FB6D";
    attribute INIT_27 of inst : label is "DE9220AD920F96E2E60ADCDBBAAB344145BAE2D1BC8471FFD70C712FB2E61772";
    attribute INIT_28 of inst : label is "BB7BC76BF6CC5C499A2E3CB7C4B983656FDB3175CC86F386D97C47323437B063";
    attribute INIT_29 of inst : label is "D17AFEB21EB078C3ACF107110F1AAE6385A387E59FB6AB825BAE5C2FC1CCB682";
    attribute INIT_2A of inst : label is "9EAB58C2386424EDB3C186F646D8A6313D56B1F1F82F5CC46D83A887AD5731C2";
    attribute INIT_2B of inst : label is "123E291D2EB5423ACB3A30F865401700161A1DE945C993E1428DA0DC98147051";
    attribute INIT_2C of inst : label is "C0CF1AF75DD0AC6B62B99658BE5BC7355B42066A809BE482212438D9B7C2D4F7";
    attribute INIT_2D of inst : label is "7B094C33094264330AC87E8C02D32C01B08C5600AD4118846115B1811A59B41B";
    attribute INIT_2E of inst : label is "B70C94557644EFF0BC804593E1AA967B3933EBF22C9B88E3A68870B293C743C8";
    attribute INIT_2F of inst : label is "A000A000800037F77280044684A3C01202561734107D22D7B142F85F0543D92D";
    attribute INIT_30 of inst : label is "002A02A00000000280080000000000020000000000000000100500002000A000";
    attribute INIT_31 of inst : label is "0000000000000A8290A92AA0A290295A978528B4095A95A0EA2C0202A4A85E80";
    attribute INIT_32 of inst : label is "4E5A86E10B1B3708B914392DB8458DF873CDF570ED1D7F528CFE9E44030D5E3C";
    attribute INIT_33 of inst : label is "B083AA67311ECFAC43EBA2750D0AE1B6D0001A1130061A40A040A8A8A2883D34";
    attribute INIT_34 of inst : label is "686EA0B270C7A674C5B48B648D9A65298F61EE37025EC7B7B1C8D8C5C98B2C64";
    attribute INIT_35 of inst : label is "33B21800D463483866F6947020E840C285D15446D0BC5AD88E75D79F80082A68";
    attribute INIT_36 of inst : label is "4CC089045A6F3F571A5CAF77C68B4C50A2B8794335CD68E21031620037A08000";
    attribute INIT_37 of inst : label is "E1A17624BC10D70870EB06D903AC1B4B9D47E20AA2A4C948540B8A16ACE7EC51";
    attribute INIT_38 of inst : label is "21E81CD800603482CBA06DDB7C773A37775C23FBC39B06CEC782D412EF29C418";
    attribute INIT_39 of inst : label is "50451411450450411410040000E1E28C4234DB8B6FC37E20102061B260C78931";
    attribute INIT_3A of inst : label is "82C0C16060B030583EDDFF6FC780000140415051511454455510554415510154";
    attribute INIT_3B of inst : label is "4AFB0092267A0C0447C63635C5A2E9C5D74E2EFA717411B40F0D92E724400A01";
    attribute INIT_3C of inst : label is "5284F427A58E52C01D45CF4BBA5457B2F390E21CA0E21D28552392159EC159A7";
    attribute INIT_3D of inst : label is "D5E2880C5B04820521AD69A23C16B8AC89801535AD0C59E7B86A761603DC9873";
    attribute INIT_3E of inst : label is "7DF7DFFFECD9FF3356E7FBBEFFBFDFDFBB77FF36DB7ACB5BF766DFF366DB7DFF";
    attribute INIT_3F of inst : label is "102DD09AB6EF565D09AB2EEADBAFDE7DF7FEFF247F0C7F3EFBEFFFF6EDFEB9FE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "7FBEBD7E9BF554001D4BB01FC02E22ACEBB89900AF3FBDD700000000000A6AFC";
    attribute INIT_01 of inst : label is "D948B650976AEA76CAF46E4D5D4FA83F098A0A320CEFAE4D5B7ADEFDF41FD6FA";
    attribute INIT_02 of inst : label is "6E259F86DC657E2CECD8668ACFC12216D9FC65ADA8E4B2D33691065A2F2B4422";
    attribute INIT_03 of inst : label is "341340F91CA739CA065418C6299C6FFF0AB634AB6DE0A84A322A93942B72DFCC";
    attribute INIT_04 of inst : label is "1026BFBF29CBCE9BB2F512FFCA8506CCD796E1BC05B60BC07132E3E0B8881805";
    attribute INIT_05 of inst : label is "0F310546046012782124B0404E0C186C4009E4C8890D1FD60A04028944A033F5";
    attribute INIT_06 of inst : label is "9E753A267F3408B2522914C845A2C3ED1022C3A711D4AE142D04C906D94D9264";
    attribute INIT_07 of inst : label is "55554554555553430266409E81994F473CFFA9DFEA4486397CB2432C05CF4A99";
    attribute INIT_08 of inst : label is "C255551551555555554554555555555155155555555455455555555515515555";
    attribute INIT_09 of inst : label is "98002C4EC3D1D34AE009E04FB8036201B2678CAAFB1EF4FFC805A2C5070469AF";
    attribute INIT_0A of inst : label is "6103A2F1F7141AD4CDA9EC07EE6A0E6F9155D45575165941018C784C3F4C260F";
    attribute INIT_0B of inst : label is "61AE01CBDAA1B2C1854CDAA5E9CBDEA397A9AB19532D3AA080196D44089B39AC";
    attribute INIT_0C of inst : label is "34297541176AFD011D6C16B8B2CB3E2FFCB2FF7F7C7DF9F7E7DFBA0CB7734000";
    attribute INIT_0D of inst : label is "CFBF9C09B57780000080B676B6B68E9729100865522C96CA6FDAF6785B9BF90A";
    attribute INIT_0E of inst : label is "FE75AB517B178920A909FACA0012DC6557A1501F20302045003D080430204C55";
    attribute INIT_0F of inst : label is "61E110F8E673391C95DD7FD37DF97AEBBD4BEDC36F183768F0DCA01E7483D41C";
    attribute INIT_10 of inst : label is "2CF2CF2CB6EB4FCFEFF3CFEBB769FBD6AEEB6E2F7F77DFFE6FFFA7D0EF81EFE2";
    attribute INIT_11 of inst : label is "F6339F7DF7CF3CF3FF2FB6DBFDB2CB29B2D2F1E5D67967967B6564FEC0BCBADF";
    attribute INIT_12 of inst : label is "B6EB5F73FCCF79E79EFBEBBFFB75965DE5A69A797FC92B466CC6869F77876F19";
    attribute INIT_13 of inst : label is "61801DF632BB4EFB7EE9EDB6D96597DF7DD75D4DB6C32CBEFBEEBAEBEFBEEBAE";
    attribute INIT_14 of inst : label is "3109281818C399018318733419061C05A2D3618C31A8686E8485DC62D7F6C2D8";
    attribute INIT_15 of inst : label is "12E2056C02B016936506330B22DA180C166030A0C3E1C0C0C61CC34318E0C187";
    attribute INIT_16 of inst : label is "C53C20CFB19C2A4031020C02B25C0BA5C18508C1255702BAEBAA135FFBF7F54A";
    attribute INIT_17 of inst : label is "653590890586E7422CAADCE6162C4E3CFEA97D9FA13BF80B6E0BC0ECE6D81F08";
    attribute INIT_18 of inst : label is "771FA975CFDEEF3F99C7BC7EAEF9DFEA74D1467FBD7379EBF3D147D5ECFAFAC1";
    attribute INIT_19 of inst : label is "18E266EFC6388721B827F5DDE20D7E953FC1525CFDEEE39C29948BD1D95DFFEA";
    attribute INIT_1A of inst : label is "F94FBD2DC7E8C5200485917F0A45B00E225458883AA734714734716730128200";
    attribute INIT_1B of inst : label is "E3B1623B28B69180740CFB19C14E6353F30C7294295B7E0A0B6312328C611341";
    attribute INIT_1C of inst : label is "E8A76D868A22244983110384F77965F5A05839F8A196F9305179AC0296C86BFA";
    attribute INIT_1D of inst : label is "8B5C6ECB25DC766193BDD5C009F18CB4E4CC626E64DC89B9937226E64D026B86";
    attribute INIT_1E of inst : label is "FB50AA0FD8A0A6DD19EEFD5CCB9492A914E29608233E993007603A3834A66FE7";
    attribute INIT_1F of inst : label is "6C9EA85A4DDD493E85A49FE93748F4DBB2AA4AF56A5492FDE937D5A9526A49DD";
    attribute INIT_20 of inst : label is "B239043DB50263C48640D51A8DB9D6119C56C0E11BA0D693290678CCC8198F0D";
    attribute INIT_21 of inst : label is "10457E0FE7A058E105404DF54022C3D740FF588E75648C7C13908E75018EA06D";
    attribute INIT_22 of inst : label is "30E5967B5DD98D594B63FC6D9B507BDEF792119FFFFFE5EFBE89C1191C13509E";
    attribute INIT_23 of inst : label is "4F58D53A0F6B2D9A9F1AA78D65AB058D59EC1C9726D5C427666CF6864B936AE2";
    attribute INIT_24 of inst : label is "B9F137215373A9B954DCEA6E55373AC6A9D65A7A9F1A09A946B9508E09A99ACB";
    attribute INIT_25 of inst : label is "04407BF5510187D02842052840A308148BA53685C75FEDF7DE0BD1FB7C632564";
    attribute INIT_26 of inst : label is "F90495882B27443FAAF948BDDD075DF440157B7DDB1A2BFAA7DF4286C8458BB1";
    attribute INIT_27 of inst : label is "D5BC0171F3C486CEB22B3D62EEEFC7407502E074B3B57EEAB53552EBAAA11C82";
    attribute INIT_28 of inst : label is "EDAB9FB00A421136E3A9303105A857DDC0290815641906408910450811B3F8FF";
    attribute INIT_29 of inst : label is "75D6E496B412D04901A0120B5A0AAA1120EB2D200050EE891B6BCA220164C3A6";
    attribute INIT_2A of inst : label is "210D8AB485F49B42C920A01BA614F2FC421B15154009564A414905AD01559090";
    attribute INIT_2B of inst : label is "0905C50FD62900F6AAB08815A0034116028295429078C901B941940045075017";
    attribute INIT_2C of inst : label is "3F7DD9E4572917AE97AC8920AC9AD701206A2BD0926D3CF3037D4ED502136278";
    attribute INIT_2D of inst : label is "45B7784DB775852A630A5191952230522693194E336524F499C65A1F43254D56";
    attribute INIT_2E of inst : label is "D06C1B028E08845122C1125F527BE960BCDFABC812F8415238E97F48297C9D8A";
    attribute INIT_2F of inst : label is "0AAA0AAA0000ECD131999D81AB3D19B2E1FC02B43C1880DEEEA44924804A6232";
    attribute INIT_30 of inst : label is "AA82AA8AAABAAAA0AAA2AAAFFFFFDFF7FFFFFFFFF7FF7FFFE02A8AAA8AAA0AAA";
    attribute INIT_31 of inst : label is "2AAAAAAAAAAAE3B6D147DB67988FB131B9F926B3E5DCF75E9D887F7C5827A86A";
    attribute INIT_32 of inst : label is "926631969C0F4CB649F189E265AA010802514C14260A2445684881802083DD04";
    attribute INIT_33 of inst : label is "E0E449E9EC2619E13C090CD70C090915F02050080000F5E9E765FD7EBD7DC249";
    attribute INIT_34 of inst : label is "A8BCE1E09155A0B501A003C1289809480961C4280662D678B5BAE1C3CB82304C";
    attribute INIT_35 of inst : label is "C64BBA7B5BE440A7BB36257060EE0263BAB0B3E6D24C627270D002D2C38000B8";
    attribute INIT_36 of inst : label is "B940038209E52580D8E3797C366337243EE045D7763143C5FC0E600BC50C1B7B";
    attribute INIT_37 of inst : label is "B323F428FF00959007944802065120172190000C812F62E2309090DE20039400";
    attribute INIT_38 of inst : label is "85019287FC3FC52805048FD012771857F5C96B86A6ACFA6BBA090499AE2B8032";
    attribute INIT_39 of inst : label is "EFB0EEB82EFB0EEA82EFF000018096BF4002406EA48C2000C2201965DB5A540D";
    attribute INIT_3A of inst : label is "984DC42266137108826299BC20615554BFBC3EEB0AEF83EEB0EEB83EFB0EEBC2";
    attribute INIT_3B of inst : label is "3C9C231A54600FD7098E6C14CC082EDDF957FECBB77F02FFAEECC3971BE6CB99";
    attribute INIT_3C of inst : label is "835FDAFFC04833B06FDC4E089C1113CA7B82FDDE82BDDB0FAC1FC8D5A9C3EDA1";
    attribute INIT_3D of inst : label is "A382205480200351EBE14804221307AA0961553D2F5D7EF770A4D81D82AEC4C1";
    attribute INIT_3E of inst : label is "6596D96597DF2BB9F5F33FBFC4C2EFF9DBE5BFF4DBC7A2F7BB7BBB32569B6F4D";
    attribute INIT_3F of inst : label is "FC8DF39BB6FD76DF39BB6FEEDBDE5965B6596576CA4E5D36DB6DB6D248FE29F9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "DA29D1E5AF9E0A6D0F3E0A8896A47E7B28E52F5533A654CAAA0000000024F148";
    attribute INIT_01 of inst : label is "F1D8ECBB8A9613AAB549E3B8C475E5AAFE555865733092EF25184604324A4219";
    attribute INIT_02 of inst : label is "83FFE0FF07DF83FF7F03BDFF783FFEFBEF03CFD7FFBF7FF5EB3AED119AEEC7F3";
    attribute INIT_03 of inst : label is "FBADDD06EB5AD6B5BDFBFF7FDEFFF800FFEFFFFDDF0E03FFFDFDAF3DFC1FF07F";
    attribute INIT_04 of inst : label is "75EB7AD6B5AC552E2FCDF448BF7FFBFFB8FFBFE1FEFDF6FBBEF77C1FDF72E77E";
    attribute INIT_05 of inst : label is "3C7C935F7D6B9EDC313DF876B5AF5ECEB3EA8DB6FADED49D8EC773B9F85B5527";
    attribute INIT_06 of inst : label is "1DCB53EAA459B2EE773B1D8FE7F590CB0FEB9C5C65A66D36B37DEB8FB8DFD4FB";
    attribute INIT_07 of inst : label is "FFFFEFFEFFBFB7DDF9FC53B5373D5B9876ED76A24F57E10760EE7F59F2308662";
    attribute INIT_08 of inst : label is "AFFFFFBFFBFEFEFFFFEFFEFFBFBFFFFBFFBFEFEFFFFEFFEFFBFBFFFFBFFBFEFE";
    attribute INIT_09 of inst : label is "D576C9982AAA0ADC4AF7DD9A256CD5D66DDC9DCF5684FBA0B3BBFBE2DC3963AA";
    attribute INIT_0A of inst : label is "63676FE52276BDFB9DF3DFD9DFFDB1D77B6DBFFBFDF7DBFB692A284F0BA42794";
    attribute INIT_0B of inst : label is "0B5D9ADE9FD3B783D7B15F2F5ADE9BD7BD6CF573E7707FDDA7FA8F8D6DE57FCA";
    attribute INIT_0C of inst : label is "FB739978D6A7529ED92BB83BCF3CCEF353CF2AAA8ACFDF3B74BD6DE3EBFFBD55";
    attribute INIT_0D of inst : label is "9DCCE2076FDB14F554544B3B4B033FD3BB1D9E8E771E5DCFCC2F41746C5416FC";
    attribute INIT_0E of inst : label is "DCEEDF74E93C8F9DCF77AD679DFA70CF119D269B9A97BFB875B6EF8917BFB3CB";
    attribute INIT_0F of inst : label is "3F3EFDE0532994CA7FCFC58CE9B0E8CF363F567779BD3C59D0F1F7BDE72F67B9";
    attribute INIT_10 of inst : label is "000000002B54020824C924001A6480066666EEEEEE666666EE66E6EBF6FBFEFC";
    attribute INIT_11 of inst : label is "6548280080082002082082082002082AD50001001040001001011A2000000000";
    attribute INIT_12 of inst : label is "2B540202A4004100004104104004104004000056A8041CDCE9D334CE397DFDDB";
    attribute INIT_13 of inst : label is "90F6D4A8218DAA4D000000100004000104004120020800820800820020800820";
    attribute INIT_14 of inst : label is "C997F5D5AF6AE49575ED5CA9D5EB57D6D92DB967F057858751DA2275294D5DA3";
    attribute INIT_15 of inst : label is "24CC32B95925DEE45755CC9789AB44E94413A64ABF118EAD7B5721A9CE8EBAD5";
    attribute INIT_16 of inst : label is "39C73E85410FA5DADE94AB554DAFD59E157BE6BC4F3C5550414568ABFF8AEF95";
    attribute INIT_17 of inst : label is "D07B9FCEA7D35E63BE316B99489C4E41F00DE2272938E6C5BF3F33C127DFBCEB";
    attribute INIT_18 of inst : label is "A62B6FE3B64D3CF1BE8AD8AC560AA1C7A3639EACD8EEE77795639E4AD6C1C3A9";
    attribute INIT_19 of inst : label is "444689B62917CA0BBF8EDAA6C5B7B57AF6BBAF3B64D34758BB1D874984AC21C7";
    attribute INIT_1A of inst : label is "D59F5AB716D3BD1AF73FBDEBAEC2CAFFEAAF05EA774B60B60B60B6263C9E4300";
    attribute INIT_1B of inst : label is "FF5C92E79309AA52F56DB2A41FFBFCFECCF7CDFFFFEFC0E077DEFFDF77F8DD83";
    attribute INIT_1C of inst : label is "BFFEFBFD82208276FDA48D3BAB26FBA2CD4ACADB3A8B8CC19782273F6F9A84BF";
    attribute INIT_1D of inst : label is "32BB153319B9E16B6B5B31AABFBFFF5BFFFFFFF79FEF3FDE7FBCFF79FE0FF77B";
    attribute INIT_1E of inst : label is "CDADC2CF66BCDB6AE7376A8DF9DD873B8B185DCFEC41A7CAD65674F1F4CCCCCB";
    attribute INIT_1F of inst : label is "7FFB56E7EBA4FD756E7EBA5FAE91E56C58F73387B72FD5EB9FE6BEDCBF57F9AE";
    attribute INIT_20 of inst : label is "EFDFBFF7EFBEDF7F7BF73FFF7ED79F8C63896FDFED7BDC36BD60E7631AA5F472";
    attribute INIT_21 of inst : label is "DE3BB5B50E7B039BB09A33A2FDFB9F69BF80E7FDDBBF77E63EEFFDDBFEFDDFBB";
    attribute INIT_22 of inst : label is "FFDFEDEFF6F6FBF7FDFC07F76EF70000007FFF6000001800007B3FFFF2050E9B";
    attribute INIT_23 of inst : label is "BE7FE7F3FBCFD6F3FBFCFEF9FADE3F7FB7BFF7EDFBBF7BF8FBDBDFFBF6FDDFBD";
    attribute INIT_24 of inst : label is "C08FFBC07FBC3FDE1FEF0FF787FBC3FF3F9FADF3FBFC7F3E7FDE1FFC7F3F73F5";
    attribute INIT_25 of inst : label is "7F566C923DEB69281F2DB3E5A07CB699CE4ECDA5FFF9B6DB6C97EC23DFBFFFFB";
    attribute INIT_26 of inst : label is "91C7BC8E792E15DDF39DCA74F0F6B14E4F1E6DA6B6F5FD6DDA6D8CAB6E5FFDEC";
    attribute INIT_27 of inst : label is "6B3D74CEFFD72BFDFABCE09D9CC9FFFB3E9F9EC9FE2DC88CECE5C8B971FA8EF7";
    attribute INIT_28 of inst : label is "CF5E69EB77F58CCBFFF3FF85CB7EBE4A8DDFD67BF5B17C77EA5CBFD7666A55B9";
    attribute INIT_29 of inst : label is "CBAE777547659D95DD3BABB0B3BBDFACFD97D1CBDBBFD4B3CEC6A7CB97F5B65B";
    attribute INIT_2A of inst : label is "96D6DD427BA765FDB1EE2CAD7EF99F592DADBABA7BA7BF57EF15DC59DDEFD67E";
    attribute INIT_2B of inst : label is "1BD6F4FD60A13C6E3CFA08A9BAD4A62F52A31FA973BEB1EED6FDC517F146851A";
    attribute INIT_2C of inst : label is "C0EB8B7FF3B94E8CF77EAF39E4AE5C844B93F743399B7FF4BFB63D6FF3D7DD72";
    attribute INIT_2D of inst : label is "FFDBDFB7DBDF7FF7BFFFEEFFEFDFFC7FFBFDFFFBFFD7FB9FE77FFDFBFFFBBFB9";
    attribute INIT_2E of inst : label is "164D2DD5549D692C8A54EDBA2DD5B6FEE33AB6176DD1972EBFFFCDB7F7EBF7FF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFE2BF7D5557EFF6F7FEFF7F02B43AA662E57A74E57397399CA29B";
    attribute INIT_30 of inst : label is "AA80A80AAABAAAA82AA2AAAEAAAA0AA0AAABAAAA82A82AAAF1147FFFFFFFFFFF";
    attribute INIT_31 of inst : label is "2AAAAAAAAAAAEA2AFB4F80AA1947D40D42FC27BBFEA1FA1EC984790214A7DA6A";
    attribute INIT_32 of inst : label is "7FFFFFEB7FFBFF5BFFBFFFBFFADFFFFFFFFFFFFFFD4C3B7B34767ED4C096F3EA";
    attribute INIT_33 of inst : label is "F5C543E78C1FEAC9AF9D19E6A258860EC2AA8B061D57531112728882A80ABFFF";
    attribute INIT_34 of inst : label is "DCDEF514FCA300D8FA380FF1A7E3453768CE73E7535D59D75E57EE47E08FF6E8";
    attribute INIT_35 of inst : label is "FFC0BF5FA1FBAC4E66E733C41F73E993E7D5E6BEF1BFFCE34FE7CB0F32DAAADC";
    attribute INIT_36 of inst : label is "6BFA56AAC3E69E25A3EED29D68F76E3174CA94BCE9A3867EAE83557FFFFBEDFF";
    attribute INIT_37 of inst : label is "E4F08B4EE3B26F3CD57953D27DE54F13A042D4AC176058C9505EDC4003473F1E";
    attribute INIT_38 of inst : label is "7BFEFDF803E0E5DE0BF776EBDA9423BB9EE7AE5FDB17DDF9D31C99D5797774CF";
    attribute INIT_39 of inst : label is "EAFFBABFEEAFFBABFEEBFFFFFFEACE94ABC2006C03781BD53D7A67FB7EEFFBFF";
    attribute INIT_3A of inst : label is "7CBF3E5F1F2FCF97ECBB66D7EFAFFFFFBFEFEBABFBEAFEFAFFFEBFFFAFFFEBBE";
    attribute INIT_3B of inst : label is "3F2C515FF693CFE3D9FD1E52FEF43C2A69E1534F0A9A9FB13C5375BCAD17F21C";
    attribute INIT_3C of inst : label is "19C88E442C58EB342C3AEC566367C5A0B5D3C8AD2BC8ACB13FC912F9EB4A912F";
    attribute INIT_3D of inst : label is "000072CA583DE8B59EC835374ADFF779DCFDEEF8FB96AD7FCD86BEDBF23EF78E";
    attribute INIT_3E of inst : label is "00104100056A80413B4028D000890C80105A495B6D00000002024905A36DA000";
    attribute INIT_3F of inst : label is "1F64D18B966B72CD18B966AE59D001040041015AA81000820800820A34400040";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "BFF9DF7D7DF777570BF7B01FC03F2FF6FFBEDBFFF3BBFF7F00000000009B76BC";
    attribute INIT_01 of inst : label is "F77FBFD5A7FBF97DEFFF87EE7F2FB8979B9FFD9FFBBFD0B3AFEEFBBF5C17F7AF";
    attribute INIT_02 of inst : label is "FCFFFF3FF9FFFCFFFFFC7FFCFFCFFF1FFFFCF7EF3FFFE7FBF7DDF4FEBEFADD7E";
    attribute INIT_03 of inst : label is "FC5FE2FF1CE739CE5FFC1CE7FFFE7FFFF3FFFCFFFFF1FC7FFE3FDFDE3FE7FF9F";
    attribute INIT_04 of inst : label is "F9236B5A96B56EDBAFDF9BF7BEE7E7FFFF3FFFFE3FFE0FFC7FF8FFE7FF8F1CBF";
    attribute INIT_05 of inst : label is "4499A8C7443B35CD65EBDAC5FF9F3E7ED50DE5CD97BFEB77BAFD7EFF5FA01AFD";
    attribute INIT_06 of inst : label is "DDB7BF777BB4A9AFD7EFF7FAFDFEE7EFE226F72711FCDD5C3644CBEEBEEFD9FD";
    attribute INIT_07 of inst : label is "FFFFFFFFFFFFFFFFC46369DFD798FFEF7E7BC5E5FAFD6BFEFDAFDFEE88EBFE6D";
    attribute INIT_08 of inst : label is "CEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_09 of inst : label is "9C00EDD169FA3EDCA1BF7BFFF801FC00FFEF86DBAFCAFFFB780DE6AD3704D99F";
    attribute INIT_0A of inst : label is "F302E4F92E6E24DC41BA4B03D26E0BDFF9E79F79E79E79F70D86DC6F1F6E379F";
    attribute INIT_0B of inst : label is "1F3B4113DEE134EA4DC49B89F913DAE027E3BA0B744F7EE0AA136DD57BE77BEC";
    attribute INIT_0C of inst : label is "BDFBBDB99EB4DA8311203D797DF73E5E737DFFFFFCFDFBF7EFDF84C4C3E790C1";
    attribute INIT_0D of inst : label is "BDDF592D7AFF83280181A44BEBD7DEBE6FF7FFA7D6C9B7BADF93F3FCFAFFBB7F";
    attribute INIT_0E of inst : label is "FD7EF7DE7F77F975FADDFF904FF79E7BDEF1DB9E6038606BC03F185EF8606F6B";
    attribute INIT_0F of inst : label is "6FEF34FBDFEFF7FBF1F87BD37DFA7EFBF79BF7DFCFFE677FDD9DBD9E7DEF7DFA";
    attribute INIT_10 of inst : label is "FF7FF7FF5CFBFEF75EBFFFFFE7DFFFFF7777FFFF77FF7FFF77777F74F3E9FFE7";
    attribute INIT_11 of inst : label is "DAF7DFDF7DF7FFFFFFFFFFFFDF7DF7D53AFBBFFFFFFFFFFFFFFEA757F9FF7FF7";
    attribute INIT_12 of inst : label is "D4EBECFD9FFFBFFBFFBEFFEFBEFBEFBEFFEFBEB9F5D9EFA75EE6DBFAEBCF7F6C";
    attribute INIT_13 of inst : label is "B9F0066BFE537DFBD7FFFFFFBFFFEFBEFFEFBFFF7DFFDF7DFFFF7FFFDFFFF7FF";
    attribute INIT_14 of inst : label is "323BFBFCB38D19FFD671A33FFE2C6809269247BFCD3BF83CF387F77FFFE7FCFF";
    attribute INIT_15 of inst : label is "3FB7824FFBFDE677FFFFF339FFFCF1FDFBC7F4FFFCE39FE59C68DA7671BFEB1A";
    attribute INIT_16 of inst : label is "FF7FEB66D7BE3B2E21DFFF03F3FC1FBF7FE7DFFF6DF707FFFFFE1E77557DDAF4";
    attribute INIT_17 of inst : label is "7FBFF5FAFDFE67DFEBFEDEE423FFFF1FFFEE7CFFFDFBEF132EFBC6E7FFDDDFFF";
    attribute INIT_18 of inst : label is "7FFBBE79F7FFAFBFDD77FFEFBF6DFFDF7CADF77F5FDBFDFDFBADF7F7FFFCFEBF";
    attribute INIT_19 of inst : label is "CFF7BFF7D3FDB5F1FF27FFEFE709FF7AF7E1F69F7FFABB9C6FF7F3F1D37EFFDF";
    attribute INIT_1A of inst : label is "FCEFFF99CFF87A3CCF8FDF7E9BDD20EFFFFDFFB43EEF66F66F66F67FB84E97BF";
    attribute INIT_1B of inst : label is "FFF1ED7BCCFFE106FF8335FFC3FFF3FFF3FFF3FE7F9FFF1F8BFF07FF8FE14A7F";
    attribute INIT_1C of inst : label is "F9FFFFFE7FFFF4CD7C1B27EEFF12EFFDE53A7FBDEB66FA74F7FBBF27F7CCFFFD";
    attribute INIT_1D of inst : label is "BBF697FBFDADB3E1FBFDFDC00FFFCFFFE7CFF3FFE7FFCFFF9FFF3FFE7FF3FFFF";
    attribute INIT_1E of inst : label is "FDF7EDCD7CDCFBFDBDEFFFDEEF37F3EB66F7B7FAFC4566C007353F71766EEC69";
    attribute INIT_1F of inst : label is "7C9FFBF3FFFC7FFFBF3FFFCFFFD4FFEF223E9AF1FE87FE7DCFFFD7FA1FF3FFFE";
    attribute INIT_20 of inst : label is "F3FFC7FFFFC7FFFCFFF8FF9FFD99F5FBDEF482BAD6E6F5976B73FF89F6112686";
    attribute INIT_21 of inst : label is "B2EFFE1FBEFCCFBF076E4DF87FE6B7FF63FFF9FFFFFF8FF9FFF1FFFF9FFFE7FF";
    attribute INIT_22 of inst : label is "F3FFFFFE7FFFFC7FFFF3FFFFFFF839CE739F9F9FFFFFE7FFFF9FCFF9FDD371FE";
    attribute INIT_23 of inst : label is "FF9FF9FCFFF3FFFCFFFF3FFE7FFFC78FFFF9FFFFFFC7FFE7FFFFFCFFFFFFE3FF";
    attribute INIT_24 of inst : label is "FFF1FFFF9FFFCFFFE7FFF3FFF9FFFCFFCFE7FFFCFFFF8FCF9FFFE7FF8FCFFCFF";
    attribute INIT_25 of inst : label is "A66E7FFFDF7B27E4EFE4BDFC93BF92CF63FB34C724912492499BFEBBFE7F3FFF";
    attribute INIT_26 of inst : label is "F77DF7BBEF7F437FBEFB7F3FDF779DFC6337EF2CB5EF8FAFDAFFE7E65AFDB5A1";
    attribute INIT_27 of inst : label is "6AFC037BFFDD6ED93BEFBF77D9D9FFB06736FE7FB62679D997EC7D8FA53BB9BE";
    attribute INIT_28 of inst : label is "FD23EBA51377B136FFD9B6937B4EFBFED44DDEEA7719AE632F37B9DC1F774F7F";
    attribute INIT_29 of inst : label is "7FABCD6FBD6EF5BB5FEB76BFCEB753BB74FE677BA89A76F64CD49BA6F67793FC";
    attribute INIT_2A of inst : label is "F27DCFF1DFFF9B7FFB5ACCDB3FFD9BFDE4FB9FDFD6BEA773FFDB5BEF5FA9DDBA";
    attribute INIT_2B of inst : label is "47A8963542388CEBEFB0AD9FBA81B3AE013391E43AFEFF5B987FD99A6667DB9F";
    attribute INIT_2C of inst : label is "3F7DCDEE5E6FE7EFBE4EFBEFBDFBC7D0F833EBF9EA69BFF5FFFF4FFFFEBF4DD2";
    attribute INIT_2D of inst : label is "E7FFFFCFFFFF9FFFFF3FF1F3FF3FF3FE7FF3F9FFF3FFE7FF9FFE7E7FE7E7CFFE";
    attribute INIT_2E of inst : label is "59551B332CBF86DF21D5ACFFDF7F93CDBCDFDBCD67FCF7DF3FF57C9E7F7CFF3F";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFEAAAA2AAAB81FFFF3FFFFF7C13B415F4FD4BCBBFDECD6CF667B6";
    attribute INIT_30 of inst : label is "FFFFFFFFFFFFFFF7FF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "5555555555557F75FFFFD75FFDDFFFFFFFFFFF75F55D55DFFFD57D555557D5FF";
    attribute INIT_32 of inst : label is "F3E7F9FFFCFFCFFFCFFFCFFE7FFE73CF9E73CF9F3E1BE6EAECCDFE003ACD9FA4";
    attribute INIT_33 of inst : label is "E0E5DDF9FEE7E7F6FBB7DF770C07C7CFF83074EF687FFFF97D755557D7FFC3CF";
    attribute INIT_34 of inst : label is "3F3FE0ED125CFD3701C727FA389BD1CAA770F7F807F7F4BDFD0FF193F727F84E";
    attribute INIT_35 of inst : label is "CFCFFFFF4BF6C0B7BBB8C6707FF9023BFABE587FF24FF77DEF77F6BBD6007D3F";
    attribute INIT_36 of inst : label is "FEE007AE8DFD77A1FDF767BC7F77F76B7EE043FBF67EF7FDAC0F77FFCFFFFFFF";
    attribute INIT_37 of inst : label is "FD61DC2FF700FFE0E499025202640933690980184B405DD958A3A0CE1147AF00";
    attribute INIT_38 of inst : label is "FF9FF3E7FFFFC73381FF9FF7B7EF79BBB7D2F3B6FBCDAF6F2EF64F5F8E7ED05F";
    attribute INIT_39 of inst : label is "AABFAAAFEAABFAABFEABFFFFFFC1ADFFC209257E96D4B6808FF01FFFFFFE7FCF";
    attribute INIT_3A of inst : label is "FF7FFBBDFFDFFEEF5A4691B8CF8FFFFFBFAFEAABFAAAFEAABFEAAFFAABFEAABE";
    attribute INIT_3B of inst : label is "BDA7BBFBB9BD5D5BF9F1381EE254DF6EFEFB77F7DBBF037EAEFEC3670EBBFB9F";
    attribute INIT_3C of inst : label is "E23FB1FD813977FA5F7DDF09981B13CE7FC2F5FF82F5FF06BD9FD4DCEFF27EDF";
    attribute INIT_3D of inst : label is "FFFFC033E67A41B1FDE1CF072191B4BABBF2D7BB7FDFDEFFC1997D3FCE4EE2C8";
    attribute INIT_3E of inst : label is "FFFFFFFFE99B7F5E26FFD13FFF37D1FFEF67FF66DBDF7F7FDDE5FFF26CDB7EEE";
    attribute INIT_3F of inst : label is "4360040C0003800040C000300027FFFBEFBFFE66DFC7CFFDF7DF7DFCCDAF8FDE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
