-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "AFFA9D6DD80586DA1654207BE37F964C49A17FE1254207BE37F964C49A17FCF5";
    attribute INIT_01 of inst : label is "0140521510440413FBFEAD13436381DAF75C0E94BBA506C50662693D75802046";
    attribute INIT_02 of inst : label is "30A2C2058140C9D8DB5BB6E8C1C2C01030A74853410A0A290C42816214C102C4";
    attribute INIT_03 of inst : label is "DCD4AF74AE5F6AFB47BAD9C325E2CFA615D1EB7BDEDBE85B25AED67BBC2A1806";
    attribute INIT_04 of inst : label is "C39D8B180008B9C02A40DAC28AAC4E0AB33941EBB4A2F016025C00546000C495";
    attribute INIT_05 of inst : label is "870F418ABCDB3B7D9BED1E3879AA1EE94812AACD4247D8206436A486E106E103";
    attribute INIT_06 of inst : label is "F974479CCFAA88AD6269D1416321A55449E4D04F66022A8488B01EBBDD543416";
    attribute INIT_07 of inst : label is "1E5BD268AB211DE67223A87F5DC355795FF3FDF0D0C09995BC20A16764606561";
    attribute INIT_08 of inst : label is "CFDCDC473333FF4FC1471A177515B690D553522743555C6F997EF2673FDE8881";
    attribute INIT_09 of inst : label is "139B59F7578FEBF9767AD2FD9F0E5FC9E2657302F454573E233E5F63966AE2D9";
    attribute INIT_0A of inst : label is "E68E6EEDCFEF91F37A6B2D04765358F7E3480FA22C74284141477CAC20D52B96";
    attribute INIT_0B of inst : label is "7A0E6FFF0730A4A7E8DF0D022A2A606F7FD99B0769D9A776958F29586683FF23";
    attribute INIT_0C of inst : label is "8ECECAC62DA6151AEB0CCE8620577F6E7F79AF61E4EDF5A4EE5FB73FBC5EF22F";
    attribute INIT_0D of inst : label is "38105C72A0250A39692C3B7BD7FC69CA2772A4650DE105771E6354DE2B2B2D37";
    attribute INIT_0E of inst : label is "ABA7B84AAAAD1134E9D6E6E8880C7BDA8B7D8A63F2E4AA311548284501CE6EEC";
    attribute INIT_0F of inst : label is "3BEEB6137B9A4D91515951113FB3A6A55E0E7377AFB464C1E86BA85D734F0492";
    attribute INIT_10 of inst : label is "05C0ED7FBF5BECB121663E7C2DB35159515136A22D535565F2F407C9BB046351";
    attribute INIT_11 of inst : label is "0670DE036C8D7B0208E0128008871FEFC42781036C841C2307B17FB00049BE02";
    attribute INIT_12 of inst : label is "6A12C431A8E6A52C4504BBDC509F6B80301FE11002407F000DB50D0708059402";
    attribute INIT_13 of inst : label is "01084410A81DD813006FC1807D07007C025A5DE818C3F758D4210C4B1884352D";
    attribute INIT_14 of inst : label is "20009D528684AABA635C12492409058C1700D8A860B027C78683A416002000BE";
    attribute INIT_15 of inst : label is "4002123676A06681431ABD88004201E840EC400A81909294553A1F80004086A1";
    attribute INIT_16 of inst : label is "80EE1270880108010A0090D0595698D78006000C243B10D64BE4C0001090D028";
    attribute INIT_17 of inst : label is "898CC8E5984E6FE6010085CA43843FDC4E4C0183005384021883EFCA81AB46F0";
    attribute INIT_18 of inst : label is "57E682A7F1CD39FBFC6FF4DB48B44A55937CEB760CBD00B0F71B18001820641C";
    attribute INIT_19 of inst : label is "C1CBEF828BC1133DCE72B27B5C10052AA2D82108610897845AA552D556AB5555";
    attribute INIT_1A of inst : label is "E4878144F2F0D29EFAC83F0C208ED40409102410A954E2F86348014F6E037086";
    attribute INIT_1B of inst : label is "77FC5908D21806B41D1006A9D43096BDA78874484C2DD09833F185815F9D2738";
    attribute INIT_1C of inst : label is "8A957E097511C0928949E010969E9255DA0363B842A0AB9ECE7DB52078860442";
    attribute INIT_1D of inst : label is "26A398BDF4A489124295C909AE3C4C04FCD656CAB25295A72AF835F5453F6FF2";
    attribute INIT_1E of inst : label is "9F56E4013C77653131F6622BC9F7A39E17BBC01A8EF086AA22C79AD352341852";
    attribute INIT_1F of inst : label is "84D1CBB5572B229D134ADA2D89D79FB205DF4E786FC0C77248B78CF33CEEF85F";
    attribute INIT_20 of inst : label is "EDEAA6344D6C30C48CCC42080521336220001185093CB29E566295DA1C0EAD12";
    attribute INIT_21 of inst : label is "9515951B3826493B6C2FE8102E0936864C406484D9246F4969D0593F6D93A736";
    attribute INIT_22 of inst : label is "795BCF39E6283E4DD9C9C0139B1EF556FB921E9E87127FD098B004805069E905";
    attribute INIT_23 of inst : label is "FD69D48D59E47C69ACEE0A7A59F5454516CA7881CE6EEC8221D5ED5645159F25";
    attribute INIT_24 of inst : label is "EF3EE5C4DA7DE12A75F44E882F544515058E834058B202A8DAC517A0F650F2B5";
    attribute INIT_25 of inst : label is "6F3CF3709624BD9325B6A1023A02A16967FB02AF958F868D316215004708284A";
    attribute INIT_26 of inst : label is "136010E81565A101A19B428AA88FD3A6FD3A62D5D0204351995D55738A62E64D";
    attribute INIT_27 of inst : label is "8B73FBC7AE79549FDB2E37791AC9B66839720DA27586E01B11813D78D08A0F58";
    attribute INIT_28 of inst : label is "FFEAFA0007FFAA00001FFF57EAF27ABF7AAA08028B803BC71D04196403C323E5";
    attribute INIT_29 of inst : label is "50540AF555550ABFFFFFFFFFFE57E0000000101FFEAD4AF201FFF52AAF20157F";
    attribute INIT_2A of inst : label is "7F044444444441B6AEB7AE005140438E44400401984504115114257C61010721";
    attribute INIT_2B of inst : label is "1FFFD00002FEFEAEAFBB3FBEF3DD98F9CEBAA6EFF3F7E7F9C035B580C763FD07";
    attribute INIT_2C of inst : label is "9249289010060000000100890492492492492890100600000003066000000000";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "500F179801DA5DB3791CBC809B7A5D990044C03701CBC809B7A5D990044C03E3";
    attribute INIT_01 of inst : label is "FFFDEFF77B7E9044361EDF5A30BC7647E9A3B23D02104BC890950D8252D2E4C8";
    attribute INIT_02 of inst : label is "72FDC96F926CC32D65EE491CD1D1220502C1C492099B2C6F38EECDC677982F0C";
    attribute INIT_03 of inst : label is "BC91805DCBEFF77FA28F957A6FF1870D6CF6B28C034504A493784D2698B6B92D";
    attribute INIT_04 of inst : label is "D742D4514AE6251D8D292F161417959DC0003A94427163962BACA523B4E56983";
    attribute INIT_05 of inst : label is "DEF5BD1349DCD8A2E51569972EFD840CB526CBBC9C9A23D5114BCBD10ED10AD9";
    attribute INIT_06 of inst : label is "C610A8003831111EE4D2AA92E5FB489AB24E3A9695D5F1F97DDFA944E6BA8AA1";
    attribute INIT_07 of inst : label is "2197A4B1526FEA10004CF2A4A2020053954590FBF7F92EE2A96AFBB498AA816C";
    attribute INIT_08 of inst : label is "B2CA33BACECEBE96AF887461D2A7DD276098746A9D8230F55FC369C20067F358";
    attribute INIT_09 of inst : label is "A574F258E87035D6B9C78FF3AB5DEA9C55D8D6A440988ACA4CC8FE9D249D550E";
    attribute INIT_0A of inst : label is "2B37955975BFFC1CB6B77BE8CCAD873BF4975515C9DF5DEAEAEEEB4B55BAD2EB";
    attribute INIT_0B of inst : label is "F6FAB593E9D549DA810FBF74CC44D4D2F12526E9D2A7488D2AF57B8EAF356251";
    attribute INIT_0C of inst : label is "9117777B50F4A224A4C9851DDA9ACACBADFF75F64ABFBE8DBCF2E5D6FFB5A55E";
    attribute INIT_0D of inst : label is "5365000E64DA5C52B643DCBF632492271007200A52CA528E600E196B544DCA42";
    attribute INIT_0E of inst : label is "4D7AC2931556EE6FDEAF012B7750B5645C8A77B097B9754FBBFF5DBAEA001129";
    attribute INIT_0F of inst : label is "5BEE66B5DE239EE6A26E22A6104C4DF275500089DB87A012023E9E8711D05944";
    attribute INIT_10 of inst : label is "510F86CB61329966B7915394FC68A26E2A66EC59523D824F6789A8004460B486";
    attribute INIT_11 of inst : label is "9C0E334E52508850C14D211CB2B5C5A03900573E1A1525869672046D296C68D8";
    attribute INIT_12 of inst : label is "BDAF29DEF3494E7692CB0FB12D69CE1486CCAB4949E900A7394B39B1AF234A9F";
    attribute INIT_13 of inst : label is "52521AC96B41A487E91B0FD4EF33B900E4BDE13DA5680FB92B4AF2BDAD295AD2";
    attribute INIT_14 of inst : label is "B5A7EAE1692F1329DDA0ACB25C9B52D88D971392C464989C5CD8B68C52E5E600";
    attribute INIT_15 of inst : label is "8E59295DCB4E14D694EFF2D1CB252535AC168E4554452EA97685201C95AC1CD7";
    attribute INIT_16 of inst : label is "FF00A5DA53B5A4E5BB596D252E64776869C9A73095ACE54920000A5AC94A1AD2";
    attribute INIT_17 of inst : label is "677623204B95840872F64D2D5AD98B639000A435E52828E5BDE79055AE53F907";
    attribute INIT_18 of inst : label is "9C018360F20B41B0036F49C5AFC9A56308D215C9CD504EB5D8E5A69C83D51161";
    attribute INIT_19 of inst : label is "69D4445D601CFDC89CE724B4715A5BC4C4274E52F7FD29C06B2994E667339999";
    attribute INIT_1A of inst : label is "D50294EB27EF2D60F9FDB2514A51796A97BE5EA976E95752BCB394A2F0E88569";
    attribute INIT_1B of inst : label is "32CAEE99A4572D22476B3FF8EF4BA0F55AB5AF75DA97EBB5BAEB523A03DE04FA";
    attribute INIT_1C of inst : label is "B659F929767779DBAF83DFC9DB3F4488ACD52BBAB4F6F1311FFE46439148E4A7";
    attribute INIT_1D of inst : label is "8075E8FF5F8A202FBD4A0065958191526804CA385A8B0641B3E4ADCBDB3C9CED";
    attribute INIT_1E of inst : label is "2AA417EF8577084EAD0D1C448C6D8A45E40476EC7449F0CDDC958E002B428BC8";
    attribute INIT_1F of inst : label is "5919D5F26EF24FEA6B29B47212AE2A1EBFC2628A90EB5774DD01E86D66810DE4";
    attribute INIT_20 of inst : label is "012376A2B209861D3031E6D2DED6368452F0B6169449592DE4AB07A1F59440AB";
    attribute INIT_21 of inst : label is "E2A6EAA4BD19966CB388B6E494D78BCAB214AB6926590040132532499658B0C9";
    attribute INIT_22 of inst : label is "B28269E29155400222129B66402D48B9142D84C72A731FCE7206D93CEC9432D6";
    attribute INIT_23 of inst : label is "15C6FDF2AE3AB326C584A5A093E98888A87195EA00112930D2831A659A26ECDA";
    attribute INIT_24 of inst : label is "11C9CB1313D2EB41A7F09567441888B8E895359A8D2CBC856848BA1D2C3B6507";
    attribute INIT_25 of inst : label is "4BAE8BF5A0E8FC655C9076B0534B5B9A4E46D7727A532BD6DB8F32B59597FFA5";
    attribute INIT_26 of inst : label is "AFAF5C2A8E684C9649B42B13311178B0578B1CB90ED60C62EEA2665AD08DCAE0";
    attribute INIT_27 of inst : label is "365D6FF974B2F9B2F4C95B8FECB7ECD54E7B5044A9A154A069322A911B9C1EEA";
    attribute INIT_28 of inst : label is "FABF9AAA07EAAA0002BFFEAFFF8AAAA6C6084251BF64A4DF7EC931D8A627A4CF";
    attribute INIT_29 of inst : label is "BAEFC80666664908445111444503A7ECFB3E8AAAFFF81F8AABFFFFD5F8AABFFF";
    attribute INIT_2A of inst : label is "3C5777777777740980199151A6FBBBFBDB3BF3AEF6BB6FAEA6CD6ACBB67670E5";
    attribute INIT_2B of inst : label is "07FF420002EEEFEFEFB9FFBDC0E5555A01ABEEA7FBF741CCDF9F1F3FE73790BD";
    attribute INIT_2C of inst : label is "9A4D3A9C128F000000000809869A69A69A4D3A9C128F0000000F8FF000000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "15050A9550D23E925BC40C1245BA002240007FE52440C1245BA002240007FC21";
    attribute INIT_01 of inst : label is "042B5AE558F5869038C2D74220FC16210DA4B54902204081128D23911430A140";
    attribute INIT_02 of inst : label is "60A980C3014A430B086280A67CF161A70723F9211028008251040408A1104A90";
    attribute INIT_03 of inst : label is "D094A162CFBF9DFCE11FD17247F1E08AEC14881284C02120003C0E170005300A";
    attribute INIT_04 of inst : label is "7720B74472D2840541D80B0ECFC6DC45694ADB811C9A99C98E8A734DE733C8AC";
    attribute INIT_05 of inst : label is "1BF0F4A9580F5C3C38E326CD9AFC2541471A30E96C6841AAAA50D0D406140211";
    attribute INIT_06 of inst : label is "C93974A575199AAF979B38F396CE6EDE1B6E62CF42CF9F0DEF6DB811B0E6A9B7";
    attribute INIT_07 of inst : label is "40FCE4F99BE3B8D294A252F408A8AAD1B543D787938DBBBB9D62A283ECE6C3BA";
    attribute INIT_08 of inst : label is "8E59DAEE307790DB0EC356204335E9B500D356ACD4031C7C029A328841787850";
    attribute INIT_09 of inst : label is "76B6BFEC1EBF8FDEED34E9F53817B8DCCD48C662A8CCCE38676CBFC6928FC5BB";
    attribute INIT_0A of inst : label is "CFD8733FFEFF1B66DCF87C6F370C04EC76DA5CF77FF1410B1B0B0D7DE10D5B1C";
    attribute INIT_0B of inst : label is "9D34FC3C6C276DFE51F474B666668C0805BFFC6C9B366ED9BB5294F5D5970BF7";
    attribute INIT_0C of inst : label is "1BF9D98C5B36B7727FD444C4E2CE38FF77F9B65B7CCBE20FC6FE7FBBFC633E35";
    attribute INIT_0D of inst : label is "5261521AC473163FDD5CEF4F01DC6A89AF7BDEF318B7B429A4AD5DF87FE7736E";
    attribute INIT_0E of inst : label is "67B861D19EDE36337635A96A6E5A9C3CE6DAECB48FFDC5622E7173CF2B52956A";
    attribute INIT_0F of inst : label is "13EE733DFF2B9BB7F73B773B7CD3FC773C5A94AB5A96A12B043758A130509854";
    attribute INIT_10 of inst : label is "3503D2E970381C20A5BD7EDA3E29F73B7737D6E8DF1C076FB7CD2D5255028426";
    attribute INIT_11 of inst : label is "8E8612C74BA8B09082530D0430A45BEF5874150F0B8509E284A46EAB5A1CBA1E";
    attribute INIT_12 of inst : label is "AD2118521108D210800203D801406A8C30FE0600C00840231D251D214B097580";
    attribute INIT_13 of inst : label is "30140200505A282D780B823C751C28406129A084210C04300842948D210A56B5";
    attribute INIT_14 of inst : label is "A521F7FA924D99B85C082024140010070468A880302264441E90C5A4312263A0";
    attribute INIT_15 of inst : label is "86000A5742E78210847B6010C001608420008234AAA9402112F11F8C04282414";
    attribute INIT_16 of inst : label is "9D052152108529202A5052493B36170248412115A521629349EE86020052C210";
    attribute INIT_17 of inst : label is "0170F94DF98F7D3C10B005415218B7F58EE86085210B08617B8708E7DA062803";
    attribute INIT_18 of inst : label is "E40F82E6F92F254000B740A16B416B4380E80C50675043D5C821648431AAAA6A";
    attribute INIT_19 of inst : label is "5CD0F615A8043F7ED6F5F6FA10521366668242B48C2903007C2E1747843D1E1F";
    attribute INIT_1A of inst : label is "C0820C24AFE8AF9552EB2842461058D79A5A6979856D8580A524842C586A0108";
    attribute INIT_1B of inst : label is "4D34B08854A148A49A4A48D30A6A54221C25438510F84A21C096B40B41CE225A";
    attribute INIT_1C of inst : label is "8904042429708E50A2A3A6C0403BF6C155BA2912D691DAB45BD31219E0467B23";
    attribute INIT_1D of inst : label is "A015C8FC76806871CC40BB225528A0D1169580483EC00122081090B6C4821A53";
    attribute INIT_1E of inst : label is "A5B6558B95AA29EDA3853AE7FCB7034C20116E281F7F32E7F7D7CA500B61CAC1";
    attribute INIT_1F of inst : label is "D504F5A40FDF69F71A4A9E589088A5772FCFE679DB8B5226CDB7A5B718044B90";
    attribute INIT_20 of inst : label is "443252B0DB2F90C5A9442A1042109600101C03848D1FEAAFBEEA05C07124A97A";
    attribute INIT_21 of inst : label is "F773BB3109C004A024A1F4E0A6D4EA4F8484F84AA012EE3B854954A004A9F220";
    attribute INIT_22 of inst : label is "DE0B5C71D2616A92AA14086294A7094DB515A4CD4A5B3AB414A218056824841F";
    attribute INIT_23 of inst : label is "D87B08DB34D6FADA00F839D44BFCCCCF2DDE6B4B52956A2014A9A336AF73BE8C";
    attribute INIT_24 of inst : label is "44BD8F8DCC3FCF7EDBFF1D1B7A8CCF2F6F19CEE6F5B56F71B7AF2DC5F78DBC1C";
    attribute INIT_25 of inst : label is "0DF661E5BF437F8743EC90A0924262F12B6B95D8DB5C1C5A22C154A5841CE729";
    attribute INIT_26 of inst : label is "886E5802A808000494B0599B9B9BA9F29A9F3AA512141077FBFB73FBDA818EE5";
    attribute INIT_27 of inst : label is "DFFBBFC4D66F29FB977FE239B1DB0ECD6C02404030296C000AA45852928C0272";
    attribute INIT_28 of inst : label is "57E01254001FD40005400002A0022227031082112C4C20DB6E831090622BCA6F";
    attribute INIT_29 of inst : label is "10054CDDDDDDCD4C44591164457BA80E0380BD5F81FFE0025550155400254A81";
    attribute INIT_2A of inst : label is "105DDDDDDDDDDD4DCC55C52A5921C00425C22C8900648218792B405114DCD15D";
    attribute INIT_2B of inst : label is "81FD0A000155550103B93FBA409C0038001154EFF03741D9C0151500C700F846";
    attribute INIT_2C of inst : label is "65B64D2E1B86000001E1B0D6FB6C92CB65B64D2E1B86000001EFC7FFFF000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "15199CCE0052929012D9A49647FA548944544281259A49647FA5489445442821";
    attribute INIT_01 of inst : label is "3DE739E888D29AC11C051958F446D28EC636947C288BC9EC0F30EB744212046C";
    attribute INIT_02 of inst : label is "52A1EA5AD9022541402892A60C404AA41301C00455338E8A5504A1A8A5504CD2";
    attribute INIT_03 of inst : label is "91708729A6BFDDFEE172C15245F44220F446981605C02020002402010AA4B949";
    attribute INIT_04 of inst : label is "07241B225B54002E516941AC8EA55C867B185B35520902803884E632B5EF7B90";
    attribute INIT_05 of inst : label is "7994DDAD11097C9083860AD1EB48804A1528D2A4A5A874AAAA4040C15691529A";
    attribute INIT_06 of inst : label is "D1F9D18C11088BCB122F12D1121ABC54AB35CEFBDE9EBA95AC37B355B64E41B2";
    attribute INIT_07 of inst : label is "586C7078895AB476302398C1AAFDFD06481EF5576D6CB15954505ABFC442F682";
    attribute INIT_08 of inst : label is "55154AD558334179B8E1A721A19CE2FB6071E74C6D81D6BA430E1EE308763850";
    attribute INIT_09 of inst : label is "B28F0B2E03DCD74AC618781BB572346BA4A8A926484445552A249FFFFE6BA595";
    attribute INIT_0A of inst : label is "55AEBFE4D26FE922EC7EAEAF53CD884C277DDAB2B76F19EBCBC9D7F7F1A539AE";
    attribute INIT_0B of inst : label is "AF1C7AAFAF21BC2D10D97B56222244C2D6F6F6AE2F18BC62F18F5AD869B6ADFA";
    attribute INIT_0C of inst : label is "4AAEE98C1923319B490C434A6EC51426937C9255BF4263C6CB591349BE435FA1";
    attribute INIT_0D of inst : label is "C32E1435866B524AC848CA106249C0E0923FC47B187FE2B7B03794F52AABA5E5";
    attribute INIT_0E of inst : label is "233A75908EC872E732B9E053E7DC8D14C2F0CDD000F5C6262E3773FFABC60453";
    attribute INIT_0F of inst : label is "E0003FA97B83319DDDD5119534D2A44D1E5E30230BF6E92B47424986F9B4CB84";
    attribute INIT_10 of inst : label is "11427030188E4600812E2E4A0A67DDD5911572AA554D852592C42FC01101BDA2";
    attribute INIT_11 of inst : label is "131B9349C98020F0828D30089631DE7B7BAE1519C9A263693AB3F6C14B5BB216";
    attribute INIT_12 of inst : label is "AD694A42115A4214860A0AD863416C88F0B78218433904202724240D2D313690";
    attribute INIT_13 of inst : label is "02B00324407C0C4CF9C9C2DCB62DB904042122842B4845290A5694AD2948C210";
    attribute INIT_14 of inst : label is "840B19929248C890A9AC29008400104508A29982284534CA120697C40244A582";
    attribute INIT_15 of inst : label is "C0648A54885B9A10A52512980C91A6842025C440AAA9060A93692E8084282914";
    attribute INIT_16 of inst : label is "191D2842148529612842524991122A6B088C2224B18DEDB75975C0432453C215";
    attribute INIT_17 of inst : label is "06A7D957B5BF7FF62219246918CBBCF7B75C0784210F5C05292C92376050814B";
    attribute INIT_18 of inst : label is "FFE8822260AB150BF8FF48643D0C2100C120051260596744C9283188D4AAAA48";
    attribute INIT_19 of inst : label is "0C653351C2AD62267219965E9A428232222F7FFBF7B56B007FC017F8043FE01F";
    attribute INIT_1A of inst : label is "9FE3043E80EE81D129949A52521A0AEE1CB872E1FFACE5E48534843F1D60A94A";
    attribute INIT_1B of inst : label is "071EBE93C0BF6624CE4B5EF1ED6B84B99B25BF758FB6AB1FA26F63490661FF83";
    attribute INIT_1C of inst : label is "99158CBEFB32EF4A64F1635A471412D4D5DA22A84611189D4F7B52E1884963A6";
    attribute INIT_1D of inst : label is "0212B0BFBD88003DAD4AC9240188BAC794211468D658834B2B32F3FCCC065E7F";
    attribute INIT_1E of inst : label is "8F13F0EC7C55E13EEC9CFA227393993DD515F6A613270E2222534DC10B70D340";
    attribute INIT_1F of inst : label is "00644513899969194D31875A97CF8F22B1F99F1CD9E9C55661934C978C85618F";
    attribute INIT_20 of inst : label is "4C70489449E77459804422164A538AAA125D8BB69045602332D882E279288039";
    attribute INIT_21 of inst : label is "55D555D584812029008376ACBB40A21C1121C10A0480B62DB229628120276E01";
    attribute INIT_22 of inst : label is "4CBD65964E297E008E96892CC5235945E19E00BA386AEFD022224B8460838215";
    attribute INIT_23 of inst : label is "482B58CB1452CB0EC32161A5F9FC44442CA8A32BC60453A0158899931DDD52C4";
    attribute INIT_24 of inst : label is "56044CB04A4B2D2839F41E276084446D6D08A6D2C498BF2FB2852CA5D3459974";
    attribute INIT_25 of inst : label is "1496429495233D470D2690A0B25042D7E92A30DA099A58484EE114A4B192B4AC";
    attribute INIT_26 of inst : label is "04417C6000C0524494154AA8888CC76E0C76E8095214165511991121B8A04C5C";
    attribute INIT_27 of inst : label is "A9349BE49B4F8CD93634F815BD4C66A574C5C200C30004A10AA7527364CE5050";
    attribute INIT_28 of inst : label is "02AA80000000000000000002AA8075FBC2014675C474C71860FD3C1FA7A94DB5";
    attribute INIT_29 of inst : label is "44414D4444444C4C4451114445792EFABEAFF80A80A80A8000A80000A8000A80";
    attribute INIT_2A of inst : label is "105555555555544DD544CD7E4D50179B64940D10D415C5050D4D401111111015";
    attribute INIT_2B of inst : label is "A1FD2A0003ABAABABBB93FB84084001800EBABA3D07741CCC015150063009004";
    attribute INIT_2C of inst : label is "01040E071B8001C003F1B0C4F000041201040E071B8001C003FFCFEBAF000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "55450280114A50E5A490B4841498D122851692DA010B4841498D122851692D3A";
    attribute INIT_01 of inst : label is "8D6358E229D09610914314C872A6D6A00B36B5001819CA88E0200F054212448B";
    attribute INIT_02 of inst : label is "CA4989431BB7402524ACD9974E80BA98936139B39DB3AC0E7014E980E7000102";
    attribute INIT_03 of inst : label is "A41DE9780CA09504AC08879FC01008F965039094254136B6DB42311886952528";
    attribute INIT_04 of inst : label is "4FE25240C2728417C54925143E3D58BF67396B11104995A9488928208C2149A2";
    attribute INIT_05 of inst : label is "5304C489192C6E110082B0C18B08910C8528D300A4BA22FFFF4949D40A540E5F";
    attribute INIT_06 of inst : label is "E17C439CC419989017ADB4F3178EB6DCEB6006C2209EF875B636B11196C685B6";
    attribute INIT_07 of inst : label is "09DCF349DBD6B5DE72AA5AD08888AAAA0AA088070739B33B0DD45A90CCC6DFA6";
    attribute INIT_08 of inst : label is "4D04D8CD34F2516B68D346E8A3B4FAD728D3468EDCA31D3A766B3A8005301940";
    attribute INIT_09 of inst : label is "72861B6D769DA798CC31E001345634C024BAA524A0CCCD34666C00C480A9A5B3";
    attribute INIT_0A of inst : label is "C498622D96C04B625D4A29EC3F6CA1EC4769DA166F51052B1B0B0C6C6F451B1C";
    attribute INIT_0B of inst : label is "9C87DA48EC84B5B5418474F66667A4A8099D9DEDADB6B6DADB02D4C2D1B69336";
    attribute INIT_0C of inst : label is "5FBBBDEF5BC6BF7FFF598AD2C6FD746C3601D79364F2DA00B611365B02E73373";
    attribute INIT_0D of inst : label is "43255281064212DCD116E54B60DD8A0497694ED298928220B4614E957EFEF5AD";
    attribute INIT_0E of inst : label is "665262D19958424E6481E443015A993DA6F082C20495B465ADAD6B1C6BCE4441";
    attribute INIT_0F of inst : label is "541120B94A9D13B777777733EFB66B53105E72221208C51F03C147A204904934";
    attribute INIT_10 of inst : label is "550A3E170F87C2C2DA496AFB02E077777FFF166C5BACAB653AAE2F4811429482";
    attribute INIT_11 of inst : label is "11F766C8F14A593800592C18923080808900D228B11A31451102890463786054";
    attribute INIT_12 of inst : label is "B5AD6B4AD2595AD3B2C80CB32F01A410C2A46B4D698951A423CC22DA873E2D99";
    attribute INIT_13 of inst : label is "62540A49716304FE79B10B1CA82A395085BDAB34A53D1A35294A529CA7295AD6";
    attribute INIT_14 of inst : label is "BD8D3B37FFF9D9B0A988ADB64ADB724AC8CB109256467880D16D63F863062528";
    attribute INIT_15 of inst : label is "88492B4A197BBCD694BD067109252734A8128C71FFFD272022596010B4A00452";
    attribute INIT_16 of inst : label is "BD59A49AD295EDA5B3DBFFFFB3362A622988A628B186250402000C4A495B1AD2";
    attribute INIT_17 of inst : label is "32A7139A289926906252482D184901289000C715AD6C2885BDB43AD780D7034F";
    attribute INIT_18 of inst : label is "FFE2C3405A98539402931B2CBD19ED50780E159B7607F7DCF9A4A298E2FFFF51";
    attribute INIT_19 of inst : label is "2E807791AA15A66EF7B1B613215EDE776684F39CE73123007FEFE04007C1001F";
    attribute INIT_1A of inst : label is "148235A3300F37E70395B5134A51297ADCEB73ADE63EC5C2B5B6B5B218AA0729";
    attribute INIT_1B of inst : label is "4F3DBC9BD4F97EA6DE636E738C6B94D35E31EBE59A9E8B35F2A30238412951C1";
    attribute INIT_1C of inst : label is "198CC496A822CE4922902AC1410006C481D80440C653197C5B531A5DE10FFB25";
    attribute INIT_1D of inst : label is "A8D52803718E2A39CC58BF2E45A8B17196110048244021A3199252A08C624251";
    attribute INIT_1E of inst : label is "95363DB80888033ACD981066F0375B01DF11472CDFE781FEEFFECC146BE6FE58";
    attribute INIT_1F of inst : label is "D50E81822B1B653B682387D892CE8576E003823ADBDF088641B785B719C44D8F";
    attribute INIT_20 of inst : label is "5CFA4BB0490E00C19145ACB25296D08C427D8BB0954E6A8636EA04987004A93A";
    attribute INIT_21 of inst : label is "7FFF7FF1EC61B6CDB6A9D1A4BEC6813C9333C93A86DBFEBF862972A1B6E0C020";
    attribute INIT_22 of inst : label is "DC032CB2C0617A408A320B2650A65B4DE1D6100068780A8326A2C935E590127F";
    attribute INIT_23 of inst : label is "D8636B4B34DAD94E5068A9D0040CCCCD2D9A694BCE4441005021B3B73777764C";
    attribute INIT_24 of inst : label is "448CAD94D819CD201801D8296A0CCD6D2D5DA6D2D1B9BF65B68D6DA5B745B804";
    attribute INIT_25 of inst : label is "5CB2C124910B00368F6CD280034952C00B64589A3B9A2B585ECD66B49094A52C";
    attribute INIT_26 of inst : label is "413A5C32058804964E806BB9999980C0980C0A151A5000773333BB637A8CAE41";
    attribute INIT_27 of inst : label is "1B65B02DD6D9AD972F6E6071B4CAA49D61AB53059620248029002600095DD056";
    attribute INIT_28 of inst : label is "FD557FD405557E00055FD5FD557FA8822558A6710404858A2805280425214065";
    attribute INIT_29 of inst : label is "10055D4444444C4400100040012D4D4A5294AD5FD555557FD555555557FD5FD5";
    attribute INIT_2A of inst : label is "FCD555555555545DCC55D5511470D1555053718D5471471C745D444551111054";
    attribute INIT_2B of inst : label is "ABFFAA000050505051BDF7BD4CBD775BB74115E41F3619D9DFDB5B7FE73FEBFA";
    attribute INIT_2C of inst : label is "00208041000003C003F048000009201000208041000003C003FFCFF404000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "5B3A0D06D94ADC1DBD848480181EC599C076E75B0048480181EC599C076E753B";
    attribute INIT_01 of inst : label is "8D6B18FAA9F0965264969D4920A416226924B550811B48A8D82186C5221254AB";
    attribute INIT_02 of inst : label is "4A69AB535BB6E96D6DA45BB6CDCBABF03BC702080C91A46738C668C67389260E";
    attribute INIT_03 of inst : label is "801398524980C4062049583252138288E61253245962D6A5B278AC562A942578";
    attribute INIT_04 of inst : label is "C636D26A565A949775496D14248419A469024A3764DBF08F18B0212484290980";
    attribute INIT_05 of inst : label is "1A9294316BFC5CD0008302C58209832E8522C3A884892299BBDB5BD48A548A59";
    attribute INIT_06 of inst : label is "851990811491135804D234D6048B48C903C302A48C8412018430A3762202D1A4";
    attribute INIT_07 of inst : label is "3496E0919A42B48204EDA019BB0002AA0AA93241494923234956D29C8E8293E3";
    attribute INIT_08 of inst : label is "49049AC920555E9308C65C2CA6214D252D861C38D4B649524A1330C248A25149";
    attribute INIT_09 of inst : label is "23A412496411045AD860A9153416358624ABA525E48CCD24546D20844C8D2DB2";
    attribute INIT_0A of inst : label is "A910400934901A5496921528250CB0AFC69052444BB5694B4A5B4B4B49075349";
    attribute INIT_0B of inst : label is "5680021928144949492414946666848941252428D23348CD2300109405148254";
    attribute INIT_0C of inst : label is "1111118C5B063A24925542DA4289244924811432488686E1442924924094A44A";
    attribute INIT_0D of inst : label is "59254A4B4E5290569174F5792E95AB0DB5494A96931292C2A2A0492444445A4D";
    attribute INIT_0E of inst : label is "441942C91240D243525500890052549D2481208051418C2C6C61614922409C89";
    attribute INIT_0F of inst : label is "5C115171AD01B6E222222222492640422A5204E45E48A09B624555B280964952";
    attribute INIT_10 of inst : label is "548B93C9E0F2781ADBD85B929ACC2222A222074A524CB266B34D290272669592";
    attribute INIT_11 of inst : label is "1C120A4E0709D61649A12C989294A4004980532E071429C6100244A52936295C";
    attribute INIT_12 of inst : label is "94A529DA572B5AD2964927116524E610AAE98ED9DB4948A438157AD14520E490";
    attribute INIT_13 of inst : label is "62526B6D5551248429060EB4C579694885A92C16AD2D9C25694AD6B5AD7B5AF6";
    attribute INIT_14 of inst : label is "B5CD22A44B691521ACB0ADB6DCB2D65418808BB2A8C5045C5D68A282622C6724";
    attribute INIT_15 of inst : label is "886DA95D5B43B072BDA926510DB52416ACB28C7266EF6EACB2C9201094A49F56";
    attribute INIT_16 of inst : label is "0B68ADCA52D5ADA5BB5B496D22A46B2C2988A63894A52748B4100C6B6D4A8E52";
    attribute INIT_17 of inst : label is "66B2B14164948008625B6D2D4A4948249100C554A72A2884A90539A748CC2325";
    attribute INIT_18 of inst : label is "FC00FE18440881000303DBADA118E52F22C8B48B6E7443F68DADA2988299BBF3";
    attribute INIT_19 of inst : label is "6DC654912B15A44AB4212524B15ADA444490421484212DFF8810084007FFFFE1";
    attribute INIT_1A of inst : label is "408114B12125292551220F094A536942100840212D682D2294929CA950AA452B";
    attribute INIT_1B of inst : label is "6924A49B56E168B6D26B6A525A4B16E21C35C3A5D0BA4BA1C302122C4BBD9D49";
    attribute INIT_1C of inst : label is "100CB8F824230A49252882494A891288509AD91044535085C9D26259F14E7C25";
    attribute INIT_1D of inst : label is "A455484042C1A9290A4B1227DCA491523E52892C6FC902A41963E891889C7441";
    attribute INIT_1E of inst : label is "0F370448C7228A04C5098844B6250A6080760524555619544495E5122B42CA62";
    attribute INIT_1F of inst : label is "F4ADC6A2AA124D226A295453120C0F502222B020920B322605B681A4161D8500";
    attribute INIT_20 of inst : label is "80265EACC28ACCB54CC8A7927392B2CC531DC3BC956B4CB424B92336689B2779";
    attribute INIT_21 of inst : label is "22AA22A69A85B6EDB6A49CA49549A4083760837EB6DB4B12C771372DB6ECD9AD";
    attribute INIT_22 of inst : label is "96E269A69851481392D24926D6953AC902A402E26B398A9866924914EDB636DA";
    attribute INIT_23 of inst : label is "9E4ACE432CB293D25C59B9F33608CCCB6D96598A409C89125365B3B7322224C8";
    attribute INIT_24 of inst : label is "D9090D3C9E12182C0B0718795A4CCB6E2A11E4F2B139CF71370A2DE5278DADC8";
    attribute INIT_25 of inst : label is "68A2A184060F41849A485292794976A4DB67105989162CC0E285329C949CC625";
    attribute INIT_26 of inst : label is "1C76D92A39AA76D24D96291111110CD8D0CD9A648A524F2222AAAA42124D0B31";
    attribute INIT_27 of inst : label is "924924092492502A84C9562DEEB72A416D92522CA6A8C4A228921C712DDD5E3B";
    attribute INIT_28 of inst : label is "AAA02A80000AAA00000000A8002AF7C48F379A57EF24ACCF3C65244E2466E642";
    attribute INIT_29 of inst : label is "51405CD555554D551114445111291D4751D4200A80AAA02A8000000002A80000";
    attribute INIT_2A of inst : label is "D0C4444444444544C444DD7B0C151051319159444D10D1450C45104015455504";
    attribute INIT_2B of inst : label is "AAFEAA0003EFEEBAB9BF37BAEDC4AA897ABFAE843676BFCCDFF1F1FF6308CA02";
    attribute INIT_2C of inst : label is "00041A0C12800180E3F168845241000000041A0C12800180E3F70FFEBF000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "0FFD5EAC542106B482DA363662590A4444D23FC825A363662590A4444D23FDE8";
    attribute INIT_01 of inst : label is "3CE739E88C32CB29C8CF0CA4A8625247C716967E4CC963E61211309298D93267";
    attribute INIT_02 of inst : label is "390CE619C8926090D2113462448868909771FDF7E64C931296192231296090E2";
    attribute INIT_03 of inst : label is "FFFCE56B6DB09D84E199F3360A18C18166298CD334E9321A6D0E2713CA409CC1";
    attribute INIT_04 of inst : label is "43490B23DEE14240902C90C1B3965E3779086BC9D39606B07BCDAD9295A52CFF";
    attribute INIT_05 of inst : label is "D328DDE8DC298DA7AF3D2912240E0C9A118D9E3E3634984466A4248A610A6109";
    attribute INIT_06 of inst : label is "D63B4A845A088EC1621B124162306C448B6A5AD91232CEC5B536BC9D98DE43B2";
    attribute INIT_07 of inst : label is "805CE0D88B18B27211BBD0D64E8A0002A016516D6D68B1116D0B88C2C45AF124";
    attribute INIT_08 of inst : label is "24B25AC4922730DB2AD926D2111261B29049264C4A416599C23B3142133B5C20";
    attribute INIT_09 of inst : label is "9226DB6D82C8B39AC596C503B256B2D4961490B010444492222C20DDB29D9591";
    attribute INIT_0A of inst : label is "CD89266DB6D06B66DCD95CAC9622466C56D959222DF6CF7B6B7B6D6D65245B65";
    attribute INIT_0B of inst : label is "9E6CD92DAEC06C6CA092D25622221614659998AE1B186C61B176D67259D64B36";
    attribute INIT_0C of inst : label is "8888898C5916B916DB3FC1714AE4936D3681B65164CAE245C6BCB69B40E73273";
    attribute INIT_0D of inst : label is "A4B0A52D7F5AD71AC6C2C098924F1679622D645EDCDAD93C4C3B85B222222364";
    attribute INIT_0E of inst : label is "225478208B4B1B0A6509A374915D1A19B2DEB10185E59530ACE56528A3422774";
    attribute INIT_0F of inst : label is "30227DF4FF038191111111116DB621413B5A113B519B0244896493493A692C88";
    attribute INIT_10 of inst : label is "0A60C462311A8D68482E2E58512911119191B6231162417FB5C4AD409DC14A4B";
    attribute INIT_11 of inst : label is "C69AA363519428DD0405924E594A164B2C27088351C98C70CEF936518C849707";
    attribute INIT_12 of inst : label is "42108421088421084D2490CCD09211C61832A536B66CA6118D428E44318A32C6";
    attribute INIT_13 of inst : label is "390821241C0CBA218C51E046328C8CA6320D10C21082619C8421094252842108";
    attribute INIT_14 of inst : label is "6378119726C08CBA7E4E1B6D2369092CA613DC496D31BEE3072218A938D1B1D3";
    attribute INIT_15 of inst : label is "63248421A41A43284205590C6490B0C218486709119A92108B658DC64210410C";
    attribute INIT_16 of inst : label is "288E122108431B13663624D811969F9384E61386CA50B1B24964E72124206508";
    attribute INIT_17 of inst : label is "89F85D2CB6C2C96739092298A52C2CB2C64E71C2108186320562C4152B20AC90";
    attribute INIT_18 of inst : label is "041F83E7FBFF7FFFFC4B245205661099A96A422624CC1A90DB12184E3844668C";
    attribute INIT_19 of inst : label is "848966F596C3022CC6B5B6488C31B02223495A5694AD93C4FFEFF7FFFBFFFFFE";
    attribute INIT_1A of inst : label is "8101C20DC511C5B82CAF5D24210C840A992A64A9B5AD9D98424842049E053084";
    attribute INIT_1B of inst : label is "8596B6CE6D8DC36D89CEC149396E6D8458E70B3702F36E059ECA5981A5293373";
    attribute INIT_1C of inst : label is "C6E2091B56382B6492815AE4211572E2F0DEBAA857085DD746AB9B258C6160B0";
    attribute INIT_1D of inst : label is "530148405AD214AD2964C9B02652CC08D528613D0FE408D0C424654AE3848CA5";
    attribute INIT_1E of inst : label is "8516756A97552376F1A52C22C4B6A34E199D95B30668D33222C6926987784868";
    attribute INIT_1F of inst : label is "0A6488F9835B7811C794675CD92C8534AA0B24925969755615926CB64F27702A";
    attribute INIT_20 of inst : label is "64335A36492C96599A7610594A59913B18531A66C2CD6366B6F408416E4050EC";
    attribute INIT_21 of inst : label is "119111998A5B6D9B6C52C232C602E10EC930EC834DB624C93C8D98D36D899252";
    attribute INIT_22 of inst : label is "590B8E38D22D6A04ED292CB329468365BD980C4FD49135769D4B2CC25044C901";
    attribute INIT_23 of inst : label is "5B7B6B4B165ADC65232E0D88CE0C4445AC8B256B422774C10891E117E1111704";
    attribute INIT_24 of inst : label is "66CD4DC659D9AB3BB20C9D8D6D0445ACAC88B2DAD8BF3C2CB244AC95B629B212";
    attribute INIT_25 of inst : label is "CC30DF5F9DF84367E127084114240ECB2370549C295B834B1EF08842CA52B4B3";
    attribute INIT_26 of inst : label is "46EB78614680D24924C98088888DA9931A992D0A610820111111116B5D394EA6";
    attribute INIT_27 of inst : label is "8B69B40DD6D928BB672F6993B0CA6E19768244925A0A362985C9B3D4E44B40B0";
    attribute INIT_28 of inst : label is "AAAA8A0000000000000A80AAAA8A02195088F32D3496539A691D9B25B3F2D36B";
    attribute INIT_29 of inst : label is "EBAECFFFFFFFCE66AAB2AACAAB7BBFEBFAFEB80A80000A8A00A80A80A8A00A80";
    attribute INIT_2A of inst : label is "BFCEEEEEEEEEED66E67FFF7BEFBEBAFBBEBBFFEEEFBEFBEFAFE73ABAB2AAB7FC";
    attribute INIT_2B of inst : label is "AABAAA000000001011BD37B85E8D775AFD5054E81F7619DCC0515140E77F87C1";
    attribute INIT_2C of inst : label is "2492412004000000F3E00032092492492492412004000000F3E007F140000002";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "0FF80C055010861016DC343242581800D0007FC125C343242581800D0007FCA1";
    attribute INIT_01 of inst : label is "1CE739C000228C21C8DD4AC0E0D2D0CECE928234088041445211289240500006";
    attribute INIT_02 of inst : label is "10AC401880020148090882020440E0801201000040000200040C0420004000C0";
    attribute INIT_03 of inst : label is "8010853365301980C09540201A00C3834674181615E0A009002C269308008801";
    attribute INIT_04 of inst : label is "03048B03DE8100020068488096BAC91739082905521003902924A51295AD2880";
    attribute INIT_05 of inst : label is "D9B059885009DC86AD353BB76E050400310E189434381000221212A840284028";
    attribute INIT_06 of inst : label is "D6384A8458088889620916E963382665D92A5A490236DA6CB5669055305E0392";
    attribute INIT_07 of inst : label is "0848404889189672102380402AA8AAAA8AB2512D25289111270A0C82444A7000";
    attribute INIT_08 of inst : label is "65964A45922560496A5972E031173097005972E45C0124CBC03B11C2091B4800";
    attribute INIT_09 of inst : label is "B722C925E2D8B64A45964D0696D29654B43831A000444596222620499394B491";
    attribute INIT_0A of inst : label is "44892664A2507122484B55A592640644124B4B2225A3072929392727256E492C";
    attribute INIT_0B of inst : label is "0A4C4B25A6C024258096D6D22222343024B0B1A709182470992652D2CCD2C962";
    attribute INIT_0C of inst : label is "88888884C9129912490443834A459725128082012C40400142AD928940421621";
    attribute INIT_0D of inst : label is "C0A0842E7D5AD20A46068194024830210225244E4A4A50BC6413849622222125";
    attribute INIT_0E of inst : label is "225830008B5E9A0B361CA158914C0C3896529380B54CB769E5ED2D28A1421558";
    attribute INIT_0F of inst : label is "24115DA6A509C1911111111124922341A94A10AA5511A006119492802C3028C0";
    attribute INIT_10 of inst : label is "0840C060301A0D00016E264CD00911119111B2211124012A9544A54055018C0A";
    attribute INIT_11 of inst : label is "869A9343499064D0004D100C518C36C968662503498B04618A5132614A44B206";
    attribute INIT_12 of inst : label is "0000000001000000000002580000088410321080002884410D230C0529093282";
    attribute INIT_13 of inst : label is "30000000180CA0218848C0C4170D888420058180000044880080000040000000";
    attribute INIT_14 of inst : label is "0020119202408C951C2C000094048005C036880026009446260294A43060A1C2";
    attribute INIT_15 of inst : label is "42000205C01A0684000D50084000A1800000460000884A081B65048400000000";
    attribute INIT_16 of inst : label is "2C04094080000008080000481193470B00C4030EAC61A196CB2CC60000105080";
    attribute INIT_17 of inst : label is "54705D64B6865B2630000700C6286DB682CC608008410420053080142A00A800";
    attribute INIT_18 of inst : label is "07E0820040080103F84B00400D450841A5692110201C8E08C809100C1000221A";
    attribute INIT_19 of inst : label is "444522D490800224429492C81800002233095AD294A50BC4FFEFF7FFFC010000";
    attribute INIT_1A of inst : label is "2101A105850184B0AA2D2810008A401ACB6B2DAC94A49C9000002104CC142012";
    attribute INIT_1B of inst : label is "859696A0600D03000B0803597B28602CD1841A1406A1280D085AD10394422262";
    attribute INIT_1C of inst : label is "22D10BEB56042B5208004A921105565150529AA8D2844A8444A95A250A5140A8";
    attribute INIT_1D of inst : label is "4A8040401AC812AD2952C9A81042880454A4D11CA9920448A22FA5481185F4A4";
    attribute INIT_1E of inst : label is "8512716A9355213680C12C224492C148115594A2822853322243206547344064";
    attribute INIT_1F of inst : label is "094444D101492011051A734AD1288525AA092596C928355234924C92C815606A";
    attribute INIT_20 of inst : label is "64335016DB24965C81550AD15AD582A294D03A02A2052102924204414C0448A2";
    attribute INIT_21 of inst : label is "1111111580080020004A4622A306A325A0125A01000024491105404000091241";
    attribute INIT_22 of inst : label is "4A090410522D2A02AE302AA02103112CA58C054918052553410AA8A140048001";
    attribute INIT_23 of inst : label is "4B296B59165A486E032C0D004A044445A48B2D29421558800080811281111204";
    attribute INIT_24 of inst : label is "564564864B4B2A6B3205CB4D2C0445A5A588964A58941C2592C5A49492289412";
    attribute INIT_25 of inst : label is "06185A9535A041725126800012921E592122D5C86B49015E8E6854228C5294A9";
    attribute INIT_26 of inst : label is "064B78600700400004154088888CA9130A91249950000211111111294CA164A6";
    attribute INIT_27 of inst : label is "89289404824B002962252997945ECA33330000004C00140100811350C08B00A0";
    attribute INIT_28 of inst : label is "0000028002A02A00000AAA00000282B9420442301814631042090980A1C88B2A";
    attribute INIT_29 of inst : label is "AEBACFFFFFFFCD5D55555555550100140501400AAA02A0028002AAAA00280AAA";
    attribute INIT_2A of inst : label is "90CEEEEEEEEEED44DD44C5041041450441440011104104105045090817EFF7FD";
    attribute INIT_2B of inst : label is "AABAA8000155554545BD37B84C842208300004C0147619C64051514073088200";
    attribute INIT_2C of inst : label is "0000000000000000618000000000000000000000000000006180038000000000";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
