-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "800424D84A3520F8AEBC5719BA6CD6CEC36141FFFFFE00A0C1FEA7A3D3F3EDB5";
    attribute INIT_01 of inst : label is "1C640055319604D58A6C25108EB3AED2531D954AAB2B0B8802200841281E3C12";
    attribute INIT_02 of inst : label is "EFF4FDFE930F1BE3FC9B4494135A75841BE7445AA86A13B5340531A3546CA70C";
    attribute INIT_03 of inst : label is "23E2AE6FBBE6C90D74C0002410480DD2B57E8747EE11EC54D2E9FCD1D9DD7FA7";
    attribute INIT_04 of inst : label is "34E14853353C444443FB4417BFEEC522AA4E33CF44EDD1897111BAA98F43EC2D";
    attribute INIT_05 of inst : label is "2A64E2981509AB80EBA4BAE9B5E17B84E3DE8E53BDB5565AD2E64DC0ABDCC71C";
    attribute INIT_06 of inst : label is "14514C4470002E0005C0003800170000E0005C0003800170000E000DD6976DC6";
    attribute INIT_07 of inst : label is "5545545545155145545545545545545545155545555545555545545555155545";
    attribute INIT_08 of inst : label is "4514514515515515515514554554555554515514555514555554514514554554";
    attribute INIT_09 of inst : label is "5455455455451551455455455455455455451555455555455555455455551555";
    attribute INIT_0A of inst : label is "A2F8D883A5145155155155145545545555545155145555145555545145145545";
    attribute INIT_0B of inst : label is "B69E8F7B30C4E0D4ACD2606A574D18981A8B669383516E9A7AF17290CF4FE196";
    attribute INIT_0C of inst : label is "6B4BC9F6DD8F7E6342C549A4267A17E8ED43E52E9436E2A98AD2F76AA579E8ED";
    attribute INIT_0D of inst : label is "03F2221208C10045A3ABBFE1E579F7CFBC282410492BFF7B333333335D76D4D2";
    attribute INIT_0E of inst : label is "40000036480000075A84399B2D8D34A828050908928924005588B5B42D16891B";
    attribute INIT_0F of inst : label is "DCCF9742DAD4C145C68A3655455C8BFDEFE7999FC0FF00004000000040000000";
    attribute INIT_10 of inst : label is "59B372526D708010C208400840D81001102C31A4BB7D6A60AE345B99B997C6E5";
    attribute INIT_11 of inst : label is "5C941A20616D44AFC5C4D13A2D27FDCBE37265F2A991ABB76F9811B057CF94D8";
    attribute INIT_12 of inst : label is "EA074EAA2216C890FAA4C30F751224644D72250AA001AD68D19E12AA5FA422D7";
    attribute INIT_13 of inst : label is "0170ABE7482F326D9F5D69152114B7E64DB3E5368229056C5A8262E89185468E";
    attribute INIT_14 of inst : label is "880000000004020100020400014082C1680002011C09028002204400440826AB";
    attribute INIT_15 of inst : label is "40080160A00080000000800000050001400000028140A15000540B0080000800";
    attribute INIT_16 of inst : label is "040000162A000000000008000000500010000100A8140A05080540B008000080";
    attribute INIT_17 of inst : label is "C000000002010080000000080000000000000800080000010080000210000000";
    attribute INIT_18 of inst : label is "06E466345440AA293C9921055245A7A956FF49FFB2D637398973A3F7F6646A05";
    attribute INIT_19 of inst : label is "429B7636754618B91A881545A7932814DBD519B1B3AAA0C5D1B28D942CC5C4CE";
    attribute INIT_1A of inst : label is "C7709AD893CA333316C2C9678B7E48D439B9662BAAADEFD491B024089B4FE2F5";
    attribute INIT_1B of inst : label is "49DB2A4ED9413061801205A3DEEB75DAD74A6F4B3DF66F5EB53A8BBA959F59A5";
    attribute INIT_1C of inst : label is "06EF313FFB16FED33593B24CDF68E5A13BE9F9BEE9B7CAC311276CA93B6504C4";
    attribute INIT_1D of inst : label is "86455F0F09ED4B1A6426984484EF2A3E19154F0F3244A6DF991E4DB9F65F66F4";
    attribute INIT_1E of inst : label is "7F8D24D3055477EFDC9C006CB488CF288AAF7770CB4DCD388F64771A925BCA8F";
    attribute INIT_1F of inst : label is "DB5924FA6AAB9277BF724461D187C7447445B7DFB15B12CB0270510130983785";
    attribute INIT_20 of inst : label is "6356B6FEFEF94F2025DC8D7EE7B936F3D652BD722832D3BB84C841040841043E";
    attribute INIT_21 of inst : label is "8AF93C8D6D93985447A5A77B0DF5C755043A0874175C71E404B8FCF1AEF73DCB";
    attribute INIT_22 of inst : label is "EFFD54CB4EEE1317055D777D7FBEEBABAAAAAAA91E9A34104172EFDF9D1ADFFB";
    attribute INIT_23 of inst : label is "46B3FB82F93D8D655EBFA5A77B098D1FA6942CBBF7E746BF05F7026E79F27D1A";
    attribute INIT_24 of inst : label is "AF5FF2D3BB84D64000000000000000000000000000000000000274D09CBBF7E7";
    attribute INIT_25 of inst : label is "7BE7D6628ECCF2F3F59B49330CC3BB529434EF84CC5D647DBEC3CD34DC9F46BE";
    attribute INIT_26 of inst : label is "7336426CD909ACC9D2C29A62E6A208AE3D9098CCDB4BEFF249FAD57F6A2BD7CC";
    attribute INIT_27 of inst : label is "D1CFF0C7BFE4B9D11D1412AB473FC31EFF92C69D42885C49029B54C1319B2131";
    attribute INIT_28 of inst : label is "F8EE74474544AAD1CF70C7BF64B1764FEFC6F66FC434DDFE079F2D34474504AA";
    attribute INIT_29 of inst : label is "17163A23A2224568E7D863DD25CBD1D11D1412AB473FC31EF92C68A85530707B";
    attribute INIT_2A of inst : label is "8698299B6BB7B6C4A4ACA2C74542A98383DCC972F474474504A2D1CF70C7B64B";
    attribute INIT_2B of inst : label is "B3BB484D25B45659F677690E0CB67184D690BAEB5159DDA42690D84E89889586";
    attribute INIT_2C of inst : label is "11A68060A28300100229E18C6C02899D159DDA42627817481D61A1A60A647962";
    attribute INIT_2D of inst : label is "E18C68028871800038E69B00100000641104000000009001A784098000240698";
    attribute INIT_2E of inst : label is "9811A68060A28204100229E18C6C028809800020069811A68060A28304000229";
    attribute INIT_2F of inst : label is "B9CC79652A16524FCE8ACEED213132A2B3BB484C4CA8ACEED213520980002006";
    attribute INIT_30 of inst : label is "39B9B93909CDCC1400501420EE803D40447EA4648A135F55A1A438576351D1AB";
    attribute INIT_31 of inst : label is "B00E60069A3185346864C97C42258D8C910C431891421400310C621886218921";
    attribute INIT_32 of inst : label is "0800100100100019040104000000244100E00A58069E28068E01504100100100";
    attribute INIT_33 of inst : label is "21E29B0102C001B04068A78E39B04044101004100400014101101300501C6400";
    attribute INIT_34 of inst : label is "100B00000600A28044008A29800901E00014020E29E2400010162C049E01F004";
    attribute INIT_35 of inst : label is "7D3E9F4FA7D3E9F4FA9E38E28258E18E01638100040104100400104041E70248";
    attribute INIT_36 of inst : label is "A7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA";
    attribute INIT_37 of inst : label is "FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4F";
    attribute INIT_38 of inst : label is "4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4";
    attribute INIT_39 of inst : label is "45145145145145145145157D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F4FA7D3E9F";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE51451451451451451451";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "7A3C0056875E9D6036D01B6C289D5401DA064CFFFFF8592DCAFBCD6603E38D93";
    attribute INIT_01 of inst : label is "7A824F0A6B466061D02B41C5B6DB77FE8440A78FBCB71F6D2B04476C99BAEE81";
    attribute INIT_02 of inst : label is "7F3D4FE7A8C2803C5524D0559149D27589EB8EC5FF3EE96ED2C9FBCC72AB849C";
    attribute INIT_03 of inst : label is "11F790A023039B4405004104800000544753F7E22C7AB348FFA364971069F9EA";
    attribute INIT_04 of inst : label is "AD05C4925B07EBEBE91405410044500518C417FF2DFD8CAE35DC9FF3D21A0931";
    attribute INIT_05 of inst : label is "674D01D807857A0965887BE276879002C3D8140197E03F478C4AAD401BBC9720";
    attribute INIT_06 of inst : label is "00000DB8F000160003C00058001F000360003C00058003F00076000BDB4F6E06";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000010000010000000000000000000";
    attribute INIT_08 of inst : label is "1001001000000000000001000000000000000000000001000000040000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000100000100000000000000000";
    attribute INIT_0A of inst : label is "F7F9EED860000000000000010000000000000000000000010000000400000000";
    attribute INIT_0B of inst : label is "376D290C8408592C77242C963BB2510B2587B92164B0F76514AA155A957FE5BD";
    attribute INIT_0C of inst : label is "993952924555310B308D90DFB4E8B322E2079C4E2072113090A61B3099FB9169";
    attribute INIT_0D of inst : label is "7AC2FBA8718B221AB014001ED4800D9E7B4C96C900060003BBBBBBBC2A18A26D";
    attribute INIT_0E of inst : label is "9F00E0381000000B0ACD03F1923A403AB09DC678421004A49DF19292B9DEE537";
    attribute INIT_0F of inst : label is "7776206F20195D9C10D0A00D8A00A3D21019E1E01FFFFFF01C00001F9D801FFF";
    attribute INIT_10 of inst : label is "8C4D2CE5024080100200400801451D50D8C3C4000C900CAEC08680CCEEE9002F";
    attribute INIT_11 of inst : label is "9558434CE8918A725B1C164364D1672C178FF8141FB41660B12A800181326200";
    attribute INIT_12 of inst : label is "AEFD1FAED2A012C4006A516622D0D5A5C298D3B90F6DFCA2163E47BBE616E01A";
    attribute INIT_13 of inst : label is "F8141E4BF0804800BD754622B697E4090017ADE0BC45BFB003ABED4C22A0FC5F";
    attribute INIT_14 of inst : label is "0011200408200280002050000540A391C104A000141C4805028955AA512A8002";
    attribute INIT_15 of inst : label is "10A051C9F4AA552A954A2552A850AA542A8140A3D3EBF4FAD51E9E4A25528040";
    attribute INIT_16 of inst : label is "100A051C9F4AA552A954A2552A850AA542A8140A3D3EBF5FA551E9E4A2552801";
    attribute INIT_17 of inst : label is "440A25528954AA552A141AA1528140A000000C0AA550A830AA0542824AA54280";
    attribute INIT_18 of inst : label is "50989B458DAB0C5F89124A586C880C8C732D34598D3978E7336C080383ED0530";
    attribute INIT_19 of inst : label is "EE000B448CB4920221B5618BF12245700032D25A24652C9005002A419225AA0F";
    attribute INIT_1A of inst : label is "2001292B68294A45A004624FB4B3E00EA6C7DB5F80007256200E96944122D548";
    attribute INIT_1B of inst : label is "72ADB2B56582C4B24D2D464D605AC077BC749875132C81BC01AA42D8FB649292";
    attribute INIT_1C of inst : label is "6B21064B180B3B66D924A49B6DB542D64B0ABAB7110981504DCB966ADC920B16";
    attribute INIT_1D of inst : label is "A8AEAF70CA3EB5228BA926D5170755DEA2BA9F70F7A948A041E4AA0094BD85EC";
    attribute INIT_1E of inst : label is "5316A6DB5D35DDA3420372298A335D611337DD77F29429EF281940A5A381D577";
    attribute INIT_1F of inst : label is "4156590F3112014E8D13F1AAE6A8388B888E93468082248225734D61B2DAD316";
    attribute INIT_20 of inst : label is "3C6A0304BCBA91C5413A300202140767E4EC062A8A9CA480221A00001A000038";
    attribute INIT_21 of inst : label is "9CB4133019373FBFAD794904C416D92DB25B64BDB16C9238A8249A66034084A8";
    attribute INIT_22 of inst : label is "27D555F292188034C00822282AAAAAAAAAAAAAA83B64FA5B2C8092934E603012";
    attribute INIT_23 of inst : label is "98041294B41030014ABFF9490C40331AD9350024A4D398080E251429CD682460";
    attribute INIT_24 of inst : label is "A55F9CA48020090AABBBBBFF57EBBAAEAEAAEEEFFFD7FBBAAAAAF690A024A4D3";
    attribute INIT_25 of inst : label is "4800601310102C959B6A900000208294E269012222471A8A0920A4121E089800";
    attribute INIT_26 of inst : label is "4B41110D044012D23B26259D5454C7DCA044032D4812514D2467189B89AF2975";
    attribute INIT_27 of inst : label is "2520C6142A8102C2E222ACFC94821050AB041923A664C0A963FFEDD36DA08803";
    attribute INIT_28 of inst : label is "0280B8B889EB37252044142A010349E303B839831880F077982C8038B888AB3F";
    attribute INIT_29 of inst : label is "34B1C45C44F49FB290230A001C10CE22E223A4DD9480105010E191152B75AD48";
    attribute INIT_2A of inst : label is "46D9A5ADA2DA45C7F7CD2C3889AB5BA56A4207043B88B888A91F6520C4140838";
    attribute INIT_2B of inst : label is "44829201F2418892DB905242553905220CF9A49E6622414900FB2817AFD9A196";
    attribute INIT_2C of inst : label is "11A6D461A39255451638E19869469C76622414910D92490DD46591B66968B3CC";
    attribute INIT_2D of inst : label is "E19869469C71D51068A78A55451451600451550451448551A38409D51471468C";
    attribute INIT_2E of inst : label is "8C11A6D461A39351451638E19869469C09D51471468C11A6D461A39251551638";
    attribute INIT_2F of inst : label is "C7398370D0801C963F31120A4882CFCC44829220B3B31120A4882E09C5547146";
    attribute INIT_30 of inst : label is "CACA4A4AD252522AF0BFABFE277BC3D19F21D5B0BBFC0000333CDA14EB3A993D";
    attribute INIT_31 of inst : label is "A51A21429A30C100852D3F90A4C21292FB5EB7B5E3BFEBCF6A56F5B52B7A5E6B";
    attribute INIT_32 of inst : label is "0951451451451458011451415551211451A50A49439E28428B50051451451450";
    attribute INIT_33 of inst : label is "60E39A50079401E51429A69A38E51441451001451551411451050051051C7144";
    attribute INIT_34 of inst : label is "451A50051350A28411448A39C41C51B55401470E69A61401451629418F50A510";
    attribute INIT_35 of inst : label is "28142A05028142A1509A68E68619A09B50279455401451450151451401A71209";
    attribute INIT_36 of inst : label is "028140A150A8542A150A8140A05028140A05028140A050A8542A15028140A050";
    attribute INIT_37 of inst : label is "5028140A05028140A05028140A05028140A05028140A050A8542A15028140A05";
    attribute INIT_38 of inst : label is "05028140A05028140A05028140A05028140A05028140A05028140A05028140A0";
    attribute INIT_39 of inst : label is "000000000000000000000128140A05028140A05028142A150A8140A05028140A";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "03454050C042026414320A19C340CC0596058B3FFFF811D543F94D7719E99B81";
    attribute INIT_01 of inst : label is "122B6A0310C00060102861C5946B45F686DDB5C994270709080A004908038E80";
    attribute INIT_02 of inst : label is "7F3DAFE7B142A5D4552C8405000A60A508957280EB8400AA008FDBC370A80400";
    attribute INIT_03 of inst : label is "FFFD8228A22812414440000000000110B30C2121A2480A5419935C954849F9ED";
    attribute INIT_04 of inst : label is "7C93F9211735AEFBAFEA5003AEEEBB81008615A00DF0542D15A48553F65A2D30";
    attribute INIT_05 of inst : label is "2EDC93B40598E2414332A0CD009393563795CCFB336B9CFDECC82C4161D08792";
    attribute INIT_06 of inst : label is "00001A576800850009A00134003280065000DA001B40042800C5001199141927";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000010400000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000040000001001000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000104000000000000000000000000000";
    attribute INIT_0A of inst : label is "B2F99445E0000000000000000000000000000000000000400000010010000000";
    attribute INIT_0B of inst : label is "6DBDA522150E334CFFFF09A67EDB49C2698FFFF8CD31FDB634AA5690847FC5BC";
    attribute INIT_0C of inst : label is "95A8DB3149D9044A308F804F3420F102C766006C76710E3E33A71A1B89FBA1D9";
    attribute INIT_0D of inst : label is "B8CA918E399FFE03300400AAFD71B586180020904003FE7BBBBBBBBDC47F4024";
    attribute INIT_0E of inst : label is "5FF803C85000000B49A90DB9DF0B740A86B8C73A9385B46C1900A49481C0E11C";
    attribute INIT_0F of inst : label is "76763C4BF2005C171002A004528A23D91001FE005FFFFC0FDC00000FDDFFFFF0";
    attribute INIT_10 of inst : label is "C5993B3B619740E89D03A0744E0C8844EF6618200EF900AA1880188ECCEFB63E";
    attribute INIT_11 of inst : label is "85C3400868F85220C5069063C537977D27148854210005BCD9BA8D8FC660DAC7";
    attribute INIT_12 of inst : label is "46010C06052000940020514624802435637C948A01212832501E43AFE624BA03";
    attribute INIT_13 of inst : label is "FA140B6FE6A01200B9E7E784A494B60240173F72AF0925DB40A8496038A0414C";
    attribute INIT_14 of inst : label is "0A41028040A01000000804028040828148140A051E8D4200008914AA15229156";
    attribute INIT_15 of inst : label is "00A0516AB40A05428140A05028000A00028110AAD168B45A05168B40A0400050";
    attribute INIT_16 of inst : label is "010A85168B40A85428140A05028000A00428100A2D168B45A05168B40A040000";
    attribute INIT_17 of inst : label is "4000285028140A05028100A45028140A04001810A156A8742A05028740A05028";
    attribute INIT_18 of inst : label is "540E0D05042F829B8D90E87C61E1080E61934DE58B5A714213692A03204001D4";
    attribute INIT_19 of inst : label is "22800D04252410878085F05371B20B1400949068212928841500A805000FA2A5";
    attribute INIT_1A of inst : label is "67A1B9B9B14A104F8636424F1BDAE6C473656D0B910C5F7E3D8080A7D96F22E1";
    attribute INIT_1B of inst : label is "7FF7FBFFB7D7E6BA6D7F53E7ECF79FBCEF7FDF7CA5BEF93905A29294D1B6DBA1";
    attribute INIT_1C of inst : label is "7DBDF7EAD75DADF36FF6FECDB6FD2767EA21B2B5990CF9906DFEFF4FF7DB5F9E";
    attribute INIT_1D of inst : label is "BC974F7C4F010E3BC33D005DDD87061EB24D1F5C77C046577FFFCF176FE6CF3A";
    attribute INIT_1E of inst : label is "4D9BA08241456E4489DE766829BBACA3B99FF57D5AD8A5B5A4371201FFE1C387";
    attribute INIT_1F of inst : label is "935FED0BA19BFF51123D4DD2F7482CCECCCB6C89103F3EBF3F71554020120D9B";
    attribute INIT_20 of inst : label is "76683786F4AAD867FD45BFE0428137B7FEE9B022A016B691205B6DB6DB6DB6FE";
    attribute INIT_21 of inst : label is "97CBED3FEBA9E150042D6D224090430C0018001DB30C140CFFA8E5F7FF52040B";
    attribute INIT_22 of inst : label is "D020025ADA458925200822282AAAAAAAAAAAAAA81924BECDB68EA3DCB77FD01B";
    attribute INIT_23 of inst : label is "DFF81B9FCBEE3FFAB0142D6D22C494976DAD23A8F72FDFF40B371FCAEB97DA7F";
    attribute INIT_24 of inst : label is "580A56B695624A8AAAAAAAAA00000000000000000002AAAAAAAB492793A8F72D";
    attribute INIT_25 of inst : label is "21ABF221987436DECDFADC19064116F7BA6D87A040E5D237F7CBED36C1F71FFD";
    attribute INIT_26 of inst : label is "5203D0280FC494835BB437F7327FEF7090FC49487AC96DFF7D3D8CCECAA9EDD9";
    attribute INIT_27 of inst : label is "B4AAE45295A39383B333F6D6D2AAB94A568E4A35B476848231F42DD6A901F892";
    attribute INIT_28 of inst : label is "3624E0ECCDBD9DB4AA6E529523925066868C68C68CB4B8C71A38AD3CECCCFDBD";
    attribute INIT_29 of inst : label is "2503667666FFDEDA5532290908998B33B337FE76D2A8B9484844A19F3B74E929";
    attribute INIT_2A of inst : label is "2410A90F7F65BAAE8E88286CCCF9DBAF4948822662CCECCCFFBDB4AA6E521211";
    attribute INIT_2B of inst : label is "661ADE25A284CCFF6CC35BE47ABD34A04ED129DF33330D6F12D1439F5A357124";
    attribute INIT_2C of inst : label is "100014500500514514514004014514173330D6D0240B6D2F504909042A41DBE6";
    attribute INIT_2D of inst : label is "4004054514004514510000514555514410514515554510514510004554514514";
    attribute INIT_2E of inst : label is "1410001450050051451451400401451400455451451410001450050051451451";
    attribute INIT_2F of inst : label is "8A109379D2891C0F0B99986B681202E6661ADA0580B99986B681220055145145";
    attribute INIT_30 of inst : label is "C141C1C14A0A0B2080180030EA02008DCC3C49F6ABB0000005095A04723E9C29";
    attribute INIT_31 of inst : label is "451450000000020CD3210D26BE5AD4D4D0C251842503000819CA338CE5094208";
    attribute INIT_32 of inst : label is "0055451451451451045451451451441451451451451451000451451451451450";
    attribute INIT_33 of inst : label is "5000005140145005145145144005141145041145005544145045145105001145";
    attribute INIT_34 of inst : label is "4500505514504514514514404404500514514514514514454500114514514514";
    attribute INIT_35 of inst : label is "28140A05028140A0509451451040040051455451411451451455451450001055";
    attribute INIT_36 of inst : label is "028140A05028140A05028140A05028140A05028140A05028140A05028140A050";
    attribute INIT_37 of inst : label is "5028140A05028140A05028140A05028140A05028140A05028140A05028140A05";
    attribute INIT_38 of inst : label is "05028140A05028140A05028140A05028140A05028140A05028140A05028140A0";
    attribute INIT_39 of inst : label is "000000000000000000000128140A05028140A05028140A05028140A05028140A";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0603502260C780741C5A0E291140558DDEC40F3FFFFC11D7C8FE64D6D8F8F289";
    attribute INIT_01 of inst : label is "40892423108C5253000131C12A61E0C1D31DB1A050A381214A92009049010608";
    attribute INIT_02 of inst : label is "AFD5B5FAB184232FA9926E24D8C37089C93EF9538D400303508F51963241109E";
    attribute INIT_03 of inst : label is "33F4929C852000131810000000000810D84C3089CCE28A5A0C511F53C8C37EAD";
    attribute INIT_04 of inst : label is "AC55C0045112505404150554410151211A05999F042C431EC3DE919980D5E5E9";
    attribute INIT_05 of inst : label is "277C51D01D046F41C590236507D5C18A9352060B1F720DE3866807408391760A";
    attribute INIT_06 of inst : label is "000013FFA0011C00168002D0004A000940013800270000E0005C0002CF0468A4";
    attribute INIT_07 of inst : label is "28000A28000028A00000000000000000000028A28A28A28A28A28A2802800000";
    attribute INIT_08 of inst : label is "000000000000000000000000028028A28028A00A28000A00A00000000000000A";
    attribute INIT_09 of inst : label is "0A28000A28000028A00000000000000000000028A28A28A28A28A28A28028000";
    attribute INIT_0A of inst : label is "AEF4554B600000000000000000028028A28028A00A28000A00A0000000000000";
    attribute INIT_0B of inst : label is "48B1CE7F185676792AFF2B3C957FB8C2CF2D45B8D9E5A8B62A131252990BF313";
    attribute INIT_0C of inst : label is "48B29D3218ED2765618B1DB159EA53692C8D0D12C8D21FC3AC73256499BD9895";
    attribute INIT_0D of inst : label is "C886458A9425DE22554460A27CA1E49A690082094012A183BBBBBBB87FC44492";
    attribute INIT_0E of inst : label is "0000000000000000116411B11F2931223A5AF7BFFC9B68B21298918203CE2528";
    attribute INIT_0F of inst : label is "54441093F09419C404A220166280A97240000000000000000000000000000000";
    attribute INIT_10 of inst : label is "08030424043702E01C0382700E1014553500C1280AF84A0CE025018AA88F907D";
    attribute INIT_11 of inst : label is "419D128020FA62A858542306C5ECFC1806148A00210024B0DAD484120008280A";
    attribute INIT_12 of inst : label is "46FBA446F518245000A00000308038F5C37010AA00A68CF563DF3A1EC4292895";
    attribute INIT_13 of inst : label is "B2C02BB6C20A9A00B1C7C124C8D6AC5340162D61B24A45D9122341AA12017AE4";
    attribute INIT_14 of inst : label is "164882CAE082104482540C12CAE482A15C101E221F0CA342A0D1A6A51C34E555";
    attribute INIT_15 of inst : label is "845229E1A0336A855508E783C042A050A8080453ABE1E0D0501C1BC1E08050F0";
    attribute INIT_16 of inst : label is "8845229E1A0336A855508E783C042A050A8080453ABE1E0D0501C1BC1E080508";
    attribute INIT_17 of inst : label is "4E8F4783D1E0F0783CDE2F0583DDF6FB088452210182C042300804068100986C";
    attribute INIT_18 of inst : label is "5124A45DD564131B16C732206649001FE2BF7B3F0118E14A590C220208400961";
    attribute INIT_19 of inst : label is "2A802451C43186292AAC826362D8E1540110C7228E21EC3151008804006AC8E2";
    attribute INIT_1A of inst : label is "7FF5B1B9B1CB185220504144FDDAC20BA765744B00409F7D5411A8C50159F5CC";
    attribute INIT_1B of inst : label is "CB176658B33B726923B6EB6B27B5B6AC62FBF6BE6D9E6C304682C0749CB2CBE1";
    attribute INIT_1C of inst : label is "65C62374626DC4B5BC9F13D6F25EFB7B79C55D5EAB576AEF232C5D3962C8EDCC";
    attribute INIT_1D of inst : label is "CE935F9B33ACA6F4D50F6169E9C7863F3A0C4F9B22C05F799B32C3192262731A";
    attribute INIT_1E of inst : label is "64FBBD550B74CF468C8889D180AAA8B08CCD757F5A58CD91CF7C03413CF1E9AF";
    attribute INIT_1F of inst : label is "487492E0988A920D1A3C6552D543C444446B268D1CC9B6493702DD3D53A864BB";
    attribute INIT_20 of inst : label is "BAE1EDF262837E2C6434ADA91AD7E9985346D6880A36973BC05A49248A4924AA";
    attribute INIT_21 of inst : label is "D769252DA0C48415506D2E770090C105248A4934110C35C58C85B4D5B708C6B4";
    attribute INIT_22 of inst : label is "528000DA5CEE0169800822282AAAAAAAAAAAAAA81EDB192000721996955B57C9";
    attribute INIT_23 of inst : label is "56D1C9D769242DA940152D2E73009612924D2C8665A756D15B93D64126D2485B";
    attribute INIT_24 of inst : label is "A00A969739804B0AAAAAAAAA00000000000000000002AAAAAAAA76D9AC8665A7";
    attribute INIT_25 of inst : label is "73E1823CCCDC16564CB25A11C4511DEF3825EDC046A34C816C818000089216D4";
    attribute INIT_26 of inst : label is "9A76E029DB00969B1890126266E26C313DB00969B7EFB6924999C466DB2C8CDA";
    attribute INIT_27 of inst : label is "B9CF3C67152019A111161642E73DD19C54804BB190120CC7771084E0453B6016";
    attribute INIT_28 of inst : label is "D80668444485B0B9CFF46715E0169C66A616616617EF1DC30898FFCC444585B0";
    attribute INIT_29 of inst : label is "69C6222222C2D85CE7FE33DF00CBA111111616C2E73FD19EE804B8DEB938C673";
    attribute INIT_2A of inst : label is "7679ED3FFDBFDBBCF8E9E6C446F5C9C6339FC032E844444585B0B9CFB467BA01";
    attribute INIT_2B of inst : label is "2332580532EC444B2C664B06490E61C0669B4E6B9111992C029973D83068819E";
    attribute INIT_2C of inst : label is "38820A48270200000659620808071B51111992E031C9264B10269D9E7B4E4962";
    attribute INIT_2D of inst : label is "620808071A20801C71A08200000000640A00000800018A01C70820800068A596";
    attribute INIT_2E of inst : label is "9638820A48270200000659620808071A20800068A59638820A48270200000659";
    attribute INIT_2F of inst : label is "0A52C112D2001DCDA8888CC9701CEA2223325C063A8888CC97018E20800068A5";
    attribute INIT_30 of inst : label is "414141414A0A0AF110011022EA0060ABC6026BE517980000C9CA702C94A6390F";
    attribute INIT_31 of inst : label is "401C608208208233590399A7975AD6529842508435023001094A338CE719C708";
    attribute INIT_32 of inst : label is "0200000000000019028000020000628001C69659659659020800000000000000";
    attribute INIT_33 of inst : label is "60820828820A00828A59659608200000A28E28000200020A28A0020002882007";
    attribute INIT_34 of inst : label is "A28828A00628E58228A31C682408002000200696596480680002100196296290";
    attribute INIT_35 of inst : label is "0000000000000000009659658200808200658A28A28000001A28A28A20820A18";
    attribute INIT_36 of inst : label is "528140A05028140005028140A05028140A05028140A050280000000000000000";
    attribute INIT_37 of inst : label is "0502954AA552A954AA5528140A05028154AA552A954AA05028140A0502954AA5";
    attribute INIT_38 of inst : label is "A05028140A05028140A05028140A0500000A05028154AA552A9540A05028140A";
    attribute INIT_39 of inst : label is "A28A28A28A28A28000028B28140A0502A954AA552A9540A05028140A05028140";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE28A00028A2CA28A28A28";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "4B8F2072094EC432A0B9505878158FC007E2C23FFFF855A908F96C444DEDBBA2";
    attribute INIT_01 of inst : label is "5232480B84596076513904C2AF264408F13543A41090902F2806012695030E02";
    attribute INIT_02 of inst : label is "C0E1B81C3108F24C7F36E828800101208A9540120D54002A12ADD834A231B8D7";
    attribute INIT_03 of inst : label is "1010A2088821524100410000002084A278093B8134E0D28F6400106269D8070D";
    attribute INIT_04 of inst : label is "614B39B3BA011144411141405501154DAF890A1A402996EFBDCB855B85B96C06";
    attribute INIT_05 of inst : label is "40E1483EEE1187280B824A6054C9005820399A242989A04988A088C111A405A9";
    attribute INIT_06 of inst : label is "145140543C00EF800DF001BE0037C006F800CF0019E0033C0027801CC0494E93";
    attribute INIT_07 of inst : label is "51E51479479E79479479E51479E51479E79E79E51479E51479E51E51479451E5";
    attribute INIT_08 of inst : label is "E51451451479479451451479451E51E51E51451E79451479E51451451451479E";
    attribute INIT_09 of inst : label is "9E51E51479479E79479479E51479E51479E79E79E51479E51479E51E51479451";
    attribute INIT_0A of inst : label is "CB02054A651451479451451479451E51E51E51451E79451479E5145145145147";
    attribute INIT_0B of inst : label is "EC9185F1108FA2726C97D139364B09F44E5D64BE89CBAC96BA7722A731A00A00";
    attribute INIT_0C of inst : label is "D0BEDC3479E14579D2BA176950AF953E3A1C0FC3A1D41002F8F625D0AA8411DD";
    attribute INIT_0D of inst : label is "D8945584D000228B149534BFA8865514514936DD8504AB28000000023BBBBBB6";
    attribute INIT_0E of inst : label is "00000000000000000EC826B32112440E04DAD6B49115B0C200132495A5D22A79";
    attribute INIT_0F of inst : label is "CDCCA8241204F80A1004A218CB55F42280000000000000000000000000000000";
    attribute INIT_10 of inst : label is "850360214118110220440981306376664AC00348C909027C108010999B90A42C";
    attribute INIT_11 of inst : label is "4F82C005C008CADF0A0A0245400944AC365DDBD0120037480B6D890D84091285";
    attribute INIT_12 of inst : label is "B87BEFB85A84126410F0419402C060B8CCD2529005A549B1C260AC3FCC925207";
    attribute INIT_13 of inst : label is "735034DACCA09408B3CFCE8292A2DC9281166F651D04960A40E085C02881BAAF";
    attribute INIT_14 of inst : label is "584D144BA572687C940B0B91010122D974AE400F1DCFE6E058F9B2FF33A31EAB";
    attribute INIT_15 of inst : label is "64F0F9DDBE6C45069E4D557ABCFEFA7D3FC9E1F3FBDDFEDF7F9FDA0450F93844";
    attribute INIT_16 of inst : label is "364F0F9DDBE6C45069E4D557ABCFEFA7D3FC9E1F3FBDDFEDF7F9FDA0450F9383";
    attribute INIT_17 of inst : label is "456AE552B954AA552A55EAA752B548A12F8299E1A353A8F66A2D028FC4A0C910";
    attribute INIT_18 of inst : label is "C21A190898AB065B3B0248586CA20915A26C0251253B65CE7B0F486A60800D94";
    attribute INIT_19 of inst : label is "A502090088A0C282831560CB67604528102282488445C6142511288904354276";
    attribute INIT_1A of inst : label is "7069B1B1B1D1114484244B0C1C0ACC8F8426890D3108C17CE902B29650129F08";
    attribute INIT_1B of inst : label is "9B37BCD9B5E364B24A37E36625738D9DEF724E1C0128A0B31884405299B6DB45";
    attribute INIT_1C of inst : label is "768C6B68C68D8CBB2D9632ECB65C336364B611859E4CE1B64A6CDE7366D38D96";
    attribute INIT_1D of inst : label is "4E9B5898832136B0D50D4D9595C4B6B13A6D589888DB57433836E357E6665F78";
    attribute INIT_1E of inst : label is "8DFB50801E38C9060992AA41A1998C21DDDD5FDF9CD887B585F8226DB2D12DAC";
    attribute INIT_1F of inst : label is "0050000CB199B61C18386CC233000CCCCCFB6E0C1D9BB71BF6868E2C0600CDFB";
    attribute INIT_20 of inst : label is "1AE92786D6EF68766C719B61485133B0570FF400008736F8845EDB6D8EDB6DB8";
    attribute INIT_21 of inst : label is "77A3FD1B69858550010E6DF108BC71CF6D8EDB3403C71C0ECD8E71B36F085210";
    attribute INIT_22 of inst : label is "C020029CDBEA1121A00822282AAAAAAAAAAAAAA80A4938000006330E3336C01B";
    attribute INIT_23 of inst : label is "CDB01B77A3FD1B6945410E6DF10896169247618CC38ECDB4EB3676C3EF47F836";
    attribute INIT_24 of inst : label is "A2A08736F8844B4AAAAAAAAA00000000000000000002AAAAAAAA5249E18CC38C";
    attribute INIT_25 of inst : label is "2FE5022DDBDCBEE6EDF4D851547113DEF34DBC0443561C020821A49249FE8DB4";
    attribute INIT_26 of inst : label is "1C5E82317A0897147BA4248623C6547017A089710010412400358CCCF1458D98";
    attribute INIT_27 of inst : label is "B0A75042D5041493333A3746C29D410B54104B47A4248230EFB0802A4E2F4112";
    attribute INIT_28 of inst : label is "8845A4CCCE8DD1B0A75042D5041219FA5A5DA5DA5F24124F6869691CCCCE8DD1";
    attribute INIT_29 of inst : label is "218C66666746E8D853A8217820A69333333A3746C29D410BC104B1DCB80ACC2F";
    attribute INIT_2A of inst : label is "D4D3462012400414C0F1C58CCEE5C056617D482DA4CCCCCE8DD1B0A71042F441";
    attribute INIT_2B of inst : label is "66F4D84432D0CCDB6CDE9B05D99DE08444990CC233337A6C2299643528440134";
    attribute INIT_2C of inst : label is "69C59E31E29E514512202716794284673337A6C221A249D5184D3430D188DD46";
    attribute INIT_2D of inst : label is "271679428459C50A00E51E51451451239E51451C51449E50A01C59C51439E202";
    attribute INIT_2E of inst : label is "0269C59E31E29E51451220271679428459C51439E20269C59E31E29E51451220";
    attribute INIT_2F of inst : label is "2E73F318D4821D2033999BD36110CCE666F4D844333999BD36110E59C51439E2";
    attribute INIT_30 of inst : label is "7676767677B3B2A290312243104E4AB9E24959F9138900001218F339B626AD0D";
    attribute INIT_31 of inst : label is "050A116716716766025949ECE46397729E739CE766262269DEF79CE739CE72CE";
    attribute INIT_32 of inst : label is "9E51451451451448E79451471451279450A10220220220459C51451451451451";
    attribute INIT_33 of inst : label is "11671679E71451679E20220279479E79E79A79451479E59E79E5165145167142";
    attribute INIT_34 of inst : label is "451679E51279A21451440A11E39C51479E59E10220231E11E79E41448850278E";
    attribute INIT_35 of inst : label is "7D3FDFEFA7D3E954AA8220221479C51E51221451451E79E78451451451671461";
    attribute INIT_36 of inst : label is "F552A954AA552A9F4AA552A954AA552A954AA552A954AA552A954AA552A9F4FA";
    attribute INIT_37 of inst : label is "AF57BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEAF57ABD5EAF57ABD5EA";
    attribute INIT_38 of inst : label is "EAF57ABD5EAF57ABD5EFF7FBE9F4FA7D3E954AA552BD5EAF57ABD5EAF57ABD5E";
    attribute INIT_39 of inst : label is "451451479E79451E79E5157D3E9F4FF7FBFDFEFF7FBFD5EAF57ABD5EAF57ABD5";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE51479E51451451479E79";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "4B4BE0E2094A846080904048000007C017E00A3FFFFAD5FB5BFE82666BEB9F8B";
    attribute INIT_01 of inst : label is "42EB686A8C7B60DEC07105C8A60406B9C027C384549494253936C9B6DD241612";
    attribute INIT_02 of inst : label is "50A94A152211B044556C89A0A699453CBC04420A4405039436AFB860B6A1F0D5";
    attribute INIT_03 of inst : label is "1010C4DB364C5B5B6DC00000000005247168350D2943028A908811C2526A854A";
    attribute INIT_04 of inst : label is "2001000030001450514151550404140DB8952E3A6E1D5C2D198BDAA0CD1F0855";
    attribute INIT_05 of inst : label is "00C00010E4000608090000400183000000300000030000408000004000800400";
    attribute INIT_06 of inst : label is "8A28A04560006C00058000B000160002C00058000B000160002C000580000800";
    attribute INIT_07 of inst : label is "28A28A00A00000000A00A28028000A00000000000028A28A00000000A28A28A2";
    attribute INIT_08 of inst : label is "A28A28A28A00000028028000A00000000000028000A28A28A00000000000028A";
    attribute INIT_09 of inst : label is "8A28A28A00A00000000A00A28028000A00000000000028A28A00000000A28A28";
    attribute INIT_0A of inst : label is "D9070DC8628A28A00028028000A00000000000028000A28A28A0000000000002";
    attribute INIT_0B of inst : label is "7D210104600AE5311D2562988E920158A624E92B94C49D24C0021EC615481E88";
    attribute INIT_0C of inst : label is "969950D9C54399CB144A944954B899A2A284CC5A28599002B0A04D14CC861178";
    attribute INIT_0D of inst : label is "01847794556FFE6B72D49368ACDC539E7924924DC077D24BBBBBBBBDC4444224";
    attribute INIT_0E of inst : label is "000000000000000009AE4391099B74931698C631B795B4D64B13B6D73BDD6C7B";
    attribute INIT_0F of inst : label is "444439B69A48108E724EA4CEEA08281360000000000000000000000000000000";
    attribute INIT_10 of inst : label is "9525A4E54EE0E01C0380700E005411006FC924E118452408539252888884F4A4";
    attribute INIT_11 of inst : label is "010B4925A346EA6A4C8E5249CCDB043C9E0EA8E0936495094C20BD2E94923A96";
    attribute INIT_12 of inst : label is "1251541257C892740251861862A26CA0C4105299242508A45220ED1A441B7A48";
    attribute INIT_13 of inst : label is "6021980A47A44E0191454392DAA26409C03225231726D34F49310504F90CD014";
    attribute INIT_14 of inst : label is "FA1D3EDFEFF77AFDD4AA5D3A954AA552A954AA5723D1E8E5526CFC5A6D1E93FF";
    attribute INIT_15 of inst : label is "4EA552A954AA552E9F4FF7FBFDFEFA7D3E9D4AA552A954AA552A954AF5FBF9B4";
    attribute INIT_16 of inst : label is "F4EA552A954AA552E9F4FF7FBFDFEFA7D3E9D4AA552A954AA552A954AF5FBF9F";
    attribute INIT_17 of inst : label is "DF4FB7FBEDFEFF7FBF9F4FF3FBE9F4FB7FAA854BF6F97DBCDF7FABD16AF5F3E9";
    attribute INIT_18 of inst : label is "605E5D288CAD37590172E96965E74826A56136C1053960E73007E80624D925D4";
    attribute INIT_19 of inst : label is "A7804D2C8CACB2979195A6EB202E453C0232B26964654594B527A13D40AF8F2C";
    attribute INIT_1A of inst : label is "C0A9A5A5A311680E94B4C260584E469425330D27132908D42D229AD753360248";
    attribute INIT_1B of inst : label is "0205F01027BA46BA6AA42A45385AC956B4F48AD2934190B139B45A50C9A69AE8";
    attribute INIT_1C of inst : label is "69294A4A94A928220904A08824120A4A4825D0751448912E68081740409AE91E";
    attribute INIT_1D of inst : label is "6D5B60DF6B1D9636C86C25FDFD88B6C1B56D80DF6E994C0220A49A22543425AD";
    attribute INIT_1E of inst : label is "193A51860E28A089313A22D96531365F1312A000D09100A101080465BEE22DB0";
    attribute INIT_1F of inst : label is "49349205931164CA24C1299DA2341998889AC91260B2343234838A244220591A";
    attribute INIT_20 of inst : label is "917E6D04BC3A904449291254A52B6D203525235FF5F4248408AA4924AA49249A";
    attribute INIT_21 of inst : label is "B4924A925D0507EAABA8490C1151451D24BA495095545008892549224BE52944";
    attribute INIT_22 of inst : label is "BFD555D09210222CE00822282AAAAAAAAAAAAAA82A497C92490492A92A24A812";
    attribute INIT_23 of inst : label is "892E12B4924B9256AFFEA8490C11131E925C0124AA4A892E9A25749945249524";
    attribute INIT_24 of inst : label is "57FF5424860889CAAAAAAAAA00000000000000000002AAAAAAABD24A8124AA4A";
    attribute INIT_25 of inst : label is "29030655D84134D4C9AC90721C8726B5AA4923089AF248F49262A4925125C92B";
    attribute INIT_26 of inst : label is "C8518441461112163935B6E400406412046111214DB4DA4DA621088A91450D5E";
    attribute INIT_27 of inst : label is "3030C082BFC8368322220640C0C2020AFE20C963B5B694A6F7008C304428C222";
    attribute INIT_28 of inst : label is "4009A0C88881903030C082BFC832C8F212092092086DAA4769681B68C8888190";
    attribute INIT_29 of inst : label is "2CE866644440C8181860414E41B4833322220640C0C2020A620C9116AB0C8408";
    attribute INIT_2A of inst : label is "40414429A49B69366651450888B558642043104D20CCC88881903030C0829883";
    attribute INIT_2B of inst : label is "448490889250CCDA68929B0FC3E908088A4964852222424844C92BB438620410";
    attribute INIT_2C of inst : label is "79C51451451479E79C51671451E514322224248444A36D1701041010510895A4";
    attribute INIT_2D of inst : label is "671451E51451679451E51479E79E79C51479E79679E71479451C51679E514516";
    attribute INIT_2E of inst : label is "1679C51451451479E79C51671451E51451679E51451679C51451451479E79C51";
    attribute INIT_2F of inst : label is "0739B81ACE805CA41911121242224644448490889191112124222651679E5145";
    attribute INIT_30 of inst : label is "7676767677B3B32290392273BA4A448AEC104AFD93B000005B5EC168B2AE4CA5";
    attribute INIT_31 of inst : label is "451E79E71459E73650596CC8E5731392CEF7BCEF23272269CE739CE739CE72DE";
    attribute INIT_32 of inst : label is "1479E79E79E79E71451E79E59E79C51E79451679C51679E79C51451451451451";
    attribute INIT_33 of inst : label is "79E71451459E79E79E79C51679451451451451E79E79E79E79E51651451459E5";
    attribute INIT_34 of inst : label is "451451479C51451451451E79E79C51451451451679C51451451479E71451679E";
    attribute INIT_35 of inst : label is "2A940A0552A9540A059679C51451679E51679E79E79E79E79E79E79E79E71451";
    attribute INIT_36 of inst : label is "0028140A0502814AA552A954AA552A940A05028140AA552A8140A0502814AA55";
    attribute INIT_37 of inst : label is "0000140A05028140A05028140A05028140A05028140A00000000000000000000";
    attribute INIT_38 of inst : label is "00000000000000000005028140A0502A9540A050280000000000000000000000";
    attribute INIT_39 of inst : label is "00000000000000000000012A954AA5028140A050281400000000000000000000";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00028A00000000000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "31032240E001801F7F6FBFB3FFFFF83FF81FFCFFFFFF23A9E5FF46E2C9F9C9B8";
    attribute INIT_01 of inst : label is "0920012010C92212412073C0AE6707B4570C19111444C6108491309244DA6D68";
    attribute INIT_02 of inst : label is "50ADAA15B90499C3D480471A7C6438826CC98BE37910578A591D516639509845";
    attribute INIT_03 of inst : label is "3210DB04C131C0208240000000208E09208D9111E084582600011E698868856D";
    attribute INIT_04 of inst : label is "9FFCFFFFEFFE40550154015405501570C8459C35955EE4151699D5D1C509AC1C";
    attribute INIT_05 of inst : label is "FFBFFFEF1BFFFDF7F6FFFFBFFE7CFFFFFFEFFFFFFEFFFFBF7FFFFFBFFE7FF3FF";
    attribute INIT_06 of inst : label is "9E79E5989FFF9BFFFB7FFF6FFFEDFFFDBFFFB7FFF6FFFEDFFFDBFFFB7FFFE7FF";
    attribute INIT_07 of inst : label is "79E79E79E79E79E79E79E79479451451451451451479E79E79E79E79E79E79E7";
    attribute INIT_08 of inst : label is "E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E51451451451479E";
    attribute INIT_09 of inst : label is "9E79E79E79E79E79E79E79E79479451451451451451479E79E79E79E79E79E79";
    attribute INIT_0A of inst : label is "9C0398E1279E79E79E79E79E79E79E79E79E79E79E79E79E79E5145145145147";
    attribute INIT_0B of inst : label is "25B1EF37D04681845DB750C22EDBD8D43082EDBA06105DB730201F2949140F2F";
    attribute INIT_0C of inst : label is "0D48D83B49C1B7050184CC041A481A616003A406003B43FD84E2AF20D04748C8";
    attribute INIT_0D of inst : label is "0C8123C30398032019C3BFEA2E432D04109249244491FF7BBBBBBBBFFFFFFE00";
    attribute INIT_0E of inst : label is "00000000000000001884989104400A484858C630004A4A07298C58D8C0E47291";
    attribute INIT_0F of inst : label is "4444069055204261892229222020809D00000000000000000000000000000000";
    attribute INIT_10 of inst : label is "62D9BB38B000000000000000012233330036D823082290212C492D8888820B64";
    attribute INIT_11 of inst : label is "04242492562A2102E56129346324BC0A42248C1A489041B620B862D06B62C168";
    attribute INIT_12 of inst : label is "0310154332934D1149236D271831026A4131084411B39E602981F9CA44490522";
    attribute INIT_13 of inst : label is "009B432E405322A4914540484809946454D2252040924C20A484703204DA1115";
    attribute INIT_14 of inst : label is "A572A9140A0583816AF572AD5EAF57ABD5EAF578BC1E0F17AB954AA552A972AA";
    attribute INIT_15 of inst : label is "AB57AB54EAD53AB940A20000010005028156AF56A954AA752AB54EAF0702854A";
    attribute INIT_16 of inst : label is "4AB57AB54EAD53AB940A20000010005028156AF56A954AA752AB54EAF0702854";
    attribute INIT_17 of inst : label is "50A05028140A05028140A05428140A04503D5EAE552A954AA552BD5EAF572A95";
    attribute INIT_18 of inst : label is "012120826200D10905898404F311049430B2C92F10942252913020921224100A";
    attribute INIT_19 of inst : label is "10A920837203094C4C401A2120B1308569C809041390104A506C836412651224";
    attribute INIT_1A of inst : label is "6824B0B0B94498184B4340841B22416038886099089425543290484028C96866";
    attribute INIT_1B of inst : label is "4B972A5CB1017061001701631E73AD9CE676EC1964964E1086C1253175B6DBB2";
    attribute INIT_1C of inst : label is "6DC621746205CCBB2D9732ECB6597171796319EC8DC6D883012E5C0972C005C5";
    attribute INIT_1D of inst : label is "6C6388DC33C24630E00C920585B4C711B18E08DC3CE425B996B6C39B66666738";
    attribute INIT_1E of inst : label is "A5D31CF3208216E5CC8000041088C514CCCA8008DC5CCEB5EF241390B2CD31C4";
    attribute INIT_1F of inst : label is "003000F1488C9223972DC4609183C444447B25CB9A4BA74BE6082097399925F3";
    attribute INIT_20 of inst : label is "260801F6D428DE35668C8B68421001B437B1B8A2AA37179B8248000008000018";
    attribute INIT_21 of inst : label is "76D96D0B61B1B000016E2F330698618C00180030030C31C6ACD02CB16C400000";
    attribute INIT_22 of inst : label is "D2AAA8DC5E6E09A2000822282AAAAAAAAAAAAAA81800180000734B059116D7DB";
    attribute INIT_23 of inst : label is "45B1DB76D96C0B6005556E2F3304D816000C0CD2C16445B5ABB6364471B2D816";
    attribute INIT_24 of inst : label is "02AA97179B826C0AAAAAAAAA00000000000000000002AAAAAAAA40008CD2C164";
    attribute INIT_25 of inst : label is "79219334CE4436C6CDB058D9364D9AD6B105E5827659E1192D8080000CB605B0";
    attribute INIT_26 of inst : label is "2532C134CB04D94B908200036752D539BCB04D94B6596C96DBB5C46CC411AD99";
    attribute INIT_27 of inst : label is "BDE3727795609B81111A9752F78CC9DE54826CB902004D6021B617333299609A";
    attribute INIT_28 of inst : label is "9826E04446A5D4BDE3327795209A264E2E06E06E04003DC61CB8800C4446A5D4";
    attribute INIT_29 of inst : label is "A21622222352EA5EF1993BC906DB8111111A9752F78DC9DE5836C8CC1DCCF379";
    attribute INIT_2A of inst : label is "0F3C12925B6CB2CB8F8412C44660EE679BCDC1B6E0444446A5D4BDE33277920D";
    attribute INIT_2B of inst : label is "23905826EB24445B6C720B26CC8F25826F7512D71111C82C1375985D8B1993CF";
    attribute INIT_2C of inst : label is "00228A28A28A28A28A28808A28A28B81111C82C13648030106F3C3CF04A45BE2";
    attribute INIT_2D of inst : label is "808A28A28A28A28A28028A28A28A28A28A28A28A28A28A28A28228A28A28A288";
    attribute INIT_2E of inst : label is "8800228A28A28A28A28A28808A28A28A28A28A28A28800228A28A28A28A28A28";
    attribute INIT_2F of inst : label is "12948130E2093E4BC0888E41609B302223905826CC0888E41609B228A28A28A2";
    attribute INIT_30 of inst : label is "0B0B0B0B18585910E01E11BC4433BD01F5BEA1E34FD60000C8CA50A2622B2A5B";
    attribute INIT_31 of inst : label is "000A28A200000080402CBF36B45AD8F97318C6319819D19E6318C6318C631963";
    attribute INIT_32 of inst : label is "8A28A28A28A28A28A28A28A28A28A28A28A28800000228A28800000000000000";
    attribute INIT_33 of inst : label is "28A20000000000000000000228000000000000000000000000028828A28A28A2";
    attribute INIT_34 of inst : label is "A28A28A28A28A28A28A28000000228A28A28A28800000000000000000000228A";
    attribute INIT_35 of inst : label is "57ABD5EAF57ABDFEFF8800000000000028800000000000000000000000008A28";
    attribute INIT_36 of inst : label is "F552A954AA552A954AA552A954AA552BD5EAF57ABD5EAF57BFDFEFF7FBFD5EAF";
    attribute INIT_37 of inst : label is "FF7FABD5EAF57ABD5EAF57ABD5EAF57ABD5EAF57ABD5EFF7FBFDFEFF7FABD5EA";
    attribute INIT_38 of inst : label is "EFF7FBFDFEFF7FBFDFEAF57ABD5EAF57ABDFEFF7FBFDFEFF7FBFDFEFF7FBFDFE";
    attribute INIT_39 of inst : label is "E79E79E51451E79479479F57ABD5EAF57ABD5EAF57ABDFEFF7FBFDFEFF7FBFDF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE79E79E79E79E79E51451";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "01210048C4A5B04000200010000000000400027FFFFEA30091FE0391C8F8C0B1";
    attribute INIT_01 of inst : label is "08A0000010D00014002462B062200124571CB101160404800000B40008020C21";
    attribute INIT_02 of inst : label is "1008A201110299C380804D38540861842CC98B4141145780051910624454AA04";
    attribute INIT_03 of inst : label is "2200C280A2A9C0104540040001000D0431459008E0C258060890C8A0C8408045";
    attribute INIT_04 of inst : label is "4002000020015500015554015000156828020E25419554150689D080570AA41C";
    attribute INIT_05 of inst : label is "0080002000000000020000800100000000000000000000800000000001000800";
    attribute INIT_06 of inst : label is "14514D99C0000800010000200004000080001000020000400008000100000000";
    attribute INIT_07 of inst : label is "51451451451451451451451E51E79E79E79E79E79E5145145145145145145145";
    attribute INIT_08 of inst : label is "451451451451451451451451451451451451451451451451479E79E79E79E514";
    attribute INIT_09 of inst : label is "1451451451451451451451451E51E79E79E79E79E79E51451451451451451451";
    attribute INIT_0A of inst : label is "12031041251451451451451451451451451451451451451451479E79E79E79E5";
    attribute INIT_0B of inst : label is "009CCF371046010050931080284998C4201084980402109230200C210B180C2A";
    attribute INIT_0C of inst : label is "200888384881870700208C001C281961A010040A011803FD84402920CA020880";
    attribute INIT_0D of inst : label is "00800102031A20002183BFEA8451604104000000D003FF7C4444444000000649";
    attribute INIT_0E of inst : label is "0000000000000000180411910D08080808508420020A4C0C28CAD4C4A0944A44";
    attribute INIT_0F of inst : label is "44440002D400404400060004008080B140000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0201800080000000000000000111000100000160286200202000218AAAA60864";
    attribute INIT_11 of inst : label is "0404000160680022C444310513649C0802000050054801B068B8021108000108";
    attribute INIT_12 of inst : label is "420045023011203100304104301004684170000801A2B4603141C10A44002402";
    attribute INIT_13 of inst : label is "00100B2E504206029145440000003440C0122520080001688080602000804145";
    attribute INIT_14 of inst : label is "05028140A05028140A05028140A05028140A05028140A05028140A0502817000";
    attribute INIT_15 of inst : label is "A05028140A05028140A05028140A05028140A05028140A05028140A05028140A";
    attribute INIT_16 of inst : label is "0A05028140A05028140A05028140A05028140A05028140A05028140A05028140";
    attribute INIT_17 of inst : label is "40A05028140A05028140A05028140A05028140A05028140A05028140A0502814";
    attribute INIT_18 of inst : label is "002020004402400905910012E20342500892D9270010200000C1600201520008";
    attribute INIT_19 of inst : label is "03842004440411080880480120B2201C011015002A2000887001800C49608220";
    attribute INIT_1A of inst : label is "2825919191405010094940031363512569A1600300122C543258000024C92054";
    attribute INIT_1B of inst : label is "193320C991033061003203229E212488426264496DB24C100F20163144924960";
    attribute INIT_1C of inst : label is "C4E72336720CE59964B3966592C863233B61981C8C0648850064CC0326400CC4";
    attribute INIT_1D of inst : label is "644100CC198002124024004080900201910400CC0C4005999292491922C2E210";
    attribute INIT_1E of inst : label is "A4D10C7100001654AC8000080088A494C88AAAA24CCAEE94CF24030010440080";
    attribute INIT_1F of inst : label is "003000E1088C924152AD04501143C444447924A95849E349E2000013118824F1";
    attribute INIT_20 of inst : label is "020000F260004E35270489200000049423A09002AA933399814A492488000018";
    attribute INIT_21 of inst : label is "F2C9240920A8A8000166673702B0C30400080010010411C6A4E0249124021080";
    attribute INIT_22 of inst : label is "400000CCCE6E01A4300822282AAAAAAAAAAAAAA80800180000738984911247C9";
    attribute INIT_23 of inst : label is "4491C9F2C9240920055566673700D0D200040CE261244491A993324821924A12";
    attribute INIT_24 of inst : label is "02AA93339B80682AAAAAAAAA00000000000000000002AAAAAAAA40008CE26124";
    attribute INIT_25 of inst : label is "792182B4CE4412626490C81504415842110CE4814600401B649080000C920490";
    attribute INIT_26 of inst : label is "44B240B2C900D12B10810003775695653C900D12B25B6596D994C4644000A488";
    attribute INIT_27 of inst : label is "99E3716795601B81111AB356678DC19E558068B101002D604225033A8259201A";
    attribute INIT_28 of inst : label is "9806E04446ACD599E3706795601A444E2E06E06E0400ADC210B800244446ACD5";
    attribute INIT_29 of inst : label is "A416222223566ACCF1B8B3CB02DB8111111AB356678CC19E481688D830CE4279";
    attribute INIT_2A of inst : label is "0A2802564964B2CA0A0202C446C1867213CCC0B6E0444446ACD599E330679205";
    attribute INIT_2B of inst : label is "2390C8068A244449247219065AA721816B4522559111C864034518594298828A";
    attribute INIT_2C of inst : label is "28A28A28A28A28A28A28A28A28A28B11111C8640B448030402A2828A00944AA2";
    attribute INIT_2D of inst : label is "A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A";
    attribute INIT_2E of inst : label is "8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28";
    attribute INIT_2F of inst : label is "000010C08620384B88888E43205A22222390C816888888E43205A228A28A28A2";
    attribute INIT_30 of inst : label is "090909090848491880989830EF023C00801E20A6870000008180080000282063";
    attribute INIT_31 of inst : label is "A28000008A28A29248249412944A505141084210918318282108421084210921";
    attribute INIT_32 of inst : label is "8A28A28A28A28A28A28A28A28A28A28A28A28A28A28800000228A28A28A28A28";
    attribute INIT_33 of inst : label is "00008A28A28A28A28A28A28800A28A28A28A28A28A28A28A28A28A28A28A28A2";
    attribute INIT_34 of inst : label is "A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A288000";
    attribute INIT_35 of inst : label is "552A954AA552A954AA8A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28";
    attribute INIT_36 of inst : label is "F7FBFDFEFF7FBFD5EAF57ABD5EAF57AA954AA552A954AA552A954AA552A954AA";
    attribute INIT_37 of inst : label is "FF7FABD5EAF57ABD5EAF552A954AA552BD5EAF57ABD5EFF7FBFDFEFF7FBFDFEF";
    attribute INIT_38 of inst : label is "EAF57ABD5EAA552A954AA552A954AA552A954AA552BD5EAF57ABDFEFF7FBFDFE";
    attribute INIT_39 of inst : label is "E51451E79E79E79E51E79F552A954AA57ABD5EAF57ABDFEFF7FBFDFEFF7FBFD5";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE79E51479E79E79E79E79";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
