-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_1L is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_1L is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_1L_0 : RAMB16_S2
	generic map (
		INIT_00 => x"A4809E409E8E69A49A481C209C2085763D217D078EE7890B7B3B8E073C2821A5",
		INIT_01 => x"9C9C6741649107269E8D589A05655BC24EF08E2192238260E49A49A481CE6898",
		INIT_02 => x"425554026C3826820835156EE257589AB59CF0A3B8E65E9C1C6741A49107279E",
		INIT_03 => x"5E43C2CEE3B5A28DC08D1E694269E635642571D989549A59041249787A108D64",
		INIT_04 => x"8D642571D989549A5989A359095C76625526966E6F4E622E628DBB8905555555",
		INIT_05 => x"45C8D050E25A6F99AF89A555555563514539AE9C6BA4119095C4642552696626",
		INIT_06 => x"B9698D69205234AEE38D4228F095554D58DCD4857D35E3735A34905526966341",
		INIT_07 => x"314E680E0E8D8D82238EF4E4E4121BD190BF897945519649188D142219491909",
		INIT_08 => x"04EA71941241D07681CF0A0865555451414DC993514102494463812910BC2068",
		INIT_09 => x"75D64D270825E561541408965C2391C50AE2490555555554A029C650590749DE",
		INIT_0A => x"398D39E9D939B8B16A36A8D989907D88D45555554125947770B9539555550777",
		INIT_0B => x"020E58E5A464164ADA1416DBBDA496810B8249D7945559649FD2E63CE4893929",
		INIT_0C => x"224BE5A46412298160AE48264A4B62359266E4BA7640E5A4652F520580B8E9D9",
		INIT_0D => x"2690B1988D64969204E5A565A6370114D15154AE562592249099573692056259",
		INIT_0E => x"CF08082CA185392919093969196B169A04E63635A481555541C70D0396966A18",
		INIT_0F => x"5639872B6B63B9ACB396B157A20E595C524A4224A5E2C27B009E4F0A324A63C2",
		INIT_10 => x"69259E49AD515B79665054DA49446908655561541408985C24A1C502E2490555",
		INIT_11 => x"515518D105165555049651DDC2C552555A49A68149225492248024B192155796",
		INIT_12 => x"A952692692692692692681555552A79689652A79689671542052A55546351663",
		INIT_13 => x"5825509506962249AA7949A25957095825509A588926A9E52689655C256081F7",
		INIT_14 => x"2E65C7DA79C22D2622E59265C7DCBD88547DC9D73E29C582255549AA7949A259",
		INIT_15 => x"B8A73A6928614F219945042779C6E60A94EA4299A5575369541C799C547D259C",
		INIT_16 => x"27639A7E2F6277FEBDC649FFAF7277FE9DCE69FFAF7277FEBDC649055519F6ED",
		INIT_17 => x"239290E64547D259C09DA4151F727621909026719511625F564A3C99B4957BBE",
		INIT_18 => x"4D246424547D259C2E4E4A65C7DA79C22D2462E59265C7DA79C19DE4971F72F6",
		INIT_19 => x"9254219565C60C126371469E69E6399151830498DC512592598265575A55071E",
		INIT_1A => x"445F71F0C1C0C1409229F26892D22E5925F49B7976935957545A79E599414966",
		INIT_1B => x"8A0F9B9F8A8646464646464444475A55071E4DC65F71F0C1C0C1409229F27992",
		INIT_1C => x"9889B8A9B8A9B8A9B8A9B8AF81F80F8DF8CF8DF8CF81F80F89F88F85F84F9B1F",
		INIT_1D => x"0C843FFFFCC840EFFFFCC840EFFFFFCC843FFFFFCC843BBAA9988BBAA9988AA9",
		INIT_1E => x"400000000FFFC048C06FFFC40C842FFFC7CC842FFFFFCC842FFC048C04BFFC84",
		INIT_1F => x"001D7CE73F9DB0C30000000000000000000000000000000000000000000804C8",
		INIT_20 => x"88EF08EC6061505552524A32B254985458501524156E6974AC62BC234ECA3B82",
		INIT_21 => x"22649559162D9556B55716E15B5D2BA8AE64A264A664A26493595555535053DB",
		INIT_22 => x"62D95555615559D5B5D4F56BE52EA82649559162D955555554F955B5D4BAB935",
		INIT_23 => x"392944506F7E56525D264D227089C022508E35D9B37A94A08E0E984ACA9AE251",
		INIT_24 => x"79939A5A7DB855D264D224662424E4A401B66E89245B62661444169B1B194A49",
		INIT_25 => x"6A654455545557EF0BEEE4169B192426F5D264D227E4A76662671A45BA99B719",
		INIT_26 => x"9699909EB36A15F6B815D264D225642401B76E89245B627615E6994D46427A7E",
		INIT_27 => x"2E91A51B15246C971B421818D0626494EA76498BA57089C022508E06D6929593",
		INIT_28 => x"7B4EE9926DE4E95A7914EF9E753B47154AE4518043C924138A18228D67195114",
		INIT_29 => x"9551D955D935925924904509925A4E4D397793BE6646424E7A4A666DBF62C111",
		INIT_2A => x"769E8916149B9A9445EDBF6EE4254A62DC84254A62DC84254A62DC8551D9551D",
		INIT_2B => x"69F5A717D266D2565256A6719627899A9489A249212B9AE5434A796DBF6249A5",
		INIT_2C => x"4271941190919C652A2E6989DD6198B062E1925B9AC1AB249ABC2AB180001A79",
		INIT_2D => x"81ECB1A65D2264662424E4A511413929CBE62726722506A2C6493489034898B6",
		INIT_2E => x"6056D9226DFADD94A62426D6602762241E627617E66976F515D89049B5DD9506",
		INIT_2F => x"0000000000000000000000000000000000000000000000000004DE09B6489B42",
		INIT_30 => x"D9CBE18525605E67E24D5345534D53533322C959588763F3BE624174AF98905D",
		INIT_31 => x"F995A9947272C9E1855434259520D914A2715C99C89C82C8E7FFDE6D64DB936D",
		INIT_32 => x"97D21EEED55AC5A3EDA9B158CB62AA72C992C828A72C892C8E565FD97A997C65",
		INIT_33 => x"99CE4E698939291909A854AA655F574D57D477642C4559F2C5B5E56448905D55",
		INIT_34 => x"1B6798986626E2E9AAE94D36E74993489BDBBA49284D66615999AAE614646488",
		INIT_35 => x"F89D49B9115155563A66F0BA6F29BBC25D264D22565E4652425E1E04AEC925D4",
		INIT_36 => x"E9546421076231B0AE6E0BD99E1504208AD82425E5D86709E185F59B42DA541E",
		INIT_37 => x"896662401A194909C65046427194AFBE62726722529EBA986D89169B7AA66199",
		INIT_38 => x"09081D651242E194203490490B825263243741E2643741E22547151A990999D4",
		INIT_39 => x"924ABAA204E9C1890628AA3922E26AA3EA6A3BAAE205289961614AF0B4D35826",
		INIT_3A => x"28559A9C12820525A70810824902C262A7E266AA28AA7922E28D4A7062498AAA",
		INIT_3B => x"00000000000000000000000000000000000000000000000000001DA345E98585",
		INIT_3C => x"13D0F92E739124F18B5E00000000000000000000000000000000000000000000",
		INIT_3D => x"893B93E4F9391393E4000009394E4339CCE71390CE7339C0E403904F403900E4",
		INIT_3E => x"000000000000000000000001B4D6208E00003E4E00003E4E000002C402013213",
		INIT_3F => x"175D73DD00000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1L_1 : RAMB16_S2
	generic map (
		INIT_00 => x"3B90E0F8E26F89C718600C3436348B4D9A22CB3ED0310D9D198C520C18A83387",
		INIT_01 => x"348CCD883C762314884B38C24303118A80628233AC3100383B945104002F8878",
		INIT_02 => x"05DDD888361043A3088B1067D3C438C23E70E2A8C521C8348CCD883C76231488",
		INIT_03 => x"C4938AA314B843CBFECBC60323081D2D1D1EF0474734F3C71CFB17232802CBB0",
		INIT_04 => x"331F1EF0C7C734F3C702CC8787BC21E1CD3CF1C471F3CE33CE4B1BCF4377560C",
		INIT_05 => x"C464B434F3C4308C608C2775600CC0B10F079A6C249900707BC01C1CD3CF1CEF",
		INIT_06 => x"C7C74B71C0312D431490C33862A00CC74830748BBC1D20C1D215A40D3CF1F2EA",
		INIT_07 => x"86DC3267DE4BCB831498CDAA18FF7337AB728CF3637077D740D76E8337379797",
		INIT_08 => x"01CBF33887C0A23480062A0CE7756DD8D4F32F70D8C0CDF74D440010C238A3ED",
		INIT_09 => x"CC73C73D8EC353471EB98C0F3E37B82B6FD3C883775600CCC9AFCCE21F0288D2",
		INIT_0A => x"174B3737F7C740D7712D4CB50CF8D74CB8377560C73C76CCD8FCF79D803364CC",
		INIT_0B => x"83EFB8DCDCDCFF27A80C0AB69A888AAC8C41CF4F3437077D7728D198AA082727",
		INIT_0C => x"499A1F1C1CFB30CF3CF3B88343B9A35DF5D8388DFDE8DCDCDE8CEA3FD8C637F7",
		INIT_0D => x"3880D760D77D7A2800DDDDDD1F2CAFAC3010FBB1E499A499B0CF1DCA2802499A",
		INIT_0E => x"6E1A8C2CB18B07070707373737A30A24031F2D2D4500600CEF5CA7A37B2C8870",
		INIT_0F => x"83371CB2D2E0C6270BFBB7DDE3AFB98CCDF1E8DC1C03EB09ABC2AE1B8DD1E986",
		INIT_10 => x"4264224225D7AADF5D75EAB7D707AA0CE580C71EB98C0D3E3BB42B6FD3C88375",
		INIT_11 => x"E38038F3224E15831CF1DB3363F3EE7628A2480082036820333473A0EE8E0426",
		INIT_12 => x"B8E882C920A24B2882C9147580E07D7B1F5E83C790F1DBB6320EC375BC3E38F3",
		INIT_13 => x"B23EE8FB2F4EA38283C792C3C7EC8FBA3EC8FD3A8E880F1EC90F1FB23EE8C4E1",
		INIT_14 => x"31A79F3BE7E3DC1E63CDF5E79F32EB3A79F32EBEE4EA07633E03A203C7B243C7",
		INIT_15 => x"E01D3F8F11C7D10ACF1E113AF427F29F423F28CFD15ABCEB1C78FCA279F3BE7E",
		INIT_16 => x"3AD27BC03ADBAC22EB49EF08BAD3AC22EB49EF083AD3AC20EB49EF0180071F07",
		INIT_17 => x"E3737C33F7DF3FF7E1F52A9E7CCBACE3737C73F7DF7DC281C7FCB9CF1DF62C40",
		INIT_18 => x"33CCDCDE79F3BE76318DCDE79F3BE763DC1FA3CDF5F7DF3FF7E1F52A9E7CCBAC",
		INIT_19 => x"F5D433A0238DB99CCEF3DBFDEF9D8CF8E36E6733BCF6FF7BE7673D5ABAC71E3F",
		INIT_1A => x"9E7CC893A29BAB98F4637149F1F63CDF5E1DF1CF1CF1CF8175EBE77D75D7AF9D",
		INIT_1B => x"DD0FCCCFCCC98A9BA8B98A9B9B9ABAC71E3F339E7CC893A29BAB98F4637149F1",
		INIT_1C => x"DEDDDDDCCCCFFFFEEEEDDDDFC4FC4FC8FC8FC0FC0FCCFCCFE0FE0FDCFDCFDD0F",
		INIT_1D => x"95554FFFFD99994FFFFD99994FFFFFD1111FFFFFD1111CFCFCFCFFEFEFEFEEDE",
		INIT_1E => x"000000000FFFD111155FFFD551111FFFDBD9999FFFFFD9999FFD5555998FFD99",
		INIT_1F => x"0063C92C3C124B24000000000000000000000000000000000000000000008400",
		INIT_20 => x"0C062824E0F0B21B02E100F393D4E486323E733D7332CB0C84E238AFC04E08CA",
		INIT_21 => x"4F3CB10F022EC0004C00000C25F83128E73CEB3CE33CCF3CB30F001003020022",
		INIT_22 => x"22EC0000119991825F4007293C04A8F3CB00F022EC0000000100025F0112A36C",
		INIT_23 => x"37379E7032F1C1C1D797D797CADF6CB7EA4A9FC219D48C8180C221C88A2B3020",
		INIT_24 => x"E19D77E1EF3179797D797E1F5C1D1D1D871C2FC73C0C15C45C88F7213975C617",
		INIT_25 => x"CF1CCC81EC01DCEE28C4A8FF11385C1F2D797D797F1F1D1C637DB1CB00CF4D75",
		INIT_26 => x"7870747319C48D42CC09797D797C1C1E871C2FC73C0C15C85E6C76C385C5F1E1",
		INIT_27 => x"60760761FC9D86F805CA030A710C5DFA38D5DF38050ADF6CB7EA4A8FC0737374",
		INIT_28 => x"C1D6FD77C73D41E1EB2DC7F9DF799EF0D0A0EFEBD447BDC71C71C0873E79E79C",
		INIT_29 => x"94119502071CF2CF1CF21048F3E1CDDB171DF59FC1C5C5C1C1CDDDC7C1D70975",
		INIT_2A => x"1C5DC70080A47475D707C1DD3CB46F2B4EC1B8AC3B82D2BCED0BC6E0191D815D",
		INIT_2B => x"87CE1F387D7C77D1E1D033E79CE41CFA700DEB080C210F1CE0C5C5C7C1F1C0C0",
		INIT_2C => x"C1E79C02727475D71985DF60C71CF698D859F5E20D88491EF438A413800021F7",
		INIT_2D => x"CF751381D7997C5D5C1CDCDE79C0272759DF3F57D97E3DD84E175E5FA5E5F413",
		INIT_2E => x"E1787E13F873C4F91D5C1C73C81D273C74D5D05DC3CF9842747C710FD26BD23D",
		INIT_2F => x"000000000000000000000000000000000000000000000000000871CF1F84FD15",
		INIT_30 => x"7EC5118B1C222D7C57E72AEB2AEB2AC9B982284F8CEC3B3A9DF3E3D2477CF8FC",
		INIT_31 => x"80780CFAA8A228118B8E0C1E5E3B0D2EA1F22E5F65FE4E64A80028E38E34E5F1",
		INIT_32 => x"E0E0AEF34563DE8E3F0857A385C200D1E5F1E4E00D1E5F1E4A81E80790CFA01E",
		INIT_33 => x"FB00C2B0CF17171717B17B0CA8B02C8C2C0B9BAB22818E43C910DD7AD4F8FC80",
		INIT_34 => x"71E0232B1F5C4C6A1C68C30065E5F5E5FCBA3F8F1F177E05E232AE4ABC0C298C",
		INIT_35 => x"3C7C001A322001DE08E2E2B1E007B98A9797D797F1F1D5C5C1C0C23FEE47BF88",
		INIT_36 => x"B3788C8E028BF2928CCE12983406206306A0CCE8DC7E3C8F118B5CF5CA817877",
		INIT_37 => x"4F81D5E8F74717079E7009C9D75C681DF3F57D97E37B8FFDC7C703FF2233FC77",
		INIT_38 => x"8CAD975D73CBDDF2B65D75CF2F77CDC1FD1AF8D97D1AF8D97E0C83E0CFF0FEC0",
		INIT_39 => x"BC70208C4323503210E00EC1C08288FD08CAD928434BC3CF9208F0E2BA438CDD",
		INIT_3A => x"100F3A340184238D8D18030AC1CC8E84BC041F2C6106C1C48613F8D000800800",
		INIT_3B => x"00002AAA8A8AA0A0800022A2BFEAAAAAAA829DDDF311003F4015E4CB8B2E4822",
		INIT_3C => x"23F0FFEA9955400000002AAAA8A88080A8A8A0200888A8A8A222020200002222",
		INIT_3D => x"0A940300C00014030019551FEACFF23AC8EB33FC8EB23ACCFC33F08FC33F0CFC",
		INIT_3E => x"00000000000000000000000187981082000183C2000183C20000000000210003",
		INIT_3F => x"0000093C00000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1L_2 : RAMB16_S2
	generic map (
		INIT_00 => x"30F8C7F8C76F0C2082082232F632C0B080302031C732CDDF2D8C878090B230E0",
		INIT_01 => x"6C171B002C950910E0C390CB0B29B10B0042C030C333C33230C6186182AF0EC2",
		INIT_02 => x"03EE404F313CF3233E4706C7E3EC90CB8202C2C8C87B216C171B002C950910E1",
		INIT_03 => x"CBCB0B2321CCB3C332C3CB2F232C3F0C3435790D0D9840C320C70F2F2C06C370",
		INIT_04 => x"B03C3DF90F0FB8404180EC0F0F7E43C3EE10106433736C336CC183CD09B99026",
		INIT_05 => x"C12C30B2F3CB380CB80CBB9901A6E450680D38DE4E3410F0F7E43C3EE10106D3",
		INIT_06 => x"0DCD410820A9060321C6430C42C1A6CD2F98D2F57534BE634BC2D0661030F0E5",
		INIT_07 => x"CA073323C7C1C16321C670622CC719C188890EDC0BB0D04180E0A0730D0DCDCD",
		INIT_08 => x"0653DC6020409090C1242C8C3B990A02C66C14D302C2C34990618238A2F0B31E",
		INIT_09 => x"64F34F358F2B098F3F748C51B231C2D723E3C10BB9901A6CCC8F718081024243",
		INIT_0A => x"0D410D0DCD0DB0E091068C190DD82820109B9902C80C3DEEC8EEF1EC069B92EE",
		INIT_0B => x"232F0C343534C773C274206A102410B08C87512DC1BB0D041902D880B08A0D0D",
		INIT_0C => x"310E363574CB0CCC32730C33230E4380106131C37344343534270231E8CB0DCD",
		INIT_0D => x"71E8E080E00410820834343477056C80C086F0D74300C300F8DD76408208310C",
		INIT_0E => x"2C1D8CF6B2C01D1D1D1D0D0D8D0B208209340404618281A6EC806810D0C31DD7",
		INIT_0F => x"230D34404048C83B48D0CD36C32F0E2F0343443534F33B3C5FCF2C1E43534A0B",
		INIT_10 => x"1C31C31C334D418924D35062496F0A8C391ACF3F748C51B230C2D723E3C10BB9",
		INIT_11 => x"2406600E205AA40B2030F7BB238BC3B0820820821C3381C332F332C8C38061C3",
		INIT_12 => x"EECE38A28A18608208E3AAB91ACE2CB28B2CA2CB28B2F772304B9BB909024080",
		INIT_13 => x"723DC8F76E6E432862CB1822CBDC8F723DD8F8B90C208B2CE38B2F723DC8C1C2",
		INIT_14 => x"32CD35C2492320764370104D35C2C118D35C2C148C6A1D23746B38E2CB28A2CB",
		INIT_15 => x"E874BF11075D5ACBD17514B06223988EE63898CDAA420B283CF92AA0D35C2492",
		INIT_16 => x"B048D369B04B06A0C1234DA8304B06A0C1234DA8304B06A0C1234D05061D378D",
		INIT_17 => x"60D0D6334D35C24934D03534D70B0460D0D6334D34D34A03C370800D3CD06668",
		INIT_18 => x"AC903434D35C249632C3434D35C249632076C370104D35C24934D03534D70B04",
		INIT_19 => x"925830C24D34B0BD859C045149268CD34D2C2F616701145249A336420A0F3E4A",
		INIT_1A => x"34D7080B080B3748D4B6E20C512C3701043CD3CD3CD3CD24D3514524934D4514",
		INIT_1B => x"004F000F000332211100033221120A0F3E4AAC34D7090B090B3748D4B6E20C51",
		INIT_1C => x"21211111111000000000000F04F04F00F00F04F04F00F00F14F14F20F20F004F",
		INIT_1D => x"44444FFFFC88888FFFFC88888FFFFFC4444FFFFFC44442222222212121212121",
		INIT_1E => x"000000000FFFC888888FFFC888888FFFCFCCCCCFFFFFCCCCCFFC4444444FFC44",
		INIT_1F => x"00A2CA243C820B280000000000000000000000000000000000000004C4840000",
		INIT_20 => x"CF042F0C38157055123CB51D33500051B39C30BC303D34C3CC3F30BC30C3C0C3",
		INIT_21 => x"53348D8D33373333B73373F70C3EC30F03370337033713348C8DCCFCCECDC000",
		INIT_22 => x"3373333333FFFFB0C32E1DD3778C373348E8D3337333333333BB30C32D30FCC3",
		INIT_23 => x"0D4D34D0A04343434DC34DC36FCD1BF34F4BE32D3F00A46187C7D3C686D3B183",
		INIT_24 => x"6C3D964D38E1D0D034D03435747434365D370FCC740F87787400C7D30DD7461D",
		INIT_25 => x"6C367846549A670C2F0C30CBD30C747604DC34DC3437343757378D20D0CDF1D7",
		INIT_26 => x"D8D0D0DD3F00E438EC20D034D03436355D370FCC740F877474F34E2003C3F343",
		INIT_27 => x"21DD1DD3D0774DD047430F0F00822491C1B1450B002FCD1BF34F4BF321D0D0D0",
		INIT_28 => x"6370FD965D77074D3C834CDC30C3C3C771F7741D3CE0D0A2CB2CB0DD74D34D34",
		INIT_29 => x"BB3B77700D75D21D31D03EF1D74D03701D75DC33434747474743434DE37385D7",
		INIT_2A => x"3432CC00A3C1D1D75D8DE37234721F87E1F97A5E9769DA729CB7EDFB333FF3FB",
		INIT_2B => x"34B0D2C0FC34F343E3FC334D346D0CD0D3CFD33CFCF3CD767643524DE37300DB",
		INIT_2C => x"474D3420D0D0D75D1B875DE39D2DDE3C382C1040CD0AF3834F30BF30C0000D2C",
		INIT_2D => x"CC7C30C34D0E347474743534D3420D0DC3531043403431F8C31D340D1344DD37",
		INIT_2E => x"59D0DD157AE3ADD0347475D754779375DE077877075D34EB09DCC01DD8F8F431",
		INIT_2F => x"0000000000000000000000000000000000000000000000000001D2DD37011E87",
		INIT_30 => x"DD4422C030B0003603748D348D348D2DCCC23E9D0C380E2E35313CDB8D4C4F36",
		INIT_31 => x"41DC4DDCDFD23A22C0276435243C0F570361440D40D00B00B2AA834D34D64378",
		INIT_32 => x"F0BCFCFB26004BBC071812DF01C619B140D280B19B140D280B07741DD4DDD077",
		INIT_33 => x"DC07C7F0CD0F0F0F0FD1DD4C32C2B045B0ACCFFC23FA0F839E32523E004F3A08",
		INIT_34 => x"D3700F0C35743C3E4C3F0C083340D340D81F3F551D9D770740F0F4C3C03C3F2C",
		INIT_35 => x"8CCC800CE1022667CC38C2F3740DC30B0DC34DC343634747474FCF32FCE0D321",
		INIT_36 => x"E0D03C3D27D7E0E0C3C30AD66C190420C3F03C3035DA779D22C075D743F1D083",
		INIT_37 => x"55034744C70D1D1D34D083435D746F353104340340DE4CD34DCC00DCB537720D",
		INIT_38 => x"4F7C4D24DF332CDDF134937CCCB3434B34BE312035BE312034745DD4DDD1DDD8",
		INIT_39 => x"B4F3A3860BD2C019046386F3CE8E037C03C3C30C33D5C4CD014E70C2F0000C34",
		INIT_3A => x"182FFC6C51861BBE1B185186C3C6860B3C0B0F4CB38AC3CE8E32D4B00A4128E2",
		INIT_3B => x"8FCFE02000002B2B2EEEEC2C000000000000130C7351400C40110CC6D74C0538",
		INIT_3C => x"23ACFFC0000000000000155566664F0F2E6E6EEEC30322222CECDCDCCFCFE8A8",
		INIT_3D => x"AAAAAB00D5400003AA8C4C4AAA8EA23A88EA23A88EA23A88EB23AC8EB23AC8EB",
		INIT_3E => x"0000000000000000000000008F8C6CF3000043F3000043F30000000021000003",
		INIT_3F => x"30C30E3200000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1L_3 : RAMB16_S2
	generic map (
		INIT_00 => x"3800E000E00F82082080003900390F0C1E03C73C240A000EA00CE43C1E003A03",
		INIT_01 => x"7803DE001C140108074F1CE8A3A31DE0CF780F3A2009280038208208000F8130",
		INIT_02 => x"00FFFC240092400390F3007331C71CE83C307800CE41C77803DE001C14010807",
		INIT_03 => x"E841E0033916808F404F28A003A00F3E0E0CFC8383FCF1C73CF003A0A0004F00",
		INIT_04 => x"2E0E0CFC8383FCF1C72CCB83833F20E0FF3C71C731C1CB31CB4F3FC7A3FFFFFF",
		INIT_05 => x"C004FA30F1E801CE81CE8FFFFFFFC3301303000F0000003033F00C0FF3C71CB3",
		INIT_06 => x"0303CF8200013C733924F3A3783FFFC7A1307A133C1E84C1E85A003F3C71F3F0",
		INIT_07 => x"32E40003248F8F0FF9243E4034F090F900D3CFDF83F031C70CC72E4003034343",
		INIT_08 => x"00B34F7001C0C0180047810E8FFFF0E0E4CF0033E0C040C70E490080083E03C0",
		INIT_09 => x"CC71C71C0DB30FC71F000C02003904C30371C083FFFFFFFC000D3DC007030060",
		INIT_0A => x"03CF0303C3030CCF2D3CF4F2CC70C304F83FFFFFCF1C7C0CC0C4C93FFFFFC0CC",
		INIT_0B => x"030F800C0C0CF007601C0870DE0008100CC0C77DF83F031C70E0D01E08080303",
		INIT_0C => x"03800E0C0CF0A00F000382800380331C71CF3800F0C00C0C0E03E03C00CD03C3",
		INIT_0D => x"3800CF1CC71C7820000C0C0C0F3D0F2CF020C800E038203810C70C3820020382",
		INIT_0E => x"07800E40B80F03030303030303838820000F3F3E0800FFFFC33C0B0038208030",
		INIT_0F => x"F0030C23E3C0CE03C0B8030CF30F83F3C0C0C00C0E8003A000E8078000C0C1E0",
		INIT_10 => x"8208208201C721C71C71C871C709800E8FFFC71F000C0300380CC30371C083FF",
		INIT_11 => x"C3FF0CFB12033FFF3C71F033032320FFE08208008200F8200A003A00E03FF820",
		INIT_12 => x"04E4924924924924920800FFFFE01C78071E01C78071F030302813FFC33C7C33",
		INIT_13 => x"3030C0C3008C339241C79241C70C0C3030C0C230CE49071E08071C3030C0C03A",
		INIT_14 => x"33471CF1C703340CB37C71C71CF04F9071CF04F33A42C3031FFF9241C79241C7",
		INIT_15 => x"540C3D0700C35002470C0013C403000CC03300C723FCB3CB1C70C42C71CF1C70",
		INIT_16 => x"13C0B1C013C13C0B4F02C702D3C13C0B4F02C702D3C13C0B4F02C703FF031D07",
		INIT_17 => x"40303031C71CF1C70876001C73C13E40303031C71C71E4F1E1F01C071C7FF440",
		INIT_18 => x"0F2C0C0C71CF1C703340C0C71CF1C703340C737C71C71CF1C70876001C73C13E",
		INIT_19 => x"71FF3A3FC71C1C25E5CF5071C71C0C71C707097973D41C71C7031FFCB2C71C31",
		INIT_1A => x"1C73C1C1C1C1F000D6479080704B37C71F1C71C71C71C7FC71C1C71C71C7071C",
		INIT_1B => x"330F330F3309999999999888888CB2C71C310F1C73C1C1C1C1F000D647908070",
		INIT_1C => x"33333333333333333333333F00F00F00F00F00F00F00F00F30F30F30F30F330F",
		INIT_1D => x"44444FFFFC44444FFFFC44444FFFFFE6664FFFFFC44443333333333333333333",
		INIT_1E => x"000000000FFFC444444FFFC444444FFFC3E2220FFFFFC0000FFC4444444FFC44",
		INIT_1F => x"002C32C33F0C33CF000000000000000000000000000000000000000400000000",
		INIT_20 => x"00B780BA84F33033F3D20701E1FC00083933CB01CB01C32C3A80DE02CBA82CE8",
		INIT_21 => x"331CF00708C0C88840880840B0C83E90F31CF31CF31CF31CF3072202232223F9",
		INIT_22 => x"8C0C888880CCCC4B0CC1C31E1C7A4031CF10708C0C888888884C8B0CC0E9033C",
		INIT_23 => x"03031C7233C0C0C0C7F1C7F1F1C70C71C1E01CC0E2C28ECB2C2C0E6C2C0E1B30",
		INIT_24 => x"C2E471F3CB1C3C731C731C0C0C0C0C0C031C7F4F1C0100C70CCCF00EA071EC03",
		INIT_25 => x"C00FEC0FCCCFFC37803A4CF03EA00C0F3C7F1C7F1C0E0C0CFF1C33D32CC70C71",
		INIT_26 => x"30303033E2C24F4F86CC731C731C0C0C031C7F4F1C0100C70F1CF2D3C0C0C0C0",
		INIT_27 => x"C031C31E0C0C787E31ECB0B0BB241C702DE1C790F3F1C70C71C1E01C40303038",
		INIT_28 => x"C1CBF471C71CF0F3C74C7870C31E2CF1C791C303C3932E4924924B071C71C71E",
		INIT_29 => x"0080000B031C73C73C700C3CB1F3C0CF031C73E1C0C0C0C0C0C0C0C741E01071",
		INIT_2A => x"1CF34F024A303031C70741E31C0C020080200802008020080200401084400800",
		INIT_2B => x"CF3F3CFC7F1C71D0D0CF31C71E43CC703A00B3A28289000FF0C0C3C741D3C033",
		INIT_2C => x"C0C71C80303031C7B0B2C72E873072E0CB3471F903E00E4CB0DE00EA000033CF",
		INIT_2D => x"0F00EA00C73F1C0C0C0C0C0C71C803030E7D3D31D31F3C0BA8031CC701CC72E1",
		INIT_2E => x"C03C7401C41C487C0C0C0C71C00C731C31C0C70C72C7C38CBC74F0071387333E",
		INIT_2F => x"000000000000000000000000000000000000000000000000000C73071D007100",
		INIT_30 => x"7442380F3E80361C61CBF1CBF1CBF1F11113C0C7C00300E0E7D3C32039F4F0C8",
		INIT_31 => x"3030CC700303CC380FFF0C0C3F03C30CF2E034C74C74E04E0C0031C71C7471D0",
		INIT_32 => x"0B8787F17FF05C770590171DC16491E04C704E091E04C704E0C0C3030CC70C0C",
		INIT_33 => x"70EC2C3CC7030303030C33CE4F3CCF00CF3332233D23C0B0C2EF7FD2C0F0C8FC",
		INIT_34 => x"31CB90900C0E4241CE43CF0241CC71CC78F1FD0703071CB0F90903A43EC2C3CC",
		INIT_35 => x"14F00093B0033FFCF2CF7800CF033DE0C7F1C7F1C0C0C0C0C0E8283C0B932CCC",
		INIT_36 => x"2C3EC6C400735B1B2424B31F780C02CB2C1EC2CC0C7C2F0B380F1C71EC0C3CF5",
		INIT_37 => x"07C0C0C0F00303031C7200C0C71EC3E7D3D31D31F032CC70C74F00730B31CC03",
		INIT_38 => x"0330072C3C03307CC01CB0F00CC1C0D21D21C8331D21C8331F1C070CC70CB400",
		INIT_39 => x"0399092410F784900249243E6424E403E4243E9240C33CC70024CF783000C00C",
		INIT_3A => x"B001C7780B2C0071DEB00B2C2E6C2CE401E430CE49241E6424970DE224009249",
		INIT_3B => x"703025657575646461212161400000000004030C3300000C00003802C0B80093",
		INIT_3C => x"0300EA800000000000003CC32121307065252121347465656121212130302565",
		INIT_3D => x"A55557AAEAAA8003AA404040000C003002C083000C00B020C083022C083000C0",
		INIT_3E => x"000000000000000000000000390338200000F1E00000B1E00000000000000003",
		INIT_3F => x"0B2CB1CC00000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
