library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic39 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic39 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"12",X"12",X"12",X"7E",X"7C",X"00",
		X"00",X"34",X"4A",X"4A",X"4A",X"7E",X"7E",X"00",X"00",X"24",X"42",X"42",X"42",X"7E",X"3C",X"00",
		X"00",X"3C",X"42",X"42",X"42",X"7E",X"7E",X"00",X"00",X"42",X"4A",X"4A",X"4A",X"7E",X"7E",X"00",
		X"00",X"02",X"0A",X"0A",X"0A",X"7E",X"7E",X"00",X"00",X"34",X"52",X"52",X"42",X"7E",X"3C",X"00",
		X"00",X"7E",X"08",X"08",X"08",X"7E",X"7E",X"00",X"00",X"42",X"42",X"7E",X"7E",X"42",X"42",X"00",
		X"00",X"7E",X"7E",X"7E",X"40",X"40",X"30",X"00",X"00",X"42",X"24",X"18",X"08",X"7E",X"7E",X"00",
		X"00",X"40",X"40",X"40",X"40",X"7E",X"7E",X"00",X"00",X"7E",X"02",X"7C",X"02",X"7E",X"7E",X"00",
		X"00",X"7E",X"20",X"18",X"04",X"7E",X"7E",X"00",X"00",X"3C",X"42",X"42",X"42",X"7E",X"3C",X"00",
		X"00",X"0C",X"12",X"12",X"12",X"7E",X"7E",X"00",X"00",X"40",X"3C",X"62",X"42",X"7E",X"3C",X"00",
		X"00",X"44",X"2A",X"1A",X"0A",X"7E",X"7E",X"00",X"00",X"34",X"72",X"4A",X"4A",X"4E",X"2C",X"00",
		X"00",X"02",X"02",X"7E",X"7E",X"02",X"02",X"00",X"00",X"3E",X"40",X"40",X"40",X"7E",X"7E",X"00",
		X"00",X"1E",X"20",X"40",X"20",X"3E",X"1E",X"00",X"00",X"3E",X"40",X"38",X"40",X"7E",X"3E",X"00",
		X"00",X"42",X"26",X"1C",X"38",X"74",X"62",X"00",X"00",X"06",X"08",X"70",X"08",X"0E",X"06",X"00",
		X"00",X"42",X"46",X"4E",X"5A",X"72",X"62",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",
		X"00",X"00",X"18",X"24",X"24",X"18",X"00",X"00",X"00",X"00",X"42",X"66",X"3C",X"18",X"00",X"00",
		X"00",X"00",X"00",X"18",X"3C",X"66",X"42",X"00",X"00",X"00",X"24",X"18",X"7E",X"18",X"24",X"00",
		X"00",X"00",X"3C",X"46",X"4A",X"52",X"3C",X"00",X"00",X"00",X"40",X"40",X"7E",X"42",X"44",X"00",
		X"00",X"00",X"64",X"4A",X"52",X"62",X"44",X"00",X"00",X"00",X"34",X"4A",X"4A",X"4A",X"42",X"00",
		X"00",X"00",X"08",X"7E",X"08",X"08",X"0E",X"00",X"00",X"00",X"30",X"4A",X"4A",X"4A",X"4E",X"00",
		X"00",X"00",X"30",X"4A",X"4A",X"4A",X"3C",X"00",X"00",X"00",X"06",X"1A",X"32",X"62",X"06",X"00",
		X"00",X"00",X"34",X"4A",X"4A",X"4A",X"34",X"00",X"00",X"00",X"3C",X"52",X"52",X"52",X"0C",X"00",
		X"00",X"00",X"60",X"F8",X"FF",X"F8",X"60",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"00",
		X"3C",X"42",X"81",X"81",X"81",X"81",X"42",X"3C",X"00",X"18",X"3C",X"66",X"66",X"3C",X"18",X"00",
		X"00",X"3C",X"42",X"5A",X"5A",X"42",X"3C",X"00",X"00",X"00",X"06",X"09",X"51",X"01",X"02",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"00",X"40",X"12",X"4B",X"A7",X"14",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"C0",
		X"80",X"50",X"2C",X"54",X"A3",X"04",X"10",X"40",X"00",X"00",X"00",X"00",X"C0",X"FF",X"C0",X"00",
		X"AB",X"55",X"23",X"0C",X"04",X"10",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"C0",X"00",X"00",
		X"00",X"00",X"C0",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"10",X"04",X"0C",X"02",X"AA",X"5D",
		X"00",X"C0",X"FF",X"C0",X"00",X"00",X"00",X"00",X"1D",X"23",X"48",X"0C",X"00",X"00",X"00",X"00",
		X"C0",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"80",X"11",X"2B",
		X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"FF",X"7F",X"7C",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"7C",X"7F",X"FF",X"FF",
		X"7F",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7C",X"7F",X"FF",X"FF",X"FF",
		X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7C",X"7F",X"FF",X"FF",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7E",X"FF",X"FF",X"FF",X"7E",X"78",
		X"78",X"7E",X"FF",X"FF",X"FF",X"7E",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"FF",X"FF",X"FF",X"7F",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7C",
		X"FF",X"FF",X"FF",X"7F",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"7C",X"7F",
		X"FF",X"FF",X"7F",X"7C",X"78",X"78",X"00",X"00",X"00",X"00",X"00",X"78",X"78",X"7C",X"7F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"03",X"0E",X"03",X"00",
		X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"03",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"30",X"E0",X"30",X"00",
		X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"30",X"E0",X"30",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"FF",X"FF",X"03",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",
		X"FF",X"FF",X"03",X"03",X"07",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"03",X"03",
		X"03",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"03",X"03",X"FF",X"FF",
		X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"03",X"03",X"FF",X"FF",X"03",X"03",
		X"0C",X"0C",X"FC",X"FC",X"0C",X"0C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",
		X"FC",X"FC",X"0C",X"0C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"0C",
		X"0C",X"0C",X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"0C",X"FC",X"FC",
		X"38",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"0C",X"FC",X"FC",X"0C",X"0C",
		X"06",X"0F",X"1F",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",
		X"1F",X"1F",X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",
		X"0F",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",X"1F",
		X"07",X"05",X"02",X"02",X"02",X"07",X"00",X"00",X"00",X"00",X"06",X"0F",X"1F",X"1F",X"0F",X"06",
		X"00",X"18",X"3F",X"3F",X"18",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"03",
		X"3F",X"3F",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",
		X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"18",X"3F",X"3F",X"18",X"00",
		X"30",X"30",X"F0",X"F0",X"30",X"30",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",
		X"F0",X"F0",X"30",X"30",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"30",
		X"30",X"30",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"30",X"F0",X"F0",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"30",X"F0",X"F0",X"30",X"30",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"00",X"00",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7B",X"87",
		X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"09",X"01",X"01",X"09",X"0E",X"00",X"00",
		X"22",X"22",X"03",X"03",X"22",X"22",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",
		X"04",X"08",X"0F",X"0F",X"08",X"84",X"87",X"7B",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"FF",X"FF",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",
		X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"FF",X"FF",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"78",X"7C",X"7C",X"7C",X"7C",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"7C",X"7C",X"7C",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7C",
		X"7C",X"78",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7C",X"7C",X"7C",
		X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7C",X"7C",X"7C",X"7C",X"78",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"C0",X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"F0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"30",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"80",
		X"1E",X"1F",X"1F",X"1F",X"1F",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",
		X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",
		X"00",X"00",X"08",X"04",X"08",X"14",X"08",X"00",X"00",X"00",X"08",X"26",X"10",X"26",X"0C",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"2C",X"00",X"4D",X"20",X"14",X"00",
		X"07",X"07",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"07",X"07",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",
		X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",
		X"1F",X"1F",X"1E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"1E",X"1F",X"1F",X"1F",X"1F",
		X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"14",X"20",X"05",X"2A",X"00",X"32",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"C2",X"C0",X"F0",X"3A",X"38",X"0C",X"46",X"0C",X"80",X"FC",X"FF",X"F0",X"82",X"F0",X"38",
		X"05",X"1C",X"78",X"F2",X"F0",X"C4",X"98",X"72",X"3F",X"3D",X"2D",X"66",X"26",X"43",X"12",X"20",
		X"3B",X"3B",X"75",X"EE",X"F5",X"3B",X"7B",X"9F",X"20",X"09",X"2C",X"84",X"44",X"ED",X"6D",X"7F",
		X"E2",X"80",X"0C",X"1E",X"1E",X"8C",X"00",X"00",X"F8",X"78",X"B0",X"60",X"F3",X"DB",X"D8",X"30",
		X"0C",X"1E",X"0C",X"80",X"C0",X"C0",X"64",X"B2",X"77",X"27",X"03",X"20",X"00",X"08",X"1C",X"08",
		X"EF",X"F9",X"77",X"37",X"7C",X"DF",X"EB",X"7D",X"20",X"41",X"04",X"31",X"7B",X"71",X"33",X"6F",
		X"00",X"00",X"04",X"00",X"24",X"0E",X"04",X"00",X"00",X"06",X"16",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"68",X"00",X"00",X"00",X"60",X"F4",X"60",X"00",X"20",X"00",X"00",
		X"B8",X"FC",X"4C",X"F8",X"F0",X"C8",X"C0",X"80",X"FC",X"3E",X"D6",X"DB",X"FB",X"F7",X"FE",X"DC",
		X"C0",X"E8",X"E0",X"70",X"F8",X"F4",X"2C",X"F8",X"9F",X"BF",X"77",X"F7",X"E6",X"FC",X"F0",X"E2",
		X"C0",X"E2",X"B8",X"9E",X"E7",X"97",X"D7",X"DF",X"E3",X"F3",X"7E",X"1E",X"0C",X"00",X"30",X"30",
		X"00",X"C2",X"C0",X"18",X"3C",X"3E",X"62",X"C3",X"EB",X"FF",X"5F",X"DD",X"C3",X"B2",X"BE",X"1C",
		X"1C",X"BD",X"E7",X"E3",X"D9",X"FD",X"FF",X"CF",X"30",X"FC",X"BE",X"3E",X"6E",X"DC",X"70",X"E0",
		X"7E",X"77",X"B7",X"B7",X"77",X"EF",X"BE",X"BC",X"B0",X"E8",X"3C",X"9E",X"EE",X"EC",X"E8",X"FC",
		X"7C",X"CF",X"F7",X"FE",X"6E",X"0F",X"0F",X"06",X"1F",X"7D",X"FB",X"B7",X"F3",X"D9",X"6F",X"3F",
		X"0F",X"07",X"1C",X"7D",X"6B",X"3F",X"7F",X"3F",X"00",X"00",X"00",X"02",X"10",X"00",X"2E",X"0F",
		X"6F",X"37",X"1F",X"14",X"0F",X"2F",X"07",X"03",X"37",X"7E",X"DF",X"DB",X"DB",X"69",X"3C",X"6F",
		X"03",X"03",X"2B",X"1E",X"1E",X"25",X"3F",X"3B",X"F3",X"F3",X"F9",X"DF",X"6F",X"27",X"9F",X"0F",
		X"0F",X"1F",X"3F",X"67",X"ED",X"D9",X"DB",X"FB",X"03",X"6E",X"F3",X"E7",X"F1",X"FE",X"1F",X"03",
		X"B1",X"59",X"0C",X"24",X"02",X"00",X"00",X"00",X"77",X"CF",X"BB",X"80",X"EF",X"77",X"FA",X"3E",
		X"01",X"00",X"02",X"04",X"7D",X"59",X"B7",X"FE",X"CB",X"F7",X"FF",X"FF",X"6C",X"9F",X"F3",X"7C",
		X"6E",X"7F",X"07",X"FB",X"FD",X"BD",X"9F",X"DF",X"FF",X"FF",X"FE",X"63",X"CB",X"9D",X"FF",X"F3",
		X"3C",X"FE",X"CF",X"BD",X"BD",X"F3",X"7E",X"18",X"19",X"3C",X"7E",X"5E",X"66",X"7E",X"9C",X"00",
		X"06",X"00",X"78",X"7C",X"65",X"3C",X"00",X"02",X"00",X"01",X"18",X"3C",X"3C",X"18",X"02",X"40");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
