-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "47474746FDB82AA24071DDBD7FD3BECEFF7F7FC55CFD82FA54D5749A94C9495D";
    attribute INIT_01 of inst : label is "D51595DFFFA566BFCFC558C75845F5D3FB7935D53625FFFAFFF5FDBA7B7F474F";
    attribute INIT_02 of inst : label is "A0F155BDFA82BE1C71564FDCAEE0AAF0653F59134B7551B5677937DA55C041DC";
    attribute INIT_03 of inst : label is "37FD36DB3A2BA24FD7D777F2BBFB22263337FE8538ABB4F9F8585F7FF851D0F1";
    attribute INIT_04 of inst : label is "D15167BBC4D6DF5BACB2DB6B69F70EDB2D3EB4DB7F5AFA7A7D7D7D7D7A16D261";
    attribute INIT_05 of inst : label is "678DFE4F2F7D34D930F5E08B545460CACF077F7BB174EDE72EF1CB6D7BCEF3F2";
    attribute INIT_06 of inst : label is "77777777EFBEEAA8F7D54FDF3EBA38E373CF187362D14061DF9D5F556EC8E571";
    attribute INIT_07 of inst : label is "77575DFDBBEBEFFBDDDFFC5344CFF913C91F75247DD17B4193FD21CBA193CC13";
    attribute INIT_08 of inst : label is "DD9DD5B1679EA9ADB5D56B70F5F55576D5F56FA1BEBEBEBEDD7D55555051F4D7";
    attribute INIT_09 of inst : label is "59155D57B8273ED867B95D7515293DFC316590EF34D0D87BB7E3BC71EE3361D3";
    attribute INIT_0A of inst : label is "3FF9EFCFE33376C25DE747072EABABAB020CDDC7429F96F3CC0A0C5352D555D5";
    attribute INIT_0B of inst : label is "FF91B6419DAD24F97CC5EC4D9FFE5FA790FF34FD74FA30F2335A49F3B075F445";
    attribute INIT_0C of inst : label is "7F6E6F7DFEC434D4A5F575F5C36C67EF15D485D57870BBDA97E2649127C8F215";
    attribute INIT_0D of inst : label is "7DDE236EF914E925657575D6524B7F7B587D55FFE248BEB426B6A565F1F7DE53";
    attribute INIT_0E of inst : label is "F97679D6A4514A52B16C591F1FFCF3377DD98DC8964B72D0D7D635D576E809F1";
    attribute INIT_0F of inst : label is "4000445C201FFFFBCCCE9DE7F3CF3CBAA0A0A0DD74F2D972775DFFC751624067";
    attribute INIT_10 of inst : label is "657D65D7D7DFF7F5A95BFDF7A56ECCC799F57B78E213B4EE4E7BECB19992D679";
    attribute INIT_11 of inst : label is "2EAD757DBD69C7B48D7D78D711FBF5697DBBBA074DE65864DFD39BA2F59F0DBF";
    attribute INIT_12 of inst : label is "A65E655B9BFB3FFFFFFF7FFADB2FCFBD4D58C5575956FB7BFC9A78D7DA89F24B";
    attribute INIT_13 of inst : label is "587F5D97B2C4DF367094256DC9659442CFDEBDD53955F555F151F151F555F19E";
    attribute INIT_14 of inst : label is "4FED6D1D5A90B335D595665E8ECFAF2A4F4DEFED1D18FB387B60509E7B8D8CF0";
    attribute INIT_15 of inst : label is "D7F17DC456DF9B4758D2692FD163348359C6D517D648D6F865FB3E7C977D5F46";
    attribute INIT_16 of inst : label is "70CCDF33999626E87CCC311FCFBAB3131B44CDF61351FDF6D713135E5E5EB64D";
    attribute INIT_17 of inst : label is "73690BDCBEE6686F9F45A0382B02E92B07FF05FF06F204F3957CE14DD15B1B34";
    attribute INIT_18 of inst : label is "D78D6945A042536ADCD55AD1289096B95359555EDCD8BF49F5230718B8C9A42C";
    attribute INIT_19 of inst : label is "9B7C3FBC98A57DB08DCAD36E42C6C918D3BB7DD722497DD84EC2D15F76E03EB9";
    attribute INIT_1A of inst : label is "7565C5F7988888D2779679E5BCEBD9DD77D7DDE5DAB25151600D4CFD2DB6AE69";
    attribute INIT_1B of inst : label is "B77745DEA6BB122A77747FF4690FBDFB88FEC5F5D2F4D2F4C11D54033138EBEB";
    attribute INIT_1C of inst : label is "76F535F0D9F193B24B68A36DFFF4D27BEF9136DB5348D756C5F535F7E8D9D972";
    attribute INIT_1D of inst : label is "3455E1F519B27E33747BEDDDD32FDCD37DF77F5DFFFFD8FA6C94755F2262FA72";
    attribute INIT_1E of inst : label is "377F1027EC5B0AA0FEDDDDBFBB3369D427D092FA29DF4FE975DBB8C44892F5DA";
    attribute INIT_1F of inst : label is "83775C539B6EAAB9D5345FDDAFAE6DBAC1575CF1F93258D2F5FCFF5DDCD35F7E";
    attribute INIT_20 of inst : label is "90593EE212612B83A652247BB6C14E21EA93683D17FFFED05F64AD5F559E96E9";
    attribute INIT_21 of inst : label is "AEC795ADEEED9249C5D5699737C147ECB6D5DFF5B80C35D4CB3CDC95D2FBF0DA";
    attribute INIT_22 of inst : label is "1CDA5E7EAA7FEA1DF727EB5F86EA96E2FFFFDD66CADEDE79BB9F7F7DD5417F5F";
    attribute INIT_23 of inst : label is "B7F72F13FFAFBFAA0533F80D2EF0BBE25B6D5FDC9E7C41519B57045F5A6C5E59";
    attribute INIT_24 of inst : label is "77FDBDDCF1D403DEE6F6C7EF4D83CDFFF1B5B9F5CA57DBD6EF0997D07BEACBFE";
    attribute INIT_25 of inst : label is "75F77D6DDF4735D1DD75FF5D1CF1E73CF3CC4C4C49C9C9EA91CF1B671BD3CFF3";
    attribute INIT_26 of inst : label is "5ED50545D6F0BFBA56197C45EEC9AEBA5FD75CDF76DA5D77DF7D75775D73DC58";
    attribute INIT_27 of inst : label is "D7DDB56EFBEDAFBA7717FDB77BDFB7FA96A35F7334FF545A627B15D4F8D4D0D1";
    attribute INIT_28 of inst : label is "7DCD9F76933791CEDDB5DDB5733B7DBB6DDC7DDB5EDE529B76DFF6FBBF777272";
    attribute INIT_29 of inst : label is "C4C63C89265ABA6E16BBBA9079F35ECF1D5ED35E32C2BC7B891E7CCD7EC019C9";
    attribute INIT_2A of inst : label is "E35B2F1DFAD267F677D3CD32F8AF99FFEDD4C1A5B8D40159DF6FDF35719ED6CB";
    attribute INIT_2B of inst : label is "5493EDBBFFCAAABE94F596D7AD5EFCAE5293EDFB45DADC24F75DFD577E3972B5";
    attribute INIT_2C of inst : label is "F1D7888FE4E6E5EDF10EEE4639DF11C70EE9908F1596147E553C6D47D236635F";
    attribute INIT_2D of inst : label is "71E134F42E64982C6F3D45F5F54E07B17471EE52DC5DE1158ADB77C6236487DB";
    attribute INIT_2E of inst : label is "EF5ED5D3B8E67F9FC31344FCA74F39EEC7FEC777EBA318BCFCF2785B17161716";
    attribute INIT_2F of inst : label is "C000000055555555F131E5CC8E8CE3A3E7B731772FAA5C03475DBF77727A70E0";
    attribute INIT_30 of inst : label is "ECF4E775FDA7D5A7369BC549AB34ABC42334DCF3A75C3B9F5FC735D8D97852FB";
    attribute INIT_31 of inst : label is "677555E823B574ACC5C5F3D5E932AC7D475D71F1FAF8DA7D6EB9D5577A71FBF7";
    attribute INIT_32 of inst : label is "FE77905E92AAF1C0DCADA54BE6C22A0C5E57F79507CF9B255EBFDF55D0D5CA62";
    attribute INIT_33 of inst : label is "F5EDEDFE5136E60437FFFF559F81FBD25937F7FF5F5F5DDBCD5F5FD7B2FAFE7E";
    attribute INIT_34 of inst : label is "90A02130E0000E60808011321470610841242090CB20028A00A9F5D1B7B2FD7F";
    attribute INIT_35 of inst : label is "D7FFFFFF9C53A657FF5420808431D0FC3841261B38600A18326822869FA22280";
    attribute INIT_36 of inst : label is "F57D577702B762B57FF55D5FBFFEFAEB7FFFFFFF787DF851DDDF5FFFD2757BD1";
    attribute INIT_37 of inst : label is "41F77C17AABEEABF7FDC1DFF8EBAAE9777D7F3FDD753B2FBBFDFDFE0D3CB7B7D";
    attribute INIT_38 of inst : label is "D07C971534872942975FD15FDDAA3B6A7FEBDDDFF35BDD5D8F7DDF6BD587507A";
    attribute INIT_39 of inst : label is "F777FD764A5E703DCBFFD772504C6A29F7FD8DD55CDAD8D615757D75F35A734C";
    attribute INIT_3A of inst : label is "1DDD3FDFFFFFAAFAFFD5DFFFFEBFFFBFD55F57555E7DA0D441F5CFFFF2FAF9B8";
    attribute INIT_3B of inst : label is "F758365B6BBEEE107DFDFF63ABE6AEAE5F5B5F5F5A52565E535F00000FAFA751";
    attribute INIT_3C of inst : label is "F5F5F5F5F6BB76A6555751DD1366FED8F5DD57F5833EFEFBF5FFF7777E5EFFD3";
    attribute INIT_3D of inst : label is "5F51D55A3FCE6F22FFC7FD4BE21BA4E9FF3DD58D7C85DFFBD7DFDDF416F8F6F0";
    attribute INIT_3E of inst : label is "877968F3643BE07BFFD5B5DBBBEFFAEE27DFDF5D5876235A75F47554BFF1BF5E";
    attribute INIT_3F of inst : label is "AED971EAAF1FC1BB17DB7A572FDB00F2F94BA50D0EDCF35FF57F7F3554DFDF5F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "2D652D60469A1BBE3E3F7D0095F3A2024C4C4C295A1484A493283EFEFCE6697D";
    attribute INIT_01 of inst : label is "632D7C054702E335A16C92E44086B4608C39BBCDB9F268965165911C08B72767";
    attribute INIT_02 of inst : label is "CE5769DBA9CF9FBC52F786BDD53BFF73F76777AA083840DA8DC165B8A1B15228";
    attribute INIT_03 of inst : label is "2046492592DCED32C484F161E6223113828646993E7BEEDB9DFDBB06443AB8E6";
    attribute INIT_04 of inst : label is "6E049223292C901A167889C5432B249002182B24AAA088880000000088F1351D";
    attribute INIT_05 of inst : label is "D2547BCAEA8208083F6E6D846CBD0D94C251B254740961C3803986060CE6A0DD";
    attribute INIT_06 of inst : label is "04040400CC104003697564B1BB7FB36B649FAD67E9B39D6DD4C8F6C3FCDF50C4";
    attribute INIT_07 of inst : label is "55514544CDB2343D50444EC900F8A423A89A04924A3304DB29313DA1B430B1C4";
    attribute INIT_08 of inst : label is "396D7DC59249C2422A4FC740455F5958184522813C3C3C230F5F1F5E55511144";
    attribute INIT_09 of inst : label is "4D2F088248CA492C964A0E7B1A463219761F68329F471C547DEC0638E6243C74";
    attribute INIT_0A of inst : label is "028877A694665BCF322C672793FFFFFFF5F1B3E7E490E924B20000420D36D20E";
    attribute INIT_0B of inst : label is "37C07702526ACB6A744DF419564D7A97E19C92B055B896DCA6DF9CD4C72DE4A6";
    attribute INIT_0C of inst : label is "1D040642C48D3E6B6969790E1442412044458B4B36395875D2A567C0E6782170";
    attribute INIT_0D of inst : label is "42C579049312F2D37A7E68D1F048111356964486971823312CEB5A6A647091A6";
    attribute INIT_0E of inst : label is "4E085F772979E97A7C3F0F13649905AA483D7E5C2E51006024105171020899D1";
    attribute INIT_0F of inst : label is "BFFFD5E5D7C2626240488DE16CB25B5FFFFFFFB4D060B0E0D000741BC5649810";
    attribute INIT_10 of inst : label is "6917298584449EA910950B4214C6464186244268A266618E4826406185894B09";
    attribute INIT_11 of inst : label is "41167A428531486ED652518D10C2D8C3522224802261192985C1008AB0F31862";
    attribute INIT_12 of inst : label is "E61C09D0C02A8335F5557FE6B84D96A07CBA89F483D628E26527BD656019D289";
    attribute INIT_13 of inst : label is "0FC61C632CBBF66D1784E02BBFB248B2444F0C5540C6961632B2921236B69E03";
    attribute INIT_14 of inst : label is "237B6392D99BAB2CDBAF1435CC8F131064697B7799855897E26011850FADCC0F";
    attribute INIT_15 of inst : label is "847911C65CC3184B53C45699124C28800BAD61266D318D1C57FC131788DCDA66";
    attribute INIT_16 of inst : label is "4584D9905C79718D62416018BF4BEA4D87D8EAD6E223FB5D768989919191C5E8";
    attribute INIT_17 of inst : label is "0358664035B9389DC201E398A06CD249E125E125E420E42299916D191B62E05F";
    attribute INIT_18 of inst : label is "4FFBDC332D8D8C4A7B874F84036B6E18618A7BC0DB88CAECC4F8586E64096199";
    attribute INIT_19 of inst : label is "601F830221CB0238C9A48019979312B28020168D963B978280678CE4E14A231C";
    attribute INIT_1A of inst : label is "1E3918664C4C4C0471871C616B2CB0004164283035C1AB7B1EF1E485D366F384";
    attribute INIT_1B of inst : label is "36E2112873236C816E2716224A4C4B24BCBB55612064306434DC74F89043F1B1";
    attribute INIT_1C of inst : label is "2B23B9378DBBD19824726802646C9811CC4EB92E421585B93823B9328DB8844A";
    attribute INIT_1D of inst : label is "6D2E5E00B791B5792B1687B2C7169EB943282412488C376497944B925717236E";
    attribute INIT_1E of inst : label is "9DD964F51EEFD77FC8DB8942E646DD0391172A3F99268909C1631031A8D9907D";
    attribute INIT_1F of inst : label is "7E67D997E3498BEFD944199FCE739D6227BEE51059BB3CBB7B0732C82C629302";
    attribute INIT_20 of inst : label is "9A160FCD406B419B79553E506E2B442B1BCF72746A0AA1AAAA55AFFAFEE8A1DA";
    attribute INIT_21 of inst : label is "7386C4571CC3D962130B00692878C0497B7B6A6936497139ED00B2C525411D96";
    attribute INIT_22 of inst : label is "61C7271961E290E66831177E7E89E44999190039345C1D9BC017465669A39BB0";
    attribute INIT_23 of inst : label is "8801E405FB67881105440481677772DD98684BABF9010740F817C0076802450E";
    attribute INIT_24 of inst : label is "6FBC404F8BEB296100C001D433006458C0220A6D2640C87DF254BE650898090B";
    attribute INIT_25 of inst : label is "294C02538841289A122B4C42045945141E0606060404048D8CADA1859A94A630";
    attribute INIT_26 of inst : label is "C1721CF6BC92FEA7823D80988A14CB2589728978C462B9C06798C1C6B80818B8";
    attribute INIT_27 of inst : label is "7B9CB1DD0498D80D5D7B98A182424026E5C2B24B8412B1B2FE8C339DD4A2A471";
    attribute INIT_28 of inst : label is "41A64C689129923E963B96BB07301330224311C019CA10C668C45D002262065D";
    attribute INIT_29 of inst : label is "25245211AB04B97186A12085B65818556392C7AA25A3DB1C11EB67C249D88A88";
    attribute INIT_2A of inst : label is "69059611526333F2614D089363F7D0A1F5F5ED19F8FAF6DB0BFC0F4247293929";
    attribute INIT_2B of inst : label is "AC622887FF8DF97CF25C7EC9A81CB8999665EA71B155139FF20020001290E690";
    attribute INIT_2C of inst : label is "EE16B2058F71A240EA6068297C4C6052F0203E0BF52D6591FDDC4C405B344071";
    attribute INIT_2D of inst : label is "75FA196E788DC2241C85D000000B6D193E649618621369CB225531AA880CE4CE";
    attribute INIT_2E of inst : label is "E7423439E5A4EACBA688AA6AB979A5C0A81E97F566B70009E6BA62BD94849496";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFF961B8E5EA93D8A4F663379BD78F0C992666913F7F7A7A7560";
    attribute INIT_30 of inst : label is "597883344F8123818D652CA16AC6D36D4BE4DB0D50E5EEC89FC8DE0D9085EEC0";
    attribute INIT_31 of inst : label is "551F45DC405A09032A254797386C4CCB420AB06062632E1D7784E6294F123E62";
    attribute INIT_32 of inst : label is "40809DAEC82A2BCB8C99A076D1E99268CAE6F39E87F4D6CB5D6D342F9DF926A3";
    attribute INIT_33 of inst : label is "8006B8ABE14209D19FD2794060741441001F12580000807B664C58701A0A2121";
    attribute INIT_34 of inst : label is "B0B96BB7FFDF6EE7BC9033B4B4F17D6FE1A77C28EABEFA9AFFBED00A9AE7FFB4";
    attribute INIT_35 of inst : label is "520000000800020000206FBCD77567F6BEFBA73BBDF7FF7BB4F168CEBBB362CE";
    attribute INIT_36 of inst : label is "01A880AA828AB26AF957FD4002748A69A4000000E02000408010008410304000";
    attribute INIT_37 of inst : label is "E4010C5A074C5F13ABE40BEA6F8924D6156E157A00F0AF08EA35CA61BF984242";
    attribute INIT_38 of inst : label is "5A5E570D26030842175EE955F70A7D4275EF125C217895389DB14C2BA892E8BE";
    attribute INIT_39 of inst : label is "D72B56EA05CA083FCEB359B37E0FF709A0A71CB4B85AE3E440E2E968B17BA145";
    attribute INIT_3A of inst : label is "1500D60C910AAF8515400115C00004043510F0B420E030AF65DEB5FE247F1AFF";
    attribute INIT_3B of inst : label is "4BFC239E93E50E9FBA0000D404650D0900464443404040406561A0A0A0A0009E";
    attribute INIT_3C of inst : label is "0000000006CD675F59B7F76F42BFFFF5B5EAA9E5146D1505414AD2A2B4AD052B";
    attribute INIT_3D of inst : label is "5FF95FC235C26592A3D5B62AF52BBC49A315E688ED936BA0876CA0065A2FE6FD";
    attribute INIT_3E of inst : label is "0B34E002B3E57D92CC05DA953C00402434024A2E008E330977FD57F2BF02FF14";
    attribute INIT_3F of inst : label is "C12A6AE597EE6BA3A6BDECBAC4E50C256A204A2847CD4282300A25740A380000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "CA8A82CC64EA7B96E279BB35FF4283F7E5A5A5B7280CFB0AF4F97FDBD6AFB3EC";
    attribute INIT_01 of inst : label is "A77FAAF770A4A7A72A60D8EAE9D5D5A8FCF3B1E73FA157154B8C1B2A321D8DCD";
    attribute INIT_02 of inst : label is "BE88B88F89A6FF8CEB32D38E69AD14B5E37C026FBD5A4FB7A6B6389F5FAEAD19";
    attribute INIT_03 of inst : label is "B73B2CBA3F65F6E68E8C60BE6999B332B198396D0F5FDE9D7EDEDD7DDF6ABFBC";
    attribute INIT_04 of inst : label is "725BE6A8EBEEBFD9FBFEAAFEEBFFB6FAEA21AEB18F23E36B666E66EE6331F6AC";
    attribute INIT_05 of inst : label is "87B980DA7F332C9260A6609BD7E7F1B688E1986CF3ECB8A728E8C93DBC44CA0B";
    attribute INIT_06 of inst : label is "EAAEEAAEBBEFBAFDEEF3C1BE371E39737BC9889EFD660D7F1BF5BBDCDEE964D6";
    attribute INIT_07 of inst : label is "EEBBBAEE9CE67308BBFEECBA00559C01AB85F2BE35EC3F8CD2CC6AE2EF2FCF0B";
    attribute INIT_08 of inst : label is "E5B4E439D7EDE363FF3C78B1B0F0FE6861F83DD0FFFFFFF37CE6F3B9EBEABEBB";
    attribute INIT_09 of inst : label is "5D7368D36D6B6FF4C7BF5718BD6753EFF22CB7CB8BDE6096A48A3EEAC626CCE6";
    attribute INIT_0A of inst : label is "3336E54D766428B4BAABA3E352ABABAB5E5FB06326EF1F36EF0517BB5BFE3B47";
    attribute INIT_0B of inst : label is "8973854BD9CD865B88BE70E493C92D1043628C9652478A35B99B084733D75EEB";
    attribute INIT_0C of inst : label is "33EC28F97CCC6CFFB1A1A3E6DB6D77CF646C9CBE63108FCBABC20882A1EDDEB2";
    attribute INIT_0D of inst : label is "FB7BB6E8ED8E4DE7F6F6F5AEDB63FC69E938EDBF3E1EAEB63A23A6F6F1EAAB8A";
    attribute INIT_0E of inst : label is "3A4BBC8E64C301C027CBFA6E1D8EB9B133EFC849DE09CA8A871BA3D36CFDCDF5";
    attribute INIT_0F of inst : label is "C000399B6FC9DD91004ECE6138E39CCCA0A0A0AAADA6ABDF32EBE971E3FC697D";
    attribute INIT_10 of inst : label is "E19CF984F790F7B114B02B5285E466678DAEFEF8E6A56DEF2B36CC38E9E9CAFD";
    attribute INIT_11 of inst : label is "22E8F6FB3FED7AF6C8E8C48F5DF95D6DE9A1A93EA3E69FF684F390B3FFAA2189";
    attribute INIT_12 of inst : label is "AEB13CC85A732668F5F5DFFA879CC2064DF71CCEFE0CE1AB7CDF3C8E874DF74E";
    attribute INIT_13 of inst : label is "1ABFE6B131E6B7AD328CA4E3EE71D04D21BE4EF1D1B767E7C3C3C34367676E6E";
    attribute INIT_14 of inst : label is "431B1828327072F50EF31B9B89C98F8F0203191D282BABEB72F6B4A6FB8EBECF";
    attribute INIT_15 of inst : label is "84E633DDEADEF9EFEC93283BF3E3F5D77A030745CA5BC8E8E20311BC8743424E";
    attribute INIT_16 of inst : label is "BAD4A1737DD6F04F814EB42065CB99A2B30D60391921BC62A830204E6A4AB29C";
    attribute INIT_17 of inst : label is "D36858F46DCB4A5B8CBBA5BAD3065919496E496E4D6A4D6A2E6E466E87521A91";
    attribute INIT_18 of inst : label is "51F4FD74C8CCC6CB65A477557233B694141F338DBEFAC9EBEDA74B6D8A48A466";
    attribute INIT_19 of inst : label is "1B9BBA8C7DDDCDE5DC48F3803B3B8561D3A314ADEE5DB5C8E87AD42430F2BFAF";
    attribute INIT_1A of inst : label is "E76B6D994DD55D9819871CF366658991618793EDBEB3075DCBFEEE67477BE9F3";
    attribute INIT_1B of inst : label is "EEFFB96B266690C9E7FF9E7CD9B66B260D9A791B931F931F83CAC7FB0F057969";
    attribute INIT_1C of inst : label is "E333A1BCCFD5FDC64C69B7CDF2B6BFFCABB331A6D21FC18E2B13A19CBA9EAB5E";
    attribute INIT_1D of inst : label is "A32AD244FD77A2F6E1B8F99DAF2DBED179E6461CFE37F9E8ECD082B8EE3FAAEB";
    attribute INIT_1E of inst : label is "3F3939B4D350C579EBF9BA4C37B8CC4E3B36923A4D974ECDFB9A38CCCEC990EE";
    attribute INIT_1F of inst : label is "42C73ABB87D88B399B279B1C8D320F229B326C1E4C406481B81A3EDB96871F6C";
    attribute INIT_20 of inst : label is "8B99462277764993A593771DEEF9E48D669E6DB316DEFBEBA1A81AA3AF9EFF21";
    attribute INIT_21 of inst : label is "4EDB876C7C6F9241A1A0A4F6ADD846F535A9FA63A30832E4A31CA286C3FEFE9C";
    attribute INIT_22 of inst : label is "34D74F363A5266DDEEA35B5504970A6AC682AF66D6C6C69F39C8283C5C6A9A3F";
    attribute INIT_23 of inst : label is "AFB313EEABA5C3BEFEAEFAABE5412A741F4F6FFEAF5F507B6CE8133A1B451DDB";
    attribute INIT_24 of inst : label is "3EEBA1387E7B49E7E590AF3906D2A1F1F17EE1DC4CB412BF678D958C9A6AF3BB";
    attribute INIT_25 of inst : label is "E1EEF861BFD565B69CE326BCF5FCF1E5AF86CA8609CD89EE9D4A324226344DCA";
    attribute INIT_26 of inst : label is "8E6E6DA366B0549DD5B9EFCD08471E3859C7780EEFCE1BEF871EEBCE1FC739BF";
    attribute INIT_27 of inst : label is "EBBFA38030CF09B1F3EBBFA3A787B07221F63AF36533169E3F7A76DECFE7F36E";
    attribute INIT_28 of inst : label is "EB8DECE6D5B7D75EBDA3BDA3D7BBFDFBE8E7B3BA3EBF3C6BE68666D3BFEB4AF6";
    attribute INIT_29 of inst : label is "65636E00674D536E2D53B2B07DF25E83999CBF84A36BA81F0004ECB8ECFBEFFD";
    attribute INIT_2A of inst : label is "EAEAEBEDF9CA656ADAFFDFD2B8CAC52AAABA4A4DDA594ADF5BA52F793B5BD3ED";
    attribute INIT_2B of inst : label is "4DB577B7002B58D622AE8F24C1BE04767B3161D26E9DE78F5557DD7F4FC8BC4B";
    attribute INIT_2C of inst : label is "59EEB2817DFFC47279949CCBA13995A146E39AF6AEFFABFB9D526A61FDF742BB";
    attribute INIT_2D of inst : label is "803CA49A81EA07D1E3BCA0A0F5EFBECE9A860CF9686F99C7A19A4FF2AF78A796";
    attribute INIT_2E of inst : label is "48A86BF2554211C5082BAA881D559DA6E6E0C8AAA9A9183FBCD34DEB93938393";
    attribute INIT_2F of inst : label is "80000000555555549B320A2C575755D5688881A89F5DBB9839BEE080258FAEEF";
    attribute INIT_30 of inst : label is "C7BD627BBEB45EBCD89C3C900051563B04D5D50229AD5AB1EA1BD6F472FBECDA";
    attribute INIT_31 of inst : label is "DBFEB6A143C8792D66F3B24CFD1468D6E3776FBDBAB9F87F8251F421D3CC7CAE";
    attribute INIT_32 of inst : label is "D54F5CFD91C4A8895CB59371A7A23AAC95452F54D213891A6A3EFD3EDC507FAC";
    attribute INIT_33 of inst : label is "60ACB8AA57C39C84355887E0352156C86E35B8F75F5E1CD4CD99175AB5A5FE7E";
    attribute INIT_34 of inst : label is "D5E4C319F471F719C63A9B1A4B0EC2F5CB0CE68244105135552AC384B7E05537";
    attribute INIT_35 of inst : label is "A9F5F5F5F7FDFDFDE5F4F1C674F2D80F10630C971EEADBFC1A6AC3ADD26DCCBA";
    attribute INIT_36 of inst : label is "56F7DF7D02BDDA778A08889FEA21AF1C8F5F5F5EEF9F4FEF3F7FDF5F7F9FDF6F";
    attribute INIT_37 of inst : label is "FF5BF5A3A9F893BC1FF5B2F9A558E8FEFE038EA47C50AEC7B98E9AD68BD0828A";
    attribute INIT_38 of inst : label is "29C2B0B4FC7595E5F055949FFDF073F474FEB48B2B00EFFEF9C4B4FEBAEEF81A";
    attribute INIT_39 of inst : label is "A2C2ABCDFEF785DC7BB0AF9ECDFFEFFDF46FEF95FAAFF1B2BE77F4B5BFA8ADAA";
    attribute INIT_3A of inst : label is "7071C31EAAAAFEA8FFEBFEFBEF2C8AEABEBF5A1E9F5F68597B7ECA561F991FA7";
    attribute INIT_3B of inst : label is "1C52FDF7ACA54B8A29FBFF0BEBE5E0E65F555A1E1C1C1E1E1F1FA0A0AFA5F873";
    attribute INIT_3C of inst : label is "F5F5F5F5C3FDF5D5AFFEA422FD49BBA5447DFC11BA5D0407011F07FDC4F50179";
    attribute INIT_3D of inst : label is "95F4B5FFB5DFFDF7F062E7FBD17FDDF5EDE07FFD38FEABF0A0AB415DA67BA2CB";
    attribute INIT_3E of inst : label is "F99A5E5216FA71D9467F3EBF82EAC3207D173CD55FFDEF5F22AE2AAFBFA7EFAF";
    attribute INIT_3F of inst : label is "67FDC547BB21404A9ECFCFBD3B8A08B35D661797DB2615D5E5FDCB22550D5F5F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "6363636CC02FACC34E9F93913F266208555F55CF1E596BE515117C9811364ACE";
    attribute INIT_01 of inst : label is "7F37F1559E529C47CED579678B29042DD8D3136F145B1C35C904291FB6906060";
    attribute INIT_02 of inst : label is "2191326CDF044F5C51892B4CDF352DF563055099EF785295CF1D39B7A451B339";
    attribute INIT_03 of inst : label is "99971C713F7EE7426464595833332226193464730412013230F0E6E67A4D90B7";
    attribute INIT_04 of inst : label is "47F1C7510B1842249E5959670A0A40021F945E71FA50D050DFD75F57D81F5CF7";
    attribute INIT_05 of inst : label is "C73F7C65B585F0779096D76722184C01650114FD99D7DC611C5945FF316052D3";
    attribute INIT_06 of inst : label is "55555555BBEFFFE95659E95C339EBCF371C1931CD46DF6681533B956F0E66BD4";
    attribute INIT_07 of inst : label is "55555555AAAAAAAA5555563858E49D63670FF1BE3BC2B612D9DC5461D12520D0";
    attribute INIT_08 of inst : label is "636E6FBB6DA63325D596E11EFBBBB8D1D7F6576BC6C6C6D5FFDFFFFFFFFBFFFF";
    attribute INIT_09 of inst : label is "D3D06D5B252936DB6DB1CDB6C61825FC5D7142ED967A69BBCF4514104D9BE0DB";
    attribute INIT_0A of inst : label is "3932CD69333270D05DC1C909EEABABAB575DD4C9D92F96DB6C0004BDFF7095E9";
    attribute INIT_0B of inst : label is "D53B54E3DAB22AE9D4CF4EF5D2CF3EA6B9F53E9678F533D7BD645453507A5A63";
    attribute INIT_0C of inst : label is "9DE6E6F33102023293D9DBE599133CDC2EEF4AF4C79DFFCBD96565595650D992";
    attribute INIT_0D of inst : label is "F37691E662040464DC5CDF75C899E6E2F7364F3569479998561694DC5CDF7588";
    attribute INIT_0E of inst : label is "9D569D077A49284A82E2B924FD9BE64C936314F432F2CE6667B69173CDC7245C";
    attribute INIT_0F of inst : label is "800067CE803AEEEA6666245B6DB2DB8800000077DB7DF6D97DF7FF7B5A7EE44F";
    attribute INIT_10 of inst : label is "D1BDD96D32E3648A01B41354C0BBBBBE7DCED8D9601D5C60E658DE502D3F5CD3";
    attribute INIT_11 of inst : label is "AF8ED679D8CD1E137CDC706FA41D2C9CDD119C37E1DEB7DD6D73B361DD489349";
    attribute INIT_12 of inst : label is "CC9AF625BB2982205FF55551D70DF7BC67D8F6B79D91440C76B137CDC702FC43";
    attribute INIT_13 of inst : label is "95314FC979CE87B1B56D5E59D8E3D9F06913467F0734F4F4F1F1F1715454590C";
    attribute INIT_14 of inst : label is "E1191F9F852508495E5ACB9B21205A5AE7E1191F92845325D0C6B927D2426255";
    attribute INIT_15 of inst : label is "6C57917E36080FB4CD77FF936DB61967D06347FBFB617B667DDB94B17D4341E5";
    attribute INIT_16 of inst : label is "D06E57B9D88767FD5EE419877F8F1F4719B64774B44C12B9D5191954D575B8E3";
    attribute INIT_17 of inst : label is "71F7545C29A67ACA654B587803BECF8E0BCD0BCD0BCC0BCD9F74CBC5FAFB193A";
    attribute INIT_18 of inst : label is "4124434946424CB4266FD0D25190918F571501522230A640445381FDC965D772";
    attribute INIT_19 of inst : label is "99167BB65B16F0510F4671DD2B3325645999916CAC65945FC62A596551AF19B6";
    attribute INIT_1A of inst : label is "F6E1E55DDCCCCCC4936DB65B7938BCCCD14F336D5E931644442C5C07A61F0C4A";
    attribute INIT_1B of inst : label is "884C6B7220222A5C84C498564A92BD6B54B5EB7B767B767B79B67C07BB94F8DC";
    attribute INIT_1C of inst : label is "C49B01110664040446F491C7998860E2613194D2D56B5D5A139B011726361ADD";
    attribute INIT_1D of inst : label is "9656C46E40C9DD89C69322330A2158C8F3CCC5347132D081C156CDB32D69CD89";
    attribute INIT_1E of inst : label is "B5233055A94A0B627221312E42EA4BB3133551BD2471E6625B79994C60B0915E";
    attribute INIT_1F of inst : label is "00473699D6588E6D71ACB13C98E359626911C6B2D4D0F5314C1D3CF311453CCC";
    attribute INIT_20 of inst : label is "62BD8DE79F929C269E97969D8BDAB95AF0785E55355C44505F28A55B557E3593";
    attribute INIT_21 of inst : label is "A46167AF05D864947461E1A658253EB49ED1D0DB49D21AD74F1E5467CEA7BD34";
    attribute INIT_22 of inst : label is "FC78C4963B52EE4D571BE9FDA9E3A3231B99C564F79D9F10F9EE66785B4D183B";
    attribute INIT_23 of inst : label is "314DA9EEAAFAFFAEBBFEBAB96EEF32C412445184B2C64E6629E54C794447DA54";
    attribute INIT_24 of inst : label is "5A5F115CAB0238C661B0EFCDBB01C0B19067B175455290D9B7CDBF5B73C26941";
    attribute INIT_25 of inst : label is "5367DC412F904167BDD3E7FC73259451306C6464EFEBEB60396B91C3805960D2";
    attribute INIT_26 of inst : label is "34F0C34B80E1BC9A2CCD6677CBE58E3853DD56D67BCC3279CD16F9C5126436B6";
    attribute INIT_27 of inst : label is "C13799997D558DBDF981379977D7B67E3C2938F1B9B1B5FDE0FB2F12462B2B51";
    attribute INIT_28 of inst : label is "C145AC5E08580888179117112A05A005C45E9179117012205C40D1B998582172";
    attribute INIT_29 of inst : label is "E6E8242B41574530AC188ABA67806CA997127BC68343B0122B664666C04E6042";
    attribute INIT_2A of inst : label is "EAF97181DF8622B69E5BD778BACFCA6ABECB61A538C42147B105259772171F48";
    attribute INIT_2B of inst : label is "D49366BB555FCFEA86CF84BC9D5FD5B77091675362FEEE661FFFFF7ECD62FAAF";
    attribute INIT_2C of inst : label is "76E7188B510446BA79048CE4AD3807AF0CE3B3B7F0273F57751A43657C5F47F5";
    attribute INIT_2D of inst : label is "9E41BE1C52895FCAC1059FFFAA542DD696994EF0DD61867999B0C5DE62624431";
    attribute INIT_2E of inst : label is "6948F5330C3600C36D33CC8493134C2AC556C1D06889BF9EEE70DD67BBBABAB9";
    attribute INIT_2F of inst : label is "0000000000000001991A6A46D2D134B469A919890005B34461B405557AF2D460";
    attribute INIT_30 of inst : label is "6C94E595F2417848303988243F95A1C6B466FE66976EE0934F613EF093F1C250";
    attribute INIT_31 of inst : label is "4B7D4621B57CA6D597FB532D74C19920659001515052E48D6A904490FD6EF690";
    attribute INIT_32 of inst : label is "7EED3264D3CAB1C166378D40E6C1620D141F399F8A6F5C526206C777933B4D48";
    attribute INIT_33 of inst : label is "75F8AAAA560A69D36075F7F460740A76CFC5185550506C14795D755F45057171";
    attribute INIT_34 of inst : label is "BAA22310F4516C41A28A13101E78626DCB2E221A4D01038E000BFFD567AD07F8";
    attribute INIT_35 of inst : label is "5555555500000000557420A29C7E40F618632E191DE68B3C1062208EBEA3238B";
    attribute INIT_36 of inst : label is "F557D5FD5AB55D7DFDD7D7D5EAAAAEBA55555555705050D05575755550505050";
    attribute INIT_37 of inst : label is "5FEFE7E1805012BA010FE000AB0000FD01400560A0F0E000E005C01F8037555D";
    attribute INIT_38 of inst : label is "F5FD7F6FBFAFEBFAFF542BDA36A00FE868F556D0FA47EA83543BE2F527D525AE";
    attribute INIT_39 of inst : label is "6FA3BE2D5B747A2BD48BD0B5734479A3AAAB52AE0EDDAE2D4AB83F4AAE4D2ED3";
    attribute INIT_3A of inst : label is "BCBDB6DFFFFFFBFFFFDFFEFFFFBDFFFFFFFFFFFFFFFFD02BD5602F582ADF8D52";
    attribute INIT_3B of inst : label is "AFF94B2C9FFAEF3F0BB7F64ABFBBBFBBFEFAF7F5F5F7F5F7FAD6FFFFF0FFF7F5";
    attribute INIT_3C of inst : label is "FFFFFFFFCF98487FABEFFCAAFBE44FF3AA8828AA8F2FAEABAAAFAB55EFFEABBF";
    attribute INIT_3D of inst : label is "CABBEABD3FDD7CEAA0EFB0D4B755C3ABABBF03D2A5D5AB89BFB8236543EDA7A7";
    attribute INIT_3E of inst : label is "8D5B6875652AE2BF5780A88FFEEC4455D5F6A025F80F5406F2AEFAAD5FA55FBA";
    attribute INIT_3F of inst : label is "FEA7AFA27C7C0D79B2730F81DB7D5757A58A9696BB8FF3777FF5FF977B787FFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "D292929141214008992675423FE028A02AF5A07A6B4000D1AB2660C8CFF6F7ED";
    attribute INIT_01 of inst : label is "3204769A16200037D1190DBCF115DC90831DC714CB2525EE1CF1D5C84C76D6D6";
    attribute INIT_02 of inst : label is "F5B04411A4D3C037B0505652309061180D45ADDC4B8A028CC9761C5201CA2CCB";
    attribute INIT_03 of inst : label is "6262492C8114519999932536A1119998E4C223008706545D41272AA226B27F68";
    attribute INIT_04 of inst : label is "8C06B027E7B5D471E5A4CDF171E7B5D464F1B3248220008888808880888001C0";
    attribute INIT_05 of inst : label is "90700A1FBFCA0CC967B96C9466DE44929457D14020292BDB6576B4064DBE314E";
    attribute INIT_06 of inst : label is "51111555CB3C8F286306FE8A2C69A698061C79CF1654848D6CD0D3115D74C406";
    attribute INIT_07 of inst : label is "0A00288A00000000A8A8AF05EA4F13A93C5F26D179BD12C925790A3C8E705114";
    attribute INIT_08 of inst : label is "9164EC4C94638080E190C0B510A0A20A604830ECE8E8E8E28080202082808280";
    attribute INIT_09 of inst : label is "0A490902E1004125B0E004123321308FE4125A1008F9E6902D80006187A05020";
    attribute INIT_0A of inst : label is "699A77A65280909C4CE98181E1575757020820C150244F0D1BB5F0924404980C";
    attribute INIT_0B of inst : label is "6EA3E20E4B720B30E0EB88F9E3890312A218BD1E461D9A679EEE1C5162777C3C";
    attribute INIT_0C of inst : label is "3441A441DCD08C0CF9F963A5A0434176A66DC75A66185305598505C971186244";
    attribute INIT_0D of inst : label is "41FAF841B7A30387FA7A6195104011F15436649F8E082EB1CA6A727AF0609246";
    attribute INIT_0E of inst : label is "1412B4056B4D374D795E5446E89A270929A9005C24514A6846364361076C9D51";
    attribute INIT_0F of inst : label is "BFFF8310B4233333000286716DB2CB4AFFFFFFAA8D0622860A208809C26C7541";
    attribute INIT_10 of inst : label is "BCE58DD184F4AC63FDFFD5F588C4E463D7738DE5BAC6BBD23D2D416EBDDA7B0C";
    attribute INIT_11 of inst : label is "7193BB04FFC4CDFC9731139110DDD4433066E4605A33E881D184E4EC26B04932";
    attribute INIT_12 of inst : label is "A24E0412808838B50000AAA28862188004E60531D4849AD0222BC97B113D161B";
    attribute INIT_13 of inst : label is "4FC21214863B4AC24CDA3586A259621E3EE27B5418E3B333B232B2B232B2347C";
    attribute INIT_14 of inst : label is "75A522F2D3F3BFE986182AFA8DDD1DBC343525A2D9F753DE6DC4D03406BC9C14";
    attribute INIT_15 of inst : label is "53484D022C53B0C1C8D106E5B0E76DC41CB251410B598BA04A8032DC9EEA4A7A";
    attribute INIT_16 of inst : label is "56D5C8776EA3BA56215DB54D4AAD926CCB85B5236A725D26B3F4E46560E01231";
    attribute INIT_17 of inst : label is "260C9BC9B28D9E6CD21D257F1C6660657F167F1E7E137E1BC7D57F58A550705F";
    attribute INIT_18 of inst : label is "602CA20A6A081C42C28D88021A0A8E9688141B1098998058667A9BABAD89726B";
    attribute INIT_19 of inst : label is "413E620038EB916D8184D8776075EC5FD0E11C879A003CD060E580073480BEA8";
    attribute INIT_1A of inst : label is "C95BF0EE555554041BCF3CF32865E820D14439BF28438565CA0E5ACE11809262";
    attribute INIT_1B of inst : label is "A6660B7A6867AD4D6770B2B60AD284289C1E298166846684740CD8860AE0EA63";
    attribute INIT_1C of inst : label is "7019719D9751911440D6F94164EC9811A87F2220FE0681011B1B639DAC9C825F";
    attribute INIT_1D of inst : label is "E808764E113AA03872BDE5959987C451C1266514489E2523B9CA723C1A0FFE62";
    attribute INIT_1E of inst : label is "88496D7094A54433BED9DC84A6200E80411132379D564B0941125B1DE80A1A20";
    attribute INIT_1F of inst : label is "BEC51CB7E618DB28C16EBB144CC3986304BB853ADEA4C495E1123249BE6233E7";
    attribute INIT_20 of inst : label is "CAF25C40157E21C879D06B54DE52C40701CD4364C32BC82EA00CB5F47F88E7C9";
    attribute INIT_21 of inst : label is "179C92071C8DD941455161ABA0614876A89FE33EB4482291D955819316E2B9ED";
    attribute INIT_22 of inst : label is "5C825E5EFA6C9D6EE6640B0AA298605288CCB94826CEC8D9956A2A257D34D243";
    attribute INIT_23 of inst : label is "D820945CFA81C0BAEA5253BC0CCDB08E421818036347222AF88CE0A1A0132C0C";
    attribute INIT_24 of inst : label is "4C06C05D4E63216114C0309D8B03C4D285A0C6AA9646C86EAC28A12422323221";
    attribute INIT_25 of inst : label is "B4B101148C4525D8E1A479610432C9042957D393D151113BDBB3E4BBC895F621";
    attribute INIT_26 of inst : label is "591D4474009CAB92034A3310A216208B0E136D1F141269851A691492489068C9";
    attribute INIT_27 of inst : label is "4FC9F586EBAAE20E058FE9F5EEE82FA84247EF5F544EDA36AEA4C1110B45471E";
    attribute INIT_28 of inst : label is "73B1A4F4D9A5D88495B995B929307730665CB191199A1226F4C84938FEF2AF01";
    attribute INIT_29 of inst : label is "0C16B890FC05F95465F8E1B1307114D47633D24CAE81483F90AD6DC6799FBACC";
    attribute INIT_2A of inst : label is "EE283638A0AC00089AEE3A330F0DCF6AC6DEEA11A100B08E0BF72F05270AC2AB";
    attribute INIT_2B of inst : label is "10C1A3DF800E0B80569847F9E41C6E860A4540515208E509C0820800050A3846";
    attribute INIT_2C of inst : label is "D36D84A313E676D9C9CA6AADB2EC8CB43B289BA86A58F2B08A556468E9A840B5";
    attribute INIT_2D of inst : label is "75E437E07951E5DC5638300000A0B5CF787182E9620C6419D294674E37E552B8";
    attribute INIT_2E of inst : label is "1EB76A41B0D2B30DAA0922E8256F30AC25985E0BA2B3CFE91AC3C68CC5C58585";
    attribute INIT_2F of inst : label is "3FFFFFFFFFFFFFFA622BAF8A4F0CD3C32E9E097E0F091A2F0E1B9FF7F7F7DEBF";
    attribute INIT_30 of inst : label is "0A2717020A012201A5A8060A1E2DE55585A0F893AC52A5C595040B012B0D9B08";
    attribute INIT_31 of inst : label is "8149E4A200224600DE0EF119864800AAB60290404441042AC8A2644E01311422";
    attribute INIT_32 of inst : label is "09BC090445080F120180C020DA05037242DC3BE3A729ECF0480440211005265B";
    attribute INIT_33 of inst : label is "00ADFDFFE28484873785000035215788C817B2F8000F187BCDA5020212AAA323";
    attribute INIT_34 of inst : label is "4D445345F65B6400575F06440A0802041E58478F144505550A5F420832F2FF50";
    attribute INIT_35 of inst : label is "30A0A0A04125D1A530015D5702029002402258044410214444535389EBE15010";
    attribute INIT_36 of inst : label is "DDF5D555D81557D5BCA008A800080000420A0A0A030E070E0A0A52020D0A0D06";
    attribute INIT_37 of inst : label is "AA6540F4460949032028AD3C0AD14D0B0164414080F004505C25420B3C41F95D";
    attribute INIT_38 of inst : label is "70541D07D074150D85FE81F2B07FA257E021F47A44E912282611C02188AA200E";
    attribute INIT_39 of inst : label is "E509D4A0E7D181C680007080B5351894000022042676AAA0A81091E828E3A8C1";
    attribute INIT_3A of inst : label is "A494984000000000A000ABA040420000000A00000E0F0F850BCA07F2A57B021F";
    attribute INIT_3B of inst : label is "088CB473255FFF64FA00219408050004010401010C000C000D01F5F5AAF0A893";
    attribute INIT_3C of inst : label is "000000001820A8D155E5F9054F70A0820B20B40A75D040010A054821D1F0003C";
    attribute INIT_3D of inst : label is "E0B1C000F5E182A50845182024A43694031580A086AA872735B0A16AA5462B2B";
    attribute INIT_3E of inst : label is "8BB8E98670E26B92ECFFC8822FBD40020DFC0A00070D08025A0C50021F0A1019";
    attribute INIT_3F of inst : label is "C2AC0480742000300A08A828152920800C050800128706A2288202E090EF8000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "6060606656819FDF69D27D14C80201F415F5550C50FED9555614408089D6490F";
    attribute INIT_01 of inst : label is "76546F0242101748E9FEF8C5D2A4BD02E5313FDDBDB821D6577DCF91CC9E6E6E";
    attribute INIT_02 of inst : label is "CB346A5ABCEB2EB855BAA65F3A6A51AAD5146F9BE2B249B9E4F0755D59C1B3C0";
    attribute INIT_03 of inst : label is "A4439E71381D431285C471FDABBB31328186564E5A8387D9052562176E9E975A";
    attribute INIT_04 of inst : label is "792182E10104B1B50020E940C1334CF084963471A82A7A7AFD7DF5F5F2B831EF";
    attribute INIT_05 of inst : label is "A237D2AA2F432D1A3A3E68A504AF00D7E4D114523C1162AA84F0C4160C8630D4";
    attribute INIT_06 of inst : label is "99999999A99267AC7D7584E43AF918C1708F7CCFE25AAFFD7796FB63FDCFD23F";
    attribute INIT_07 of inst : label is "7501440408882AA0414548C10C88BC32289B31806EC30C036A24086941BCD719";
    attribute INIT_08 of inst : label is "AFBDF7BB6DB6EA6B53ED4B6FBAAFFC1AFFF7F6E3D3D3D3DFFBEEEFBFBFFFBFFF";
    attribute INIT_09 of inst : label is "126374DDB56DB6DB6CB31E5D9D6B7B76730D30EDBFF6D2763FEB2CBA8FB6DD96";
    attribute INIT_0A of inst : label is "3A6C78CDB66347BB676EF7373BFFFFFFFDF755F7F41BB6DB6DFFFE63BBBE5377";
    attribute INIT_0B of inst : label is "8E23E08A1F090675E0FFA8F8C78C5707A2B8363C67BD3FEF3E1209F3E339F4CB";
    attribute INIT_0C of inst : label is "1F6C0EDA4C9EE6B5E1F1F3CD5349678B46EECCF42B55791AF28A0AC2A5A9BF77";
    attribute INIT_0D of inst : label is "DA2FE36C993DCD6D707472D39A4B3C5B7F3C4DA4BA0CB234B173F8606576D2CA";
    attribute INIT_0E of inst : label is "6B397D5E74186A1A69F8777398CC5267EAECC8ECC6F9A282CF35718368A97D65";
    attribute INIT_0F of inst : label is "80000FD9606FFFFFCCCCCD6138E38E1E0000002EBFEFAFAFBBBBEFF321FEFD36";
    attribute INIT_10 of inst : label is "7B9799CD844CC62F41315B56C176E6E3932EFEFBE27AFAE7A43E5671C49A7A49";
    attribute INIT_11 of inst : label is "0456EA508788543EC6D2CDAD32C8D8D7D73A371980E199998DD109933AFC186E";
    attribute INIT_12 of inst : label is "A2F9FAE5C86B23228888755AAC5DBAE909E76A65DB85E606FE23B82D23FBC6C9";
    attribute INIT_13 of inst : label is "AFE63FB92C93364DB0A4398B16B2C436E4C6445386E0B0B03435B5B5B03037A0";
    attribute INIT_14 of inst : label is "C1A9220754B4AB6CC069A090BDFDE360C08139270A04F85C7668138C43A9A80E";
    attribute INIT_15 of inst : label is "F7F9DDC7D0C71C73C0E8C7139C703EA9F8C1C12C236DE14AA9598914B06A6A86";
    attribute INIT_16 of inst : label is "F5A4BBB1DCAB729DEE456A0F08C982EE9F8EEE577A8DDD444F91915557574C6C";
    attribute INIT_17 of inst : label is "F38A667C2D8C1C8BAB713AD33044905C416C416C456C456F1FF5635F39767D57";
    attribute INIT_18 of inst : label is "FAEA9B4D16D6D740E8C716D345B5B4BD450A33DDD6CD0BCDCEB142EEEA6D37BE";
    attribute INIT_19 of inst : label is "D236DCBEFFFA7C30D7C89B6BDA557B4FDB331EC7FB0D3FC76CFFC30EB59CA239";
    attribute INIT_1A of inst : label is "38FF7CEE1199999951C71C713C39DD9973CDA0EF9EE7B5E9BEAFF6EF772B3BBA";
    attribute INIT_1B of inst : label is "74F371FD6667D2054F3336A68D8DE63CAD1E17F9C2FCC2FCC0BC700DBED5CFAB";
    attribute INIT_1C of inst : label is "3209311A9D30913B6E69E26DF364DB3CCFBDB4D47B7A9FC6A22B333FDC3CD57B";
    attribute INIT_1D of inst : label is "E6B0E8820912A612331FDD1C959F94D35B68A63CDE0F846BEEC0EC3A7B137642";
    attribute INIT_1E of inst : label is "A15BFBB0E7F1787CDDD1CD0AA39A8DEE333ADB9A799F6CC971DB33EF6D371A9E";
    attribute INIT_1F of inst : label is "824F7C9E828C9EF9D105193D8D220A32D73B44146BD7AEB769AE96DA2C8A3783";
    attribute INIT_20 of inst : label is "E716CD51E0EBD7D26D50BBD38D22567795BF4235F25311FBF51B8CA72FB0819B";
    attribute INIT_21 of inst : label is "77AC8E76A8890807574F4943621175D2FA4312793F2CFE53E436F88E0C105196";
    attribute INIT_22 of inst : label is "1FE2471768269DEE7C2197F7F6B85AD2FD9DE1452CFCDD1F5B07E77051E11690";
    attribute INIT_23 of inst : label is "CC5C241E5FDAEEAE50054005FEF5BAA6DD6D6D52395312727DEC947930755513";
    attribute INIT_24 of inst : label is "C8179455EBE3B35A07C60CC131E26C5489794BBEE6D5C90D633A027CC0E02E55";
    attribute INIT_25 of inst : label is "3B4D06CBC843A8D317A90D62BC13471C57020202C84040CB18C11960298CCE30";
    attribute INIT_26 of inst : label is "958E19A6EAB64389A219C28C9A34CB2CCB63CC5CD4639D5026BC53679800B8BC";
    attribute INIT_27 of inst : label is "C9BCBB880D44DC8C8D49BCAB1206D46D590B9ACB969B917292F81058A24141AF";
    attribute INIT_28 of inst : label is "49ECC6709B2198B49C339C33253219B208DF19C33CC632C37080CCE327716306";
    attribute INIT_29 of inst : label is "E7EE3C83E34CB3738C83301F5CDA5A07091EC84022CBCB18838367CC4CC62E89";
    attribute INIT_2A of inst : label is "EDBBC38C9FF465700FFCB6EA9F758EA09C31217D389CF7736B322F62F58FCF03";
    attribute INIT_2B of inst : label is "D9F104B8AA932ED474CE1690140145FDB7F22189F8F59BDFC75FFFFFFAD9D49F";
    attribute INIT_2C of inst : label is "ADDEB3174D79AB27B346A64513D607860B8B2805AF5BFF2BA4232321843B2EEC";
    attribute INIT_2D of inst : label is "E3C3BFF4B152C5D7FEB81FFFFF145005A0E6ECD3A1E2EC87317392A0CD4CB5E4";
    attribute INIT_2E of inst : label is "48A8AB4355C7F5DECF29AAB0B63C58764EF8FA2BCB1A3FA7BC53A1EA33333736";
    attribute INIT_2F of inst : label is "C000000000000001B123C7C8141D45078F1F20BF2FAB76CA9E7FBAAAAAAA028F";
    attribute INIT_30 of inst : label is "5AA45ED75A022A03D1791A6C3E08C11F43B42D4244083605401F06D5D5D9CA51";
    attribute INIT_31 of inst : label is "694AB695ED96AB947E8D5C7544CCC8807AC005151631D40A9997555BA5DAB7B4";
    attribute INIT_32 of inst : label is "40DC48D5E3CAFB0574C794B5F23BFACC0E8BB0C1917580B86B561EE055FDCB69";
    attribute INIT_33 of inst : label is "B40CA8AA6AAB99D43511B15460740AAA517518555040C0D4743C9870F5056161";
    attribute INIT_34 of inst : label is "DFF774FCE4104EEDD7DF7DFDBCF337497DF77767FED053DE554B20D3B7A557CA";
    attribute INIT_35 of inst : label is "440000001040204010157DD7DF7F2DE0F9E5F67BF1548856FD9776969F2675D3";
    attribute INIT_36 of inst : label is "818AA977F89F57FD3022A000028A00A250000001114110114000580802440212";
    attribute INIT_37 of inst : label is "5B9ABFE9E88080B82D75BE45202A08F414010404145CAC12A510175E8105C567";
    attribute INIT_38 of inst : label is "AAEABABEBEAFABEABA01BE8BFFA07FE82AF156AF3ABCFA2DC6BE8A31AD47ADAF";
    attribute INIT_39 of inst : label is "FA2BE8A34FD50EBFB1BFAAAC7FD7FFEBFBEEC2AFABAFF7B71AAEAEBFFEAFAEAE";
    attribute INIT_3A of inst : label is "DCC8F78F555FFFD7AFFEABAED7D77555FFFAFFFFEFEFC02FF02FFA0BFE8FAF1F";
    attribute INIT_3B of inst : label is "10129971B02FF10F47DEFB38DFFBDFDBFFFDFFFFFCFCFCFCB9BCFFFFFAFAFF55";
    attribute INIT_3C of inst : label is "FFFFFFFFD280401C067950301547FF8FBC7FF7EFEA183FECEE1785FFE57BBD5A";
    attribute INIT_3D of inst : label is "8AAE9FC43FDD6FAAFABAFA11FF75BEABAEEBAC47ADC32FB0EA2FBB194E7FE7BF";
    attribute INIT_3E of inst : label is "0B38C8C2741C6CD7EF91AB8FD22375FDC412AFB9FABFC3FAA2ABA7F10FA71FFA";
    attribute INIT_3F of inst : label is "A5BABA3679F57DD9B38B7BEFDAFD5FDEAF32FAFEAFAEAD77657DDA047162FFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "E3E3E3EC35FEFD75E6A9C662AA1555F5E0F5F5D9B4BBFAF22D849F797D3AD3D3";
    attribute INIT_01 of inst : label is "958899E5DBF775CA5334FD722CF941FC79EFE5F6FF7B9F6DAC906DAFF24CECEC";
    attribute INIT_02 of inst : label is "F6897E3F77A6039FAD3DFF5B6DA9B6F99E68C34455DF157FFE9BD3CB5A9113D7";
    attribute INIT_03 of inst : label is "5BFDF79FBBEBFEC8F8F93BFA9999E6643B28293B45D6C5467ADED5EA3D7E6F1B";
    attribute INIT_04 of inst : label is "A6F472D5949063C7ED8574F3AC94F063FD6DD5D57AFA727275757575FAFFFE7E";
    attribute INIT_05 of inst : label is "77FDF7FFCFF165B4F0E7A7B7D9B1F9775766C7BDEB76FF18FD9C37E9D62DCA2B";
    attribute INIT_06 of inst : label is "BBBBBFFFABAAEBBB8FBE7F3E19349A6B3FD4CB5D847B1F9BEBDFED5D93D1AFDB";
    attribute INIT_07 of inst : label is "FFFFFFFFAAAAAAAAFFFFF5BB0866BC016B9179AE67C66F1E9A9E5D6A963F1E5F";
    attribute INIT_08 of inst : label is "D881B9B8679C75FF96FDFD70B4E4E9F5E1B18DB59292929BF5F5F5F5FAFAFAFA";
    attribute INIT_09 of inst : label is "F7F6ECF3BD77BCD177FFE3EDCDF3CFFCC6BDE5E3F9B6DA6ED053FFDD18DECB9E";
    attribute INIT_0A of inst : label is "3D751D6974626EA6ABD7EC6C9AAAAAAA0A0E992C2D5F867BDC0E5F5D5BDA4743";
    attribute INIT_0B of inst : label is "997B9DE889278E9E9CB25EE36EA219A05A870B7D1BC70D3B18471F073949D549";
    attribute INIT_0C of inst : label is "E3FCE7FD7DF09D9CB4B4A5F5CBFDF7D75333F8B1D2EAAEDA276FE7F97B9BDBBB";
    attribute INIT_0D of inst : label is "FD3DB7FCEDEB2D2F35B5E5F457F7ECE3236D957B5EDAFEBE99B7AF35BBEAFA5A";
    attribute INIT_0E of inst : label is "F7EF65D9DEFFF9DE048123F5AA6CB8D925CFD5BFD52FF7DFDF5FBEDF7D7B4F3F";
    attribute INIT_0F of inst : label is "80001F49CBE99991EEEEB1AC9269A6BCA0A0A0DB4F1F5F5F1E5B5FD4FF370F69";
    attribute INIT_10 of inst : label is "347DDCF0F3B3A8F4A545BCE7615DDDD4ED91351579BBC63293852985524787FE";
    attribute INIT_11 of inst : label is "ABCDB5FD7959F3A5FDA9F4F3F57D367DADF18DDB993C7AD6F0F7B2FDBB102191";
    attribute INIT_12 of inst : label is "7FEDFFBA3B858EE8AAAA801F5B2268146F18DF8F9B5D57171B8F4FDA9F6F3B5E";
    attribute INIT_13 of inst : label is "D15DF9ECDB6E699AC9F27FCDE261D9EA7F5117FACF5909090D0D8D8D89898255";
    attribute INIT_14 of inst : label is "A4949C9C953536757576B3C3B9F9F9FBA7A4949C9A9AEBDB9D064912F4BABAF2";
    attribute INIT_15 of inst : label is "F1B3E4ED97BE15552DF7FD94D55634B2F863BFF3CDFBADCBF806E347ED2322A2";
    attribute INIT_16 of inst : label is "ABFE677AE80EA66E9DEAFFA362E719861A3F44283D3E463B899B9A0A0E0E7ADE";
    attribute INIT_17 of inst : label is "93BFC9A48A026862FDF47DBEAFBC6FA67752775277577757D28AE602D52D2F38";
    attribute INIT_18 of inst : label is "EAF23F9DB0F0FBF78BB0E7E7ECB4B5ECF1FFE4ECF6FEF9FFFC74C5D69A4AFA26";
    attribute INIT_19 of inst : label is "BECBB37FE5761DA4B468B7FD40C4C353B7A2E3B46EB06CBD78D1EF516BF4EEBB";
    attribute INIT_1A of inst : label is "6CFCEE8888888993E4B2CF3C86BE3B912FDFD7DAC27C3503757B29704E6F5D7B";
    attribute INIT_1B of inst : label is "BDEEB48AFCEEF8BFDFF9496DA7AB42947F42367F9F7F9F7F9A5F0F7FDF7D3F7F";
    attribute INIT_1C of inst : label is "F1FFF7F3B1DEFDEAF9DDB6FDB3B5F7ECA3F3F3CD289FE756DDFFE7F2AF7EAD23";
    attribute INIT_1D of inst : label is "F3DFAFFFEDFC73DFE346A979F17DE557EDD7D3FDF671D99B77E1BF66EEB6BFDB";
    attribute INIT_1E of inst : label is "76279E7A62389F87AAB7BA753FB8A166FD5D9E574A9B5E8F2FDF3BDEFF564FCA";
    attribute INIT_1F of inst : label is "C1BD6EEF08A66F99F6B146F5AFB822999B577A45239E4B66105FD957D7DF5D7D";
    attribute INIT_20 of inst : label is "B149922EFAA478B4A76FF4691D8C5DCD7CBD9DD1BCFD7A905FECDA0B017E7773";
    attribute INIT_21 of inst : label is "E6F5B1E9FD7CBED4F5E4E5DFDDD777BCA59CD7A5D2E3AB86727935B1DAABE648";
    attribute INIT_22 of inst : label is "C6BEDAE6931862CD8FECFAD58E4BA67BC6C69C64CFC7C3C62F9939292ECDC77B";
    attribute INIT_23 of inst : label is "37FF7FAFFFFBBAEFAABBEB7DADCFB0625E9690CDDE4DBD0D83CB7E7AC7CE7B5B";
    attribute INIT_24 of inst : label is "9B73D7B0F794DC23596DED39D6F4B38846DAF3C5ECB876971BFE34B3BB7AD37A";
    attribute INIT_25 of inst : label is "F5F6FDE5FFF5F5F5F9E5F7F9F537F5D574E4E4E4EBEBEBE6E023B123A66E2D5A";
    attribute INIT_26 of inst : label is "EEDBFF2FEC73EB17BDC6F9FF61C3AEBB578F5B4F6FDF5F6F9E5B7F1F5F774F5F";
    attribute INIT_27 of inst : label is "946FFF5D326FABDAB6946FFFAB79B8983DFF5D2F7F7F5ECA7F7A6D2A1B2D2B7F";
    attribute INIT_28 of inst : label is "FCF9D3B5F7F6F5C56DF56DF5F157EDD7FDF54CB7F6BEFAD1B7F3FBFEADBBFAB6";
    attribute INIT_29 of inst : label is "6C63FEA0B47956FEDF5FB23BEDABFFA3996FBF349B69736BA0F5D1B9F6B98BBB";
    attribute INIT_2A of inst : label is "DB3FFDEF82B0469A5FABE7FC0CA8A4CB9ACBD24F4F85CDA265DF354D7E4383E6";
    attribute INIT_2B of inst : label is "4BBD927D2871F46A7FF7992A81DC075A693B54560D6F5C926F5F5F5E34DD57D7";
    attribute INIT_2C of inst : label is "18DBE2B4E9D75F3D71B898EC41B9B1EDC283B9F87A8BFE6AC474D5DEE8CCDEEA";
    attribute INIT_2D of inst : label is "94532596C17D27F9F3AC65F5F5A1D9EE9EDC66DA9AFC9AB6A1C356E7EBBB7F54";
    attribute INIT_2E of inst : label is "E9E8FF9B987299876D934C960F6798246EC659DEEDBC5FF74E583F571B1B1B18";
    attribute INIT_2F of inst : label is "0000000055555551939A6B66C7CE71F3E98DBB2DB0F3C6DDF9CAC7FFFFFF5BEF";
    attribute INIT_30 of inst : label is "3BD42786BD7CD57CF1E5C94DB5B6E1DDE8EA23FFD74FE32A65E8FEE6A92FCB3A";
    attribute INIT_31 of inst : label is "B7FFE177D599FB7425CCBFF0CFB5F7BF87BFF3F3FEFB8BD6DDF4A3B0EBBCBFDD";
    attribute INIT_32 of inst : label is "AB4FFE0B139381E1E33E7FFF4EFE15866028081E785BFB55974BDB250F4E4D7D";
    attribute INIT_33 of inst : label is "75E1EDFE420AE5D305055DF435754200FB9FB2FF5F5E7C7FC62FDF5F1FAFFE7E";
    attribute INIT_34 of inst : label is "5F438619022A9B18422ADB194B0E82984B0FD2DA440505250A2B57D187B55552";
    attribute INIT_35 of inst : label is "F5F5F5F5F5F5F5F5F5F4D9422A8A98031D570FDF174C01D41946873F554D8D21";
    attribute INIT_36 of inst : label is "00AAAA00A2A008AA8A02AABFAAAAAAAA5F5F5F5F5F5F5F5F5F5F0F5F5F5F5F5F";
    attribute INIT_37 of inst : label is "DEBFFDEA3FFDDEABFABDFFAF0BDDDDC9E97FF96FEB0F5FBC4FF17BBF7FF70785";
    attribute INIT_38 of inst : label is "559565516559D67565A0F56BFC55FF95BFD5F45BAC6EA0BEF7F56FF5FEFFFFFF";
    attribute INIT_39 of inst : label is "F5EBD4F7BFF8F57FF5F95FB5FFA7FFD7FBFBF3FBFA5FBFFAFFEFE57FF87FF852";
    attribute INIT_3A of inst : label is "CBDBEFBFAAAAAAAAFFFFFEFBA8AAAAAA5F5F5F5F5F5F5F3FFE3ED50BB94FFC5F";
    attribute INIT_3B of inst : label is "ED51679ECFF515A2BB6FFE63AAAFABAD5E5B5F5657575757521E5F5F0A5A0A82";
    attribute INIT_3C of inst : label is "F5F5F5F5EDFDF5FDF1BFFDF5FF4FFFFFFFEAABFFAF8FFFFFF5EAF2AABFAFFFAB";
    attribute INIT_3D of inst : label is "7FE57FFDFFF8FFF5FFB5FFF5FFC1FFD7BAD7FDF7FE7BFFFAA5FFFEBDEEBFFFBE";
    attribute INIT_3E of inst : label is "F5DB7BE9189BE47077AABFFEA803FDF05A4ABFFF55FF5FFF5FFB5FFF4FFC5FFD";
    attribute INIT_3F of inst : label is "3CA1F5F2EFAFE1DB575567F57EEF84D3B5FBD7F3DFEA7D57D7FFDFA355455F5F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "06060604A174EE73C4909BE02A37C434200000F9EC0F22EA91A295D3D4C922A1";
    attribute INIT_01 of inst : label is "E7C8ECA51FE776FF625129062C7948F504D5D165DEDBC61879C509A1B2300808";
    attribute INIT_02 of inst : label is "20FF1785C8828D247A1B638D26909250510E0D224FCF23EC67DCD6335D604037";
    attribute INIT_03 of inst : label is "A338638E918558032F2ECE8833330006467C6C369306099C630304E649253050";
    attribute INIT_04 of inst : label is "548413C8347512008C1009A25902A516083001840220888008880888084CC832";
    attribute INIT_05 of inst : label is "12FA0325405094891192D7629044F109861B36C418DA9D04184002253E08C25A";
    attribute INIT_06 of inst : label is "EEEEEEEE01140116724B61CA920892492E99131C425916659F1A940056984C02";
    attribute INIT_07 of inst : label is "2888222000000000AA22AE67A20DB2888650E01967846B244388A08A200DCB4A";
    attribute INIT_08 of inst : label is "BCB68174632C9138D4B08935F5F5F1B105F17D28D6D6D6D0A575957470D8D262";
    attribute INIT_09 of inst : label is "CDC5DC770933BC9167B9D4B4D131E8E885F5D0D390A2880044A69A40482043C0";
    attribute INIT_0A of inst : label is "3B342D6D60025C80DDE14909295757570A0ADC090987547BCD1E4C155BD43054";
    attribute INIT_0B of inst : label is "DC40918B01AE08B65C2D3C0594523BB0D3D786A092D38B670954164122D8814B";
    attribute INIT_0C of inst : label is "91E4E6F9392A1939938181E4B19536D6CA4B61BDF9F0A2C2A3ACE331CB36D199";
    attribute INIT_0D of inst : label is "797991E4244E20EE9444C52484B0E0A2E300C51F1D929C885A918E9448DA20C8";
    attribute INIT_0E of inst : label is "1CB308C35A386B3A300C00C6055AA87B21C75CB65368EE0E4F1319116567624C";
    attribute INIT_0F of inst : label is "400075C6850BBBB344466CD969861A9AA0A0A09450401246471E4DC14A70065D";
    attribute INIT_10 of inst : label is "5331696571B23350E011ABE2741B1B3574ECF2F86DCB0F2DA6C27A890324E5B7";
    attribute INIT_11 of inst : label is "EDB050697C7A93D374F47325C51D4F10F184B4C08ADA32626530E36609E231C0";
    attribute INIT_12 of inst : label is "4CBA326F936DA66800002005F61DA2B8121F9243C9336F250109374F4C125842";
    attribute INIT_13 of inst : label is "9F980CDB698A5695BF67D8F384D309A0411946CC893B1B1B1E1E9E9E9B9B9407";
    attribute INIT_14 of inst : label is "89C140302444549100C186367272EC6C8C8941403228A328FAF73C4CB93626CC";
    attribute INIT_15 of inst : label is "26C49930560CC5365A65B429CD138420C1064CE686EB6663702DD21766D4F488";
    attribute INIT_16 of inst : label is "3528F20140A806C4C8854834C04DB0081132087C486D9A699C08080506044C03";
    attribute INIT_17 of inst : label is "E0B638782D95024B6C01D87806B81E9893649364916491654087885F8069616B";
    attribute INIT_18 of inst : label is "2A83A1B5B43474BFF924ECEDA58593ADC5349331602242E261D08376CAC2C9B2";
    attribute INIT_19 of inst : label is "909A36BC112455807D4030FDD05772027081872184B82A6D40E127409B340CB2";
    attribute INIT_1A of inst : label is "7472E7D588088889B16DB2C9605D3800494F91C9CC4F30186EA0082406061873";
    attribute INIT_1B of inst : label is "C81980332020688C819A28DCD683A55A77AC0271177115710A564EA3194C1A5A";
    attribute INIT_1C of inst : label is "913991A364646449E0B191E5909125E423A18182201564D2313991A372226408";
    attribute INIT_1D of inst : label is "517E0CC660E485C4922734006EFB3BCEE9C64494703198C0C7208F220480DC88";
    attribute INIT_1E of inst : label is "A63231CAE2289F0E3322224E108951AA1923180C475842060A1818CA4243ADC4";
    attribute INIT_1F of inst : label is "42EF261807548F0832AC2B9C8E301D5259146A30B8D1C421581D9851930C1C64";
    attribute INIT_20 of inst : label is "6C142C7D99D53527C63D9035FBE53BA0E932F4E5DE27AA3AFE6403FD7AC60661";
    attribute INIT_21 of inst : label is "B5216D84FC686DB0A1A0B48E618637BD14F9E2D141E11BE28238C06CCBFAA09B";
    attribute INIT_22 of inst : label is "C4788CB430968A6EF21B61D42CE22C7093D7CC1E0ED6D2982BDD7D6C6C1B951B";
    attribute INIT_23 of inst : label is "E3A7E15DEBFFBCFA5500036B0EE672C932D0C38CA60CCB45C7D649770C180C41";
    attribute INIT_24 of inst : label is "EEE721F5F7C001B77505AD2D448081E50DC1E3409800122B98125097CB4201AA";
    attribute INIT_25 of inst : label is "D1A4B4F17D9445659151E4D4C1A498E1F380008001898928640610A6120600C2";
    attribute INIT_26 of inst : label is "7D05F611C9E140BD64662832DB0008211B0C3616494C164F45124B4417EF1717";
    attribute INIT_27 of inst : label is "AB9719E6A0448B88A12B9719A2B2A0204C091C5C19741E08400E1916485C5821";
    attribute INIT_28 of inst : label is "68240A50264424FB940094003E65C06580020920A824A2025022BFE98E59E0F0";
    attribute INIT_29 of inst : label is "C1C23CA11701449F8349920F45A8CCA091342504AA4BE103A145842060644322";
    attribute INIT_2A of inst : label is "8AFB65354038CC025E8F772B8C9A44014A6D0A065AC90FB35B560A4E11469EC6";
    attribute INIT_2B of inst : label is "86993779224B42C0C8DD83E1A3682E421C1E290A4508451D5F5D5D5F664F3306";
    attribute INIT_2C of inst : label is "340810A3A00E5F9D700CCCC224B111ED02C1919D00C344AA55362F0B74882808";
    attribute INIT_2D of inst : label is "94172110046C3220B21C50A0A01408B8540D2472BF0787258196CED227E6C810";
    attribute INIT_2E of inst : label is "4C0C80D33C429B44450822548425BC2E8DD25C8680118FE446723F0B13120212";
    attribute INIT_2F of inst : label is "8000000055555551D12149488E84E3A1C50531652FAAA640B1A8800A00000AC0";
    attribute INIT_30 of inst : label is "6450143225C4B5C521F8BC8CB5C22BA8BF6CF46CA2936BD380BDAB11101F16EA";
    attribute INIT_31 of inst : label is "472A0D0491B12C44D093D5AD61F13F7BD410240424098B8031B6C5E5B9F8DD54";
    attribute INIT_32 of inst : label is "F6DFBA8EBBA8326BAF7B286ECC88922C332E5F5D0F1A4F4D504DC4703E170048";
    attribute INIT_33 of inst : label is "1F514555E28E24864520A1FE212008220B2D18520F0F4294620A0A5D2D052E2E";
    attribute INIT_34 of inst : label is "CFF786C9E7BEDF99E32ECEC96B8E86D93EDBF24F34CF2D25AAFE2279C010550A";
    attribute INIT_35 of inst : label is "20A0A0A04125D1A520A0F9E33EFE0912CD36DBCEC70C21C4C90687FBCF7D8DF3";
    attribute INIT_36 of inst : label is "757F7F5F080A00025FD7FFE800000000020A0A0A020E070E0A0A0A020D0A0D04";
    attribute INIT_37 of inst : label is "A1E5E20380000146A38A088ABE0000400BC20BC20B0F030D0A0FCA080F02D2D7";
    attribute INIT_38 of inst : label is "AAEAFA16ADA3E8FA7AA132A5F5A5B5A980D42081FA02FA38D4328455F84022DA";
    attribute INIT_39 of inst : label is "6A55A8C50554761551D484F461C071E9F0F5C4751A8A7ABB11F47215FA2A0A86";
    attribute INIT_3A of inst : label is "86F9E39FAAA2AAAAE55FFFF5A8A8AAAA5F5F555D5F5F571F740548065E840F5E";
    attribute INIT_3B of inst : label is "F4F8BBEFBDF545D5D9FFB703AAA4AAAC1D1B1F5B585A5A52131700000F55018C";
    attribute INIT_3C of inst : label is "F5F5F5F5CEF4C1A0575551F51BE5F450A59574E1DFBAFAAAA0F5F5557A5AAAD2";
    attribute INIT_3D of inst : label is "B5E295D575FC60AAF4AAF07585F5B4E994A985551A504A1AAA35D1B502F8AAC3";
    attribute INIT_3E of inst : label is "9FE7B3F5801BC6F8FBFF291FD0A2A020564E4657585F530AAD52A557405F505E";
    attribute INIT_3F of inst : label is "AFFBFB7BFE20085E164D769F1FE2A62F4F5A5D474B107975E555DF204E4ADF5F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
