library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity joust_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of joust_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"00",X"08",X"BD",X"E0",X"0C",X"BE",X"5E",X"E9",X"BD",X"E0",X"15",X"86",X"02",X"BD",X"E0",
		X"37",X"BD",X"3B",X"2E",X"8E",X"D2",X"24",X"BD",X"E0",X"15",X"BD",X"3B",X"5E",X"CC",X"6C",X"55",
		X"8E",X"1C",X"BD",X"BD",X"4A",X"53",X"10",X"8E",X"12",X"11",X"BD",X"5E",X"E6",X"8E",X"CC",X"00",
		X"BD",X"3B",X"31",X"4D",X"27",X"23",X"CC",X"F7",X"33",X"8E",X"1F",X"AB",X"BD",X"4A",X"53",X"C6",
		X"CC",X"34",X"10",X"8E",X"CC",X"00",X"BD",X"3B",X"31",X"35",X"10",X"85",X"F0",X"26",X"02",X"8A",
		X"F0",X"BD",X"4A",X"56",X"86",X"F8",X"BD",X"4A",X"53",X"86",X"01",X"BD",X"E0",X"37",X"8E",X"D1",
		X"5B",X"CC",X"11",X"FF",X"BD",X"E0",X"09",X"8E",X"D0",X"ED",X"CC",X"10",X"FF",X"BD",X"E0",X"09",
		X"CE",X"D3",X"5D",X"7F",X"BC",X"1E",X"A6",X"C0",X"B7",X"BC",X"1F",X"A6",X"C0",X"B7",X"BC",X"0A",
		X"EC",X"C1",X"FD",X"BC",X"08",X"4F",X"E6",X"C0",X"F3",X"BC",X"1E",X"FD",X"BC",X"00",X"4F",X"E6",
		X"C0",X"FD",X"BC",X"02",X"4F",X"E6",X"C4",X"27",X"11",X"F3",X"BC",X"1E",X"FD",X"BC",X"04",X"4F",
		X"E6",X"41",X"FD",X"BC",X"06",X"BD",X"D2",X"A8",X"20",X"DB",X"33",X"41",X"E6",X"C0",X"27",X"02",
		X"20",X"C9",X"A6",X"C0",X"27",X"05",X"B7",X"BC",X"1F",X"20",X"C0",X"DE",X"2E",X"86",X"6F",X"A7",
		X"4D",X"86",X"0A",X"BD",X"E0",X"37",X"6A",X"4D",X"26",X"F7",X"CC",X"00",X"40",X"BD",X"E0",X"0C",
		X"10",X"8E",X"A0",X"10",X"CC",X"FF",X"FF",X"ED",X"A1",X"CC",X"00",X"00",X"ED",X"A1",X"ED",X"A1",
		X"ED",X"A1",X"ED",X"A1",X"ED",X"A1",X"ED",X"A1",X"A7",X"A4",X"7E",X"5E",X"E3",X"CC",X"FF",X"FF",
		X"ED",X"4D",X"CC",X"D2",X"2C",X"ED",X"C8",X"10",X"86",X"02",X"BD",X"E0",X"37",X"9E",X"1E",X"EC",
		X"4D",X"2A",X"0C",X"10",X"AE",X"C4",X"A6",X"22",X"81",X"11",X"27",X"3B",X"CC",X"00",X"10",X"27",
		X"23",X"C3",X"FF",X"FF",X"ED",X"4D",X"26",X"2F",X"10",X"AE",X"C8",X"10",X"31",X"28",X"10",X"8C",
		X"D2",X"54",X"25",X"04",X"10",X"8E",X"D2",X"2C",X"10",X"AF",X"C8",X"10",X"10",X"AF",X"C8",X"12",
		X"86",X"08",X"A7",X"4F",X"10",X"AE",X"C8",X"12",X"AE",X"A0",X"10",X"AF",X"C8",X"12",X"6A",X"4F",
		X"26",X"05",X"CC",X"00",X"57",X"ED",X"4D",X"DC",X"1C",X"DD",X"1D",X"DC",X"1A",X"DD",X"1B",X"DC",
		X"18",X"DD",X"19",X"1F",X"10",X"D6",X"17",X"DD",X"17",X"20",X"9D",X"6F",X"C8",X"15",X"8E",X"00",
		X"0F",X"10",X"8E",X"00",X"10",X"86",X"08",X"30",X"01",X"8D",X"30",X"8C",X"01",X"2E",X"25",X"F7",
		X"30",X"10",X"31",X"2F",X"31",X"21",X"8D",X"40",X"10",X"8C",X"00",X"F2",X"25",X"F6",X"31",X"30",
		X"30",X"1F",X"8D",X"17",X"8C",X"00",X"66",X"26",X"00",X"8C",X"00",X"00",X"22",X"F2",X"31",X"3F",
		X"8D",X"26",X"10",X"8C",X"00",X"10",X"22",X"F6",X"7E",X"E0",X"0F",X"4C",X"84",X"0F",X"8A",X"08",
		X"AF",X"4D",X"10",X"AF",X"4F",X"ED",X"C8",X"11",X"C6",X"10",X"8D",X"46",X"31",X"21",X"4C",X"84",
		X"0F",X"8A",X"08",X"5A",X"26",X"F4",X"20",X"1B",X"4C",X"84",X"0F",X"8A",X"08",X"AF",X"4D",X"10",
		X"AF",X"4F",X"ED",X"C8",X"11",X"C6",X"10",X"8D",X"29",X"30",X"01",X"4C",X"84",X"0F",X"8A",X"08",
		X"5A",X"26",X"F4",X"EC",X"E1",X"ED",X"C8",X"13",X"6A",X"C8",X"15",X"2E",X"0A",X"86",X"03",X"A7",
		X"C8",X"15",X"86",X"01",X"BD",X"E0",X"37",X"EC",X"C8",X"11",X"10",X"AE",X"4F",X"AE",X"4D",X"6E",
		X"D8",X"13",X"34",X"36",X"86",X"00",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"1F",X"10",X"44",X"56",
		X"1F",X"98",X"E6",X"65",X"1F",X"01",X"86",X"0F",X"E6",X"E4",X"25",X"06",X"58",X"58",X"58",X"58",
		X"86",X"F0",X"A4",X"84",X"26",X"04",X"EA",X"84",X"E7",X"84",X"86",X"01",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"35",X"B6",X"00",X"00",X"07",X"3F",X"05",X"FF",X"E8",X"E8",X"00",X"01",X"03",X"05",
		X"07",X"05",X"03",X"01",X"00",X"08",X"18",X"28",X"38",X"28",X"18",X"08",X"00",X"00",X"40",X"80",
		X"C0",X"80",X"40",X"00",X"00",X"09",X"1B",X"2D",X"3F",X"2D",X"1B",X"09",X"00",X"09",X"52",X"A4",
		X"FF",X"A4",X"52",X"09",X"34",X"10",X"30",X"01",X"FC",X"BC",X"1A",X"B4",X"BC",X"09",X"34",X"02",
		X"B6",X"BC",X"1A",X"A4",X"84",X"26",X"0F",X"E4",X"84",X"EA",X"E0",X"E7",X"84",X"1E",X"01",X"5C",
		X"1E",X"10",X"26",X"E4",X"34",X"02",X"35",X"92",X"86",X"40",X"B5",X"BC",X"16",X"26",X"08",X"FC",
		X"BC",X"00",X"83",X"00",X"01",X"20",X"06",X"FC",X"BC",X"00",X"C3",X"00",X"01",X"FD",X"BC",X"00",
		X"39",X"7D",X"BC",X"16",X"2B",X"08",X"FC",X"BC",X"02",X"83",X"00",X"01",X"20",X"06",X"FC",X"BC",
		X"02",X"C3",X"00",X"01",X"FD",X"BC",X"02",X"39",X"7F",X"BC",X"16",X"FC",X"BC",X"00",X"B3",X"BC",
		X"04",X"76",X"BC",X"16",X"2A",X"05",X"43",X"53",X"C3",X"00",X"01",X"FD",X"BC",X"12",X"FD",X"BC",
		X"10",X"FC",X"BC",X"02",X"B3",X"BC",X"06",X"76",X"BC",X"16",X"2B",X"05",X"43",X"53",X"C3",X"00",
		X"01",X"83",X"00",X"01",X"FD",X"BC",X"14",X"7F",X"BC",X"0B",X"43",X"53",X"4F",X"F3",X"BC",X"12",
		X"24",X"03",X"7C",X"BC",X"0B",X"FD",X"BC",X"0C",X"20",X"03",X"BD",X"D2",X"78",X"FC",X"BC",X"10",
		X"F3",X"BC",X"14",X"FD",X"BC",X"10",X"34",X"01",X"7F",X"BF",X"FF",X"7F",X"C9",X"00",X"FC",X"BC",
		X"00",X"47",X"56",X"1F",X"98",X"F6",X"BC",X"03",X"1F",X"01",X"C6",X"F0",X"24",X"01",X"53",X"1F",
		X"98",X"53",X"FD",X"BC",X"1A",X"B4",X"BC",X"08",X"E4",X"84",X"34",X"04",X"1F",X"89",X"EA",X"E0",
		X"8C",X"98",X"00",X"24",X"34",X"E7",X"84",X"7D",X"BC",X"0A",X"2A",X"03",X"BD",X"D2",X"54",X"86",
		X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"FC",X"BC",X"0C",X"83",X"00",X"01",X"26",X"08",X"7D",
		X"BC",X"0B",X"27",X"17",X"7A",X"BC",X"0B",X"FD",X"BC",X"0C",X"35",X"01",X"25",X"9C",X"BD",X"D2",
		X"91",X"FC",X"BC",X"10",X"F3",X"BC",X"12",X"20",X"9A",X"32",X"62",X"35",X"81",X"44",X"00",X"11",
		X"11",X"02",X"50",X"03",X"64",X"08",X"74",X"0C",X"7A",X"14",X"7F",X"1E",X"7F",X"26",X"7A",X"2A",
		X"75",X"30",X"64",X"30",X"50",X"00",X"01",X"00",X"22",X"22",X"1C",X"5C",X"1C",X"55",X"1E",X"50",
		X"20",X"4B",X"00",X"01",X"00",X"11",X"11",X"20",X"4B",X"23",X"56",X"23",X"5E",X"00",X"01",X"80",
		X"11",X"33",X"0E",X"56",X"0E",X"5F",X"11",X"68",X"16",X"70",X"1B",X"70",X"21",X"68",X"24",X"5E",
		X"00",X"01",X"80",X"22",X"44",X"1C",X"5C",X"1D",X"62",X"21",X"68",X"00",X"01",X"80",X"11",X"44",
		X"0E",X"5F",X"0E",X"56",X"11",X"4C",X"15",X"44",X"17",X"42",X"1A",X"42",X"1C",X"44",X"20",X"4A",
		X"00",X"01",X"80",X"11",X"33",X"03",X"64",X"02",X"50",X"08",X"42",X"0E",X"3A",X"16",X"36",X"1E",
		X"36",X"25",X"3A",X"2C",X"42",X"30",X"50",X"00",X"01",X"80",X"22",X"44",X"20",X"35",X"2B",X"3A",
		X"00",X"00",X"05",X"00",X"11",X"11",X"09",X"6D",X"0C",X"6E",X"16",X"7A",X"20",X"7F",X"29",X"7E",
		X"2F",X"7B",X"34",X"79",X"00",X"01",X"00",X"22",X"22",X"2E",X"7C",X"46",X"75",X"00",X"01",X"80",
		X"11",X"44",X"45",X"74",X"41",X"64",X"40",X"50",X"00",X"01",X"80",X"11",X"44",X"34",X"79",X"3A",
		X"70",X"3A",X"50",X"3C",X"48",X"41",X"3B",X"00",X"01",X"80",X"22",X"44",X"41",X"3B",X"47",X"41",
		X"00",X"01",X"00",X"22",X"22",X"1E",X"4C",X"2C",X"4C",X"00",X"01",X"80",X"11",X"44",X"1E",X"4B",
		X"2C",X"46",X"00",X"01",X"80",X"11",X"33",X"1E",X"4B",X"1E",X"46",X"41",X"3B",X"00",X"01",X"80",
		X"11",X"33",X"2C",X"46",X"2C",X"68",X"2A",X"6C",X"24",X"6F",X"1F",X"6E",X"1B",X"6A",X"18",X"64",
		X"17",X"5F",X"16",X"5D",X"15",X"5F",X"09",X"6D",X"00",X"01",X"80",X"22",X"44",X"16",X"5D",X"24",
		X"5B",X"26",X"5C",X"28",X"63",X"2C",X"64",X"00",X"00",X"6E",X"00",X"22",X"33",X"01",X"76",X"0D",
		X"6B",X"00",X"01",X"80",X"11",X"44",X"01",X"75",X"07",X"64",X"00",X"01",X"00",X"11",X"44",X"0A",
		X"58",X"0A",X"62",X"0C",X"6A",X"00",X"01",X"00",X"11",X"44",X"0D",X"6B",X"13",X"75",X"1A",X"7C",
		X"22",X"7E",X"2C",X"7E",X"33",X"7C",X"36",X"7A",X"00",X"01",X"00",X"22",X"33",X"36",X"7A",X"38",
		X"7F",X"00",X"01",X"00",X"11",X"33",X"39",X"76",X"38",X"80",X"3F",X"7E",X"44",X"7E",X"4C",X"80",
		X"00",X"01",X"80",X"11",X"44",X"35",X"79",X"39",X"76",X"00",X"01",X"80",X"11",X"33",X"4A",X"7E",
		X"47",X"72",X"46",X"54",X"00",X"01",X"80",X"11",X"33",X"1A",X"50",X"1A",X"58",X"1C",X"60",X"1F",
		X"66",X"24",X"69",X"2A",X"6A",X"30",X"68",X"35",X"64",X"38",X"5A",X"39",X"4D",X"3A",X"42",X"00",
		X"01",X"00",X"11",X"11",X"08",X"34",X"0C",X"3E",X"00",X"01",X"00",X"22",X"22",X"0C",X"3F",X"14",
		X"3E",X"00",X"01",X"00",X"11",X"11",X"4E",X"32",X"48",X"40",X"46",X"54",X"00",X"01",X"80",X"22",
		X"44",X"27",X"2C",X"2A",X"58",X"2C",X"5C",X"2E",X"58",X"2E",X"3C",X"36",X"2C",X"00",X"01",X"80",
		X"11",X"44",X"36",X"2C",X"38",X"36",X"39",X"42",X"39",X"4D",X"00",X"01",X"80",X"11",X"33",X"36",
		X"2C",X"3C",X"2D",X"4E",X"31",X"00",X"01",X"80",X"11",X"44",X"1A",X"50",X"1C",X"46",X"22",X"36",
		X"27",X"2C",X"00",X"01",X"80",X"11",X"33",X"0A",X"58",X"0C",X"4F",X"10",X"44",X"14",X"3E",X"1F",
		X"30",X"00",X"01",X"80",X"11",X"44",X"0D",X"3E",X"14",X"36",X"1F",X"30",X"00",X"01",X"80",X"11",
		X"33",X"09",X"33",X"11",X"2F",X"1A",X"2D",X"27",X"2B",X"00",X"01",X"80",X"22",X"44",X"00",X"3A",
		X"10",X"44",X"00",X"00",X"AA",X"00",X"11",X"33",X"38",X"76",X"30",X"7C",X"28",X"7F",X"19",X"7B",
		X"12",X"7A",X"00",X"01",X"00",X"22",X"44",X"12",X"7A",X"0C",X"72",X"00",X"01",X"80",X"11",X"33",
		X"13",X"79",X"14",X"71",X"14",X"66",X"00",X"01",X"80",X"11",X"44",X"14",X"66",X"12",X"5A",X"00",
		X"01",X"80",X"22",X"44",X"0C",X"55",X"13",X"5A",X"00",X"01",X"80",X"11",X"33",X"12",X"5A",X"22",
		X"6A",X"29",X"6C",X"2C",X"68",X"2C",X"63",X"00",X"01",X"80",X"11",X"44",X"2B",X"62",X"28",X"5E",
		X"14",X"52",X"10",X"4E",X"0F",X"46",X"00",X"01",X"00",X"22",X"44",X"38",X"76",X"44",X"7B",X"00",
		X"01",X"80",X"11",X"44",X"37",X"76",X"3B",X"6D",X"00",X"01",X"80",X"11",X"33",X"3A",X"6C",X"38",
		X"63",X"32",X"58",X"20",X"4C",X"1E",X"46",X"00",X"01",X"00",X"22",X"44",X"24",X"4E",X"38",X"52",
		X"00",X"01",X"80",X"11",X"44",X"37",X"51",X"30",X"48",X"25",X"42",X"20",X"42",X"1E",X"46",X"00",
		X"01",X"80",X"11",X"33",X"37",X"51",X"37",X"3F",X"2C",X"39",X"24",X"36",X"1C",X"35",X"17",X"38",
		X"10",X"40",X"10",X"4E",X"00",X"01",X"80",X"22",X"44",X"0D",X"3F",X"15",X"3A",X"00",X"00",X"DE",
		X"00",X"11",X"33",X"0F",X"7A",X"15",X"7E",X"20",X"7F",X"34",X"7D",X"3C",X"66",X"00",X"01",X"00",
		X"11",X"33",X"1E",X"60",X"28",X"4E",X"00",X"01",X"00",X"11",X"33",X"30",X"44",X"41",X"37",X"00",
		X"01",X"00",X"22",X"44",X"28",X"4E",X"3C",X"4C",X"00",X"01",X"00",X"11",X"33",X"3C",X"4C",X"40",
		X"48",X"00",X"01",X"80",X"11",X"44",X"29",X"4D",X"2D",X"4B",X"3C",X"4B",X"00",X"01",X"80",X"11",
		X"44",X"0F",X"79",X"0A",X"6F",X"00",X"01",X"80",X"11",X"33",X"0B",X"6E",X"0B",X"68",X"0E",X"60",
		X"15",X"51",X"20",X"48",X"00",X"01",X"80",X"11",X"33",X"3B",X"67",X"34",X"70",X"28",X"74",X"20",
		X"70",X"1E",X"6A",X"1E",X"60",X"00",X"01",X"80",X"22",X"44",X"3B",X"66",X"2F",X"63",X"2A",X"66",
		X"24",X"6A",X"1E",X"6A",X"00",X"01",X"80",X"22",X"44",X"01",X"5A",X"0B",X"4F",X"00",X"01",X"80",
		X"11",X"44",X"0B",X"4F",X"1A",X"4A",X"1F",X"49",X"00",X"01",X"00",X"22",X"44",X"04",X"50",X"07",
		X"51",X"00",X"01",X"80",X"22",X"44",X"04",X"41",X"09",X"3E",X"00",X"01",X"80",X"11",X"33",X"09",
		X"50",X"09",X"3E",X"1A",X"40",X"25",X"42",X"32",X"3A",X"40",X"37",X"00",X"01",X"80",X"11",X"33",
		X"30",X"44",X"3F",X"48",X"00",X"00",X"00",X"00",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",
		X"29",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",
		X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F3",X"0F",X"A3",X"0F",X"A4",X"7E",X"6E",X"C4",X"86",X"01",X"97",X"B0",X"6F",X"C8",X"34",X"39",
		X"6D",X"C8",X"34",X"27",X"08",X"6A",X"C8",X"2F",X"26",X"03",X"6C",X"C8",X"2F",X"6A",X"C8",X"33",
		X"39",X"6D",X"C8",X"34",X"27",X"02",X"86",X"8A",X"A7",X"C8",X"2F",X"39",X"25",X"03",X"86",X"CE",
		X"39",X"6D",X"C8",X"34",X"27",X"0F",X"EC",X"47",X"83",X"01",X"0B",X"2E",X"05",X"83",X"FF",X"9A",
		X"2E",X"03",X"86",X"88",X"39",X"86",X"7F",X"39",X"A7",X"C8",X"33",X"6D",X"C8",X"34",X"27",X"0C",
		X"67",X"C8",X"11",X"66",X"C8",X"12",X"67",X"C8",X"11",X"66",X"C8",X"12",X"39",X"6D",X"C8",X"34",
		X"27",X"02",X"CB",X"02",X"E7",X"C8",X"2E",X"39",X"FC",X"B3",X"00",X"C3",X"FF",X"FF",X"2E",X"12",
		X"FC",X"B3",X"02",X"10",X"83",X"05",X"00",X"22",X"06",X"C3",X"00",X"01",X"FD",X"B3",X"02",X"CC",
		X"00",X"01",X"FD",X"B3",X"00",X"86",X"01",X"7E",X"E0",X"12",X"ED",X"A8",X"1C",X"CC",X"07",X"08",
		X"FD",X"B3",X"00",X"FC",X"B1",X"B0",X"FD",X"B3",X"02",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A6",X"0B",X"81",X"A9",X"25",X"03",X"0C",X"8A",X"39",X"81",X"51",X"25",X"03",X"0C",X"89",X"39",
		X"0C",X"88",X"39",X"E6",X"C8",X"13",X"86",X"60",X"3D",X"1F",X"89",X"4F",X"83",X"00",X"60",X"E3",
		X"C8",X"11",X"ED",X"C8",X"11",X"96",X"32",X"48",X"AB",X"C8",X"14",X"2D",X"08",X"81",X"08",X"2E",
		X"0B",X"A7",X"C8",X"14",X"39",X"81",X"F8",X"2D",X"03",X"A7",X"C8",X"14",X"39",X"AD",X"D8",X"24",
		X"4D",X"27",X"07",X"6F",X"4F",X"4D",X"2A",X"02",X"63",X"4F",X"6C",X"C8",X"13",X"26",X"03",X"6A",
		X"C8",X"13",X"BD",X"8E",X"8E",X"DC",X"32",X"39",X"DB",X"48",X"1D",X"E3",X"C8",X"11",X"ED",X"C8",
		X"11",X"E3",X"4B",X"AB",X"C8",X"23",X"6F",X"C8",X"23",X"81",X"20",X"22",X"14",X"6C",X"C8",X"23",
		X"EC",X"C8",X"11",X"2A",X"07",X"43",X"50",X"82",X"FF",X"ED",X"C8",X"11",X"CC",X"20",X"00",X"20",
		X"00",X"81",X"E6",X"24",X"14",X"ED",X"4B",X"A6",X"C8",X"14",X"EC",X"86",X"EB",X"C8",X"16",X"E7",
		X"C8",X"16",X"89",X"00",X"1F",X"89",X"7E",X"DD",X"D2",X"8E",X"EF",X"CB",X"A6",X"42",X"81",X"89",
		X"27",X"03",X"8E",X"EF",X"9A",X"BD",X"E0",X"2D",X"BD",X"8E",X"4D",X"BD",X"D8",X"EB",X"86",X"03",
		X"BD",X"E0",X"37",X"BD",X"8E",X"8E",X"BD",X"D8",X"EB",X"A6",X"42",X"2A",X"1C",X"E6",X"07",X"C1",
		X"03",X"27",X"16",X"84",X"7F",X"A7",X"42",X"CC",X"00",X"00",X"ED",X"C8",X"1E",X"ED",X"C8",X"1A",
		X"8E",X"00",X"00",X"10",X"AE",X"4D",X"AD",X"B8",X"10",X"6C",X"4B",X"A6",X"4B",X"81",X"F4",X"25",
		X"C7",X"86",X"1E",X"BD",X"E0",X"37",X"AE",X"4D",X"6E",X"98",X"0E",X"8D",X"07",X"EC",X"C8",X"1E",
		X"27",X"1B",X"30",X"16",X"A6",X"07",X"88",X"04",X"AB",X"05",X"81",X"E0",X"25",X"0F",X"A6",X"05",
		X"81",X"E0",X"25",X"0A",X"86",X"F0",X"A7",X"04",X"CC",X"04",X"04",X"ED",X"06",X"39",X"40",X"8B",
		X"E0",X"88",X"04",X"A7",X"07",X"39",X"6F",X"C8",X"22",X"6F",X"C8",X"23",X"6F",X"C8",X"14",X"1D",
		X"F3",X"B3",X"02",X"E3",X"C8",X"11",X"ED",X"C8",X"11",X"10",X"83",X"FE",X"80",X"2D",X"43",X"E3",
		X"4B",X"ED",X"4B",X"81",X"E6",X"25",X"1D",X"AE",X"C4",X"A6",X"02",X"81",X"16",X"26",X"05",X"CC",
		X"6A",X"8D",X"ED",X"05",X"9E",X"2C",X"CC",X"6A",X"EE",X"ED",X"05",X"CC",X"D8",X"58",X"ED",X"C8",
		X"30",X"7E",X"D8",X"99",X"EC",X"47",X"10",X"83",X"00",X"08",X"2E",X"03",X"CC",X"00",X"08",X"10",
		X"83",X"01",X"16",X"2D",X"03",X"CC",X"01",X"16",X"ED",X"47",X"1F",X"32",X"BD",X"6A",X"A1",X"26",
		X"01",X"39",X"A6",X"42",X"2A",X"07",X"86",X"50",X"AE",X"4D",X"BD",X"E6",X"B1",X"AE",X"C4",X"A6",
		X"02",X"81",X"16",X"26",X"05",X"CC",X"6A",X"8D",X"ED",X"05",X"9E",X"2C",X"CC",X"6A",X"E3",X"ED",
		X"05",X"86",X"01",X"A7",X"04",X"CC",X"D8",X"58",X"ED",X"C8",X"30",X"EC",X"C8",X"11",X"E3",X"4B",
		X"ED",X"4B",X"39",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"B0",X"02",X"A4",X"A9",X"EA",X"97",
		X"26",X"10",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"37",X"27",X"03",X"BD",X"DA",X"3E",X"86",
		X"01",X"39",X"81",X"08",X"25",X"0C",X"27",X"22",X"81",X"20",X"25",X"24",X"85",X"20",X"26",X"26",
		X"20",X"2A",X"81",X"02",X"27",X"08",X"22",X"0C",X"C6",X"44",X"E7",X"4B",X"4F",X"39",X"C6",X"50",
		X"E7",X"4B",X"4F",X"39",X"C6",X"80",X"E7",X"4B",X"4F",X"39",X"C6",X"89",X"E7",X"4B",X"4F",X"39",
		X"C6",X"A2",X"E7",X"4B",X"4F",X"39",X"C6",X"D2",X"E7",X"4B",X"4F",X"39",X"96",X"A0",X"26",X"3B",
		X"96",X"96",X"26",X"37",X"A6",X"42",X"81",X"89",X"27",X"04",X"81",X"8F",X"26",X"2D",X"0C",X"96",
		X"86",X"15",X"E6",X"43",X"8E",X"69",X"DD",X"DE",X"2C",X"BD",X"E0",X"30",X"DE",X"2E",X"EF",X"A8",
		X"24",X"6F",X"A8",X"10",X"CC",X"00",X"D6",X"ED",X"2A",X"EC",X"47",X"C3",X"FF",X"FE",X"ED",X"27",
		X"CC",X"00",X"00",X"ED",X"A8",X"1C",X"86",X"01",X"A7",X"A8",X"2D",X"E6",X"4B",X"39",X"1F",X"89",
		X"9A",X"4B",X"97",X"4B",X"5D",X"10",X"2B",X"00",X"D6",X"C1",X"08",X"25",X"11",X"10",X"27",X"00",
		X"8C",X"C4",X"70",X"C1",X"20",X"10",X"22",X"00",X"E3",X"25",X"18",X"7E",X"DA",X"C5",X"C1",X"02",
		X"27",X"56",X"10",X"22",X"00",X"C6",X"10",X"AE",X"9F",X"00",X"00",X"CC",X"FF",X"E0",X"8E",X"00",
		X"45",X"20",X"0B",X"10",X"AE",X"9F",X"00",X"08",X"CC",X"FF",X"E0",X"8E",X"00",X"8A",X"34",X"20",
		X"BD",X"DB",X"F9",X"24",X"30",X"10",X"AC",X"E1",X"26",X"14",X"A6",X"04",X"2B",X"0D",X"A6",X"08",
		X"2B",X"09",X"A6",X"0C",X"2B",X"05",X"A6",X"88",X"10",X"2A",X"03",X"7E",X"DB",X"BF",X"A6",X"24",
		X"2B",X"7A",X"EC",X"A4",X"E3",X"22",X"A3",X"84",X"A3",X"02",X"D3",X"34",X"D3",X"34",X"10",X"2B",
		X"00",X"C4",X"7E",X"DB",X"85",X"32",X"62",X"39",X"10",X"AE",X"9F",X"00",X"02",X"CC",X"00",X"FC",
		X"8E",X"00",X"45",X"20",X"23",X"10",X"AE",X"9F",X"00",X"0A",X"CC",X"00",X"CA",X"8E",X"00",X"81",
		X"BD",X"DB",X"F9",X"24",X"E2",X"E6",X"4B",X"C1",X"93",X"22",X"2D",X"20",X"17",X"10",X"AE",X"9F",
		X"00",X"0A",X"CC",X"00",X"CA",X"8E",X"00",X"81",X"34",X"20",X"BD",X"DB",X"F9",X"24",X"C6",X"10",
		X"AC",X"E1",X"26",X"14",X"A6",X"04",X"2B",X"0D",X"A6",X"08",X"2B",X"09",X"A6",X"0C",X"2B",X"05",
		X"A6",X"88",X"10",X"2A",X"03",X"7E",X"DB",X"BF",X"A6",X"24",X"2B",X"10",X"EC",X"A4",X"E3",X"22",
		X"A3",X"84",X"A3",X"02",X"D3",X"34",X"D3",X"34",X"10",X"2A",X"00",X"79",X"7E",X"DB",X"85",X"10",
		X"AE",X"9F",X"00",X"0E",X"CC",X"00",X"36",X"8E",X"00",X"D3",X"20",X"1B",X"10",X"AE",X"9F",X"00",
		X"04",X"CC",X"00",X"56",X"8E",X"00",X"51",X"20",X"0E",X"32",X"62",X"39",X"10",X"AE",X"9F",X"00",
		X"0C",X"CC",X"00",X"6A",X"8E",X"00",X"A3",X"34",X"20",X"BD",X"DB",X"F9",X"24",X"EB",X"10",X"AC",
		X"E1",X"26",X"11",X"A6",X"04",X"2B",X"68",X"A6",X"08",X"2B",X"64",X"A6",X"0C",X"2B",X"60",X"A6",
		X"88",X"10",X"2B",X"5B",X"A6",X"24",X"2B",X"1D",X"EC",X"A4",X"E3",X"22",X"A3",X"84",X"A3",X"02",
		X"D3",X"34",X"D3",X"34",X"2A",X"1F",X"A6",X"C8",X"14",X"2C",X"06",X"40",X"80",X"02",X"A7",X"C8",
		X"14",X"8B",X"06",X"20",X"1D",X"EC",X"C8",X"11",X"2A",X"09",X"43",X"50",X"82",X"FF",X"47",X"56",
		X"ED",X"C8",X"11",X"20",X"1F",X"A6",X"C8",X"14",X"2F",X"06",X"40",X"8B",X"02",X"A7",X"C8",X"14",
		X"80",X"06",X"A7",X"C8",X"22",X"EC",X"C8",X"11",X"10",X"83",X"FF",X"C0",X"2A",X"03",X"CC",X"FF",
		X"C0",X"ED",X"C8",X"11",X"86",X"02",X"A7",X"C8",X"23",X"8E",X"EF",X"8F",X"7E",X"E0",X"2D",X"EC",
		X"C8",X"11",X"2B",X"07",X"43",X"53",X"47",X"56",X"ED",X"C8",X"11",X"86",X"FE",X"A7",X"C8",X"23",
		X"A6",X"C8",X"14",X"26",X"13",X"EC",X"A4",X"E3",X"22",X"A3",X"84",X"A3",X"02",X"D3",X"34",X"D3",
		X"34",X"2A",X"0B",X"86",X"02",X"A7",X"C8",X"14",X"8E",X"EF",X"8F",X"7E",X"E0",X"2D",X"86",X"FE",
		X"A7",X"C8",X"14",X"8E",X"EF",X"8F",X"7E",X"E0",X"2D",X"A3",X"47",X"DD",X"34",X"1F",X"10",X"AE",
		X"D8",X"1C",X"E0",X"C8",X"28",X"2B",X"07",X"58",X"58",X"49",X"30",X"8B",X"20",X"13",X"50",X"58",
		X"58",X"49",X"31",X"AB",X"20",X"0B",X"A6",X"84",X"AA",X"A4",X"46",X"25",X"64",X"30",X"04",X"31",
		X"24",X"EC",X"02",X"2D",X"F3",X"A3",X"A4",X"29",X"ED",X"93",X"34",X"2D",X"1E",X"EC",X"84",X"A3",
		X"22",X"93",X"34",X"2E",X"62",X"43",X"39",X"30",X"88",X"10",X"31",X"A8",X"10",X"EC",X"02",X"2D",
		X"40",X"A3",X"A4",X"29",X"3C",X"93",X"34",X"2D",X"02",X"43",X"39",X"EC",X"06",X"2D",X"32",X"A3",
		X"24",X"29",X"2E",X"93",X"34",X"2D",X"06",X"30",X"04",X"31",X"24",X"43",X"39",X"EC",X"0A",X"2D",
		X"20",X"A3",X"28",X"29",X"1C",X"93",X"34",X"2D",X"06",X"30",X"08",X"31",X"28",X"43",X"39",X"EC",
		X"0E",X"2D",X"0E",X"A3",X"2C",X"29",X"0A",X"93",X"34",X"2D",X"BC",X"30",X"0C",X"31",X"2C",X"43",
		X"39",X"4F",X"39",X"30",X"88",X"10",X"31",X"A8",X"10",X"EC",X"84",X"2D",X"F4",X"A3",X"22",X"29",
		X"F0",X"93",X"34",X"2E",X"02",X"43",X"39",X"EC",X"04",X"2D",X"E6",X"A3",X"26",X"29",X"E2",X"93",
		X"34",X"2E",X"06",X"30",X"04",X"31",X"24",X"43",X"39",X"EC",X"08",X"2D",X"D4",X"A3",X"2A",X"29",
		X"D0",X"93",X"34",X"2E",X"06",X"30",X"08",X"31",X"28",X"43",X"39",X"EC",X"0C",X"2D",X"C2",X"A3",
		X"2E",X"29",X"BE",X"93",X"34",X"2E",X"BC",X"30",X"0C",X"31",X"2C",X"43",X"39",X"FE",X"00",X"FF",
		X"00",X"FF",X"80",X"FF",X"C0",X"00",X"00",X"00",X"40",X"00",X"80",X"01",X"00",X"02",X"00",X"08",
		X"DD",X"3A",X"07",X"07",X"07",X"00",X"00",X"DD",X"3C",X"F9",X"00",X"07",X"00",X"08",X"DD",X"4D",
		X"1C",X"00",X"07",X"02",X"04",X"DD",X"4D",X"F9",X"00",X"07",X"04",X"02",X"DD",X"4D",X"15",X"00",
		X"07",X"06",X"01",X"DD",X"4D",X"15",X"00",X"00",X"08",X"02",X"DD",X"8E",X"DD",X"DD",X"E4",X"02",
		X"02",X"DD",X"9C",X"15",X"15",X"E4",X"04",X"02",X"DD",X"9C",X"07",X"07",X"E4",X"06",X"02",X"DD",
		X"9C",X"07",X"07",X"D6",X"04",X"02",X"DD",X"9C",X"07",X"07",X"CF",X"04",X"04",X"DD",X"9C",X"07",
		X"07",X"C1",X"02",X"04",X"DD",X"9C",X"B3",X"B3",X"BA",X"02",X"63",X"4F",X"CC",X"0C",X"00",X"6F",
		X"C8",X"10",X"39",X"18",X"00",X"3C",X"03",X"30",X"02",X"24",X"01",X"18",X"02",X"E6",X"C8",X"10",
		X"2F",X"2D",X"5A",X"2E",X"02",X"C6",X"04",X"E7",X"C8",X"10",X"C1",X"01",X"26",X"19",X"AE",X"4D",
		X"6C",X"C8",X"35",X"A6",X"C8",X"35",X"46",X"24",X"05",X"AE",X"88",X"24",X"20",X"03",X"AE",X"88",
		X"26",X"BD",X"E0",X"2D",X"E6",X"C8",X"10",X"58",X"8E",X"DD",X"43",X"3A",X"EC",X"84",X"39",X"C6",
		X"04",X"E7",X"C8",X"10",X"FC",X"DD",X"43",X"39",X"00",X"00",X"02",X"04",X"01",X"01",X"8E",X"DD",
		X"89",X"E6",X"C8",X"10",X"E6",X"85",X"86",X"0C",X"6F",X"C8",X"10",X"39",X"A6",X"C8",X"10",X"2B",
		X"08",X"AE",X"4D",X"AE",X"88",X"20",X"BD",X"E0",X"2D",X"86",X"FF",X"A7",X"C8",X"10",X"CC",X"00",
		X"02",X"39",X"B6",X"C8",X"07",X"8A",X"08",X"20",X"05",X"B6",X"C8",X"07",X"84",X"F7",X"B7",X"C8",
		X"07",X"B6",X"C8",X"04",X"5F",X"85",X"04",X"27",X"01",X"5C",X"84",X"03",X"47",X"82",X"00",X"DD",
		X"32",X"39",X"A6",X"C8",X"22",X"27",X"22",X"2D",X"0D",X"81",X"03",X"2F",X"16",X"CB",X"03",X"80",
		X"03",X"A7",X"C8",X"22",X"20",X"13",X"81",X"FD",X"2C",X"09",X"CB",X"FD",X"80",X"FD",X"A7",X"C8",
		X"22",X"20",X"06",X"EB",X"C8",X"22",X"6F",X"C8",X"22",X"1D",X"E3",X"47",X"10",X"83",X"01",X"24",
		X"2F",X"03",X"C3",X"FE",X"D1",X"10",X"83",X"FF",X"F6",X"2C",X"03",X"C3",X"01",X"2F",X"ED",X"47",
		X"39",X"00",X"0B",X"00",X"06",X"00",X"04",X"00",X"01",X"FA",X"86",X"44",X"33",X"21",X"FF",X"00",
		X"04",X"00",X"06",X"00",X"08",X"00",X"2D",X"FA",X"86",X"43",X"33",X"21",X"02",X"00",X"10",X"00",
		X"08",X"00",X"04",X"00",X"01",X"FA",X"86",X"44",X"33",X"21",X"FF",X"00",X"60",X"00",X"40",X"00",
		X"20",X"00",X"10",X"FF",X"CA",X"86",X"43",X"21",X"FE",X"00",X"5E",X"00",X"38",X"00",X"22",X"00",
		X"08",X"CA",X"53",X"A5",X"25",X"21",X"FC",X"00",X"0E",X"00",X"0E",X"00",X"0C",X"00",X"0B",X"FF",
		X"FF",X"FF",X"F8",X"42",X"FF",X"F0",X"00",X"F2",X"00",X"F8",X"00",X"FF",X"00",X"42",X"11",X"42",
		X"14",X"21",X"20",X"00",X"80",X"01",X"00",X"02",X"00",X"03",X"00",X"42",X"11",X"F8",X"13",X"21",
		X"20",X"FF",X"F1",X"FF",X"F2",X"FF",X"F4",X"FF",X"F5",X"FF",X"FF",X"FF",X"F8",X"42",X"01",X"10",
		X"00",X"0E",X"00",X"08",X"00",X"01",X"00",X"42",X"11",X"42",X"14",X"21",X"E0",X"00",X"03",X"00",
		X"02",X"00",X"01",X"00",X"01",X"FA",X"86",X"44",X"33",X"21",X"FF",X"00",X"0A",X"00",X"08",X"00",
		X"06",X"00",X"02",X"FA",X"86",X"44",X"33",X"21",X"FF",X"00",X"20",X"00",X"15",X"00",X"10",X"00",
		X"02",X"77",X"66",X"44",X"33",X"21",X"FF",X"00",X"0F",X"00",X"0E",X"00",X"0C",X"00",X"0B",X"FF",
		X"FF",X"FF",X"FA",X"22",X"FF",X"F0",X"00",X"F2",X"00",X"F8",X"00",X"FF",X"00",X"FF",X"FF",X"FF",
		X"84",X"22",X"20",X"01",X"00",X"02",X"00",X"03",X"00",X"03",X"80",X"FF",X"FF",X"FF",X"84",X"84",
		X"20",X"FF",X"F1",X"FF",X"F2",X"FF",X"F4",X"FF",X"F5",X"FF",X"FF",X"FF",X"F8",X"22",X"01",X"10",
		X"00",X"0E",X"00",X"08",X"00",X"01",X"00",X"FF",X"F8",X"FF",X"84",X"22",X"E0",X"00",X"03",X"00",
		X"02",X"00",X"01",X"00",X"01",X"FF",X"F8",X"FF",X"83",X"22",X"FF",X"00",X"0A",X"00",X"08",X"00",
		X"06",X"00",X"02",X"FF",X"F8",X"FF",X"83",X"22",X"FF",X"FF",X"80",X"FF",X"00",X"FE",X"00",X"FE",
		X"00",X"FF",X"FF",X"FF",X"84",X"84",X"20",X"00",X"20",X"00",X"15",X"00",X"10",X"00",X"02",X"FF",
		X"F8",X"84",X"33",X"22",X"FF",X"00",X"14",X"00",X"10",X"00",X"0E",X"00",X"0C",X"FF",X"FF",X"FF",
		X"FA",X"82",X"FF",X"FF",X"EC",X"FF",X"E0",X"FF",X"F2",X"FF",X"F4",X"FF",X"FF",X"FF",X"FA",X"82",
		X"01",X"FF",X"F0",X"FE",X"00",X"FD",X"00",X"FC",X"00",X"FF",X"FF",X"FF",X"FA",X"84",X"20",X"00",
		X"14",X"00",X"0A",X"00",X"08",X"00",X"02",X"FF",X"FF",X"FF",X"FA",X"82",X"FF",X"00",X"20",X"00",
		X"15",X"00",X"10",X"00",X"02",X"FF",X"FF",X"FF",X"FA",X"82",X"FF",X"00",X"0A",X"00",X"08",X"00",
		X"06",X"00",X"02",X"FF",X"FF",X"FF",X"FA",X"61",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"F0",X"10",X"CE",X"BF",X"00",X"7E",X"E0",X"3D",X"7E",X"E2",X"82",X"7E",X"E2",X"4D",X"7E",
		X"E2",X"0F",X"7E",X"E1",X"59",X"7E",X"E4",X"B2",X"7E",X"E4",X"C0",X"7E",X"E2",X"A1",X"7E",X"E2",
		X"B8",X"7E",X"E2",X"CF",X"7E",X"E2",X"F9",X"7E",X"E3",X"22",X"7E",X"E3",X"58",X"7E",X"E4",X"CD",
		X"7E",X"E2",X"84",X"E5",X"FA",X"E4",X"E6",X"7E",X"E1",X"57",X"7E",X"E6",X"0A",X"86",X"A0",X"1F",
		X"8B",X"8E",X"00",X"00",X"5F",X"86",X"39",X"B7",X"CB",X"FF",X"4F",X"ED",X"81",X"ED",X"81",X"8C",
		X"BF",X"80",X"25",X"F1",X"5C",X"F7",X"BF",X"FF",X"F7",X"C9",X"00",X"B7",X"C8",X"05",X"B7",X"C8",
		X"07",X"B7",X"C8",X"04",X"B7",X"C8",X"06",X"C6",X"34",X"F7",X"C8",X"05",X"F7",X"C8",X"07",X"B7",
		X"C8",X"0D",X"B7",X"C8",X"0F",X"B7",X"C8",X"0C",X"43",X"B7",X"C8",X"0E",X"C6",X"34",X"F7",X"C8",
		X"0D",X"C6",X"35",X"F7",X"C8",X"0F",X"C6",X"3F",X"F7",X"C8",X"0E",X"86",X"3C",X"97",X"8B",X"97",
		X"B4",X"CE",X"A1",X"00",X"DF",X"08",X"86",X"14",X"30",X"C8",X"38",X"AF",X"C4",X"33",X"88",X"38",
		X"EF",X"84",X"4A",X"26",X"F3",X"8E",X"A9",X"C0",X"9F",X"25",X"8E",X"AC",X"21",X"9F",X"68",X"8E",
		X"E5",X"FA",X"BD",X"E4",X"B2",X"CC",X"0E",X"10",X"DD",X"99",X"8E",X"CD",X"00",X"BD",X"3B",X"34",
		X"1F",X"98",X"81",X"20",X"22",X"06",X"84",X"0F",X"81",X"09",X"23",X"07",X"5F",X"8E",X"CD",X"00",
		X"BD",X"3B",X"3D",X"D7",X"F2",X"CE",X"A0",X"0A",X"8E",X"5E",X"D0",X"4F",X"5F",X"BD",X"E2",X"84",
		X"1C",X"EF",X"8E",X"A9",X"C0",X"96",X"27",X"2A",X"03",X"8E",X"AC",X"21",X"9F",X"28",X"03",X"27",
		X"6D",X"84",X"26",X"FC",X"30",X"09",X"9F",X"2A",X"96",X"61",X"27",X"1D",X"0A",X"61",X"26",X"19",
		X"9E",X"63",X"27",X"15",X"EC",X"81",X"2B",X"03",X"8E",X"00",X"00",X"9F",X"63",X"D7",X"61",X"C6",
		X"FF",X"F7",X"C8",X"0E",X"84",X"3F",X"B7",X"C8",X"0E",X"4F",X"5F",X"8E",X"A0",X"00",X"AF",X"04",
		X"ED",X"81",X"AF",X"04",X"ED",X"84",X"30",X"88",X"3E",X"AF",X"04",X"ED",X"81",X"AF",X"04",X"ED",
		X"84",X"30",X"88",X"3E",X"AF",X"04",X"ED",X"81",X"AF",X"04",X"ED",X"84",X"30",X"88",X"3E",X"AF",
		X"04",X"ED",X"81",X"AF",X"04",X"ED",X"84",X"CE",X"A0",X"0A",X"10",X"CE",X"BF",X"00",X"0F",X"65",
		X"20",X"11",X"DF",X"2E",X"6E",X"D8",X"05",X"AE",X"E1",X"DE",X"2E",X"AF",X"45",X"A7",X"44",X"96",
		X"65",X"26",X"1D",X"DF",X"2C",X"EE",X"C4",X"27",X"0A",X"A6",X"43",X"26",X"F6",X"6A",X"44",X"27",
		X"E1",X"20",X"F0",X"10",X"CE",X"BF",X"00",X"03",X"65",X"DE",X"66",X"26",X"03",X"CE",X"A0",X"0A",
		X"DF",X"2C",X"A6",X"9F",X"A0",X"68",X"27",X"0E",X"EE",X"C4",X"27",X"0B",X"A6",X"43",X"27",X"F0",
		X"6A",X"44",X"27",X"BE",X"20",X"EA",X"12",X"DF",X"66",X"DE",X"28",X"DF",X"68",X"33",X"41",X"8E",
		X"00",X"00",X"DC",X"00",X"ED",X"C4",X"AF",X"9F",X"A0",X"04",X"DC",X"40",X"26",X"06",X"DC",X"02",
		X"ED",X"42",X"20",X"08",X"ED",X"42",X"DC",X"02",X"ED",X"9F",X"A0",X"44",X"AF",X"9F",X"A0",X"06",
		X"DC",X"80",X"26",X"06",X"DC",X"42",X"ED",X"44",X"20",X"08",X"ED",X"44",X"DC",X"42",X"ED",X"9F",
		X"A0",X"84",X"AF",X"9F",X"A0",X"46",X"DC",X"C0",X"26",X"14",X"DC",X"82",X"26",X"06",X"DC",X"C2",
		X"ED",X"46",X"20",X"22",X"ED",X"46",X"DC",X"C2",X"ED",X"9F",X"A0",X"86",X"20",X"18",X"ED",X"46",
		X"DC",X"82",X"26",X"08",X"DC",X"C2",X"ED",X"9F",X"A0",X"C4",X"20",X"0A",X"ED",X"9F",X"A0",X"C4",
		X"DC",X"C2",X"ED",X"9F",X"A0",X"86",X"AF",X"9F",X"A0",X"C6",X"6C",X"5F",X"7E",X"E0",X"E2",X"10",
		X"CE",X"BF",X"00",X"DE",X"2E",X"EC",X"C4",X"ED",X"9F",X"A0",X"2C",X"DC",X"08",X"ED",X"C4",X"DF",
		X"08",X"DE",X"2C",X"7E",X"E1",X"5F",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",X"29",X"31",
		X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"34",X"46",X"8E",
		X"A0",X"0A",X"DE",X"0A",X"27",X"15",X"E6",X"61",X"E4",X"42",X"E1",X"E4",X"26",X"07",X"11",X"93",
		X"2E",X"26",X"0A",X"9F",X"2C",X"1F",X"31",X"EE",X"C4",X"26",X"EB",X"35",X"C6",X"11",X"93",X"66",
		X"26",X"02",X"9F",X"66",X"EC",X"C4",X"ED",X"84",X"DC",X"08",X"ED",X"C4",X"DF",X"08",X"1F",X"13",
		X"20",X"E5",X"DE",X"2E",X"34",X"06",X"10",X"9E",X"08",X"EC",X"A4",X"DD",X"08",X"EC",X"C4",X"ED",
		X"A4",X"10",X"AF",X"C4",X"86",X"01",X"A7",X"24",X"AF",X"25",X"35",X"06",X"A7",X"22",X"E7",X"23",
		X"39",X"C4",X"C0",X"8E",X"A0",X"04",X"3A",X"DC",X"2A",X"ED",X"94",X"C3",X"00",X"08",X"ED",X"84",
		X"C3",X"00",X"02",X"9E",X"2A",X"DD",X"2A",X"39",X"C4",X"C0",X"8E",X"A0",X"06",X"3A",X"DC",X"2A",
		X"ED",X"94",X"C3",X"00",X"08",X"ED",X"84",X"C3",X"00",X"02",X"9E",X"2A",X"DD",X"2A",X"39",X"E6",
		X"4B",X"D7",X"31",X"C4",X"C0",X"8E",X"A0",X"04",X"3A",X"DC",X"2A",X"ED",X"94",X"C3",X"00",X"08",
		X"ED",X"84",X"C3",X"00",X"02",X"9E",X"2A",X"DD",X"2A",X"EC",X"47",X"46",X"56",X"D7",X"30",X"86",
		X"1A",X"24",X"02",X"8A",X"20",X"5F",X"ED",X"84",X"39",X"E6",X"4B",X"D7",X"31",X"C4",X"C0",X"8E",
		X"A0",X"06",X"3A",X"DC",X"2A",X"ED",X"94",X"C3",X"00",X"08",X"ED",X"84",X"C3",X"00",X"02",X"9E",
		X"2A",X"DD",X"2A",X"EC",X"47",X"46",X"56",X"D7",X"30",X"86",X"0A",X"24",X"02",X"8A",X"20",X"A7",
		X"84",X"39",X"E6",X"4B",X"D7",X"31",X"C4",X"C0",X"8E",X"A0",X"04",X"3A",X"DC",X"2A",X"ED",X"94",
		X"C3",X"00",X"08",X"ED",X"84",X"C3",X"00",X"02",X"ED",X"94",X"C3",X"00",X"08",X"ED",X"84",X"C3",
		X"00",X"02",X"9E",X"2A",X"DD",X"2A",X"EC",X"47",X"46",X"56",X"D7",X"30",X"86",X"1A",X"24",X"02",
		X"8A",X"20",X"5F",X"ED",X"84",X"ED",X"0A",X"39",X"E6",X"4B",X"D7",X"31",X"C4",X"C0",X"8E",X"A0",
		X"06",X"3A",X"DC",X"2A",X"ED",X"94",X"C3",X"00",X"08",X"ED",X"84",X"C3",X"00",X"02",X"ED",X"94",
		X"C3",X"00",X"08",X"ED",X"84",X"C3",X"00",X"02",X"9E",X"2A",X"DD",X"2A",X"EC",X"47",X"46",X"56",
		X"D7",X"30",X"86",X"0A",X"24",X"02",X"8A",X"20",X"A7",X"84",X"A7",X"0A",X"39",X"10",X"DF",X"1F",
		X"86",X"39",X"B7",X"CB",X"FF",X"0C",X"0D",X"0A",X"0E",X"B6",X"BF",X"FF",X"8A",X"01",X"B7",X"C9",
		X"00",X"F6",X"C8",X"0E",X"F6",X"CB",X"00",X"C4",X"C0",X"10",X"26",X"00",X"A4",X"CE",X"A0",X"0F",
		X"37",X"76",X"CE",X"C0",X"08",X"36",X"76",X"CE",X"A0",X"17",X"37",X"76",X"CE",X"C0",X"10",X"36",
		X"76",X"10",X"DE",X"1F",X"96",X"90",X"2A",X"11",X"DC",X"99",X"83",X"00",X"01",X"2E",X"08",X"C6",
		X"06",X"BD",X"3B",X"2B",X"CC",X"0E",X"10",X"DD",X"99",X"96",X"8D",X"27",X"02",X"0A",X"8D",X"DC",
		X"BA",X"DD",X"BB",X"DC",X"B8",X"DD",X"B9",X"DC",X"B6",X"DD",X"B7",X"DC",X"B4",X"DD",X"B5",X"B6",
		X"C8",X"0C",X"97",X"B4",X"85",X"40",X"27",X"04",X"C6",X"78",X"D7",X"8D",X"D6",X"B4",X"DA",X"B5",
		X"DA",X"B6",X"DA",X"B7",X"DA",X"B8",X"DA",X"B9",X"DA",X"BA",X"DA",X"BB",X"DA",X"BC",X"D4",X"8B",
		X"D7",X"8C",X"94",X"B5",X"9A",X"8C",X"D6",X"8B",X"97",X"8B",X"53",X"D4",X"8B",X"C4",X"3E",X"27",
		X"30",X"54",X"34",X"04",X"64",X"E4",X"24",X"03",X"BD",X"F0",X"03",X"96",X"8D",X"26",X"07",X"64",
		X"E4",X"24",X"03",X"BD",X"3B",X"4F",X"64",X"E4",X"24",X"03",X"BD",X"3B",X"25",X"96",X"8D",X"26",
		X"0E",X"64",X"E4",X"24",X"03",X"BD",X"3B",X"49",X"64",X"E4",X"24",X"03",X"BD",X"3B",X"4C",X"35",
		X"04",X"9E",X"25",X"96",X"23",X"6D",X"84",X"27",X"4E",X"2B",X"05",X"63",X"80",X"9F",X"21",X"4F",
		X"B7",X"A0",X"23",X"B8",X"CB",X"00",X"84",X"C0",X"27",X"3D",X"BE",X"A0",X"21",X"EE",X"81",X"BF",
		X"A0",X"21",X"30",X"C4",X"27",X"17",X"7A",X"C8",X"0F",X"B6",X"C8",X"0E",X"10",X"CE",X"CA",X"08",
		X"37",X"3F",X"34",X"3F",X"EE",X"C4",X"26",X"F4",X"1A",X"FF",X"7C",X"C8",X"0F",X"B6",X"A0",X"23",
		X"8B",X"40",X"26",X"CC",X"BE",X"A0",X"25",X"6F",X"84",X"8E",X"A9",X"C0",X"73",X"A0",X"24",X"2A",
		X"03",X"8E",X"AC",X"21",X"BF",X"A0",X"25",X"10",X"FE",X"A0",X"1F",X"B6",X"BF",X"FF",X"B7",X"C9",
		X"00",X"3B",X"10",X"8E",X"A0",X"0F",X"C6",X"10",X"A6",X"80",X"A7",X"A0",X"5A",X"26",X"F9",X"39",
		X"96",X"0E",X"44",X"44",X"44",X"98",X"0E",X"44",X"06",X"0D",X"06",X"0E",X"39",X"A6",X"80",X"2B",
		X"04",X"D6",X"90",X"2A",X"10",X"D6",X"61",X"27",X"04",X"91",X"62",X"25",X"08",X"97",X"62",X"86",
		X"01",X"97",X"61",X"9F",X"63",X"39",X"8E",X"00",X"FF",X"9F",X"9C",X"CC",X"E5",X"E9",X"DD",X"B1",
		X"86",X"14",X"BD",X"E0",X"37",X"9E",X"9C",X"C6",X"44",X"B6",X"BF",X"FF",X"84",X"FE",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"E7",X"84",X"30",X"89",X"01",X"00",X"8C",X"96",X"00",X"22",X"28",X"A6",
		X"84",X"84",X"EE",X"27",X"EF",X"85",X"F0",X"26",X"04",X"8A",X"40",X"A7",X"84",X"DC",X"9C",X"86",
		X"96",X"1F",X"01",X"C6",X"44",X"E7",X"84",X"30",X"89",X"FF",X"00",X"A6",X"84",X"27",X"F6",X"85",
		X"0F",X"26",X"04",X"8A",X"04",X"A7",X"84",X"B6",X"BF",X"FF",X"8A",X"01",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"0A",X"9D",X"D6",X"9D",X"D1",X"9B",X"2C",X"A6",X"86",X"01",X"BD",X"E0",X"37",X"BD",
		X"E0",X"18",X"A7",X"4F",X"84",X"0F",X"9E",X"B1",X"A6",X"86",X"24",X"4A",X"E6",X"4E",X"C4",X"0F",
		X"CA",X"02",X"DB",X"9D",X"5C",X"1F",X"01",X"AF",X"C8",X"14",X"86",X"40",X"A7",X"84",X"8E",X"E6",
		X"92",X"BD",X"E4",X"CD",X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"14",X"86",X"04",X"A7",X"84",
		X"A7",X"89",X"01",X"00",X"86",X"40",X"A7",X"1F",X"A7",X"01",X"86",X"08",X"BD",X"E0",X"37",X"AE",
		X"C8",X"14",X"86",X"44",X"A7",X"1F",X"A7",X"84",X"A7",X"01",X"A7",X"89",X"01",X"00",X"86",X"05",
		X"AB",X"4E",X"A7",X"4E",X"20",X"9E",X"D6",X"9D",X"5C",X"ED",X"C8",X"14",X"1F",X"01",X"6F",X"01",
		X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"14",X"C6",X"44",X"E7",X"01",X"6F",X"84",X"E7",X"1F",
		X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"14",X"C6",X"44",X"E7",X"84",X"E7",X"89",X"FE",X"FF",
		X"E7",X"89",X"00",X"FF",X"6F",X"1F",X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"14",X"6F",X"89",
		X"FE",X"FF",X"6F",X"89",X"00",X"FF",X"7E",X"E5",X"44",X"1C",X"17",X"10",X"0D",X"06",X"04",X"74",
		X"78",X"7F",X"85",X"89",X"8C",X"15",X"90",X"83",X"05",X"AC",X"00",X"FF",X"70",X"58",X"0F",X"3F",
		X"51",X"E8",X"14",X"90",X"5D",X"11",X"1F",X"A4",X"0A",X"67",X"8E",X"00",X"36",X"10",X"8E",X"00",
		X"D3",X"FE",X"00",X"36",X"34",X"36",X"6F",X"E4",X"E6",X"E4",X"4F",X"4C",X"58",X"26",X"04",X"E6",
		X"C0",X"58",X"5C",X"24",X"F6",X"8D",X"58",X"80",X"02",X"A7",X"61",X"86",X"03",X"8D",X"50",X"E7",
		X"E4",X"E6",X"61",X"26",X"0C",X"84",X"07",X"27",X"06",X"AE",X"62",X"31",X"21",X"20",X"D9",X"35",
		X"B6",X"84",X"07",X"27",X"02",X"8B",X"07",X"34",X"26",X"B6",X"BF",X"FF",X"84",X"FE",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"1F",X"10",X"46",X"56",X"1F",X"98",X"E6",X"63",X"1F",X"02",X"A6",X"E4",
		X"25",X"04",X"48",X"48",X"48",X"48",X"AA",X"A4",X"A7",X"A4",X"30",X"01",X"6A",X"61",X"26",X"E4",
		X"B6",X"BF",X"FF",X"8A",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"26",X"20",X"99",X"34",
		X"02",X"86",X"01",X"58",X"26",X"04",X"E6",X"C0",X"58",X"5C",X"49",X"6A",X"E4",X"26",X"F4",X"32",
		X"61",X"39",X"01",X"72",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"AE",X"04",X"27",X"6F",X"AB",X"22",X"20",
		X"14",X"10",X"AE",X"04",X"27",X"66",X"1F",X"89",X"84",X"F0",X"C4",X"0F",X"AB",X"23",X"19",X"A7",
		X"23",X"1F",X"98",X"A9",X"22",X"19",X"A7",X"22",X"6C",X"24",X"A6",X"21",X"89",X"00",X"19",X"A7",
		X"21",X"A6",X"A4",X"89",X"00",X"19",X"24",X"02",X"8B",X"10",X"A7",X"A4",X"DC",X"97",X"27",X"3C",
		X"EC",X"21",X"AB",X"27",X"19",X"10",X"A3",X"28",X"25",X"32",X"A6",X"29",X"9B",X"98",X"19",X"A7",
		X"29",X"A6",X"28",X"99",X"97",X"19",X"A7",X"28",X"81",X"30",X"25",X"0C",X"8B",X"80",X"19",X"A7",
		X"28",X"A6",X"27",X"8B",X"80",X"19",X"A7",X"27",X"34",X"30",X"BD",X"87",X"19",X"8E",X"EF",X"67",
		X"BD",X"E0",X"2D",X"C6",X"05",X"BD",X"3B",X"2B",X"35",X"30",X"20",X"C4",X"39",X"A0",X"50",X"1A",
		X"55",X"A0",X"4C",X"24",X"D9",X"E7",X"D8",X"A0",X"4D",X"27",X"D9",X"E7",X"D4",X"A0",X"4D",X"2A",
		X"D9",X"E7",X"D8",X"A0",X"4E",X"2D",X"D9",X"E7",X"D4",X"A0",X"4E",X"30",X"D9",X"E7",X"D8",X"A0",
		X"4F",X"33",X"D9",X"E7",X"D4",X"00",X"00",X"FF",X"A0",X"4F",X"36",X"D9",X"E7",X"D8",X"00",X"00",
		X"FF",X"A0",X"5A",X"1A",X"77",X"A0",X"56",X"4B",X"D9",X"E7",X"D8",X"A0",X"57",X"4E",X"D9",X"E7",
		X"D4",X"A0",X"57",X"51",X"D9",X"E7",X"D8",X"A0",X"58",X"54",X"D9",X"E7",X"D4",X"A0",X"58",X"57",
		X"D9",X"E7",X"D8",X"A0",X"59",X"5A",X"D9",X"E7",X"D4",X"00",X"00",X"FF",X"A0",X"59",X"5D",X"D9",
		X"E7",X"D8",X"00",X"00",X"FF",X"AE",X"4D",X"30",X"88",X"2B",X"AF",X"4F",X"10",X"AE",X"4D",X"EE",
		X"22",X"10",X"AE",X"02",X"2B",X"0B",X"E6",X"94",X"AD",X"98",X"04",X"AE",X"4F",X"30",X"06",X"20",
		X"E9",X"86",X"02",X"BD",X"E0",X"37",X"AE",X"4D",X"E6",X"94",X"27",X"F5",X"6F",X"94",X"30",X"04",
		X"E6",X"94",X"26",X"D6",X"30",X"06",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"CC",X"30",X"06",
		X"20",X"C8",X"30",X"0C",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",X"BE",X"30",X"06",X"20",X"BA",
		X"30",X"0C",X"20",X"B6",X"56",X"56",X"56",X"56",X"C4",X"0F",X"86",X"17",X"3D",X"34",X"01",X"1A",
		X"F0",X"E3",X"9F",X"4A",X"68",X"C3",X"00",X"02",X"FD",X"CA",X"02",X"CC",X"07",X"03",X"FD",X"CA",
		X"06",X"10",X"BF",X"CA",X"04",X"CC",X"12",X"EE",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"1F",X"30",
		X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"01",X"86",X"01",X"7E",X"E0",X"37",X"00",X"51",X"00",
		X"00",X"55",X"00",X"00",X"50",X"00",X"05",X"55",X"00",X"05",X"55",X"00",X"00",X"55",X"50",X"01",
		X"10",X"55",X"00",X"57",X"00",X"00",X"77",X"00",X"00",X"07",X"00",X"00",X"77",X"70",X"00",X"77",
		X"70",X"07",X"77",X"00",X"77",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
		X"38",X"38",X"38",X"38",X"38",X"38",X"30",X"30",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"80",X"80",X"80",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",
		X"C4",X"84",X"84",X"84",X"84",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"8A",X"8A",X"8A",X"AA",X"AA",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",
		X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"2A",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"02",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",
		X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"A0",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"18",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"08",
		X"08",X"08",X"08",X"08",X"08",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"28",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",
		X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"32",X"22",X"22",X"22",X"22",X"22",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"24",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"84",X"84",X"8C",X"8C",X"8C",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8D",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"6F",X"4D",X"6F",X"4E",X"6F",X"4F",X"86",X"01",
		X"BD",X"E0",X"37",X"AE",X"4D",X"A6",X"81",X"AB",X"4F",X"A7",X"4F",X"AF",X"4D",X"2A",X"EF",X"B1",
		X"EE",X"C1",X"27",X"E4",X"BD",X"7A",X"75",X"20",X"DF",X"F0",X"F0",X"20",X"01",X"80",X"48",X"40",
		X"48",X"E0",X"01",X"F8",X"F8",X"28",X"01",X"10",X"F8",X"68",X"5E",X"48",X"10",X"01",X"20",X"28",
		X"5E",X"28",X"58",X"28",X"28",X"2E",X"68",X"20",X"01",X"30",X"58",X"3E",X"28",X"38",X"3E",X"28",
		X"2E",X"48",X"50",X"01",X"40",X"B8",X"4E",X"98",X"40",X"01",X"80",X"88",X"3E",X"28",X"B0",X"01",
		X"D0",X"28",X"2E",X"48",X"C0",X"01",X"00",X"10",X"01",X"F0",X"F0",X"20",X"01",X"F0",X"F0",X"20",
		X"01",X"70",X"58",X"30",X"58",X"E0",X"01",X"10",X"A8",X"B8",X"5E",X"48",X"10",X"01",X"20",X"28",
		X"5E",X"98",X"28",X"2E",X"68",X"20",X"01",X"30",X"38",X"5E",X"58",X"3E",X"28",X"2E",X"48",X"50",
		X"01",X"40",X"98",X"8E",X"78",X"40",X"01",X"80",X"68",X"30",X"2E",X"28",X"B0",X"01",X"D0",X"18",
		X"1E",X"20",X"38",X"C0",X"01",X"00",X"10",X"01",X"10",X"01",X"10",X"01",X"F0",X"F0",X"20",X"01",
		X"F0",X"F0",X"20",X"01",X"70",X"58",X"30",X"58",X"E0",X"01",X"10",X"AE",X"B8",X"5E",X"28",X"1E",
		X"18",X"10",X"01",X"20",X"28",X"5E",X"28",X"3E",X"68",X"2E",X"28",X"48",X"20",X"01",X"30",X"38",
		X"7E",X"38",X"3E",X"18",X"18",X"3E",X"38",X"50",X"01",X"40",X"18",X"28",X"38",X"28",X"18",X"8E",
		X"28",X"3E",X"28",X"40",X"01",X"80",X"18",X"4E",X"18",X"30",X"2E",X"28",X"B0",X"01",X"F0",X"F0",
		X"20",X"01",X"D0",X"1E",X"1E",X"20",X"3E",X"C0",X"01",X"00",X"10",X"01",X"10",X"01",X"10",X"01",
		X"10",X"01",X"10",X"01",X"F0",X"F0",X"20",X"01",X"F0",X"F0",X"20",X"01",X"70",X"5E",X"30",X"5E",
		X"E0",X"01",X"10",X"AE",X"4E",X"38",X"9E",X"18",X"2E",X"1E",X"1E",X"10",X"01",X"20",X"28",X"5E",
		X"28",X"3E",X"28",X"5E",X"38",X"28",X"40",X"01",X"30",X"38",X"7E",X"38",X"3E",X"18",X"18",X"3E",
		X"38",X"50",X"01",X"40",X"1E",X"28",X"3E",X"2E",X"18",X"8E",X"2E",X"5E",X"40",X"01",X"80",X"1E",
		X"4E",X"1E",X"50",X"2E",X"B0",X"01",X"A0",X"1E",X"20",X"1E",X"1E",X"10",X"1E",X"20",X"1E",X"1E",
		X"C0",X"01",X"B0",X"1E",X"10",X"1E",X"20",X"2E",X"10",X"C0",X"01",X"00",X"10",X"01",X"10",X"01",
		X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"10",X"01",X"F0",X"F0",X"20",X"01",X"F0",X"F0",
		X"20",X"01",X"F0",X"F0",X"20",X"01",X"10",X"AE",X"10",X"2E",X"10",X"3E",X"90",X"1E",X"20",X"1E",
		X"1E",X"10",X"01",X"20",X"2E",X"5E",X"2E",X"3E",X"2E",X"50",X"3E",X"2E",X"40",X"01",X"30",X"3E",
		X"10",X"1E",X"20",X"1E",X"20",X"1E",X"3E",X"30",X"1E",X"1E",X"30",X"3E",X"50",X"01",X"40",X"1E",
		X"2E",X"3E",X"2E",X"1E",X"2E",X"20",X"1E",X"10",X"1E",X"20",X"1E",X"50",X"2E",X"40",X"01",X"80",
		X"1E",X"40",X"1E",X"50",X"2E",X"B0",X"01",X"F0",X"F0",X"20",X"01",X"A0",X"1E",X"20",X"1E",X"10",
		X"10",X"1E",X"20",X"10",X"1E",X"C0",X"01",X"C0",X"1E",X"10",X"1E",X"20",X"1E",X"20",X"C0",X"01",
		X"00",X"E8",X"EC",X"47",X"10",X"83",X"FF",X"F9",X"2D",X"36",X"10",X"83",X"01",X"21",X"2E",X"30",
		X"86",X"45",X"E6",X"4B",X"C1",X"65",X"25",X"08",X"86",X"81",X"C1",X"A1",X"25",X"02",X"86",X"D0",
		X"5F",X"A0",X"4B",X"2A",X"0D",X"A6",X"C8",X"11",X"2B",X"08",X"CC",X"EF",X"12",X"ED",X"C8",X"24",
		X"C6",X"01",X"A6",X"4F",X"2B",X"05",X"86",X"01",X"DD",X"32",X"39",X"86",X"FF",X"DD",X"32",X"39",
		X"BD",X"8E",X"8E",X"86",X"3C",X"BD",X"E0",X"37",X"8E",X"00",X"96",X"AF",X"47",X"AE",X"4D",X"6E",
		X"98",X"0E",X"CC",X"EE",X"C2",X"ED",X"C8",X"24",X"5F",X"20",X"D7",X"C8",X"75",X"28",X"C8",X"64",
		X"01",X"BE",X"63",X"06",X"BE",X"EE",X"3C",X"EF",X"14",X"EF",X"1E",X"F0",X"78",X"EF",X"3C",X"EF",
		X"64",X"F0",X"F0",X"E5",X"14",X"E5",X"64",X"EF",X"3C",X"F0",X"F0",X"E5",X"1E",X"E7",X"F0",X"EF",
		X"50",X"EF",X"3C",X"EF",X"14",X"F0",X"F0",X"EF",X"14",X"EF",X"3C",X"EF",X"50",X"EF",X"3C",X"EF",
		X"14",X"EF",X"3C",X"F0",X"F0",X"EF",X"14",X"EF",X"3C",X"EF",X"50",X"EF",X"3C",X"EF",X"14",X"EF",
		X"3C",X"EF",X"50",X"F0",X"78",X"70",X"F0",X"64",X"74",X"5A",X"43",X"66",X"5A",X"42",X"E9",X"0F",
		X"E9",X"0F",X"E9",X"07",X"E9",X"07",X"69",X"5A",X"41",X"DB",X"1E",X"5A",X"1E",X"41",X"5B",X"78",
		X"32",X"63",X"3C",X"32",X"76",X"1E",X"2D",X"7C",X"1E",X"2D",X"7D",X"1E",X"2D",X"73",X"1E",X"0A",
		X"79",X"0A",X"28",X"F8",X"5A",X"00",X"01",X"28",X"69",X"14",X"28",X"72",X"1E",X"09",X"F7",X"1E",
		X"00",X"01",X"06",X"5E",X"3C",X"06",X"5F",X"3C",X"06",X"5D",X"3C",X"06",X"5C",X"3C",X"06",X"59",
		X"3C",X"06",X"58",X"1E",X"06",X"00",X"01",X"50",X"69",X"14",X"46",X"ED",X"1E",X"EB",X"FF",X"7F",
		X"A5",X"46",X"ED",X"2B",X"EA",X"FF",X"7F",X"98",X"46",X"00",X"01",X"3C",X"72",X"1E",X"14",X"F7",
		X"1E",X"00",X"01",X"0A",X"5E",X"5A",X"0A",X"5F",X"5A",X"0A",X"5D",X"46",X"0A",X"5C",X"46",X"0A",
		X"59",X"46",X"0A",X"58",X"28",X"0A",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E3",X"8D",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"7E",X"F0",X"25",X"7E",X"F3",X"42",X"7E",X"F4",X"6B",X"7E",X"F9",X"45",X"7E",X"FE",X"AD",X"7E",
		X"FF",X"87",X"7E",X"FF",X"1C",X"00",X"F9",X"07",X"28",X"2F",X"00",X"A4",X"15",X"C7",X"FF",X"38",
		X"17",X"CC",X"81",X"81",X"2F",X"1A",X"FF",X"10",X"CE",X"BF",X"00",X"7F",X"C8",X"0D",X"7F",X"C8",
		X"0C",X"86",X"3C",X"B7",X"C8",X"0D",X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",
		X"B7",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"F0",X"15",
		X"10",X"8E",X"C0",X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"25",X"25",X"F7",X"86",X"02",X"10",
		X"8E",X"F0",X"68",X"8E",X"00",X"00",X"20",X"3A",X"10",X"8E",X"F0",X"6F",X"7E",X"F2",X"90",X"86",
		X"34",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"7F",X"C8",X"0E",X"86",X"A0",X"1F",X"8B",X"10",X"CE",
		X"BF",X"00",X"BD",X"3B",X"2E",X"86",X"05",X"8E",X"30",X"70",X"C6",X"99",X"BD",X"4A",X"53",X"86",
		X"06",X"8E",X"3A",X"90",X"C6",X"99",X"BD",X"4A",X"53",X"10",X"8E",X"3B",X"10",X"86",X"07",X"7E",
		X"F1",X"D0",X"1A",X"3F",X"7F",X"C9",X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",X"8E",X"00",X"00",
		X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",
		X"56",X"20",X"02",X"44",X"56",X"ED",X"81",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",
		X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",
		X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",X"C8",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",
		X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",
		X"44",X"56",X"10",X"A3",X"81",X"26",X"43",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",
		X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",
		X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",X"C5",X"1F",X"03",X"1F",X"B8",X"81",X"FF",X"26",X"05",
		X"1F",X"30",X"7E",X"F0",X"AD",X"4A",X"1F",X"8B",X"81",X"80",X"27",X"07",X"4D",X"1F",X"30",X"10",
		X"26",X"FF",X"6A",X"C6",X"01",X"F7",X"C9",X"00",X"6E",X"A4",X"30",X"1E",X"A8",X"84",X"E8",X"01",
		X"4D",X"26",X"07",X"5D",X"26",X"04",X"30",X"02",X"20",X"AD",X"CE",X"00",X"30",X"1E",X"10",X"5F",
		X"1E",X"10",X"8C",X"00",X"00",X"27",X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",X"10",X"11",X"83",
		X"00",X"30",X"23",X"EE",X"CE",X"00",X"10",X"20",X"E9",X"33",X"41",X"47",X"25",X"05",X"57",X"25",
		X"02",X"20",X"F6",X"1F",X"30",X"86",X"01",X"B7",X"C9",X"00",X"10",X"CE",X"F1",X"90",X"20",X"54",
		X"86",X"A0",X"1F",X"8B",X"1F",X"A8",X"43",X"10",X"CE",X"BF",X"00",X"BD",X"3B",X"2E",X"85",X"C0",
		X"26",X"0A",X"86",X"05",X"8E",X"30",X"70",X"C6",X"22",X"BD",X"4A",X"53",X"86",X"07",X"8E",X"40",
		X"90",X"C6",X"22",X"BD",X"4A",X"53",X"1F",X"30",X"1F",X"98",X"C6",X"22",X"BD",X"4A",X"56",X"1F",
		X"A8",X"85",X"40",X"26",X"03",X"7E",X"F8",X"D7",X"10",X"8E",X"3B",X"10",X"20",X"00",X"86",X"20",
		X"8E",X"58",X"00",X"30",X"1F",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",
		X"26",X"EE",X"6E",X"A4",X"1F",X"03",X"86",X"02",X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"F1",X"F3",
		X"7E",X"F2",X"6E",X"86",X"02",X"10",X"8E",X"F1",X"FB",X"20",X"D5",X"10",X"8E",X"F2",X"01",X"20",
		X"5D",X"86",X"01",X"10",X"8E",X"F2",X"09",X"20",X"C7",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",
		X"44",X"10",X"8E",X"F2",X"17",X"20",X"57",X"86",X"02",X"10",X"8E",X"F2",X"1F",X"20",X"B1",X"10",
		X"8E",X"F2",X"25",X"20",X"39",X"86",X"01",X"10",X"8E",X"F2",X"2D",X"20",X"A3",X"1F",X"30",X"1F",
		X"98",X"10",X"8E",X"F2",X"37",X"20",X"37",X"86",X"02",X"10",X"8E",X"F2",X"3F",X"20",X"91",X"10",
		X"8E",X"F2",X"45",X"20",X"19",X"86",X"05",X"10",X"8E",X"F2",X"4D",X"20",X"83",X"1F",X"B8",X"4A",
		X"1F",X"8B",X"26",X"96",X"10",X"8E",X"F2",X"5A",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",
		X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",
		X"46",X"46",X"46",X"84",X"C0",X"B7",X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",
		X"B7",X"C8",X"0F",X"86",X"34",X"C5",X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",
		X"1A",X"3F",X"8E",X"F3",X"20",X"8C",X"F3",X"40",X"26",X"02",X"6E",X"A4",X"A6",X"01",X"27",X"18",
		X"A6",X"84",X"5F",X"1F",X"03",X"86",X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",
		X"1E",X"03",X"26",X"F3",X"E1",X"01",X"26",X"04",X"30",X"02",X"20",X"D9",X"A6",X"84",X"44",X"44",
		X"44",X"44",X"81",X"0D",X"25",X"02",X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",
		X"CE",X"F2",X"D6",X"7E",X"F1",X"E4",X"86",X"A0",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",
		X"CE",X"BF",X"00",X"BD",X"3B",X"2E",X"1F",X"A8",X"43",X"D7",X"D5",X"85",X"C0",X"26",X"0A",X"86",
		X"05",X"8E",X"30",X"70",X"C6",X"22",X"BD",X"4A",X"53",X"86",X"08",X"8E",X"40",X"90",X"C6",X"22",
		X"BD",X"4A",X"53",X"96",X"D5",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"C6",X"22",X"BD",X"4A",X"56",
		X"1F",X"A9",X"C5",X"40",X"26",X"03",X"7E",X"F8",X"DC",X"10",X"8E",X"3B",X"10",X"7E",X"F1",X"CE",
		X"00",X"A2",X"10",X"A9",X"20",X"50",X"30",X"FA",X"40",X"A7",X"50",X"BF",X"60",X"85",X"70",X"47",
		X"80",X"51",X"90",X"00",X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",X"3D",X"E0",X"D5",X"F0",X"77",
		X"00",X"11",X"86",X"04",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",
		X"86",X"FF",X"97",X"D8",X"BD",X"F4",X"5A",X"B6",X"C8",X"0C",X"46",X"10",X"25",X"05",X"F6",X"BD",
		X"3B",X"2E",X"1A",X"BF",X"10",X"8E",X"F3",X"6B",X"7E",X"F2",X"5E",X"86",X"39",X"B7",X"CB",X"FF",
		X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"10",X"8E",X"F3",X"7E",X"7E",X"F2",X"90",X"86",X"A0",
		X"1F",X"8B",X"BD",X"3B",X"2E",X"86",X"00",X"BD",X"4A",X"62",X"C6",X"03",X"8E",X"70",X"00",X"86",
		X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"16",X"30",X"1F",X"8C",X"00",X"00",
		X"26",X"ED",X"5A",X"26",X"E7",X"10",X"8E",X"F3",X"B1",X"8E",X"00",X"00",X"86",X"FF",X"7E",X"F0",
		X"A2",X"86",X"01",X"B7",X"C9",X"00",X"86",X"A0",X"1F",X"8B",X"BD",X"3B",X"2E",X"86",X"01",X"BD",
		X"4A",X"62",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"8E",X"9C",
		X"00",X"6F",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",X"01",X"26",X"F4",X"CC",X"A5",X"5A",
		X"DD",X"DA",X"97",X"D8",X"8D",X"67",X"BD",X"F9",X"15",X"BD",X"FE",X"4A",X"86",X"02",X"24",X"24",
		X"C6",X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",X"10",X"CE",X"F4",X"02",X"86",X"03",X"7E",
		X"F1",X"E4",X"10",X"CE",X"BF",X"00",X"8D",X"45",X"86",X"A0",X"1F",X"8B",X"86",X"03",X"C1",X"1F",
		X"22",X"02",X"86",X"04",X"BD",X"3B",X"2E",X"BD",X"4A",X"62",X"BD",X"F9",X"15",X"0F",X"D7",X"BD",
		X"FD",X"D3",X"BD",X"FD",X"DC",X"BD",X"F9",X"38",X"24",X"F8",X"86",X"3F",X"B7",X"C8",X"0E",X"4F",
		X"BD",X"F9",X"45",X"4F",X"B7",X"C8",X"0E",X"BD",X"F9",X"15",X"BD",X"F7",X"65",X"BD",X"F9",X"15",
		X"BD",X"F6",X"D1",X"BD",X"F9",X"38",X"24",X"03",X"BD",X"F9",X"15",X"20",X"75",X"7F",X"C8",X"0E",
		X"86",X"34",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"39",X"8E",X"F0",X"15",X"10",X"8E",X"C0",
		X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"25",X"25",X"F7",X"39",X"86",X"3C",X"B7",X"C8",X"05",
		X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",X"3F",X"1F",X"8A",X"86",X"8F",X"BE",
		X"A6",X"D0",X"30",X"89",X"12",X"34",X"10",X"8E",X"F4",X"8D",X"7E",X"F0",X"A2",X"10",X"8E",X"F4",
		X"94",X"7E",X"F2",X"90",X"86",X"A0",X"1F",X"8B",X"10",X"CE",X"BF",X"00",X"BD",X"FE",X"4A",X"24",
		X"16",X"86",X"04",X"8C",X"CD",X"00",X"23",X"02",X"86",X"03",X"BD",X"3B",X"2E",X"BD",X"4A",X"62",
		X"86",X"39",X"B7",X"CB",X"FF",X"20",X"F9",X"8D",X"31",X"10",X"8E",X"F4",X"6B",X"86",X"04",X"7E",
		X"F1",X"D0",X"8D",X"76",X"BD",X"F9",X"15",X"BD",X"3B",X"2E",X"86",X"07",X"B7",X"C0",X"00",X"BD",
		X"F9",X"15",X"86",X"38",X"B7",X"C0",X"00",X"BD",X"F9",X"15",X"86",X"C0",X"B7",X"C0",X"00",X"BD",
		X"F9",X"15",X"8D",X"06",X"BD",X"F9",X"15",X"7E",X"F9",X"55",X"8E",X"C0",X"00",X"10",X"8E",X"F5",
		X"2A",X"EC",X"A1",X"ED",X"81",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"C0",X"10",X"25",X"F2",X"CC",
		X"00",X"00",X"8E",X"00",X"00",X"9F",X"D5",X"30",X"89",X"0F",X"00",X"ED",X"83",X"34",X"02",X"86",
		X"39",X"B7",X"CB",X"FF",X"35",X"02",X"9C",X"D5",X"26",X"F1",X"30",X"89",X"09",X"00",X"4D",X"26",
		X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",X"DC",X"39",X"05",X"05",X"28",X"28",X"80",X"80",
		X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",X"BD",X"3B",X"2E",X"4F",X"BD",X"F7",
		X"5A",X"7F",X"C9",X"00",X"86",X"FF",X"B7",X"C0",X"01",X"86",X"C0",X"B7",X"C0",X"02",X"86",X"38",
		X"B7",X"C0",X"03",X"86",X"07",X"B7",X"C0",X"04",X"10",X"8E",X"F6",X"59",X"CC",X"01",X"01",X"AE",
		X"A4",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"01",X"ED",X"81",X"AC",X"22",X"26",X"FA",X"31",X"24",
		X"10",X"8C",X"F6",X"81",X"26",X"E9",X"86",X"11",X"10",X"8E",X"F6",X"39",X"AE",X"A4",X"9F",X"D5",
		X"A7",X"84",X"0C",X"D5",X"C6",X"39",X"F7",X"CB",X"FF",X"9E",X"D5",X"AC",X"22",X"26",X"F1",X"31",
		X"24",X"10",X"8C",X"F6",X"59",X"26",X"E5",X"10",X"8E",X"F6",X"81",X"AE",X"A4",X"9F",X"D5",X"A6",
		X"24",X"A7",X"84",X"0C",X"D5",X"C6",X"39",X"F7",X"CB",X"FF",X"9E",X"D5",X"AC",X"22",X"26",X"F1",
		X"31",X"25",X"10",X"8C",X"F6",X"BD",X"26",X"E3",X"10",X"8E",X"F6",X"BD",X"AE",X"A4",X"A6",X"24",
		X"A7",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"AC",X"22",X"26",X"F5",X"31",X"25",X"10",X"8C",X"F6",
		X"D1",X"26",X"E9",X"86",X"21",X"B7",X"43",X"7E",X"86",X"20",X"B7",X"93",X"7E",X"8E",X"4B",X"0A",
		X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",X"6D",
		X"26",X"EE",X"8E",X"4B",X"90",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",
		X"A7",X"80",X"8C",X"4B",X"F3",X"26",X"EE",X"8E",X"0B",X"18",X"9F",X"D5",X"9E",X"D5",X"A6",X"84",
		X"84",X"F0",X"8A",X"01",X"A7",X"84",X"D6",X"D6",X"CB",X"22",X"25",X"04",X"D7",X"D6",X"20",X"EC",
		X"C6",X"18",X"D7",X"D6",X"D6",X"D5",X"CB",X"10",X"D7",X"D5",X"C1",X"9B",X"26",X"DE",X"C6",X"01",
		X"F7",X"C9",X"00",X"C6",X"39",X"F7",X"CB",X"FF",X"39",X"04",X"07",X"94",X"07",X"04",X"29",X"94",
		X"29",X"04",X"4B",X"94",X"4B",X"04",X"6D",X"94",X"6D",X"04",X"8F",X"94",X"8F",X"04",X"B1",X"94",
		X"B1",X"04",X"D3",X"94",X"D3",X"04",X"F5",X"94",X"F5",X"03",X"07",X"03",X"F5",X"13",X"07",X"13",
		X"F5",X"23",X"07",X"23",X"F5",X"33",X"07",X"33",X"F5",X"43",X"07",X"43",X"F5",X"53",X"07",X"53",
		X"F5",X"63",X"07",X"63",X"F5",X"73",X"07",X"73",X"F5",X"83",X"07",X"83",X"F5",X"93",X"07",X"93",
		X"F5",X"45",X"05",X"52",X"05",X"44",X"45",X"06",X"52",X"06",X"44",X"45",X"07",X"52",X"07",X"00",
		X"45",X"08",X"52",X"08",X"33",X"45",X"09",X"52",X"09",X"33",X"45",X"F3",X"52",X"F3",X"33",X"45",
		X"F4",X"52",X"F4",X"33",X"45",X"F5",X"52",X"F5",X"00",X"45",X"F6",X"52",X"F6",X"44",X"45",X"F7",
		X"52",X"F7",X"44",X"04",X"7E",X"43",X"7E",X"22",X"54",X"7E",X"93",X"7E",X"22",X"02",X"6F",X"02",
		X"8E",X"04",X"03",X"6F",X"03",X"8E",X"30",X"93",X"6F",X"93",X"8E",X"00",X"94",X"6F",X"94",X"8E",
		X"34",X"BD",X"3B",X"2E",X"86",X"05",X"BD",X"4A",X"62",X"86",X"80",X"97",X"F7",X"4F",X"BD",X"F9",
		X"45",X"BD",X"F9",X"38",X"25",X"2E",X"0A",X"F7",X"26",X"F3",X"B6",X"F7",X"42",X"8D",X"6B",X"8D",
		X"24",X"8E",X"F7",X"42",X"A6",X"80",X"9F",X"D5",X"8D",X"60",X"86",X"80",X"97",X"F7",X"4F",X"BD",
		X"F9",X"45",X"BD",X"F9",X"38",X"25",X"0D",X"0A",X"F7",X"26",X"F3",X"9E",X"D5",X"8C",X"F7",X"4A",
		X"25",X"E2",X"20",X"DD",X"39",X"8E",X"00",X"00",X"10",X"8E",X"F7",X"4A",X"9F",X"D5",X"30",X"89",
		X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"C6",X"39",X"F7",X"CB",X"FF",X"9C",X"D5",X"26",
		X"F3",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"10",X"8C",X"F7",X"5A",X"26",
		X"DB",X"39",X"02",X"03",X"04",X"10",X"18",X"20",X"40",X"80",X"00",X"FF",X"11",X"EE",X"22",X"DD",
		X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",X"8E",X"C0",X"00",X"A7",X"80",X"8C",
		X"C0",X"10",X"25",X"F9",X"39",X"86",X"0A",X"97",X"D5",X"BD",X"3B",X"2E",X"86",X"06",X"BD",X"4A",
		X"62",X"C6",X"39",X"F7",X"CB",X"FF",X"CE",X"A0",X"F7",X"6F",X"C0",X"11",X"83",X"A1",X"00",X"23",
		X"F8",X"CE",X"F8",X"47",X"8D",X"28",X"86",X"34",X"B7",X"C8",X"07",X"C6",X"39",X"F7",X"CB",X"FF",
		X"8D",X"1C",X"86",X"3C",X"B7",X"C8",X"07",X"8D",X"25",X"BD",X"F9",X"38",X"24",X"09",X"C6",X"39",
		X"F7",X"CB",X"FF",X"0A",X"D5",X"27",X"06",X"4F",X"BD",X"F9",X"45",X"20",X"D4",X"39",X"AE",X"C1",
		X"27",X"0B",X"10",X"AE",X"C1",X"A6",X"84",X"A8",X"A4",X"A7",X"21",X"20",X"F1",X"39",X"CE",X"F8",
		X"5F",X"10",X"8E",X"A0",X"F7",X"C6",X"01",X"E5",X"21",X"27",X"02",X"8D",X"1B",X"33",X"43",X"58",
		X"24",X"F5",X"C6",X"39",X"F7",X"CB",X"FF",X"31",X"22",X"10",X"8C",X"A1",X"00",X"22",X"08",X"20",
		X"E4",X"10",X"8C",X"A0",X"FC",X"23",X"DE",X"39",X"34",X"14",X"86",X"3F",X"B7",X"C8",X"0E",X"E8",
		X"A4",X"E7",X"A4",X"E6",X"E4",X"E5",X"A4",X"26",X"27",X"E6",X"42",X"27",X"48",X"86",X"40",X"1F",
		X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"CC",X"34",X"02",X"FD",X"CA",X"06",X"BF",X"CA",X"04",X"C6",
		X"00",X"F7",X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"94",
		X"E6",X"42",X"27",X"21",X"86",X"40",X"1F",X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"A6",
		X"C4",X"BD",X"4A",X"5C",X"A6",X"41",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"BD",X"4A",X"5F",
		X"86",X"3C",X"B7",X"C8",X"0E",X"35",X"94",X"C8",X"0C",X"A0",X"F7",X"C8",X"04",X"A0",X"F9",X"C8",
		X"06",X"A0",X"FB",X"00",X"00",X"C8",X"04",X"A0",X"FD",X"C8",X"06",X"A0",X"FF",X"00",X"00",X"16",
		X"FF",X"2C",X"17",X"FF",X"33",X"18",X"FF",X"3A",X"19",X"FF",X"41",X"1A",X"FF",X"48",X"1B",X"FF",
		X"4F",X"1C",X"FF",X"56",X"00",X"00",X"00",X"1F",X"F1",X"5D",X"20",X"F1",X"64",X"21",X"F1",X"6B",
		X"00",X"00",X"00",X"1E",X"FF",X"72",X"1D",X"FF",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F2",X"80",X"20",X"F2",X"87",X"21",X"F2",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F3",X"CE",X"20",X"03",X"CE",X"F3",X"A5",X"10",
		X"CE",X"BF",X"00",X"10",X"8E",X"F8",X"EC",X"86",X"01",X"7E",X"F1",X"D0",X"B6",X"C8",X"0C",X"85",
		X"02",X"26",X"F0",X"10",X"8E",X"F8",X"FC",X"86",X"01",X"7E",X"F1",X"D0",X"B6",X"C8",X"0C",X"85",
		X"02",X"27",X"F0",X"10",X"8E",X"F9",X"0C",X"86",X"01",X"7E",X"F1",X"D0",X"B6",X"C8",X"0C",X"85",
		X"02",X"26",X"F0",X"6E",X"C4",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"06",X"86",X"01",X"8D",X"25",
		X"20",X"F3",X"7F",X"C0",X"00",X"BD",X"3B",X"2E",X"20",X"07",X"B6",X"C8",X"0C",X"85",X"02",X"27",
		X"06",X"86",X"01",X"8D",X"10",X"20",X"F3",X"39",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"03",X"1A",
		X"01",X"39",X"1C",X"FE",X"39",X"C6",X"39",X"8E",X"03",X"00",X"F7",X"CB",X"FF",X"30",X"1F",X"26",
		X"F9",X"4A",X"2A",X"F1",X"39",X"86",X"A0",X"1F",X"8B",X"BD",X"F4",X"5A",X"8D",X"DA",X"24",X"02",
		X"8D",X"B3",X"86",X"07",X"BD",X"4A",X"62",X"CE",X"CD",X"02",X"8E",X"1A",X"30",X"86",X"24",X"34",
		X"12",X"C6",X"88",X"BD",X"4A",X"53",X"1E",X"31",X"BD",X"3B",X"34",X"C5",X"F0",X"26",X"08",X"CA",
		X"F0",X"C5",X"0F",X"26",X"02",X"CA",X"0F",X"1F",X"98",X"43",X"34",X"06",X"BD",X"3B",X"37",X"6D",
		X"E0",X"26",X"12",X"85",X"F0",X"26",X"0E",X"8A",X"F0",X"85",X"0F",X"26",X"08",X"8A",X"0F",X"C5",
		X"F0",X"26",X"02",X"CA",X"F0",X"1F",X"02",X"1E",X"31",X"1F",X"10",X"86",X"6A",X"1F",X"01",X"35",
		X"02",X"C6",X"88",X"BD",X"4A",X"56",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"20",X"34",X"04",X"C6",
		X"88",X"BD",X"4A",X"56",X"35",X"02",X"BD",X"4A",X"56",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"12",
		X"30",X"88",X"10",X"4C",X"11",X"83",X"CD",X"38",X"23",X"95",X"86",X"2E",X"C6",X"88",X"BD",X"4A",
		X"53",X"1F",X"10",X"86",X"6E",X"1F",X"01",X"1E",X"31",X"8E",X"CD",X"20",X"BD",X"3B",X"34",X"D7",
		X"DF",X"BD",X"3B",X"37",X"DD",X"E0",X"8E",X"CD",X"38",X"BD",X"3B",X"34",X"D7",X"E2",X"BD",X"3B",
		X"37",X"DD",X"E3",X"1E",X"31",X"8D",X"20",X"C6",X"88",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",
		X"4A",X"56",X"86",X"32",X"BD",X"4A",X"50",X"96",X"E1",X"BD",X"4A",X"56",X"86",X"39",X"B7",X"CB",
		X"FF",X"BD",X"F9",X"15",X"7E",X"FB",X"02",X"34",X"30",X"8D",X"67",X"DC",X"DF",X"27",X"0C",X"86",
		X"99",X"34",X"02",X"97",X"E1",X"0F",X"E0",X"0F",X"DF",X"20",X"3D",X"96",X"E1",X"34",X"02",X"DC",
		X"DC",X"DD",X"DF",X"96",X"DE",X"97",X"E1",X"CC",X"00",X"00",X"DD",X"DC",X"97",X"DE",X"86",X"04",
		X"08",X"E1",X"09",X"E0",X"09",X"DF",X"09",X"DE",X"4A",X"26",X"F5",X"8E",X"A0",X"E2",X"10",X"8E",
		X"A0",X"E2",X"CE",X"A0",X"E2",X"8D",X"13",X"DC",X"DE",X"DD",X"E5",X"DC",X"E0",X"DD",X"E7",X"8E",
		X"A0",X"E9",X"8D",X"06",X"8D",X"04",X"8D",X"21",X"35",X"B2",X"34",X"70",X"C6",X"04",X"20",X"04",
		X"34",X"70",X"C6",X"03",X"1C",X"FE",X"A6",X"82",X"A9",X"A2",X"19",X"A7",X"C2",X"5A",X"26",X"F6",
		X"35",X"F0",X"CC",X"00",X"00",X"DD",X"DC",X"97",X"DE",X"DC",X"E2",X"26",X"0C",X"96",X"E4",X"26",
		X"08",X"CC",X"00",X"00",X"DD",X"DF",X"97",X"E1",X"39",X"86",X"07",X"97",X"E5",X"8E",X"A0",X"DF",
		X"10",X"8E",X"A0",X"E5",X"CE",X"A0",X"E9",X"8D",X"29",X"0A",X"E5",X"26",X"02",X"20",X"23",X"86",
		X"04",X"08",X"E1",X"09",X"E0",X"09",X"DF",X"09",X"DE",X"09",X"DD",X"09",X"DC",X"4A",X"26",X"F1",
		X"8D",X"AE",X"25",X"02",X"20",X"E3",X"DC",X"E6",X"DD",X"DC",X"96",X"E8",X"97",X"DE",X"0C",X"E1",
		X"20",X"EE",X"34",X"20",X"C6",X"03",X"86",X"99",X"A0",X"A2",X"A7",X"A4",X"5A",X"26",X"F7",X"10",
		X"AE",X"E4",X"C6",X"03",X"1A",X"01",X"A6",X"3F",X"89",X"00",X"19",X"A7",X"A2",X"5A",X"26",X"F6",
		X"35",X"A0",X"8E",X"CC",X"18",X"6F",X"80",X"8C",X"CC",X"24",X"25",X"F9",X"BD",X"3B",X"2E",X"BD",
		X"F9",X"38",X"24",X"03",X"BD",X"F9",X"15",X"86",X"08",X"BD",X"4A",X"62",X"CE",X"CC",X"00",X"8E",
		X"1A",X"20",X"86",X"30",X"34",X"12",X"C6",X"22",X"BD",X"4A",X"5C",X"D7",X"E9",X"D7",X"DC",X"1F",
		X"12",X"BD",X"FC",X"BA",X"33",X"42",X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"12",X"30",X"0A",X"4C",
		X"11",X"83",X"CC",X"24",X"2D",X"DE",X"86",X"09",X"BD",X"4A",X"65",X"0F",X"DC",X"B6",X"CC",X"07",
		X"84",X"0F",X"81",X"09",X"26",X"0A",X"86",X"6E",X"D6",X"E9",X"8E",X"70",X"3E",X"BD",X"4A",X"5C",
		X"10",X"8E",X"16",X"20",X"CE",X"CC",X"00",X"1F",X"21",X"86",X"30",X"C6",X"33",X"DD",X"F7",X"BD",
		X"4A",X"59",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"04",X"84",X"03",X"27",X"02",X"8D",X"1F",
		X"C6",X"34",X"F7",X"C8",X"07",X"B6",X"C8",X"04",X"84",X"03",X"27",X"03",X"BD",X"FC",X"22",X"C6",
		X"3C",X"F7",X"C8",X"07",X"BD",X"F9",X"38",X"24",X"D9",X"BD",X"F9",X"15",X"7E",X"3B",X"19",X"97",
		X"FB",X"91",X"F9",X"27",X"10",X"0F",X"FA",X"96",X"FB",X"97",X"F9",X"86",X"02",X"BD",X"F9",X"45",
		X"B6",X"C8",X"04",X"26",X"18",X"C6",X"05",X"D7",X"FC",X"B6",X"C8",X"04",X"26",X"03",X"0F",X"F9",
		X"39",X"86",X"02",X"BD",X"F9",X"45",X"0A",X"FC",X"26",X"EF",X"B6",X"C8",X"04",X"85",X"02",X"26",
		X"21",X"85",X"01",X"27",X"3F",X"10",X"8C",X"16",X"20",X"27",X"39",X"8D",X"3C",X"31",X"36",X"33",
		X"5E",X"11",X"83",X"CC",X"12",X"26",X"09",X"0D",X"D9",X"27",X"05",X"31",X"A8",X"C4",X"33",X"54",
		X"20",X"1B",X"10",X"8C",X"16",X"CA",X"27",X"1C",X"8D",X"1F",X"31",X"2A",X"33",X"42",X"11",X"83",
		X"CC",X"08",X"26",X"09",X"0D",X"D9",X"27",X"05",X"31",X"A8",X"3C",X"33",X"4C",X"1F",X"21",X"DC",
		X"F7",X"BD",X"4A",X"59",X"4F",X"BD",X"F9",X"45",X"39",X"1F",X"21",X"96",X"F7",X"5F",X"BD",X"4A",
		X"59",X"39",X"97",X"FB",X"91",X"FD",X"27",X"10",X"0F",X"FE",X"96",X"FB",X"97",X"FD",X"86",X"02",
		X"BD",X"F9",X"45",X"B6",X"C8",X"04",X"26",X"19",X"C6",X"08",X"F7",X"A1",X"00",X"B6",X"C8",X"04",
		X"26",X"03",X"0F",X"FE",X"39",X"4F",X"BD",X"F9",X"45",X"7A",X"A1",X"00",X"26",X"EF",X"B6",X"C8",
		X"04",X"34",X"02",X"1F",X"31",X"BD",X"3B",X"31",X"34",X"02",X"5F",X"D7",X"E9",X"8D",X"5B",X"C6",
		X"39",X"F7",X"CB",X"FF",X"8E",X"FC",X"96",X"1F",X"30",X"30",X"85",X"35",X"06",X"C4",X"03",X"C5",
		X"02",X"26",X"0C",X"C5",X"01",X"27",X"14",X"A1",X"84",X"27",X"10",X"8B",X"99",X"20",X"06",X"A1",
		X"01",X"27",X"08",X"8B",X"01",X"19",X"1F",X"31",X"BD",X"3B",X"3A",X"C6",X"22",X"D7",X"E9",X"BD",
		X"FC",X"BA",X"4F",X"7E",X"F9",X"45",X"00",X"99",X"01",X"99",X"00",X"01",X"00",X"09",X"00",X"99",
		X"00",X"99",X"00",X"99",X"01",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"03",X"20",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"1F",X"30",X"54",X"8E",X"FD",X"17",
		X"30",X"85",X"6D",X"84",X"2B",X"29",X"1F",X"31",X"BD",X"3B",X"31",X"11",X"83",X"CC",X"06",X"26",
		X"08",X"97",X"D9",X"0D",X"DC",X"26",X"02",X"8D",X"50",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"34",
		X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"D6",X"E9",X"BD",X"4A",X"5F",X"39",X"A6",
		X"84",X"85",X"01",X"26",X"1B",X"1F",X"31",X"BD",X"3B",X"34",X"86",X"0D",X"5D",X"27",X"02",X"86",
		X"44",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"D6",X"E9",X"7E",X"4A",X"5C",
		X"8D",X"B4",X"86",X"2F",X"7E",X"4A",X"59",X"81",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"34",X"76",X"8E",X"00",X"3C",X"BF",X"CA",
		X"06",X"8E",X"6A",X"48",X"BF",X"CA",X"04",X"5F",X"F7",X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",
		X"8E",X"FD",X"97",X"81",X"09",X"26",X"0E",X"34",X"12",X"86",X"6E",X"D6",X"E9",X"8E",X"70",X"3E",
		X"BD",X"4A",X"5C",X"35",X"12",X"1F",X"89",X"58",X"34",X"04",X"58",X"EB",X"E0",X"3A",X"33",X"42",
		X"1E",X"31",X"8C",X"CC",X"14",X"27",X"2E",X"A6",X"C0",X"BD",X"3B",X"3A",X"C6",X"39",X"F7",X"CB",
		X"FF",X"1E",X"31",X"31",X"2A",X"34",X"10",X"30",X"5E",X"BD",X"3B",X"31",X"85",X"F0",X"26",X"02",
		X"8A",X"F0",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"D6",X"E9",X"BD",X"4A",
		X"5F",X"35",X"10",X"20",X"CB",X"35",X"F6",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"04",X"01",
		X"02",X"04",X"00",X"06",X"00",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"01",
		X"16",X"06",X"02",X"00",X"00",X"01",X"04",X"01",X"02",X"00",X"00",X"01",X"00",X"04",X"01",X"00",
		X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"01",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BD",X"3B",X"2E",X"CC",X"FE",X"01",X"DD",X"F8",X"39",X"86",X"3F",X"B7",X"C8",
		X"0E",X"86",X"03",X"BD",X"F9",X"45",X"4F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"45",X"86",
		X"3F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"45",X"DC",X"F8",X"84",X"3F",X"B7",X"C8",X"0E",
		X"C6",X"99",X"8E",X"3A",X"80",X"86",X"22",X"BD",X"4A",X"53",X"96",X"F9",X"8A",X"F0",X"C6",X"99",
		X"BD",X"4A",X"56",X"86",X"40",X"97",X"F7",X"86",X"01",X"BD",X"F9",X"45",X"BD",X"F9",X"38",X"25",
		X"04",X"0A",X"F7",X"26",X"F2",X"96",X"D7",X"26",X"06",X"B6",X"C8",X"0C",X"46",X"24",X"1A",X"8E",
		X"57",X"80",X"96",X"F9",X"8A",X"F0",X"C6",X"00",X"BD",X"4A",X"56",X"DC",X"F8",X"1A",X"01",X"49",
		X"5C",X"C1",X"07",X"25",X"02",X"8D",X"8F",X"DD",X"F8",X"39",X"8E",X"CC",X"00",X"10",X"8E",X"9C",
		X"00",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",X"C6",X"06",X"DE",X"DA",X"10",X"9E",
		X"D9",X"8E",X"CC",X"00",X"BD",X"FE",X"AD",X"A7",X"80",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",
		X"00",X"26",X"F1",X"10",X"9F",X"D9",X"DF",X"DA",X"8E",X"CC",X"00",X"BD",X"FE",X"AD",X"A8",X"80",
		X"84",X"0F",X"26",X"24",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"ED",X"5A",X"26",
		X"CB",X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"9C",X"00",X"10",X"8E",X"CC",X"00",X"A6",X"C0",X"A7",
		X"A0",X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",X"8D",X"EC",X"1A",X"01",X"39",X"34",X"04",X"D6",
		X"D9",X"86",X"03",X"3D",X"CB",X"11",X"96",X"DB",X"44",X"44",X"44",X"98",X"DB",X"44",X"06",X"DA",
		X"06",X"DB",X"DB",X"DB",X"D9",X"DA",X"D7",X"D9",X"96",X"D9",X"35",X"84",X"20",X"4A",X"4F",X"55",
		X"53",X"54",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"20",
		X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",
		X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",
		X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",
		X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"6E",X"9F",X"EF",X"F8",X"86",X"0D",X"8E",X"FF",
		X"E0",X"E6",X"84",X"E7",X"C8",X"17",X"E6",X"80",X"E7",X"C6",X"4C",X"81",X"15",X"26",X"F7",X"4F",
		X"A7",X"C8",X"16",X"31",X"C8",X"14",X"10",X"AF",X"C8",X"2B",X"86",X"04",X"BD",X"E0",X"37",X"C6",
		X"0D",X"EB",X"C8",X"16",X"A6",X"C8",X"17",X"A7",X"C5",X"A6",X"C8",X"16",X"4C",X"81",X"08",X"26",
		X"01",X"4F",X"81",X"04",X"26",X"13",X"30",X"4D",X"E6",X"80",X"34",X"04",X"E6",X"80",X"E7",X"1E",
		X"AC",X"C8",X"2B",X"2F",X"F7",X"35",X"04",X"E7",X"1F",X"A7",X"C8",X"16",X"8B",X"0D",X"E6",X"C6",
		X"E7",X"C8",X"17",X"C6",X"E8",X"E7",X"C6",X"8E",X"A0",X"17",X"31",X"4D",X"A6",X"A0",X"A7",X"80",
		X"8C",X"A0",X"1E",X"2F",X"F7",X"20",X"B3",X"86",X"77",X"97",X"D5",X"8E",X"09",X"12",X"8D",X"34",
		X"30",X"89",X"06",X"00",X"8C",X"8D",X"00",X"25",X"F5",X"8D",X"24",X"30",X"0C",X"8C",X"8D",X"E8",
		X"25",X"F7",X"30",X"89",X"F9",X"F8",X"8D",X"1C",X"8C",X"09",X"E3",X"30",X"89",X"FA",X"00",X"22",
		X"F5",X"30",X"89",X"01",X"FC",X"8D",X"08",X"30",X"14",X"8C",X"05",X"0E",X"22",X"F7",X"39",X"CC",
		X"00",X"08",X"20",X"03",X"CC",X"02",X"0C",X"FD",X"CA",X"06",X"BF",X"CA",X"04",X"96",X"D5",X"8B",
		X"11",X"24",X"02",X"86",X"88",X"97",X"D5",X"B7",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",X"39",
		X"AF",X"77",X"37",X"1F",X"17",X"0F",X"04",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"18",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"3C",X"00",X"E1",X"01",X"DF",X"04",X"D3",X"03",X"A1",X"06",X"20",X"07",X"1A",X"08",X"4C",
		X"0D",X"D9",X"0D",X"E1",X"0D",X"E9",X"0D",X"F1",X"0D",X"F9",X"23",X"2A",X"0E",X"65",X"2B",X"A1",
		X"2C",X"1F",X"2C",X"9D",X"2D",X"5F",X"2E",X"49",X"2F",X"0B",X"31",X"0B",X"32",X"F6",X"34",X"12",
		X"34",X"18",X"34",X"1E",X"34",X"A8",X"0A",X"48",X"39",X"1B",X"39",X"1B",X"00",X"C1",X"00",X"4A",
		X"01",X"45",X"15",X"03",X"00",X"4A",X"01",X"45",X"15",X"02",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"88",X"8C",X"CC",X"CA",X"AE",
		X"EC",X"CC",X"CC",X"88",X"8C",X"CC",X"AA",X"CC",X"CC",X"CC",X"CC",X"C0",X"88",X"CC",X"C8",X"88",
		X"88",X"EE",X"CC",X"88",X"88",X"CC",X"88",X"8C",X"EE",X"E8",X"88",X"00",X"00",X"EE",X"EE",X"EE",
		X"C8",X"88",X"CE",X"EC",X"C8",X"88",X"8C",X"EE",X"E8",X"8C",X"EE",X"00",X"00",X"00",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"8E",X"EE",X"C8",X"8C",X"CE",X"EE",X"EE",X"E8",X"00",X"00",X"00",X"00",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EC",X"EE",X"EE",X"88",X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"EE",X"EE",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"02",X"0A",X"02",X"43",X"02",X"0A",X"02",X"43",X"02",X"0A",X"02",X"40",X"02",X"0A",X"02",
		X"3E",X"02",X"0A",X"02",X"3C",X"02",X"0A",X"02",X"3B",X"02",X"33",X"02",X"39",X"81",X"00",X"81",
		X"00",X"01",X"97",X"00",X"EF",X"7E",X"45",X"1C",X"03",X"00",X"EF",X"7E",X"45",X"1C",X"02",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"CC",X"CC",X"C8",X"88",X"88",X"CC",X"88",X"8A",X"CC",
		X"88",X"88",X"CC",X"8C",X"CC",X"CA",X"AC",X"CC",X"AA",X"AA",X"88",X"CC",X"88",X"8A",X"A0",X"00",
		X"0E",X"EE",X"EE",X"EE",X"E8",X"88",X"88",X"CC",X"CC",X"88",X"8C",X"EE",X"E8",X"88",X"88",X"88",
		X"AA",X"88",X"CE",X"E8",X"88",X"88",X"80",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"88",X"88",
		X"88",X"88",X"CE",X"EE",X"EE",X"E8",X"C8",X"88",X"8C",X"CE",X"EE",X"EE",X"E8",X"88",X"80",X"00",
		X"00",X"00",X"00",X"CC",X"C8",X"88",X"8E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"EE",X"EE",
		X"E8",X"8E",X"EE",X"EC",X"8E",X"EE",X"E0",X"00",X"00",X"00",X"00",X"88",X"8E",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"CE",X"EE",X"E8",X"EE",X"EE",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",
		X"88",X"00",X"00",X"08",X"EE",X"EE",X"E0",X"02",X"01",X"02",X"44",X"02",X"01",X"02",X"44",X"02",
		X"04",X"02",X"44",X"02",X"07",X"02",X"44",X"02",X"09",X"02",X"44",X"02",X"09",X"02",X"44",X"02",
		X"1E",X"02",X"44",X"81",X"00",X"81",X"00",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",X"29",
		X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",
		X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"03",
		X"79",X"01",X"ED",X"2B",X"51",X"28",X"0D",X"01",X"ED",X"2B",X"51",X"28",X"0C",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AC",X"CC",X"C8",X"EE",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"EC",X"CC",X"AC",X"CA",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AC",X"CC",X"CC",X"CC",
		X"CC",X"C8",X"8E",X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DE",X"88",X"88",X"88",X"88",X"CC",X"CC",X"CC",X"CC",X"CA",X"AA",X"AC",X"CC",X"CC",X"CA",X"AA",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"0C",X"CC",X"C8",X"88",X"88",X"CC",X"CC",X"88",X"88",X"EE",
		X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DE",X"E8",X"88",X"88",X"88",
		X"88",X"88",X"8C",X"CC",X"CC",X"CC",X"8C",X"C8",X"8C",X"CC",X"CC",X"88",X"8E",X"EE",X"EE",X"E0",
		X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"E8",X"8E",X"E8",X"88",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"8E",X"EE",X"88",X"88",X"8E",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"EE",X"EE",X"EE",X"EC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"CC",X"88",X"88",X"88",X"EE",X"E8",X"88",X"8E",X"EE",X"E8",X"88",X"8E",X"88",X"8E",
		X"EE",X"88",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"CC",X"8C",X"C8",X"88",X"88",
		X"EE",X"EE",X"88",X"88",X"8E",X"C8",X"88",X"00",X"00",X"00",X"00",X"00",X"CC",X"88",X"88",X"88",
		X"EE",X"EE",X"88",X"EE",X"E8",X"EE",X"88",X"8E",X"EE",X"E8",X"88",X"EE",X"E8",X"88",X"CC",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"88",X"88",X"EE",X"EE",X"E8",X"CC",X"88",X"EE",X"EE",X"88",X"8E",X"EE",
		X"E8",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"88",X"8E",X"EE",X"EE",X"EE",X"EE",X"E8",X"8E",
		X"EE",X"E8",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"88",X"CE",X"EE",X"EE",X"EE",X"88",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"88",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"02",X"58",X"02",X"01",X"02",
		X"58",X"02",X"04",X"02",X"55",X"02",X"07",X"02",X"54",X"02",X"09",X"02",X"54",X"02",X"07",X"02",
		X"54",X"02",X"07",X"02",X"52",X"02",X"0D",X"02",X"43",X"02",X"19",X"02",X"2E",X"81",X"00",X"81",
		X"00",X"04",X"AF",X"03",X"AF",X"01",X"8A",X"24",X"0C",X"03",X"AF",X"01",X"8A",X"24",X"03",X"0A",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"EE",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"EA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"06",
		X"AA",X"AA",X"AA",X"CC",X"C8",X"8E",X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DE",X"88",X"88",X"CE",X"AA",X"CC",X"A8",X"88",X"88",X"88",X"CC",X"CC",X"08",
		X"88",X"88",X"88",X"8E",X"E8",X"88",X"EE",X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DE",X"E8",X"88",X"C8",X"EE",X"88",X"88",X"CC",X"CE",X"EE",X"EE",X"E0",X"00",X"08",
		X"88",X"88",X"88",X"88",X"EE",X"E8",X"88",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"88",X"C8",X"EE",X"E8",X"88",X"88",X"8E",X"EE",X"EE",X"EE",X"00",X"00",X"08",
		X"88",X"88",X"88",X"88",X"EE",X"EE",X"E8",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"EE",X"EE",X"EE",X"88",X"88",X"CC",X"CC",X"C8",X"88",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"EE",X"EE",X"EE",X"EE",X"EC",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"C8",X"8E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"02",
		X"01",X"02",X"62",X"02",X"01",X"02",X"62",X"02",X"01",X"02",X"5F",X"02",X"01",X"02",X"5E",X"02",
		X"01",X"02",X"5E",X"02",X"2F",X"02",X"5B",X"02",X"33",X"02",X"5C",X"02",X"4C",X"02",X"5C",X"81",
		X"00",X"81",X"00",X"06",X"D6",X"04",X"E1",X"65",X"81",X"19",X"0F",X"04",X"E1",X"65",X"81",X"19",
		X"0F",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EE",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"EA",X"AA",X"AA",X"AA",X"CC",X"C8",
		X"88",X"88",X"AA",X"AA",X"AC",X"CC",X"C8",X"88",X"8E",X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DE",X"8C",X"AA",X"8C",X"C0",X"08",X"88",X"8E",X"EE",X"EE",
		X"CC",X"CC",X"CC",X"CE",X"88",X"88",X"EE",X"ED",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DE",X"E8",X"88",X"8E",X"EE",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"88",X"8E",X"EE",
		X"E8",X"EE",X"88",X"88",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"88",X"8E",X"EE",X"E0",X"00",X"00",X"0C",X"CC",X"CC",X"88",X"88",X"8C",X"CC",X"C8",X"8E",X"EE",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"8C",
		X"C0",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"8E",X"EE",X"EE",X"EE",X"EE",
		X"E8",X"88",X"EE",X"88",X"88",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"8E",X"E8",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"8E",X"EE",X"EE",X"E8",X"8E",X"EE",X"EE",
		X"EE",X"EE",X"E8",X"88",X"EE",X"EE",X"EE",X"E8",X"88",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"C8",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"88",X"8E",X"88",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"CE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"88",X"8E",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EC",X"88",X"EE",X"EE",X"E0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"D6",X"06",X"2E",X"7F",X"8A",X"1C",X"03",X"06",X"2E",X"7F",X"8A",X"1C",X"02",X"00",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"00",X"CC",X"C8",X"8C",X"CC",X"88",X"8C",X"AC",X"CA",X"8C",
		X"88",X"88",X"AA",X"AA",X"AE",X"EC",X"C8",X"88",X"A8",X"88",X"88",X"88",X"88",X"88",X"00",X"00",
		X"E8",X"8E",X"E8",X"88",X"8E",X"EE",X"EE",X"88",X"88",X"88",X"88",X"88",X"88",X"EE",X"EE",X"C8",
		X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"EE",X"88",X"88",X"8C",X"C8",X"88",X"8E",X"88",
		X"EE",X"EC",X"88",X"88",X"88",X"8E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",
		X"00",X"EE",X"88",X"C8",X"8E",X"EE",X"EE",X"E8",X"EE",X"EE",X"CE",X"EE",X"EE",X"88",X"8E",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"0C",X"CC",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"8C",X"EE",X"E8",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"8E",X"EE",X"EE",X"EE",X"EE",X"EE",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"02",X"3A",X"02",X"01",X"02",X"39",X"02",X"02",
		X"02",X"38",X"02",X"02",X"02",X"37",X"02",X"04",X"02",X"37",X"02",X"05",X"02",X"36",X"02",X"08",
		X"02",X"35",X"02",X"15",X"02",X"33",X"02",X"15",X"02",X"33",X"02",X"1C",X"02",X"76",X"02",X"29",
		X"02",X"76",X"02",X"37",X"02",X"76",X"02",X"39",X"02",X"76",X"02",X"3A",X"02",X"76",X"02",X"3D",
		X"02",X"4E",X"02",X"3D",X"02",X"4A",X"81",X"00",X"81",X"00",X"08",X"28",X"07",X"28",X"35",X"A3",
		X"24",X"0C",X"07",X"28",X"35",X"A3",X"24",X"03",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"88",X"CA",X"AA",X"AA",X"AA",X"CC",X"CC",X"CA",
		X"AC",X"CC",X"CC",X"AA",X"AA",X"CC",X"CC",X"AA",X"AA",X"AA",X"AA",X"CC",X"CA",X"CC",X"CA",X"CC",
		X"AA",X"CA",X"CC",X"CC",X"CC",X"CC",X"AC",X"CC",X"00",X"08",X"CC",X"CC",X"CA",X"AC",X"CC",X"C8",
		X"8A",X"AA",X"CC",X"CC",X"CC",X"CC",X"AA",X"A8",X"CC",X"AC",X"CC",X"8E",X"EE",X"88",X"88",X"CC",
		X"C8",X"88",X"8C",X"C8",X"88",X"88",X"EE",X"EE",X"00",X"00",X"88",X"CC",X"C8",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"8C",X"CC",X"CC",X"CC",X"CC",X"CA",X"AE",X"EE",X"EE",X"E8",X"88",
		X"88",X"88",X"EE",X"8E",X"EE",X"EE",X"00",X"00",X"00",X"00",X"08",X"88",X"EE",X"EE",X"EE",X"88",
		X"EE",X"EE",X"EE",X"88",X"EE",X"CC",X"88",X"EE",X"88",X"88",X"8C",X"CC",X"AE",X"EE",X"EE",X"E8",
		X"8E",X"88",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"E8",X"88",X"8E",X"E8",X"E8",X"EE",X"8E",X"EE",X"EE",X"88",X"88",X"CA",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"88",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"EE",X"EE",X"EE",X"EE",X"E8",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"02",X"40",X"02",X"01",X"02",X"40",
		X"02",X"04",X"02",X"40",X"02",X"05",X"02",X"3C",X"02",X"06",X"02",X"36",X"02",X"09",X"02",X"38",
		X"02",X"10",X"02",X"2A",X"02",X"1A",X"02",X"28",X"81",X"00",X"81",X"00",X"09",X"F8",X"09",X"3E",
		X"1B",X"D3",X"59",X"06",X"09",X"3E",X"1B",X"D3",X"59",X"06",X"08",X"CE",X"1B",X"D3",X"0C",X"09",
		X"08",X"66",X"70",X"D3",X"0C",X"09",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"88",X"88",X"8C",X"CC",X"CC",X"CC",X"C0",X"88",X"88",
		X"CC",X"CC",X"C8",X"88",X"8C",X"A0",X"CC",X"8C",X"CC",X"CC",X"CE",X"E8",X"C8",X"00",X"EC",X"8C",
		X"CC",X"EE",X"E8",X"EE",X"00",X"00",X"8E",X"E8",X"EE",X"88",X"8E",X"E0",X"00",X"00",X"88",X"EE",
		X"E8",X"88",X"E0",X"00",X"00",X"00",X"88",X"88",X"8E",X"00",X"00",X"00",X"00",X"00",X"8E",X"E8",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"88",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"8E",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CC",X"CC",
		X"CC",X"88",X"88",X"8C",X"CC",X"CC",X"0E",X"EE",X"EE",X"88",X"88",X"CC",X"CC",X"CC",X"0E",X"EE",
		X"EE",X"EE",X"88",X"88",X"8C",X"88",X"00",X"00",X"AC",X"C8",X"8C",X"CC",X"CC",X"88",X"00",X"00",
		X"EC",X"CE",X"EE",X"E8",X"EE",X"88",X"00",X"00",X"0E",X"88",X"EE",X"EE",X"E8",X"88",X"00",X"00",
		X"00",X"E8",X"88",X"88",X"88",X"C8",X"00",X"00",X"00",X"0E",X"EE",X"EE",X"E8",X"88",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"CC",X"CC",X"C8",X"EE",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"E8",X"CC",X"CC",
		X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AC",X"CC",X"CC",X"CC",X"88",X"88",X"CC",X"8E",X"ED",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DE",X"88",X"88",X"CC",X"CC",X"CA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AC",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",X"01",X"02",X"BA",X"02",X"01",X"02",X"BA",
		X"02",X"01",X"02",X"B9",X"02",X"02",X"02",X"B9",X"02",X"02",X"02",X"B8",X"02",X"05",X"02",X"B6",
		X"02",X"05",X"02",X"B5",X"02",X"06",X"02",X"B3",X"02",X"07",X"02",X"B0",X"02",X"08",X"02",X"AF",
		X"02",X"0E",X"02",X"AE",X"02",X"0F",X"02",X"AD",X"02",X"10",X"02",X"AB",X"02",X"10",X"02",X"AB",
		X"02",X"10",X"02",X"AB",X"02",X"10",X"02",X"AB",X"02",X"10",X"02",X"AB",X"02",X"10",X"02",X"AB",
		X"02",X"10",X"02",X"AB",X"81",X"00",X"81",X"00",X"0E",X"9F",X"76",X"F7",X"29",X"C7",X"B7",X"F2",
		X"F4",X"15",X"DC",X"43",X"56",X"4D",X"62",X"97",X"29",X"C7",X"37",X"D8",X"BD",X"0A",X"1A",X"50",
		X"B5",X"C4",X"8A",X"E4",X"9B",X"B6",X"AC",X"59",X"A9",X"7A",X"85",X"DE",X"56",X"96",X"56",X"B1",
		X"5E",X"31",X"93",X"96",X"52",X"EF",X"AC",X"C4",X"A9",X"25",X"2A",X"95",X"AC",X"C8",X"AA",X"52",
		X"A9",X"26",X"B3",X"4A",X"E4",X"AB",X"1C",X"3F",X"62",X"4D",X"43",X"D5",X"2F",X"50",X"AD",X"24",
		X"AD",X"42",X"B5",X"89",X"55",X"0A",X"D4",X"23",X"7D",X"4B",X"D7",X"29",X"50",X"AD",X"52",X"B5",
		X"8B",X"5C",X"AD",X"13",X"29",X"49",X"2D",X"58",X"B5",X"20",X"BD",X"63",X"DD",X"C7",X"04",X"F7",
		X"3D",X"02",X"78",X"A5",X"C9",X"15",X"3E",X"7B",X"98",X"B0",X"DA",X"54",X"2F",X"54",X"EC",X"12",
		X"86",X"D8",X"EC",X"12",X"86",X"F3",X"FE",X"E5",X"6A",X"FC",X"A7",X"8B",X"0F",X"A5",X"6F",X"94",
		X"EA",X"50",X"02",X"4F",X"C3",X"14",X"00",X"93",X"F0",X"85",X"3E",X"53",X"A9",X"4F",X"17",X"1F",
		X"42",X"FD",X"4F",X"70",X"09",X"7F",X"A8",X"7B",X"80",X"4B",X"FD",X"42",X"BD",X"4F",X"E2",X"40",
		X"F9",X"27",X"B9",X"40",X"09",X"7F",X"08",X"50",X"02",X"5F",X"C3",X"9F",X"C4",X"90",X"47",X"53",
		X"80",X"4D",X"E8",X"70",X"09",X"BF",X"29",X"F3",X"F8",X"9E",X"3F",X"9F",X"E0",X"13",X"7A",X"1C",
		X"02",X"6F",X"42",X"9E",X"22",X"01",X"3E",X"41",X"33",X"B1",X"04",X"CE",X"85",X"3C",X"44",X"47",
		X"F3",X"80",X"4B",X"EC",X"70",X"09",X"7D",X"0C",X"44",X"47",X"D0",X"E0",X"12",X"79",X"07",X"00",
		X"93",X"F3",X"11",X"20",X"04",X"D9",X"88",X"90",X"72",X"B5",X"4A",X"51",X"F2",X"D4",X"13",X"0B",
		X"51",X"62",X"B5",X"CC",X"44",X"83",X"14",X"EA",X"7E",X"E5",X"6E",X"56",X"B1",X"6A",X"51",X"4B",
		X"95",X"A2",X"45",X"38",X"4E",X"7E",X"69",X"5E",X"F5",X"4A",X"D5",X"2B",X"58",X"AD",X"52",X"55",
		X"CF",X"73",X"11",X"11",X"9D",X"E5",X"2E",X"5B",X"A5",X"CB",X"55",X"EF",X"72",X"57",X"CB",X"51",
		X"62",X"BC",X"28",X"3F",X"4A",X"49",X"EA",X"77",X"2B",X"F2",X"BF",X"2F",X"54",X"AD",X"2F",X"F7",
		X"2B",X"51",X"C4",X"44",X"67",X"A8",X"7A",X"22",X"7E",X"95",X"7A",X"15",X"E2",X"25",X"3A",X"52",
		X"4A",X"F0",X"AC",X"FD",X"AB",X"1E",X"A7",X"CF",X"F2",X"47",X"53",X"FC",X"F5",X"0B",X"54",X"3D",
		X"7E",X"85",X"3E",X"7F",X"94",X"A8",X"F3",X"11",X"10",X"85",X"2A",X"16",X"E8",X"5F",X"E1",X"2E",
		X"57",X"A9",X"4E",X"85",X"AA",X"95",X"F9",X"5E",X"85",X"3A",X"54",X"3D",X"43",X"F0",X"B8",X"FD",
		X"2B",X"14",X"B8",X"23",X"E5",X"3E",X"49",X"F9",X"4E",X"B7",X"E8",X"7A",X"47",X"CB",X"74",X"BF",
		X"CF",X"62",X"20",X"32",X"95",X"0B",X"74",X"24",X"7C",X"6D",X"29",X"07",X"EA",X"52",X"E4",X"8E",
		X"85",X"BE",X"33",X"FC",X"B5",X"4E",X"18",X"95",X"FD",X"CF",X"D0",X"1F",X"D4",X"A7",X"42",X"FD",
		X"4E",X"1B",X"A1",X"FE",X"5B",X"A1",X"DC",X"4E",X"08",X"D6",X"FF",X"2B",X"F2",X"DF",X"2B",X"F0",
		X"87",X"E9",X"54",X"FD",X"0A",X"D5",X"E8",X"7E",X"85",X"FE",X"3E",X"C5",X"B8",X"68",X"5B",X"A9",
		X"50",X"77",X"CA",X"FC",X"A7",X"5A",X"87",X"78",X"23",X"B1",X"5B",X"B8",X"9C",X"33",X"B4",X"2B",
		X"D0",X"AF",X"42",X"DD",X"02",X"77",X"3F",X"20",X"99",X"D4",X"7F",X"AA",X"7E",X"1D",X"9F",X"98",
		X"4D",X"E8",X"53",X"E5",X"AE",X"D0",X"2F",X"42",X"9D",X"4F",X"D2",X"E7",X"F1",X"38",X"21",X"11",
		X"E8",X"17",X"E7",X"B9",X"EA",X"75",X"27",X"7C",X"02",X"21",X"4F",X"9E",X"92",X"7A",X"80",X"9F",
		X"9F",X"E7",X"F9",X"27",X"E0",X"8F",X"9F",X"A9",X"5F",X"98",X"98",X"12",X"E7",X"AC",X"4C",X"E8",
		X"18",X"91",X"D0",X"95",X"D0",X"27",X"C2",X"9E",X"82",X"11",X"4E",X"59",X"EE",X"17",X"A0",X"7F",
		X"92",X"BA",X"02",X"FA",X"94",X"B1",X"30",X"21",X"4A",X"84",X"DE",X"80",X"82",X"BD",X"4B",X"77",
		X"1D",X"CE",X"3F",X"8C",X"EC",X"82",X"9C",X"3D",X"2B",X"C9",X"28",X"D4",X"21",X"C2",X"FC",X"B7",
		X"53",X"DD",X"F5",X"C1",X"3F",X"29",X"77",X"F8",X"98",X"33",X"D3",X"7A",X"8F",X"E0",X"A2",X"BD",
		X"0A",X"F7",X"19",X"EA",X"1F",X"E3",X"3B",X"73",X"D4",X"E1",X"49",X"FE",X"7E",X"26",X"5B",X"B9",
		X"4B",X"BF",X"A0",X"43",X"DC",X"17",X"D2",X"EF",X"24",X"82",X"7F",X"51",X"C5",X"82",X"7C",X"A3",
		X"EB",X"12",X"79",X"03",X"3B",X"63",X"DC",X"AF",X"52",X"DD",X"87",X"54",X"A0",X"EE",X"D8",X"F5",
		X"79",X"A7",X"F9",X"4E",X"32",X"7F",X"95",X"E2",X"27",X"E8",X"57",X"F7",X"2B",X"72",X"9D",X"02",
		X"9E",X"A8",X"6F",X"9F",X"A1",X"EF",X"CA",X"0F",X"D0",X"A5",X"8B",X"0F",X"A9",X"FA",X"92",X"B9",
		X"23",X"6C",X"7B",X"95",X"EA",X"5F",X"A8",X"CF",X"D4",X"A0",X"DA",X"54",X"3D",X"CA",X"72",X"8F",
		X"F3",X"F4",X"29",X"C6",X"0F",X"D4",X"A0",X"4E",X"59",X"4E",X"49",X"33",X"A8",X"42",X"95",X"43",
		X"7C",X"AF",X"CF",X"4A",X"04",X"75",X"31",X"61",X"95",X"F9",X"27",X"9C",X"1A",X"E5",X"7A",X"97",
		X"EC",X"10",X"AF",X"41",X"96",X"B9",X"4E",X"71",X"5F",X"81",X"63",X"F6",X"3F",X"40",X"BD",X"CF",
		X"F3",X"F4",X"2D",X"C8",X"24",X"77",X"08",X"7E",X"C1",X"FB",X"14",X"0A",X"54",X"15",X"D4",X"A7",
		X"8A",X"04",X"29",X"50",X"93",X"C9",X"1D",X"CF",X"DC",X"3F",X"52",X"FC",X"80",X"DD",X"42",X"96",
		X"F9",X"FE",X"53",X"A9",X"7E",X"A1",X"38",X"81",X"6E",X"A5",X"7E",X"50",X"2F",X"42",X"9C",X"40",
		X"BF",X"28",X"2F",X"60",X"9D",X"0F",X"D0",X"FD",X"07",X"D4",X"A0",X"5E",X"A5",X"3B",X"1F",X"C5",
		X"03",X"12",X"F9",X"01",X"2A",X"1F",X"B0",X"5E",X"C4",X"8E",X"48",X"4E",X"C0",X"8E",X"A4",X"DE",
		X"C0",X"8E",X"22",X"5F",X"A0",X"7E",X"84",X"8E",X"85",X"FA",X"92",X"39",X"C0",X"EF",X"9F",X"A8",
		X"5E",X"C5",X"7E",X"7F",X"14",X"0A",X"4C",X"E4",X"84",X"3F",X"20",X"1D",X"C4",X"00",X"9F",X"24",
		X"13",X"F2",X"9D",X"89",X"BD",X"80",X"F7",X"34",X"1F",X"F2",X"A1",X"BB",X"95",X"F1",X"80",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"0D",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"0D",X"DD",X"DD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"D0",X"00",X"0A",X"00",X"0D",X"AF",X"35",X"51",X"0A",
		X"07",X"0A",X"00",X"0D",X"AF",X"70",X"81",X"0A",X"07",X"0A",X"00",X"0D",X"AF",X"08",X"8A",X"0A",
		X"07",X"0A",X"00",X"0D",X"AF",X"3C",X"D3",X"0A",X"07",X"0F",X"49",X"00",X"EF",X"1D",X"A2",X"11",
		X"15",X"01",X"EF",X"21",X"AA",X"10",X"C1",X"00",X"ED",X"1D",X"00",X"12",X"65",X"01",X"ED",X"21",
		X"08",X"0F",X"9D",X"00",X"ED",X"1B",X"1A",X"11",X"69",X"01",X"ED",X"1F",X"4A",X"10",X"19",X"00",
		X"ED",X"1B",X"BC",X"11",X"BD",X"02",X"ED",X"1F",X"EC",X"10",X"6D",X"00",X"ED",X"1C",X"5E",X"12",
		X"11",X"02",X"ED",X"20",X"7A",X"10",X"C1",X"00",X"ED",X"1D",X"00",X"12",X"65",X"01",X"ED",X"21",
		X"08",X"0E",X"D1",X"00",X"ED",X"1E",X"34",X"0F",X"0D",X"00",X"ED",X"22",X"3C",X"0E",X"D1",X"00",
		X"ED",X"1E",X"34",X"0F",X"0D",X"00",X"ED",X"22",X"3C",X"0E",X"D1",X"00",X"ED",X"1E",X"D3",X"0F",
		X"0D",X"00",X"ED",X"22",X"B3",X"0F",X"49",X"00",X"EE",X"15",X"7D",X"11",X"15",X"02",X"EE",X"19",
		X"AA",X"10",X"C1",X"00",X"ED",X"14",X"C7",X"12",X"65",X"01",X"ED",X"19",X"08",X"0F",X"9D",X"00",
		X"ED",X"12",X"B9",X"11",X"69",X"00",X"ED",X"17",X"0E",X"10",X"19",X"00",X"ED",X"13",X"6F",X"11",
		X"BD",X"01",X"ED",X"17",X"C4",X"10",X"6D",X"00",X"ED",X"14",X"11",X"12",X"11",X"01",X"ED",X"18",
		X"66",X"10",X"C1",X"00",X"ED",X"14",X"C7",X"12",X"65",X"01",X"ED",X"19",X"08",X"0E",X"D1",X"00",
		X"ED",X"16",X"17",X"0F",X"0D",X"01",X"ED",X"1A",X"31",X"0E",X"D1",X"00",X"ED",X"16",X"17",X"0F",
		X"0D",X"01",X"ED",X"1A",X"31",X"0E",X"D1",X"00",X"ED",X"16",X"97",X"0F",X"0D",X"00",X"ED",X"1A",
		X"A3",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",
		X"0A",X"02",X"06",X"02",X"11",X"02",X"02",X"02",X"0A",X"02",X"02",X"02",X"0E",X"02",X"02",X"02",
		X"0E",X"02",X"04",X"02",X"0D",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",
		X"0C",X"02",X"0B",X"02",X"0C",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"02",X"0A",X"02",
		X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"02",X"02",
		X"0D",X"02",X"09",X"02",X"11",X"02",X"05",X"02",X"11",X"02",X"05",X"02",X"11",X"02",X"06",X"02",
		X"0F",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",
		X"08",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",
		X"00",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",
		X"0A",X"02",X"06",X"02",X"0A",X"02",X"02",X"02",X"0A",X"02",X"02",X"02",X"0B",X"02",X"03",X"02",
		X"0B",X"02",X"04",X"02",X"0B",X"02",X"05",X"02",X"0B",X"02",X"05",X"02",X"0B",X"02",X"06",X"02",
		X"0A",X"02",X"07",X"02",X"0B",X"02",X"07",X"02",X"0B",X"02",X"07",X"02",X"0C",X"02",X"07",X"02",
		X"0D",X"02",X"07",X"02",X"0E",X"02",X"08",X"02",X"0F",X"81",X"00",X"81",X"00",X"02",X"07",X"02",
		X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",
		X"11",X"02",X"02",X"02",X"0A",X"02",X"02",X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"04",X"02",
		X"0D",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",X"0C",X"02",X"06",X"02",X"0A",X"02",X"04",X"02",
		X"0A",X"02",X"04",X"02",X"09",X"02",X"06",X"02",X"09",X"02",X"07",X"02",X"0A",X"02",X"07",X"02",
		X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"0A",X"81",X"00",X"81",
		X"00",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"02",X"07",X"02",X"09",X"02",X"07",X"02",
		X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"11",X"02",X"02",X"02",
		X"0A",X"02",X"02",X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"04",X"02",X"0D",X"02",X"05",X"02",
		X"0C",X"02",X"05",X"02",X"0C",X"02",X"06",X"02",X"0A",X"02",X"08",X"02",X"0A",X"02",X"07",X"02",
		X"0A",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"0C",X"02",X"06",X"02",X"0C",X"02",X"06",X"02",
		X"0D",X"02",X"06",X"02",X"0D",X"02",X"06",X"02",X"08",X"81",X"00",X"81",X"00",X"02",X"07",X"02",
		X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",
		X"11",X"02",X"02",X"02",X"0A",X"02",X"02",X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"04",X"02",
		X"0D",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",X"0C",X"02",X"06",X"02",X"0B",X"02",X"07",X"02",
		X"0B",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"0B",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",
		X"0D",X"02",X"05",X"02",X"0E",X"02",X"05",X"02",X"0E",X"02",X"05",X"02",X"0E",X"81",X"00",X"81",
		X"00",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",
		X"0A",X"02",X"06",X"02",X"11",X"02",X"02",X"02",X"0A",X"02",X"02",X"02",X"0E",X"02",X"03",X"02",
		X"0E",X"02",X"04",X"02",X"0D",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",X"0C",X"02",X"06",X"02",
		X"0A",X"02",X"04",X"02",X"0A",X"02",X"04",X"02",X"09",X"02",X"04",X"02",X"09",X"02",X"05",X"02",
		X"09",X"02",X"05",X"02",X"0A",X"02",X"04",X"02",X"0A",X"02",X"04",X"02",X"0A",X"02",X"04",X"02",
		X"0B",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"02",X"0A",X"02",
		X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"09",X"02",
		X"0D",X"02",X"09",X"02",X"11",X"02",X"08",X"02",X"11",X"02",X"08",X"02",X"10",X"02",X"08",X"02",
		X"0F",X"02",X"08",X"02",X"0E",X"02",X"08",X"02",X"0E",X"02",X"08",X"02",X"0D",X"02",X"08",X"02",
		X"0C",X"02",X"08",X"02",X"0C",X"02",X"07",X"02",X"0C",X"02",X"06",X"02",X"0C",X"02",X"05",X"02",
		X"0C",X"02",X"04",X"02",X"0D",X"81",X"00",X"81",X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",
		X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"02",X"02",X"0D",X"02",X"09",X"02",
		X"11",X"02",X"05",X"02",X"11",X"02",X"05",X"02",X"10",X"02",X"06",X"02",X"0F",X"02",X"07",X"02",
		X"0E",X"02",X"07",X"02",X"0E",X"02",X"09",X"02",X"0D",X"02",X"09",X"02",X"0F",X"02",X"0A",X"02",
		X"0F",X"02",X"0A",X"02",X"0D",X"02",X"09",X"02",X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",
		X"0C",X"02",X"0A",X"02",X"0C",X"02",X"09",X"02",X"0C",X"81",X"00",X"81",X"00",X"02",X"0A",X"02",
		X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"02",X"02",
		X"0D",X"02",X"09",X"02",X"11",X"02",X"05",X"02",X"11",X"02",X"05",X"02",X"10",X"02",X"06",X"02",
		X"0F",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",X"0E",X"02",X"09",X"02",X"0D",X"02",X"09",X"02",
		X"0B",X"02",X"09",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"05",X"02",X"0D",X"02",X"05",X"02",
		X"0D",X"02",X"04",X"02",X"0D",X"02",X"04",X"02",X"0D",X"02",X"0B",X"02",X"0D",X"81",X"00",X"81",
		X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",
		X"0D",X"02",X"02",X"02",X"0D",X"02",X"09",X"02",X"11",X"02",X"05",X"02",X"11",X"02",X"05",X"02",
		X"10",X"02",X"06",X"02",X"0F",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",X"0E",X"02",X"09",X"02",
		X"0D",X"02",X"08",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"07",X"02",
		X"0E",X"02",X"06",X"02",X"0E",X"02",X"05",X"02",X"0E",X"02",X"05",X"02",X"0E",X"02",X"05",X"02",
		X"0E",X"81",X"00",X"81",X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",
		X"0C",X"02",X"09",X"02",X"0D",X"02",X"02",X"02",X"0D",X"02",X"09",X"02",X"11",X"02",X"05",X"02",
		X"11",X"02",X"05",X"02",X"10",X"02",X"06",X"02",X"0F",X"02",X"07",X"02",X"0E",X"02",X"07",X"02",
		X"0E",X"02",X"09",X"02",X"0D",X"02",X"09",X"02",X"0F",X"02",X"0A",X"02",X"0F",X"02",X"0A",X"02",
		X"0F",X"02",X"0A",X"02",X"0E",X"02",X"09",X"02",X"0E",X"02",X"09",X"02",X"0F",X"02",X"09",X"02",
		X"0F",X"02",X"08",X"02",X"0F",X"81",X"00",X"81",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",
		X"06",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"94",X"C4",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"09",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"D6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"D1",X"10",X"00",X"00",X"00",X"00",X"06",X"DD",X"55",X"11",
		X"D0",X"00",X"00",X"00",X"00",X"CD",X"5D",X"D5",X"15",X"60",X"00",X"00",X"00",X"05",X"85",X"51",
		X"54",X"1D",X"60",X"00",X"00",X"04",X"84",X"C4",X"55",X"8D",X"56",X"00",X"00",X"00",X"04",X"4C",
		X"CC",X"88",X"D5",X"80",X"00",X"00",X"00",X"00",X"0D",X"DD",X"D1",X"D8",X"00",X"00",X"00",X"00",
		X"00",X"DD",X"88",X"E8",X"80",X"00",X"00",X"00",X"00",X"00",X"0E",X"88",X"08",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"08",X"CC",X"CC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"CC",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"EE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C6",X"00",X"00",X"00",X"00",X"0C",
		X"10",X"00",X"00",X"00",X"00",X"00",X"6D",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"4C",
		X"40",X"00",X"00",X"00",X"00",X"00",X"91",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",
		X"00",X"00",X"00",X"00",X"00",X"06",X"D1",X"10",X"00",X"00",X"00",X"06",X"DD",X"55",X"11",X"50",
		X"00",X"00",X"00",X"CD",X"5D",X"D5",X"15",X"D0",X"00",X"00",X"05",X"85",X"51",X"5C",X"15",X"60",
		X"00",X"00",X"84",X"CC",X"55",X"8D",X"56",X"00",X"00",X"04",X"44",X"CC",X"88",X"DD",X"80",X"00",
		X"00",X"00",X"0D",X"DD",X"D1",X"D8",X"00",X"00",X"00",X"00",X"DD",X"86",X"88",X"80",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"8C",X"CC",X"E0",X"00",X"00",X"00",X"00",X"0E",X"C8",X"EC",X"C8",X"00",
		X"00",X"00",X"00",X"08",X"C0",X"00",X"EC",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"08",X"80",
		X"00",X"00",X"00",X"08",X"CE",X"00",X"00",X"80",X"00",X"00",X"00",X"0E",X"CC",X"00",X"00",X"00",
		X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"6D",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"4C",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"D1",X"10",
		X"00",X"00",X"00",X"00",X"06",X"DD",X"55",X"11",X"50",X"00",X"00",X"00",X"00",X"CD",X"5D",X"D5",
		X"15",X"D0",X"00",X"00",X"00",X"05",X"85",X"51",X"5C",X"15",X"60",X"00",X"00",X"00",X"84",X"CC",
		X"55",X"8D",X"56",X"00",X"00",X"00",X"04",X"44",X"CC",X"88",X"DD",X"80",X"00",X"00",X"00",X"00",
		X"0D",X"DD",X"D1",X"D8",X"00",X"00",X"00",X"00",X"00",X"DD",X"60",X"08",X"88",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"C8",X"EC",X"80",X"00",X"00",X"00",X"00",X"00",X"EC",X"80",X"0C",X"8E",
		X"00",X"00",X"00",X"00",X"00",X"8C",X"80",X"00",X"CC",X"E0",X"00",X"00",X"00",X"00",X"8C",X"E0",
		X"00",X"08",X"CE",X"00",X"00",X"00",X"00",X"C8",X"00",X"00",X"0E",X"88",X"00",X"00",X"00",X"00",
		X"CC",X"00",X"00",X"0E",X"EC",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"06",X"D3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"94",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"D1",X"10",X"00",X"00",X"00",X"00",X"06",X"DD",X"55",X"11",X"D0",X"00",
		X"00",X"00",X"00",X"CD",X"5D",X"D5",X"15",X"60",X"00",X"00",X"00",X"05",X"85",X"51",X"5C",X"1D",
		X"60",X"00",X"00",X"00",X"84",X"CC",X"55",X"8D",X"56",X"00",X"00",X"00",X"04",X"44",X"CC",X"88",
		X"DD",X"80",X"00",X"00",X"00",X"00",X"0D",X"DD",X"D1",X"D8",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"68",X"8E",X"88",X"00",X"00",X"00",X"00",X"00",X"0E",X"CC",X"08",X"CE",X"00",X"00",X"00",X"00",
		X"00",X"08",X"CE",X"08",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"CE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"00",X"EC",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"0C",X"C0",X"00",X"00",X"00",X"0C",X"17",X"00",
		X"00",X"00",X"00",X"03",X"D3",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"94",X"CE",X"00",X"00",
		X"00",X"00",X"00",X"09",X"18",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"61",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"06",X"DD",X"55",X"11",X"50",X"00",X"00",
		X"00",X"CD",X"5D",X"D5",X"15",X"D0",X"00",X"00",X"05",X"85",X"51",X"5C",X"15",X"60",X"00",X"00",
		X"84",X"CC",X"55",X"8D",X"56",X"00",X"00",X"04",X"44",X"CC",X"88",X"DD",X"80",X"00",X"00",X"00",
		X"0D",X"DD",X"D1",X"D8",X"00",X"00",X"00",X"00",X"DD",X"68",X"88",X"C8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8C",X"EC",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"CE",X"CE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"EC",X"EC",X"E0",X"00",X"00",X"00",X"00",X"00",X"0E",X"CE",X"CE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"EC",X"00",X"0D",X"0A",X"00",X"00",X"00",X"00",X"00",X"6D",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"4C",X"4E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"09",X"77",X"99",X"0D",X"10",X"00",X"00",X"00",
		X"00",X"6D",X"15",X"DC",X"6D",X"10",X"00",X"00",X"00",X"06",X"15",X"51",X"5C",X"D1",X"50",X"00",
		X"00",X"00",X"6D",X"55",X"15",X"D6",X"DD",X"60",X"00",X"00",X"00",X"DD",X"55",X"5C",X"58",X"68",
		X"00",X"00",X"00",X"04",X"86",X"DC",X"CC",X"CC",X"E0",X"00",X"00",X"00",X"08",X"48",X"68",X"C4",
		X"C4",X"88",X"00",X"00",X"00",X"00",X"80",X"EE",X"88",X"4E",X"CE",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"8E",X"8E",X"00",X"00",X"00",X"0D",X"09",X"00",X"C8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"04",X"D0",X"00",X"00",X"06",X"D3",X"00",X"00",X"00",X"44",X"DD",X"00",X"00",
		X"0D",X"94",X"C4",X"E0",X"04",X"48",X"84",X"90",X"00",X"09",X"18",X"00",X"00",X"00",X"CC",X"88",
		X"C9",X"00",X"00",X"1D",X"00",X"00",X"0C",X"CC",X"CC",X"85",X"90",X"00",X"1D",X"00",X"00",X"00",
		X"0C",X"5C",X"8D",X"58",X"9D",X"16",X"00",X"00",X"00",X"CC",X"5D",X"DC",X"5D",X"D1",X"D6",X"00",
		X"00",X"00",X"08",X"4D",X"D1",X"51",X"11",X"60",X"00",X"00",X"00",X"4C",X"55",X"11",X"11",X"D6",
		X"00",X"00",X"00",X"04",X"C4",X"58",X"8C",X"1D",X"C0",X"00",X"00",X"00",X"04",X"54",X"0E",X"E8",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"E0",X"08",X"00",X"00",X"00",X"00",X"0D",X"10",
		X"00",X"00",X"3D",X"60",X"00",X"00",X"00",X"00",X"00",X"0E",X"4C",X"49",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1D",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"11",X"55",X"DD",X"60",X"00",X"00",X"00",X"00",X"06",X"51",X"5D",X"D5",X"DC",X"00",
		X"00",X"00",X"00",X"06",X"D1",X"45",X"15",X"58",X"50",X"00",X"00",X"00",X"00",X"65",X"D8",X"55",
		X"4C",X"48",X"40",X"00",X"00",X"00",X"08",X"5D",X"88",X"CC",X"C4",X"40",X"00",X"00",X"00",X"00",
		X"8D",X"1D",X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"08",X"8E",X"88",X"DD",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"80",X"88",X"E0",X"00",X"00",X"00",X"00",X"00",X"08",X"CC",X"CC",X"80",X"00",
		X"00",X"00",X"00",X"0E",X"CC",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"EE",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",
		X"80",X"00",X"00",X"00",X"0C",X"10",X"00",X"03",X"D6",X"00",X"00",X"00",X"00",X"00",X"04",X"C4",
		X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1D",X"60",X"00",X"00",X"00",X"00",X"00",X"05",
		X"11",X"55",X"DD",X"60",X"00",X"00",X"00",X"0D",X"51",X"5D",X"D5",X"DC",X"00",X"00",X"00",X"06",
		X"51",X"C5",X"15",X"58",X"50",X"00",X"00",X"00",X"65",X"D8",X"55",X"CC",X"48",X"00",X"00",X"00",
		X"08",X"DD",X"88",X"CC",X"44",X"40",X"00",X"00",X"00",X"8D",X"1D",X"DD",X"D0",X"00",X"00",X"00",
		X"00",X"08",X"88",X"68",X"DD",X"00",X"00",X"00",X"0E",X"CC",X"C8",X"E0",X"00",X"00",X"00",X"00",
		X"8C",X"CE",X"8C",X"E0",X"00",X"00",X"00",X"00",X"CE",X"00",X"0C",X"80",X"00",X"00",X"00",X"08",
		X"80",X"00",X"0F",X"80",X"00",X"00",X"00",X"08",X"00",X"00",X"EC",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CC",X"E0",X"00",X"00",X"0C",X"10",X"00",X"03",X"D6",X"00",X"00",X"00",X"00",X"00",
		X"E4",X"C4",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"19",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1D",X"60",X"00",X"00",X"00",X"00",
		X"00",X"05",X"11",X"55",X"DD",X"60",X"00",X"00",X"00",X"0D",X"51",X"5D",X"D5",X"DC",X"00",X"00",
		X"00",X"06",X"51",X"C5",X"15",X"58",X"50",X"00",X"00",X"00",X"65",X"D8",X"55",X"CC",X"48",X"00",
		X"00",X"00",X"08",X"DD",X"88",X"CC",X"44",X"40",X"00",X"00",X"00",X"8D",X"1D",X"DD",X"D0",X"00",
		X"00",X"00",X"00",X"88",X"80",X"06",X"DD",X"00",X"00",X"00",X"08",X"CE",X"8C",X"80",X"00",X"00",
		X"00",X"00",X"E8",X"C0",X"08",X"CE",X"00",X"00",X"00",X"0E",X"CC",X"00",X"08",X"C8",X"00",X"00",
		X"00",X"EC",X"80",X"00",X"0E",X"C8",X"00",X"00",X"00",X"88",X"E0",X"00",X"00",X"8C",X"00",X"00",
		X"00",X"CE",X"E0",X"00",X"00",X"CC",X"00",X"00",X"0C",X"10",X"00",X"3D",X"60",X"00",X"00",X"00",
		X"00",X"00",X"4C",X"49",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"1D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"11",X"55",X"DD",X"60",X"00",X"00",X"00",X"06",X"51",X"5D",X"D5",X"DC",
		X"00",X"00",X"00",X"06",X"D1",X"C5",X"15",X"58",X"50",X"00",X"00",X"00",X"65",X"D8",X"55",X"CC",
		X"48",X"00",X"00",X"00",X"08",X"DD",X"88",X"CC",X"44",X"40",X"00",X"00",X"00",X"8D",X"1D",X"DD",
		X"D0",X"00",X"00",X"00",X"00",X"88",X"E8",X"86",X"DD",X"00",X"00",X"00",X"00",X"EC",X"80",X"CC",
		X"E0",X"00",X"00",X"00",X"00",X"0C",X"80",X"EC",X"80",X"00",X"00",X"00",X"00",X"EC",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"CE",X"00",X"0C",
		X"80",X"00",X"00",X"00",X"0C",X"C0",X"00",X"0C",X"C0",X"00",X"03",X"17",X"00",X"3D",X"30",X"00",
		X"00",X"00",X"00",X"EC",X"49",X"D0",X"00",X"00",X"00",X"00",X"48",X"81",X"90",X"00",X"00",X"00",
		X"00",X"06",X"16",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"05",X"11",X"55",
		X"DD",X"60",X"00",X"00",X"0D",X"51",X"5D",X"D5",X"DC",X"00",X"00",X"06",X"51",X"C5",X"15",X"58",
		X"50",X"00",X"00",X"65",X"D8",X"55",X"CC",X"48",X"00",X"00",X"08",X"DD",X"88",X"CC",X"44",X"40",
		X"00",X"00",X"8D",X"1D",X"DD",X"D0",X"00",X"00",X"00",X"8C",X"88",X"86",X"DD",X"00",X"00",X"08",
		X"CE",X"C8",X"00",X"00",X"00",X"00",X"EC",X"EC",X"80",X"00",X"00",X"00",X"0E",X"CE",X"CE",X"00",
		X"00",X"00",X"00",X"EC",X"EC",X"E0",X"00",X"00",X"00",X"00",X"CE",X"CC",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"0A",X"00",X"03",X"D6",X"00",X"00",X"00",X"00",X"00",X"E4",X"C4",X"91",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"D0",X"99",X"77",
		X"90",X"00",X"00",X"00",X"01",X"D6",X"CD",X"51",X"D6",X"00",X"00",X"00",X"05",X"1D",X"C5",X"15",
		X"51",X"60",X"00",X"00",X"06",X"DD",X"6D",X"51",X"55",X"D6",X"00",X"00",X"00",X"86",X"85",X"C5",
		X"55",X"DD",X"00",X"00",X"00",X"0E",X"CC",X"CC",X"CD",X"68",X"40",X"00",X"00",X"88",X"4C",X"4C",
		X"86",X"84",X"80",X"00",X"0C",X"EC",X"E4",X"88",X"EE",X"08",X"00",X"00",X"00",X"E8",X"E8",X"E0",
		X"00",X"00",X"00",X"0D",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"00",X"00",X"00",
		X"3D",X"60",X"00",X"00",X"0D",X"40",X"C0",X"0E",X"4C",X"49",X"D0",X"00",X"00",X"DD",X"44",X"00",
		X"00",X"00",X"81",X"90",X"00",X"09",X"48",X"84",X"40",X"00",X"00",X"D1",X"00",X"00",X"9C",X"88",
		X"CC",X"00",X"00",X"00",X"D1",X"00",X"09",X"58",X"CC",X"CC",X"C0",X"00",X"00",X"61",X"D9",X"85",
		X"D8",X"C5",X"C0",X"00",X"00",X"00",X"6D",X"1D",X"D5",X"CD",X"D5",X"CC",X"00",X"00",X"00",X"06",
		X"11",X"15",X"1D",X"D4",X"80",X"00",X"00",X"00",X"00",X"6D",X"11",X"11",X"55",X"C4",X"00",X"00",
		X"00",X"00",X"0C",X"D1",X"C8",X"85",X"4C",X"40",X"00",X"00",X"00",X"00",X"88",X"8E",X"E0",X"45",
		X"40",X"00",X"00",X"00",X"00",X"80",X"0E",X"88",X"00",X"00",X"0C",X"10",X"00",X"00",X"00",X"00",
		X"00",X"08",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"7F",X"50",X"00",X"00",X"00",X"00",
		X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"8F",X"00",X"09",X"70",X"00",X"00",X"00",X"00",X"8F",X"00",X"07",X"17",X"97",X"66",
		X"66",X"00",X"8F",X"00",X"00",X"69",X"76",X"71",X"77",X"98",X"FE",X"00",X"00",X"06",X"96",X"07",
		X"97",X"7F",X"80",X"00",X"00",X"00",X"97",X"96",X"77",X"79",X"00",X"00",X"00",X"00",X"66",X"98",
		X"99",X"60",X"00",X"00",X"00",X"00",X"88",X"8E",X"88",X"00",X"00",X"00",X"00",X"0F",X"F8",X"00",
		X"F8",X"00",X"00",X"00",X"00",X"0E",X"FF",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"08",X"FF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",
		X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"F8",X"00",X"00",X"00",X"0C",X"10",X"00",X"00",
		X"00",X"00",X"00",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F5",X"00",X"00",X"00",
		X"00",X"00",X"00",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"F0",X"00",X"09",X"70",X"00",X"00",X"00",X"00",X"8F",X"00",X"07",X"17",
		X"97",X"66",X"66",X"00",X"8F",X"00",X"00",X"69",X"76",X"71",X"77",X"98",X"F8",X"00",X"00",X"06",
		X"96",X"07",X"97",X"7F",X"80",X"00",X"00",X"00",X"97",X"99",X"11",X"77",X"00",X"00",X"00",X"00",
		X"69",X"97",X"77",X"96",X"00",X"00",X"00",X"00",X"06",X"88",X"88",X"60",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"8E",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"8F",X"F8",X"00",X"00",X"00",X"00",X"00",X"0E",X"F8",X"0F",X"F8",X"00",X"00",X"00",X"00",
		X"08",X"F0",X"00",X"EF",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"08",X"80",X"00",X"00",X"00",
		X"08",X"F8",X"00",X"00",X"80",X"00",X"00",X"00",X"0E",X"FF",X"00",X"00",X"00",X"00",X"0C",X"10",
		X"00",X"00",X"00",X"00",X"00",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"F5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"09",X"70",X"00",X"00",X"00",X"00",X"8F",X"00",
		X"07",X"17",X"97",X"67",X"76",X"00",X"8F",X"00",X"00",X"69",X"70",X"71",X"77",X"98",X"F8",X"00",
		X"00",X"06",X"96",X"67",X"97",X"7F",X"80",X"00",X"00",X"00",X"97",X"71",X"17",X"79",X"00",X"00",
		X"00",X"00",X"69",X"67",X"77",X"96",X"00",X"00",X"00",X"00",X"06",X"88",X"88",X"60",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"FF",X"E0",X"00",X"00",X"00",X"00",X"08",X"F8",X"EF",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"80",X"EF",X"80",X"00",X"00",X"00",X"00",X"EF",X"80",X"08",X"F8",X"00",X"00",
		X"00",X"00",X"8F",X"E0",X"00",X"8F",X"E0",X"00",X"00",X"00",X"8F",X"00",X"00",X"08",X"FE",X"00",
		X"00",X"00",X"F8",X"00",X"00",X"0E",X"88",X"00",X"00",X"00",X"FF",X"00",X"00",X"0E",X"EF",X"00",
		X"0C",X"10",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"7F",X"50",X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"00",X"09",X"70",X"00",X"00",X"00",X"00",
		X"8F",X"00",X"07",X"17",X"97",X"66",X"66",X"00",X"8F",X"00",X"00",X"69",X"76",X"71",X"17",X"98",
		X"F8",X"00",X"00",X"06",X"96",X"07",X"77",X"98",X"80",X"00",X"00",X"00",X"67",X"96",X"76",X"69",
		X"00",X"00",X"00",X"00",X"66",X"98",X"99",X"60",X"00",X"00",X"00",X"00",X"88",X"8E",X"88",X"00",
		X"00",X"00",X"00",X"0E",X"FF",X"00",X"F8",X"00",X"00",X"00",X"00",X"08",X"FE",X"08",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"F0",X"08",X"F0",X"00",X"00",X"00",X"00",X"08",X"F0",X"08",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"FE",X"00",X"00",X"00",X"00",X"0E",X"F0",X"00",X"88",X"00",
		X"00",X"00",X"00",X"08",X"F0",X"00",X"EF",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"0F",X"F0",
		X"00",X"00",X"0C",X"16",X"00",X"00",X"00",X"00",X"00",X"0E",X"88",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"7F",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"88",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"8F",X"00",X"09",X"19",X"69",X"70",
		X"00",X"00",X"8F",X"00",X"09",X"97",X"97",X"71",X"17",X"AA",X"8F",X"00",X"00",X"61",X"70",X"71",
		X"11",X"9A",X"FF",X"00",X"00",X"07",X"99",X"66",X"97",X"7F",X"F8",X"00",X"00",X"00",X"97",X"71",
		X"77",X"7F",X"80",X"00",X"00",X"00",X"67",X"1F",X"F7",X"76",X"00",X"00",X"00",X"00",X"06",X"8F",
		X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"0F",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",X"EF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"FE",X"F0",X"0D",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"7F",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"E0",X"00",X"00",X"69",X"77",X"79",X"96",X"00",X"EF",X"E0",X"00",X"09",X"61",X"19",X"77",
		X"79",X"9E",X"8F",X"00",X"00",X"00",X"66",X"07",X"17",X"77",X"98",X"F8",X"00",X"00",X"00",X"09",
		X"61",X"76",X"71",X"98",X"80",X"00",X"00",X"00",X"00",X"66",X"06",X"17",X"99",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"99",X"99",X"9E",X"00",X"00",X"00",X"00",X"00",X"E8",X"88",X"EE",X"8E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"00",X"4A",X"4F",X"55",X"53",X"54",
		X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",
		X"4E",X"43",X"2E",X"0D",X"09",X"07",X"96",X"00",X"00",X"00",X"00",X"8F",X"80",X"00",X"01",X"17",
		X"79",X"00",X"00",X"00",X"F7",X"F5",X"00",X"00",X"77",X"79",X"00",X"00",X"00",X"F8",X"00",X"00",
		X"00",X"11",X"79",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"07",X"77",X"90",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"01",X"17",X"97",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"77",X"77",X"79",
		X"08",X"C8",X"00",X"00",X"09",X"D7",X"60",X"7D",X"D7",X"9F",X"FE",X"00",X"00",X"09",X"69",X"96",
		X"6D",X"D6",X"9F",X"E0",X"00",X"00",X"00",X"00",X"99",X"96",X"69",X"98",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"99",X"99",X"9E",X"00",X"00",X"00",X"00",X"00",X"E8",X"88",X"EE",X"8E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"00",X"00",X"0C",X"10",X"00",X"8F",X"80",X"00",
		X"00",X"00",X"00",X"00",X"05",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"07",X"90",X"00",X"F8",X"00",X"66",
		X"66",X"79",X"71",X"70",X"00",X"EF",X"89",X"77",X"17",X"67",X"96",X"00",X"00",X"08",X"F7",X"79",
		X"70",X"69",X"60",X"00",X"00",X"00",X"97",X"77",X"69",X"79",X"00",X"00",X"00",X"00",X"06",X"99",
		X"89",X"66",X"00",X"00",X"00",X"00",X"00",X"88",X"E8",X"88",X"00",X"00",X"00",X"00",X"00",X"8F",
		X"00",X"8F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"80",X"FF",X"E0",X"00",X"00",X"00",X"00",X"08",
		X"FF",X"80",X"00",X"00",X"00",X"00",X"00",X"EF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"88",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"8E",X"00",X"00",X"00",X"03",X"10",X"08",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"5F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"00",X"00",
		X"00",X"F8",X"00",X"00",X"00",X"00",X"07",X"90",X"F8",X"00",X"66",X"66",X"79",X"71",X"70",X"8F",
		X"89",X"77",X"17",X"67",X"96",X"00",X"08",X"F7",X"79",X"70",X"69",X"60",X"00",X"00",X"77",X"11",
		X"99",X"79",X"00",X"00",X"00",X"69",X"77",X"79",X"96",X"00",X"00",X"00",X"06",X"88",X"88",X"60",
		X"00",X"00",X"00",X"00",X"8F",X"F0",X"00",X"00",X"00",X"00",X"00",X"E8",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"8F",X"F8",X"E0",X"00",X"00",X"00",X"8F",X"F0",X"8F",X"E0",X"00",X"00",X"00",X"FE",
		X"00",X"0F",X"80",X"00",X"00",X"08",X"80",X"00",X"0F",X"80",X"00",X"00",X"08",X"00",X"00",X"8F",
		X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"E0",X"00",X"00",X"03",X"10",X"08",X"F8",X"00",X"00",
		X"00",X"00",X"00",X"5F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"00",X"00",X"00",X"F8",
		X"00",X"00",X"00",X"00",X"07",X"90",X"F8",X"00",X"67",X"76",X"79",X"71",X"70",X"8F",X"89",X"77",
		X"17",X"07",X"96",X"00",X"08",X"F7",X"79",X"76",X"69",X"60",X"00",X"00",X"97",X"71",X"17",X"79",
		X"00",X"00",X"00",X"69",X"77",X"76",X"96",X"00",X"00",X"00",X"06",X"88",X"88",X"60",X"00",X"00",
		X"00",X"0E",X"FF",X"8F",X"00",X"00",X"00",X"00",X"00",X"FE",X"8F",X"80",X"00",X"00",X"00",X"08",
		X"FE",X"08",X"F0",X"00",X"00",X"00",X"8F",X"80",X"08",X"FE",X"00",X"00",X"0E",X"F8",X"00",X"0E",
		X"F8",X"00",X"00",X"EF",X"80",X"00",X"00",X"F8",X"00",X"00",X"88",X"E0",X"00",X"00",X"8F",X"00",
		X"00",X"FE",X"E0",X"00",X"00",X"FF",X"00",X"00",X"0C",X"10",X"00",X"8F",X"80",X"00",X"00",X"00",
		X"00",X"00",X"05",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",X"07",X"90",X"00",X"F8",X"00",X"66",X"66",X"79",
		X"71",X"70",X"00",X"8F",X"89",X"71",X"17",X"67",X"96",X"00",X"00",X"08",X"89",X"77",X"70",X"69",
		X"60",X"00",X"00",X"00",X"96",X"67",X"69",X"76",X"00",X"00",X"00",X"00",X"06",X"99",X"89",X"66",
		X"00",X"00",X"00",X"00",X"00",X"88",X"E8",X"88",X"00",X"00",X"00",X"00",X"00",X"8F",X"00",X"FF",
		X"E0",X"00",X"00",X"00",X"00",X"0F",X"80",X"EF",X"80",X"00",X"00",X"00",X"00",X"0F",X"80",X"0F",
		X"F0",X"00",X"00",X"00",X"00",X"0F",X"80",X"0F",X"80",X"00",X"00",X"00",X"00",X"EF",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"0F",X"E0",X"00",X"00",X"00",X"00",X"FE",X"00",X"0F",
		X"80",X"00",X"00",X"00",X"0F",X"F0",X"00",X"0F",X"80",X"00",X"0C",X"16",X"00",X"88",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"05",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",
		X"00",X"00",X"79",X"00",X"00",X"F8",X"00",X"00",X"07",X"96",X"91",X"90",X"00",X"F8",X"AA",X"71",
		X"17",X"79",X"79",X"90",X"00",X"FF",X"A9",X"11",X"17",X"07",X"16",X"00",X"00",X"8F",X"F7",X"79",
		X"66",X"99",X"70",X"00",X"00",X"08",X"F7",X"77",X"17",X"79",X"00",X"00",X"00",X"00",X"67",X"7F",
		X"F1",X"76",X"00",X"00",X"00",X"00",X"08",X"8F",X"F8",X"60",X"00",X"00",X"00",X"00",X"0E",X"8F",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"8F",X"80",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"EF",X"F0",X"00",X"00",X"00",X"00",X"00",X"0D",X"09",X"00",X"8F",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"F7",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FE",X"00",X"69",
		X"97",X"77",X"96",X"00",X"00",X"00",X"F8",X"E9",X"97",X"77",X"91",X"16",X"90",X"00",X"00",X"8F",
		X"89",X"77",X"71",X"70",X"66",X"00",X"00",X"00",X"08",X"89",X"17",X"67",X"16",X"90",X"00",X"00",
		X"00",X"00",X"99",X"71",X"60",X"66",X"00",X"00",X"00",X"00",X"00",X"E9",X"99",X"99",X"EE",X"00",
		X"00",X"00",X"00",X"00",X"E8",X"EE",X"88",X"8E",X"00",X"00",X"00",X"00",X"00",X"8E",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"09",X"00",X"08",X"F8",X"00",X"00",X"00",X"00",X"69",X"70",X"00",X"5F",
		X"7F",X"00",X"00",X"00",X"97",X"71",X"10",X"00",X"00",X"8F",X"00",X"00",X"00",X"97",X"77",X"00",
		X"00",X"00",X"8F",X"00",X"00",X"00",X"97",X"11",X"00",X"00",X"00",X"8F",X"00",X"00",X"09",X"77",
		X"70",X"00",X"00",X"00",X"8F",X"00",X"00",X"79",X"71",X"10",X"00",X"00",X"00",X"8C",X"80",X"97",
		X"77",X"77",X"00",X"00",X"00",X"00",X"EF",X"F9",X"7D",X"D7",X"06",X"7D",X"90",X"00",X"00",X"0E",
		X"F9",X"6D",X"D6",X"69",X"96",X"90",X"00",X"00",X"00",X"89",X"96",X"69",X"99",X"00",X"00",X"00",
		X"00",X"00",X"E9",X"99",X"99",X"EE",X"00",X"00",X"00",X"00",X"00",X"E8",X"EE",X"88",X"8E",X"00",
		X"00",X"00",X"00",X"00",X"8E",X"00",X"00",X"00",X"00",X"00",X"24",X"0A",X"00",X"F4",X"27",X"5A",
		X"24",X"B2",X"01",X"F4",X"2A",X"76",X"24",X"5E",X"00",X"F3",X"26",X"DA",X"25",X"06",X"00",X"F3",
		X"29",X"F6",X"24",X"5E",X"00",X"F3",X"25",X"5A",X"25",X"06",X"00",X"F3",X"28",X"92",X"24",X"5E",
		X"00",X"F3",X"25",X"DA",X"25",X"06",X"01",X"F3",X"29",X"12",X"24",X"5E",X"00",X"F3",X"26",X"5A",
		X"25",X"06",X"01",X"F3",X"29",X"84",X"24",X"5E",X"00",X"F3",X"26",X"DA",X"25",X"06",X"00",X"F3",
		X"29",X"F6",X"23",X"96",X"00",X"F2",X"27",X"D1",X"23",X"D2",X"00",X"F2",X"2A",X"E0",X"23",X"96",
		X"00",X"ED",X"27",X"D1",X"23",X"D2",X"00",X"ED",X"2A",X"E0",X"23",X"96",X"00",X"ED",X"28",X"1B",
		X"23",X"D2",X"00",X"ED",X"2B",X"2A",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",
		X"02",X"08",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"11",X"02",X"06",X"02",X"0A",X"02",X"05",
		X"02",X"0B",X"02",X"04",X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"04",X"02",X"0E",X"02",X"05",
		X"02",X"0D",X"02",X"05",X"02",X"0C",X"02",X"05",X"02",X"0D",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",
		X"02",X"0D",X"02",X"02",X"02",X"0D",X"02",X"09",X"02",X"0D",X"02",X"08",X"02",X"0E",X"02",X"05",
		X"02",X"0F",X"02",X"05",X"02",X"10",X"02",X"05",X"02",X"0F",X"02",X"06",X"02",X"0E",X"02",X"07",
		X"02",X"0E",X"02",X"06",X"02",X"0E",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"80",X"00",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",
		X"02",X"0A",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"0A",X"02",X"06",X"02",X"0B",X"02",X"05",
		X"02",X"0B",X"02",X"05",X"02",X"0B",X"02",X"03",X"02",X"0B",X"02",X"03",X"02",X"0B",X"02",X"03",
		X"02",X"0B",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"02",X"07",
		X"02",X"09",X"02",X"07",X"02",X"09",X"02",X"07",X"02",X"08",X"02",X"06",X"02",X"0A",X"02",X"06",
		X"02",X"11",X"02",X"07",X"02",X"0A",X"02",X"06",X"02",X"0E",X"02",X"05",X"02",X"0E",X"02",X"04",
		X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"03",X"02",X"0E",X"02",X"02",X"02",X"0E",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",
		X"02",X"0C",X"02",X"0B",X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"09",X"02",X"0D",X"02",X"09",
		X"02",X"0D",X"02",X"08",X"02",X"0D",X"02",X"08",X"02",X"0E",X"02",X"08",X"02",X"0E",X"02",X"08",
		X"02",X"10",X"02",X"08",X"02",X"10",X"02",X"08",X"02",X"10",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"02",X"0A",X"02",X"0C",X"02",X"0A",X"02",X"0C",X"02",X"0B",
		X"02",X"0C",X"02",X"09",X"02",X"0D",X"02",X"02",X"02",X"0D",X"02",X"09",X"02",X"0C",X"02",X"05",
		X"02",X"0D",X"02",X"05",X"02",X"0E",X"02",X"05",X"02",X"0F",X"02",X"05",X"02",X"10",X"02",X"05",
		X"02",X"10",X"02",X"05",X"02",X"11",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"0D",X"0A",X"00",X"00",X"00",X"B6",
		X"60",X"00",X"0F",X"F8",X"00",X"00",X"00",X"06",X"33",X"31",X"D0",X"0F",X"55",X"50",X"00",X"00",
		X"6B",X"33",X"3B",X"1B",X"0E",X"F0",X"50",X"00",X"0B",X"0B",X"BD",X"B1",X"1D",X"08",X"F0",X"00",
		X"00",X"B0",X"BB",X"32",X"BB",X"1F",X"FF",X"80",X"00",X"0B",X"6B",X"B3",X"33",X"BD",X"D8",X"F8",
		X"00",X"00",X"00",X"0B",X"3B",X"BB",X"88",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"FF",X"E0",X"00",X"00",X"00",X"0D",X"0A",X"00",X"00",X"0B",X"36",
		X"60",X"00",X"FF",X"80",X"00",X"00",X"00",X"6B",X"33",X"31",X"DE",X"F5",X"55",X"00",X"00",X"06",
		X"B3",X"33",X"BB",X"DE",X"EF",X"05",X"00",X"00",X"6B",X"0B",X"3D",X"B1",X"18",X"8F",X"00",X"00",
		X"00",X"B0",X"B3",X"32",X"3B",X"FF",X"FF",X"00",X"00",X"03",X"6B",X"B3",X"33",X"BD",X"8F",X"FE",
		X"00",X"00",X"00",X"0B",X"B3",X"8B",X"88",X"00",X"00",X"00",X"00",X"00",X"3B",X"3B",X"8F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"F0",X"FF",X"FF",X"80",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F8",X"00",X"00",X"00",
		X"00",X"0F",X"80",X"00",X"80",X"0F",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EF",X"FE",X"00",X"00",X"00",X"00",X"0D",X"0A",X"00",X"00",X"0B",X"36",
		X"60",X"00",X"FF",X"80",X"00",X"00",X"00",X"63",X"33",X"B1",X"DE",X"F5",X"55",X"00",X"00",X"06",
		X"BB",X"33",X"3D",X"DE",X"EF",X"05",X"00",X"00",X"6B",X"03",X"3D",X"B1",X"18",X"8F",X"00",X"00",
		X"00",X"B0",X"BB",X"23",X"BC",X"FF",X"FF",X"00",X"00",X"03",X"BB",X"B3",X"3B",X"BD",X"8F",X"FE",
		X"00",X"00",X"00",X"0B",X"33",X"8B",X"88",X"00",X"00",X"00",X"00",X"00",X"3B",X"3B",X"88",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"0F",X"FE",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"8F",
		X"E0",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"FE",X"00",X"00",X"8F",X"00",X"00",X"00",X"00",
		X"00",X"FE",X"00",X"00",X"08",X"F0",X"00",X"00",X"00",X"00",X"8F",X"80",X"00",X"0E",X"FF",X"00",
		X"00",X"00",X"00",X"EF",X"F8",X"00",X"08",X"08",X"F0",X"00",X"0D",X"0A",X"00",X"00",X"0B",X"36",
		X"60",X"00",X"0F",X"F8",X"00",X"00",X"00",X"63",X"33",X"31",X"D0",X"0F",X"55",X"50",X"00",X"06",
		X"B3",X"33",X"3B",X"1C",X"0E",X"F0",X"50",X"00",X"6B",X"03",X"3D",X"B1",X"1F",X"08",X"F0",X"00",
		X"00",X"B0",X"BB",X"32",X"BB",X"1F",X"FF",X"80",X"00",X"03",X"BB",X"BB",X"3B",X"BD",X"D8",X"F8",
		X"00",X"00",X"00",X"0B",X"33",X"8E",X"88",X"00",X"00",X"00",X"00",X"03",X"3B",X"EF",X"88",X"FE",
		X"00",X"00",X"00",X"00",X"0B",X"BE",X"F8",X"EF",X"80",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",
		X"0F",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"08",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"EF",X"FE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"00",X"00",X"00",X"0D",X"09",X"00",X"0B",X"22",X"36",
		X"00",X"0F",X"F8",X"00",X"00",X"00",X"32",X"33",X"BB",X"B0",X"0F",X"55",X"50",X"00",X"00",X"B0",
		X"30",X"66",X"6B",X"08",X"F0",X"50",X"00",X"00",X"00",X"0B",X"66",X"31",X"D0",X"88",X"00",X"00",
		X"00",X"BB",X"BB",X"B3",X"3B",X"1E",X"8F",X"00",X"00",X"03",X"30",X"BB",X"BD",X"31",X"1F",X"F8",
		X"00",X"00",X"06",X"3B",X"B3",X"32",X"BD",X"D8",X"E0",X"00",X"00",X"00",X"00",X"63",X"38",X"8D",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"FF",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E8",X"FE",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"E8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"8E",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"E8",X"EF",X"E8",
		X"00",X"0D",X"0C",X"00",X"00",X"06",X"B3",X"6B",X"60",X"00",X"00",X"00",X"00",X"00",X"62",X"63",
		X"36",X"B6",X"8F",X"80",X"00",X"00",X"0B",X"32",X"36",X"6B",X"B6",X"8F",X"55",X"00",X"00",X"63",
		X"3B",X"3B",X"BB",X"B3",X"88",X"05",X"00",X"00",X"33",X"33",X"B6",X"B3",X"BB",X"36",X"00",X"00",
		X"03",X"3B",X"0B",X"0B",X"30",X"33",X"B3",X"B0",X"00",X"00",X"6B",X"EE",X"E0",X"B3",X"03",X"30",
		X"33",X"00",X"00",X"00",X"E8",X"8E",X"0B",X"30",X"23",X"02",X"30",X"0D",X"09",X"03",X"03",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"20",X"3B",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"33",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"3B",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"30",X"BB",X"66",X"00",X"00",X"00",X"00",X"00",X"03",X"B3",X"3B",X"B6",X"BE",X"00",
		X"00",X"00",X"00",X"00",X"2B",X"33",X"B6",X"6B",X"BE",X"00",X"00",X"00",X"00",X"03",X"3B",X"BB",
		X"BB",X"DB",X"E8",X"F8",X"00",X"00",X"00",X"63",X"3B",X"BB",X"BD",X"88",X"F5",X"50",X"00",X"0B",
		X"06",X"36",X"B0",X"11",X"FF",X"E0",X"50",X"03",X"B3",X"B0",X"EE",X"BB",X"0D",X"8E",X"00",X"00",
		X"0B",X"B6",X"E8",X"8E",X"EE",X"8E",X"00",X"00",X"00",X"00",X"60",X"E8",X"EE",X"0E",X"00",X"80",
		X"00",X"00",X"0D",X"0A",X"00",X"8F",X"F0",X"00",X"06",X"6B",X"00",X"00",X"00",X"05",X"55",X"F0",
		X"0D",X"13",X"33",X"60",X"00",X"00",X"05",X"0F",X"E0",X"B1",X"B3",X"33",X"B6",X"00",X"00",X"00",
		X"0F",X"80",X"D1",X"1B",X"DB",X"B0",X"B0",X"00",X"00",X"08",X"FF",X"F1",X"BB",X"23",X"BB",X"0B",
		X"00",X"00",X"00",X"8F",X"8D",X"DB",X"33",X"3B",X"B6",X"B0",X"00",X"00",X"00",X"00",X"88",X"BB",
		X"B3",X"B0",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"8F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"8F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FF",X"E0",X"00",
		X"00",X"00",X"0C",X"0A",X"08",X"FF",X"00",X"06",X"63",X"B0",X"00",X"00",X"55",X"5F",X"ED",X"13",
		X"33",X"B6",X"00",X"00",X"50",X"FE",X"ED",X"BB",X"33",X"3B",X"60",X"00",X"00",X"F8",X"81",X"1B",
		X"D3",X"B0",X"B6",X"00",X"00",X"FF",X"FF",X"B3",X"23",X"3B",X"0B",X"00",X"00",X"EF",X"F8",X"DB",
		X"33",X"3B",X"B6",X"30",X"00",X"00",X"00",X"88",X"B8",X"3B",X"B0",X"00",X"00",X"00",X"00",X"0F",
		X"F8",X"B3",X"B3",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"BB",X"00",X"00",X"08",X"FF",X"FF",
		X"0F",X"F0",X"00",X"00",X"00",X"8F",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"08",X"00",
		X"08",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"EF",
		X"FE",X"00",X"00",X"00",X"0C",X"0A",X"08",X"FF",X"00",X"06",X"63",X"B0",X"00",X"00",X"55",X"5F",
		X"ED",X"1B",X"33",X"36",X"00",X"00",X"50",X"FE",X"ED",X"D3",X"33",X"BB",X"60",X"00",X"00",X"F8",
		X"81",X"1B",X"D3",X"30",X"B6",X"00",X"00",X"FF",X"FF",X"CB",X"32",X"BB",X"0B",X"00",X"00",X"EF",
		X"F8",X"DB",X"B3",X"3B",X"BB",X"30",X"00",X"00",X"00",X"88",X"B8",X"33",X"B0",X"00",X"00",X"00",
		X"00",X"8F",X"88",X"B3",X"B3",X"00",X"00",X"00",X"0E",X"FF",X"EF",X"F0",X"BB",X"00",X"00",X"00",
		X"0F",X"F0",X"0E",X"F8",X"00",X"00",X"00",X"00",X"F8",X"00",X"00",X"EF",X"00",X"00",X"00",X"0F",
		X"80",X"00",X"00",X"EF",X"00",X"00",X"00",X"FF",X"E0",X"00",X"08",X"F8",X"00",X"00",X"0F",X"80",
		X"80",X"00",X"8F",X"FE",X"00",X"00",X"0D",X"0A",X"00",X"8F",X"F0",X"00",X"06",X"63",X"B0",X"00",
		X"00",X"05",X"55",X"F0",X"0D",X"13",X"33",X"36",X"00",X"00",X"05",X"0F",X"E0",X"C1",X"B3",X"33",
		X"3B",X"60",X"00",X"00",X"0F",X"80",X"F1",X"1B",X"D3",X"30",X"B6",X"00",X"00",X"08",X"FF",X"F1",
		X"BB",X"23",X"BB",X"0B",X"00",X"00",X"00",X"8F",X"8D",X"DB",X"B3",X"BB",X"BB",X"30",X"00",X"00",
		X"00",X"00",X"88",X"E8",X"33",X"B0",X"00",X"00",X"00",X"00",X"00",X"EF",X"88",X"FE",X"B3",X"30",
		X"00",X"00",X"00",X"00",X"08",X"FE",X"8F",X"EB",X"B0",X"00",X"00",X"00",X"00",X"0E",X"F0",X"08",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"EF",X"FE",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"FF",X"08",X"00",X"00",X"00",X"00",X"0C",X"09",X"00",X"8F",X"F0",X"00",X"63",X"22",X"B0",X"00",
		X"05",X"55",X"F0",X"0B",X"BB",X"33",X"23",X"00",X"05",X"0F",X"80",X"B6",X"66",X"03",X"0B",X"00",
		X"00",X"88",X"0D",X"13",X"66",X"B0",X"00",X"00",X"00",X"F8",X"E1",X"B3",X"3B",X"BB",X"BB",X"00",
		X"00",X"8F",X"F1",X"13",X"DB",X"BB",X"03",X"30",X"00",X"0E",X"8D",X"DB",X"23",X"3B",X"B3",X"60",
		X"00",X"00",X"08",X"D8",X"83",X"36",X"00",X"00",X"00",X"00",X"8E",X"FF",X"8E",X"00",X"00",X"00",
		X"00",X"08",X"EF",X"8E",X"00",X"00",X"00",X"00",X"00",X"8E",X"8F",X"00",X"00",X"00",X"00",X"00",
		X"08",X"E8",X"F0",X"00",X"00",X"00",X"00",X"00",X"8E",X"FE",X"8E",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0C",X"00",X"00",X"00",X"06",X"B6",X"3B",X"60",X"00",X"00",X"00",X"08",X"F8",X"6B",X"63",
		X"36",X"26",X"00",X"00",X"00",X"55",X"F8",X"6B",X"B6",X"63",X"23",X"B0",X"00",X"00",X"50",X"88",
		X"3B",X"BB",X"B3",X"B3",X"36",X"00",X"00",X"00",X"63",X"BB",X"3B",X"6B",X"33",X"33",X"00",X"00",
		X"0B",X"3B",X"33",X"03",X"B0",X"B0",X"B3",X"30",X"00",X"33",X"03",X"30",X"3B",X"0E",X"EE",X"B6",
		X"00",X"03",X"20",X"32",X"03",X"B0",X"E8",X"8E",X"00",X"00",X"0D",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"30",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"B3",X"02",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"33",X"B0",X"00",X"00",X"00",X"00",X"00",X"0B",X"B3",X"30",X"20",
		X"00",X"00",X"00",X"00",X"00",X"66",X"BB",X"03",X"B0",X"00",X"00",X"00",X"00",X"EB",X"6B",X"B3",
		X"3B",X"30",X"00",X"00",X"00",X"EB",X"B6",X"6B",X"33",X"B2",X"00",X"00",X"8F",X"8E",X"BD",X"BB",
		X"BB",X"B3",X"30",X"00",X"05",X"5F",X"88",X"DB",X"BB",X"B3",X"36",X"00",X"00",X"05",X"0E",X"FF",
		X"11",X"0B",X"63",X"60",X"B0",X"00",X"00",X"00",X"E8",X"D0",X"BB",X"EE",X"0B",X"3B",X"30",X"00",
		X"00",X"00",X"E8",X"EE",X"E8",X"8E",X"6B",X"B0",X"00",X"00",X"08",X"00",X"E0",X"EE",X"8E",X"06",
		X"00",X"00",X"00",X"02",X"EF",X"2B",X"B9",X"00",X"00",X"00",X"EF",X"2B",X"EC",X"00",X"00",X"02",
		X"ED",X"2B",X"B9",X"00",X"00",X"00",X"ED",X"2B",X"EC",X"03",X"03",X"00",X"55",X"50",X"00",X"00",
		X"00",X"00",X"00",X"57",X"70",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",
		X"05",X"55",X"55",X"00",X"00",X"00",X"00",X"05",X"55",X"55",X"75",X"55",X"55",X"50",X"05",X"55",
		X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"03",X"03",X"00",X"00",
		X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"00",X"00",X"07",X"75",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"05",X"55",X"55",X"57",X"55",X"55",
		X"50",X"00",X"00",X"00",X"00",X"55",X"55",X"50",X"00",X"00",X"00",X"05",X"55",X"55",X"00",X"00",
		X"00",X"02",X"EF",X"2C",X"37",X"00",X"00",X"00",X"EF",X"2C",X"6A",X"00",X"00",X"02",X"ED",X"2C",
		X"37",X"00",X"00",X"00",X"ED",X"2C",X"6A",X"03",X"03",X"00",X"77",X"70",X"00",X"00",X"00",X"00",
		X"00",X"75",X"50",X"00",X"00",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"07",X"77",
		X"77",X"00",X"00",X"00",X"00",X"07",X"77",X"77",X"57",X"77",X"77",X"70",X"07",X"77",X"77",X"00",
		X"00",X"00",X"00",X"00",X"77",X"77",X"70",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",
		X"07",X"77",X"00",X"00",X"00",X"00",X"00",X"05",X"57",X"00",X"00",X"00",X"00",X"00",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"70",X"07",X"77",X"77",X"75",X"77",X"77",X"70",X"00",
		X"00",X"00",X"00",X"77",X"77",X"70",X"00",X"00",X"00",X"07",X"77",X"77",X"00",X"00",X"00",X"02",
		X"EF",X"2C",X"BB",X"00",X"00",X"00",X"EF",X"2C",X"EE",X"00",X"00",X"02",X"ED",X"2C",X"BB",X"00",
		X"00",X"00",X"ED",X"2C",X"EE",X"2F",X"95",X"00",X"F5",X"2D",X"21",X"03",X"03",X"00",X"44",X"40",
		X"00",X"00",X"00",X"00",X"00",X"49",X"90",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"04",X"41",X"11",X"11",X"11",X"11",X"10",
		X"04",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"03",X"03",
		X"00",X"00",X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"00",X"00",X"09",X"94",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"01",X"11",X"11",X"11",
		X"11",X"14",X"40",X"00",X"00",X"00",X"00",X"44",X"44",X"40",X"00",X"00",X"00",X"04",X"44",X"44",
		X"00",X"01",X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"E4",X"4E",X"01",X"00",X"00",X"49",X"9E",
		X"01",X"00",X"00",X"E4",X"4E",X"01",X"00",X"04",X"44",X"40",X"4D",X"00",X"4E",X"E4",X"40",X"44",
		X"00",X"00",X"E4",X"46",X"6D",X"00",X"00",X"44",X"4E",X"61",X"00",X"00",X"4E",X"E4",X"61",X"00",
		X"0E",X"4E",X"E4",X"61",X"00",X"08",X"80",X"04",X"81",X"00",X"88",X"80",X"E8",X"81",X"00",X"00",
		X"00",X"02",X"EF",X"2D",X"7D",X"00",X"00",X"00",X"EF",X"2D",X"D8",X"00",X"00",X"02",X"ED",X"2D",
		X"7D",X"00",X"00",X"00",X"ED",X"2D",X"D8",X"2F",X"95",X"00",X"F5",X"2E",X"0B",X"03",X"03",X"00",
		X"DD",X"D0",X"00",X"00",X"00",X"00",X"00",X"D4",X"40",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"0D",X"DD",X"DD",X"00",X"00",X"00",X"00",X"0D",X"D1",X"11",X"11",X"11",
		X"11",X"10",X"0D",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"DD",X"DD",X"D0",X"00",X"00",X"00",
		X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",
		X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"03",X"03",X"00",X"00",X"00",X"00",X"0D",X"DD",
		X"00",X"00",X"00",X"00",X"00",X"04",X"4D",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"DD",X"DD",X"D0",X"01",X"11",X"11",X"11",X"11",X"1D",X"D0",X"00",X"00",X"00",
		X"00",X"DD",X"DD",X"D0",X"00",X"00",X"00",X"0D",X"DD",X"DD",X"00",X"01",X"08",X"00",X"00",X"00",
		X"01",X"00",X"00",X"9D",X"D9",X"01",X"00",X"00",X"D4",X"4E",X"01",X"00",X"00",X"ED",X"D6",X"01",
		X"00",X"0D",X"DD",X"D9",X"DA",X"00",X"D9",X"6D",X"D9",X"DD",X"00",X"00",X"6D",X"D6",X"6A",X"00",
		X"00",X"DD",X"DE",X"61",X"00",X"00",X"D9",X"9D",X"61",X"00",X"09",X"DE",X"ED",X"61",X"00",X"03",
		X"30",X"0D",X"31",X"00",X"33",X"30",X"93",X"31",X"00",X"00",X"00",X"02",X"EF",X"2E",X"67",X"00",
		X"00",X"00",X"EF",X"2E",X"9A",X"00",X"00",X"02",X"ED",X"2E",X"67",X"00",X"00",X"00",X"ED",X"2E",
		X"9A",X"2F",X"95",X"00",X"F5",X"2E",X"CD",X"03",X"03",X"00",X"99",X"90",X"00",X"00",X"00",X"00",
		X"00",X"95",X"50",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"09",X"99",
		X"99",X"00",X"00",X"00",X"00",X"09",X"91",X"11",X"11",X"11",X"11",X"10",X"09",X"99",X"99",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",
		X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"05",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"01",X"11",X"11",X"11",X"11",X"19",X"90",X"00",
		X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"01",X"08",X"00",
		X"00",X"00",X"01",X"00",X"00",X"E9",X"9E",X"01",X"00",X"00",X"95",X"5E",X"01",X"00",X"00",X"E9",
		X"9E",X"01",X"00",X"09",X"99",X"90",X"9D",X"00",X"9E",X"E9",X"90",X"99",X"00",X"00",X"E9",X"96",
		X"6D",X"00",X"00",X"99",X"9E",X"61",X"00",X"00",X"96",X"69",X"61",X"00",X"0E",X"9E",X"E9",X"61",
		X"00",X"03",X"30",X"09",X"31",X"00",X"33",X"30",X"E3",X"31",X"00",X"2F",X"35",X"00",X"FA",X"2F",
		X"C5",X"2F",X"55",X"00",X"FB",X"2F",X"FD",X"2F",X"75",X"00",X"FB",X"2F",X"E3",X"2F",X"35",X"00",
		X"FB",X"30",X"17",X"2F",X"95",X"FF",X"F6",X"30",X"37",X"2F",X"95",X"FE",X"F5",X"30",X"91",X"2F",
		X"95",X"00",X"F5",X"2E",X"0B",X"02",X"03",X"02",X"06",X"02",X"02",X"02",X"07",X"02",X"02",X"02",
		X"07",X"02",X"02",X"02",X"07",X"02",X"02",X"02",X"07",X"02",X"02",X"02",X"07",X"02",X"03",X"02",
		X"06",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"02",X"02",X"02",X"06",X"02",X"01",X"02",
		X"07",X"02",X"01",X"02",X"07",X"02",X"01",X"02",X"07",X"02",X"02",X"02",X"07",X"02",X"03",X"02",
		X"06",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"02",X"03",X"02",X"06",X"02",X"02",X"02",
		X"07",X"02",X"01",X"02",X"07",X"02",X"01",X"02",X"07",X"02",X"01",X"02",X"06",X"02",X"02",X"02",
		X"05",X"81",X"00",X"81",X"00",X"02",X"03",X"02",X"06",X"02",X"03",X"02",X"06",X"02",X"03",X"02",
		X"06",X"02",X"02",X"02",X"04",X"02",X"01",X"02",X"04",X"02",X"03",X"02",X"08",X"02",X"03",X"02",
		X"08",X"02",X"03",X"02",X"06",X"02",X"03",X"02",X"06",X"02",X"02",X"02",X"07",X"02",X"01",X"02",
		X"08",X"81",X"00",X"81",X"00",X"00",X"03",X"00",X"B2",X"2B",X"00",X"0B",X"21",X"12",X"B0",X"02",
		X"11",X"11",X"20",X"02",X"15",X"15",X"20",X"02",X"51",X"55",X"20",X"03",X"25",X"52",X"30",X"00",
		X"32",X"23",X"00",X"00",X"02",X"00",X"25",X"52",X"00",X"02",X"51",X"15",X"B0",X"32",X"11",X"11",
		X"30",X"35",X"11",X"52",X"B0",X"B2",X"55",X"23",X"00",X"0B",X"33",X"30",X"00",X"00",X"02",X"02",
		X"55",X"20",X"00",X"B5",X"11",X"52",X"00",X"31",X"11",X"12",X"30",X"B2",X"51",X"15",X"30",X"03",
		X"25",X"52",X"B0",X"00",X"33",X"3B",X"00",X"01",X"02",X"02",X"00",X"63",X"53",X"00",X"25",X"36",
		X"4E",X"52",X"30",X"51",X"5E",X"63",X"51",X"30",X"21",X"52",X"E2",X"15",X"30",X"32",X"12",X"35",
		X"22",X"00",X"0B",X"22",X"32",X"3B",X"00",X"0C",X"0F",X"00",X"00",X"63",X"36",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B6",X"46",X"00",X"00",X"00",X"00",X"55",X"00",X"B3",X"3E",X"00",X"00",X"00",
		X"00",X"32",X"03",X"33",X"E0",X"80",X"00",X"05",X"00",X"00",X"B0",X"E3",X"B0",X"00",X"00",X"23",
		X"00",X"00",X"00",X"0B",X"B3",X"35",X"30",X"00",X"00",X"02",X"30",X"06",X"6E",X"31",X"30",X"00",
		X"00",X"01",X"03",X"36",X"63",X"23",X"00",X"00",X"00",X"01",X"15",X"36",X"E0",X"00",X"00",X"05",
		X"00",X"02",X"11",X"23",X"E0",X"21",X"03",X"11",X"00",X"00",X"22",X"22",X"E2",X"12",X"33",X"23",
		X"00",X"0E",X"08",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"15",X"00",X"00",
		X"6D",X"D6",X"01",X"00",X"00",X"00",X"00",X"32",X"00",X"00",X"34",X"43",X"01",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"ED",X"D3",X"01",X"00",X"00",X"52",X"00",X"00",X"00",X"03",X"3D",X"D0",
		X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"DE",X"63",X"D0",X"2D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"63",X"36",X"6D",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"32",X"3E",X"61",X"00",
		X"00",X"00",X"00",X"03",X"20",X"00",X"D6",X"63",X"61",X"00",X"00",X"01",X"00",X"00",X"00",X"03",
		X"3E",X"E2",X"61",X"00",X"00",X"12",X"00",X"00",X"00",X"03",X"30",X"03",X"31",X"00",X"00",X"00",
		X"00",X"00",X"00",X"33",X"30",X"E3",X"31",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"31",
		X"2F",X"00",X"00",X"00",X"F8",X"31",X"43",X"00",X"00",X"00",X"F8",X"31",X"69",X"00",X"00",X"00",
		X"F2",X"31",X"A1",X"00",X"00",X"00",X"F0",X"31",X"FD",X"00",X"00",X"00",X"EF",X"32",X"76",X"07",
		X"02",X"44",X"8E",X"00",X"0E",X"44",X"E0",X"00",X"04",X"80",X"00",X"0E",X"40",X"00",X"00",X"40",
		X"00",X"00",X"40",X"00",X"0D",X"00",X"00",X"0C",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"44",
		X"00",X"00",X"0E",X"44",X"00",X"0E",X"44",X"4E",X"00",X"E4",X"44",X"E0",X"00",X"44",X"E0",X"00",
		X"00",X"48",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"02",X"0D",X"00",X"00",X"00",X"40",X"04",
		X"00",X"00",X"04",X"00",X"40",X"04",X"E0",X"00",X"04",X"0E",X"40",X"E4",X"E0",X"00",X"04",X"4C",
		X"C4",X"44",X"00",X"00",X"04",X"4A",X"CC",X"4E",X"00",X"00",X"E4",X"AA",X"44",X"E0",X"00",X"00",
		X"4A",X"A4",X"E0",X"00",X"00",X"04",X"A8",X"E0",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"00",
		X"00",X"02",X"0B",X"00",X"00",X"A0",X"00",X"80",X"00",X"00",X"00",X"A0",X"0E",X"A0",X"00",X"08",
		X"00",X"A8",X"0A",X"80",X"00",X"EA",X"0E",X"A8",X"8A",X"80",X"A0",X"AA",X"08",X"AA",X"AA",X"0A",
		X"A0",X"CA",X"0A",X"AA",X"A8",X"8A",X"80",X"8C",X"AA",X"AA",X"AA",X"AC",X"00",X"EC",X"AA",X"AA",
		X"AC",X"4E",X"00",X"08",X"CA",X"CA",X"A4",X"E0",X"00",X"0E",X"4C",X"AC",X"4E",X"00",X"00",X"00",
		X"4C",X"C4",X"E0",X"00",X"00",X"00",X"44",X"4E",X"00",X"00",X"00",X"0E",X"44",X"E0",X"00",X"00",
		X"00",X"E4",X"4E",X"00",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"00",X"00",X"03",X"15",X"00",
		X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"0E",X"80",X"0A",X"00",X"00",X"00",X"00",X"0E",
		X"E0",X"8E",X"0E",X"E0",X"0A",X"00",X"08",X"EE",X"80",X"08",X"80",X"E8",X"00",X"E8",X"08",X"80",
		X"88",X"00",X"88",X"00",X"EA",X"A8",X"E8",X"80",X"00",X"EA",X"80",X"88",X"5F",X"AA",X"0E",X"80",
		X"0A",X"AF",X"FE",X"8F",X"5E",X"88",X"E0",X"0E",X"A8",X"F8",X"AA",X"AA",X"80",X"00",X"08",X"AA",
		X"8A",X"AA",X"E8",X"00",X"00",X"0E",X"88",X"8F",X"5F",X"80",X"00",X"00",X"00",X"8A",X"A5",X"FA",
		X"E0",X"00",X"00",X"08",X"8E",X"8A",X"8E",X"00",X"00",X"00",X"04",X"AA",X"8E",X"E0",X"00",X"00",
		X"00",X"E4",X"C4",X"CE",X"00",X"00",X"00",X"00",X"84",X"48",X"E0",X"00",X"00",X"00",X"00",X"48",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"03",X"16",X"00",X"00",X"00",X"00",X"AA",X"F0",X"00",X"00",
		X"00",X"00",X"8A",X"88",X"E8",X"80",X"00",X"00",X"0E",X"F8",X"EA",X"EA",X"A0",X"00",X"00",X"0F",
		X"AE",X"08",X"88",X"E0",X"00",X"00",X"AF",X"AE",X"8A",X"AF",X"F0",X"00",X"0E",X"AA",X"EE",X"EE",
		X"08",X"80",X"00",X"08",X"88",X"8E",X"8A",X"FF",X"80",X"00",X"EA",X"FE",X"A8",X"E0",X"88",X"00",
		X"0E",X"8F",X"88",X"FA",X"0F",X"08",X"00",X"08",X"4A",X"88",X"8E",X"81",X"E0",X"00",X"04",X"A4",
		X"8E",X"08",X"F1",X"E0",X"00",X"04",X"A8",X"E0",X"0F",X"8F",X"E0",X"00",X"04",X"CE",X"00",X"0F",
		X"EF",X"E0",X"00",X"08",X"CE",X"00",X"00",X"F8",X"E0",X"00",X"0E",X"48",X"00",X"00",X"00",X"00",
		X"00",X"00",X"48",X"00",X"00",X"00",X"00",X"00",X"04",X"4E",X"00",X"00",X"00",X"00",X"00",X"48",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"33",X"0E",X"00",X"00",X"00",X"F1",
		X"33",X"4C",X"00",X"00",X"00",X"F1",X"33",X"8E",X"00",X"00",X"00",X"F5",X"33",X"E0",X"00",X"0B",
		X"00",X"00",X"40",X"00",X"00",X"0E",X"44",X"00",X"00",X"04",X"C4",X"00",X"00",X"04",X"A8",X"00",
		X"00",X"08",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"80",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"E4",X"40",X"00",X"00",X"E4",X"C4",X"00",
		X"00",X"8C",X"5A",X"E0",X"0E",X"CA",X"55",X"C0",X"E4",X"A5",X"55",X"A0",X"00",X"14",X"00",X"0E",
		X"4E",X"00",X"00",X"0E",X"44",X"00",X"00",X"00",X"4A",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"EE",X"00",X"00",X"0E",X"48",
		X"E0",X"00",X"0E",X"44",X"80",X"00",X"00",X"44",X"CE",X"00",X"00",X"4C",X"A8",X"00",X"00",X"4A",
		X"5C",X"00",X"0E",X"C5",X"5C",X"00",X"08",X"A5",X"5C",X"00",X"4A",X"55",X"5A",X"00",X"01",X"14",
		X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"00",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",
		X"00",X"40",X"00",X"0E",X"44",X"0E",X"40",X"00",X"04",X"4E",X"0C",X"40",X"00",X"04",X"C0",X"4A",
		X"80",X"00",X"0C",X"54",X"C8",X"E0",X"00",X"0A",X"5A",X"C4",X"00",X"00",X"0A",X"55",X"C4",X"00",
		X"00",X"05",X"55",X"A8",X"00",X"00",X"05",X"55",X"A8",X"00",X"00",X"4A",X"55",X"A8",X"00",X"00",
		X"00",X"08",X"00",X"00",X"04",X"00",X"00",X"04",X"44",X"00",X"00",X"4C",X"48",X"00",X"0E",X"CA",
		X"40",X"00",X"04",X"AE",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"84",X"80",
		X"00",X"00",X"4C",X"CE",X"00",X"00",X"4A",X"5C",X"E0",X"00",X"45",X"55",X"A0",X"00",X"4A",X"55",
		X"AE",X"00",X"00",X"00",X"01",X"E8",X"34",X"24",X"00",X"00",X"01",X"E2",X"34",X"35",X"00",X"00",
		X"00",X"DD",X"34",X"64",X"07",X"01",X"00",X"04",X"00",X"00",X"44",X"40",X"04",X"41",X"44",X"00",
		X"44",X"40",X"00",X"04",X"00",X"01",X"0D",X"00",X"00",X"70",X"00",X"00",X"07",X"00",X"70",X"07",
		X"00",X"00",X"70",X"00",X"70",X"00",X"00",X"05",X"05",X"00",X"00",X"77",X"00",X"00",X"07",X"70",
		X"00",X"05",X"05",X"00",X"00",X"00",X"70",X"00",X"70",X"00",X"07",X"00",X"70",X"07",X"00",X"00",
		X"00",X"70",X"00",X"00",X"02",X"0F",X"00",X"07",X"00",X"07",X"00",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"07",X"01",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"70",X"71",X"00",X"01",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"01",X"07",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"07",X"00",X"07",X"00",X"00",X"34",X"CC",X"01",X"F5",X"36",X"04",X"35",X"68",
		X"01",X"F5",X"37",X"8C",X"35",X"00",X"01",X"F9",X"36",X"88",X"35",X"9C",X"00",X"F9",X"38",X"10",
		X"35",X"34",X"00",X"F6",X"36",X"E5",X"35",X"D0",X"00",X"F6",X"38",X"74",X"80",X"00",X"80",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"02",X"09",X"02",X"0E",
		X"02",X"09",X"02",X"16",X"02",X"05",X"02",X"1A",X"02",X"03",X"02",X"18",X"02",X"05",X"02",X"15",
		X"02",X"08",X"02",X"0F",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"02",X"14",X"02",X"18",X"02",X"0A",X"02",X"1B",X"02",X"07",X"02",X"19",X"02",X"05",X"02",X"19",
		X"02",X"07",X"02",X"1A",X"02",X"05",X"02",X"15",X"02",X"03",X"02",X"07",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"02",X"1B",X"02",X"1C",X"02",X"17",X"02",X"1B",
		X"02",X"16",X"02",X"1A",X"02",X"14",X"02",X"19",X"02",X"09",X"02",X"1B",X"02",X"06",X"02",X"19",
		X"02",X"04",X"02",X"1A",X"02",X"06",X"02",X"15",X"02",X"08",X"02",X"10",X"02",X"05",X"02",X"0C",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"02",X"0F",X"02",X"14",X"02",X"07",X"02",X"14",
		X"02",X"03",X"02",X"18",X"02",X"05",X"02",X"1A",X"02",X"08",X"02",X"18",X"02",X"0E",X"02",X"15",
		X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",X"80",X"00",X"80",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"02",X"05",X"02",X"09",
		X"02",X"02",X"02",X"13",X"02",X"04",X"02",X"16",X"02",X"04",X"02",X"18",X"02",X"03",X"02",X"16",
		X"02",X"0C",X"02",X"18",X"02",X"16",X"02",X"1A",X"81",X"00",X"81",X"00",X"81",X"00",X"81",X"00",
		X"80",X"00",X"80",X"00",X"02",X"01",X"02",X"02",X"02",X"02",X"02",X"06",X"02",X"03",X"02",X"07",
		X"02",X"04",X"02",X"09",X"02",X"02",X"02",X"14",X"02",X"04",X"02",X"17",X"02",X"03",X"02",X"19",
		X"02",X"08",X"02",X"17",X"02",X"0D",X"02",X"15",X"02",X"11",X"02",X"18",X"81",X"00",X"81",X"00",
		X"81",X"00",X"81",X"00",X"09",X"0E",X"99",X"99",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"44",X"F7",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"CF",X"79",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"44",X"FF",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"4F",X"79",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"94",X"CF",X"70",X"00",X"0D",X"1F",
		X"FD",X"00",X"00",X"00",X"00",X"99",X"44",X"88",X"F4",X"14",X"90",X"00",X"04",X"00",X"D1",X"1F",
		X"00",X"99",X"64",X"8C",X"FF",X"CC",X"C5",X"FF",X"CA",X"88",X"FF",X"DD",X"00",X"00",X"00",X"99",
		X"44",X"CD",X"FF",X"88",X"4F",X"FC",X"34",X"E0",X"00",X"00",X"00",X"00",X"00",X"09",X"44",X"48",
		X"86",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"1F",X"FD",X"00",X"00",X"00",X"00",X"00",X"06",X"36",X"9F",X"F1",X"90",X"00",
		X"04",X"00",X"11",X"10",X"00",X"00",X"69",X"94",X"9F",X"FC",X"F9",X"A0",X"00",X"EC",X"8F",X"80",
		X"00",X"00",X"69",X"4E",X"94",X"FC",X"D8",X"E8",X"9C",X"9F",X"FD",X"C9",X"F0",X"00",X"00",X"00",
		X"94",X"FC",X"99",X"6E",X"98",X"AD",X"CF",X"8E",X"00",X"ED",X"00",X"00",X"94",X"DD",X"66",X"0E",
		X"E6",X"88",X"E0",X"00",X"00",X"00",X"00",X"00",X"94",X"F4",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FD",X"ED",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"14",X"F1",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"69",X"86",X"00",X"00",X"00",X"0F",X"DC",X"E8",
		X"40",X"00",X"00",X"00",X"06",X"99",X"AA",X"AC",X"FC",X"A6",X"00",X"00",X"CD",X"43",X"F0",X"00",
		X"00",X"00",X"06",X"94",X"84",X"C3",X"FF",X"F1",X"8A",X"CD",X"FF",X"D8",X"00",X"ED",X"00",X"00",
		X"00",X"00",X"06",X"64",X"6F",X"FC",X"F9",X"8C",X"DC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"4C",X"78",X"66",X"8E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"4C",X"AA",X"F7",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"44",X"CA",
		X"AA",X"FF",X"D7",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"7F",X"44",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"FC",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FF",X"44",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"97",X"F4",X"49",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DF",X"F1",X"D0",X"00",X"07",X"FC",X"49",X"00",X"00",X"00",X"00",X"F1",X"1D",X"00",X"40",
		X"00",X"09",X"41",X"4F",X"88",X"44",X"99",X"00",X"00",X"00",X"DD",X"FF",X"88",X"AC",X"FF",X"5C",
		X"CC",X"FF",X"C8",X"46",X"99",X"00",X"00",X"00",X"0E",X"43",X"CF",X"F4",X"88",X"FF",X"DC",X"44",
		X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"68",X"84",X"44",X"90",X"00",X"00",X"00",
		X"0A",X"03",X"00",X"00",X"DF",X"F1",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"11",X"00",X"40",X"00",X"09",X"1F",X"F9",X"63",X"60",X"00",X"00",X"00",X"00",X"00",X"08",
		X"F8",X"CE",X"00",X"0A",X"9F",X"CF",X"F9",X"49",X"96",X"00",X"00",X"00",X"00",X"0F",X"9C",X"DF",
		X"F9",X"C9",X"8E",X"8D",X"CF",X"49",X"E4",X"96",X"00",X"00",X"00",X"DE",X"00",X"E8",X"FC",X"DA",
		X"89",X"E6",X"99",X"CF",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"88",X"6E",
		X"E0",X"66",X"DD",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"4F",X"49",X"00",X"0B",X"0F",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"DE",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FD",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"1F",X"41",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"8E",X"CD",X"F0",X"00",X"00",X"00",X"68",X"96",X"36",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"34",X"DC",X"00",X"00",X"6A",X"CF",X"CA",X"AA",X"99",X"60",X"00",X"00",X"00",
		X"00",X"DE",X"00",X"8D",X"FF",X"DC",X"A8",X"1F",X"FF",X"3C",X"48",X"49",X"60",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"8F",X"CD",X"C8",X"9F",X"CF",X"F6",X"46",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E8",X"66",X"87",X"C4",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"AA",X"C4",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0D",X"7D",X"FF",X"AA",X"AC",X"44",X"99",X"00",X"D0",X"1C",X"01",X"B0",X"2C",
		X"14",X"01",X"C0",X"14",X"01",X"B0",X"14",X"1C",X"01",X"40",X"34",X"30",X"24",X"1C",X"1C",X"01",
		X"30",X"14",X"3C",X"14",X"20",X"14",X"2C",X"01",X"20",X"24",X"2C",X"34",X"2C",X"10",X"14",X"01",
		X"30",X"34",X"5C",X"01",X"30",X"24",X"3C",X"01",X"20",X"2C",X"01",X"24",X"5C",X"00",X"D0",X"14",
		X"01",X"B0",X"24",X"1E",X"01",X"C0",X"2E",X"01",X"B0",X"1E",X"14",X"01",X"40",X"3E",X"30",X"2E",
		X"1E",X"14",X"01",X"30",X"2E",X"24",X"1E",X"20",X"1E",X"24",X"01",X"20",X"3E",X"14",X"2E",X"10",
		X"1E",X"14",X"2E",X"01",X"30",X"1E",X"10",X"2E",X"24",X"24",X"01",X"30",X"1E",X"2E",X"24",X"01",
		X"20",X"3E",X"14",X"01",X"3E",X"24",X"24",X"00",X"E0",X"01",X"B0",X"1E",X"14",X"1E",X"01",X"C0",
		X"2E",X"01",X"B0",X"1E",X"1E",X"01",X"40",X"2E",X"40",X"2E",X"1E",X"1E",X"01",X"30",X"1E",X"10",
		X"1E",X"14",X"1E",X"20",X"1E",X"14",X"1E",X"01",X"30",X"2E",X"10",X"1E",X"20",X"1E",X"10",X"2E",
		X"01",X"50",X"2E",X"1E",X"14",X"1E",X"14",X"01",X"40",X"2E",X"1E",X"14",X"01",X"20",X"2E",X"1E",
		X"01",X"1E",X"2E",X"20",X"1E",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"3D",X"36",X"7E",X"3D",X"AF",X"7E",X"3B",X"CF",X"7E",X"3C",X"57",X"7E",X"3F",X"C1",X"7E",
		X"3E",X"09",X"7E",X"3D",X"E9",X"7E",X"3D",X"BD",X"7E",X"41",X"16",X"7E",X"41",X"10",X"7E",X"40",
		X"BC",X"7E",X"40",X"E1",X"7E",X"40",X"F2",X"7E",X"40",X"F0",X"7E",X"40",X"FA",X"7E",X"41",X"08",
		X"7E",X"41",X"06",X"7E",X"41",X"4F",X"7E",X"42",X"E7",X"7E",X"43",X"09",X"7E",X"43",X"03",X"7E",
		X"42",X"FD",X"7E",X"43",X"65",X"7E",X"43",X"7B",X"7E",X"43",X"90",X"7E",X"43",X"F6",X"7E",X"44",
		X"D4",X"7E",X"46",X"4F",X"0D",X"F5",X"27",X"5A",X"CC",X"00",X"40",X"BD",X"E0",X"0C",X"86",X"04",
		X"BD",X"E0",X"37",X"34",X"01",X"1A",X"FF",X"CC",X"9C",X"D7",X"FD",X"CA",X"06",X"4F",X"5F",X"FD",
		X"CA",X"04",X"B7",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",X"35",X"01",X"8E",X"39",X"20",X"86",
		X"69",X"C6",X"11",X"BD",X"4A",X"53",X"8E",X"14",X"CA",X"86",X"6B",X"C6",X"99",X"BD",X"4A",X"5C",
		X"BE",X"5E",X"DB",X"BD",X"E0",X"2D",X"6F",X"C8",X"32",X"86",X"1E",X"BD",X"E0",X"37",X"6A",X"C8",
		X"32",X"27",X"0F",X"AE",X"C4",X"A6",X"02",X"81",X"41",X"27",X"EE",X"81",X"42",X"27",X"EA",X"7E",
		X"5E",X"D3",X"CC",X"42",X"FF",X"BD",X"E0",X"0C",X"86",X"03",X"BD",X"E0",X"37",X"20",X"F0",X"34",
		X"02",X"A6",X"80",X"1E",X"12",X"BD",X"40",X"FA",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",X"8E",
		X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",X"36",X"8E",X"3C",X"11",X"10",
		X"8E",X"CC",X"00",X"C6",X"12",X"8D",X"D8",X"35",X"B6",X"34",X"36",X"8E",X"3C",X"23",X"10",X"8E",
		X"CC",X"24",X"C6",X"34",X"8D",X"C9",X"BD",X"3D",X"0F",X"8E",X"CC",X"8E",X"BD",X"40",X"FA",X"35",
		X"B6",X"20",X"05",X"01",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"05",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"1A",X"1C",X"0F",X"1D",X"0F",X"18",
		X"1E",X"0F",X"0E",X"0A",X"0C",X"23",X"32",X"0A",X"0A",X"0A",X"0A",X"0A",X"21",X"13",X"16",X"16",
		X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",
		X"0A",X"13",X"18",X"0D",X"2E",X"25",X"29",X"BD",X"3C",X"F6",X"BD",X"40",X"BC",X"B6",X"C8",X"0C",
		X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1B",X"84",X"0F",X"27",X"11",X"7F",X"CC",X"1B",X"BD",X"3C",
		X"F6",X"BD",X"40",X"BC",X"BD",X"3D",X"98",X"86",X"40",X"BD",X"F0",X"09",X"B6",X"CC",X"1D",X"84",
		X"0F",X"27",X"0D",X"7F",X"CC",X"1D",X"8D",X"6E",X"BD",X"3B",X"1F",X"86",X"40",X"BD",X"F0",X"09",
		X"B6",X"CC",X"21",X"84",X"0F",X"27",X"1F",X"7F",X"CC",X"21",X"8D",X"5A",X"BD",X"40",X"BC",X"86",
		X"0A",X"BD",X"4A",X"62",X"BD",X"45",X"57",X"B6",X"00",X"20",X"BD",X"F0",X"09",X"BD",X"3D",X"0F",
		X"8E",X"CC",X"8E",X"BD",X"40",X"FA",X"B6",X"CC",X"23",X"84",X"0F",X"27",X"13",X"7F",X"CC",X"23",
		X"8D",X"34",X"BD",X"40",X"BC",X"86",X"10",X"BD",X"4A",X"62",X"BD",X"43",X"A7",X"BD",X"3F",X"88",
		X"B6",X"CC",X"1F",X"84",X"0F",X"27",X"0A",X"7F",X"CC",X"1F",X"8D",X"1A",X"8D",X"07",X"7E",X"F0",
		X"06",X"8D",X"02",X"20",X"51",X"B6",X"CC",X"19",X"84",X"0F",X"27",X"09",X"7C",X"CC",X"8C",X"7C",
		X"CC",X"8C",X"7F",X"CC",X"19",X"39",X"34",X"12",X"8D",X"08",X"8E",X"CC",X"8C",X"BD",X"40",X"FA",
		X"35",X"92",X"34",X"34",X"8E",X"CC",X"00",X"10",X"8E",X"CC",X"24",X"8D",X"09",X"35",X"B4",X"8E",
		X"CC",X"24",X"10",X"8E",X"CC",X"8C",X"10",X"9F",X"D5",X"4F",X"E6",X"80",X"C4",X"0F",X"34",X"04",
		X"AB",X"E0",X"9C",X"D5",X"26",X"F4",X"8B",X"37",X"39",X"8D",X"D7",X"34",X"02",X"8E",X"CC",X"8C",
		X"BD",X"40",X"E1",X"A1",X"E0",X"39",X"8D",X"70",X"8D",X"EF",X"27",X"3D",X"86",X"39",X"B7",X"CB",
		X"FF",X"BD",X"3B",X"EA",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"AB",X"86",X"39",X"B7",X"CB",X"FF",
		X"BD",X"40",X"BC",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"28",X"BD",X"3B",X"22",X"BD",X"3B",X"1C",
		X"8D",X"C7",X"27",X"1A",X"86",X"0B",X"BD",X"4A",X"62",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",
		X"0C",X"85",X"02",X"27",X"F4",X"6E",X"9F",X"EF",X"FE",X"BD",X"3B",X"1C",X"20",X"F7",X"86",X"0C",
		X"20",X"E4",X"8E",X"CD",X"02",X"C6",X"04",X"A6",X"80",X"84",X"0F",X"81",X"09",X"23",X"03",X"5A",
		X"27",X"06",X"8C",X"CD",X"3E",X"26",X"F0",X"39",X"86",X"0D",X"BD",X"4A",X"62",X"8E",X"CD",X"02",
		X"6F",X"80",X"8C",X"CD",X"3E",X"26",X"F9",X"39",X"8D",X"05",X"27",X"FB",X"7E",X"3B",X"F9",X"BD",
		X"3D",X"0F",X"34",X"02",X"8E",X"CC",X"8E",X"BD",X"40",X"E1",X"A1",X"E0",X"39",X"86",X"18",X"97",
		X"E2",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"08",X"BD",X"F0",X"09",X"B6",X"C8",X"0C",X"85",X"08",
		X"27",X"16",X"0A",X"E2",X"26",X"F0",X"10",X"8E",X"CD",X"3E",X"8E",X"3E",X"42",X"C6",X"17",X"BD",
		X"3B",X"16",X"BD",X"3F",X"88",X"7F",X"C8",X"0E",X"39",X"10",X"8E",X"CD",X"74",X"C6",X"08",X"BD",
		X"3F",X"AF",X"A8",X"26",X"84",X"0F",X"27",X"03",X"5A",X"27",X"0E",X"86",X"39",X"B7",X"CB",X"FF",
		X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"E7",X"39",X"86",X"39",X"B7",X"CB",X"FF",X"8E",X"3E",
		X"42",X"10",X"8E",X"CD",X"3E",X"C6",X"7D",X"BD",X"3B",X"16",X"8E",X"3E",X"BF",X"10",X"8E",X"CE",
		X"38",X"C6",X"B6",X"BD",X"3B",X"16",X"BD",X"3F",X"88",X"10",X"8E",X"CD",X"74",X"BD",X"3F",X"A7",
		X"86",X"39",X"B7",X"CB",X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"F0",X"86",X"0E",X"7E",
		X"4A",X"62",X"14",X"19",X"1F",X"1D",X"1E",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"21",X"13",X"16",X"00",X"10",X"91",X"02",X"17",X"1C",X"1D",
		X"00",X"04",X"84",X"93",X"14",X"1C",X"18",X"00",X"04",X"71",X"13",X"1A",X"10",X"24",X"00",X"04",
		X"61",X"75",X"0D",X"21",X"15",X"00",X"04",X"52",X"22",X"15",X"10",X"16",X"00",X"04",X"42",X"10",
		X"1A",X"11",X"0E",X"00",X"04",X"32",X"17",X"15",X"0F",X"18",X"00",X"04",X"29",X"99",X"14",X"0B",
		X"18",X"00",X"04",X"10",X"11",X"0D",X"14",X"17",X"00",X"04",X"05",X"23",X"1D",X"14",X"17",X"00",
		X"03",X"99",X"09",X"0D",X"1C",X"0C",X"00",X"03",X"80",X"01",X"1A",X"20",X"0B",X"00",X"03",X"72",
		X"10",X"11",X"21",X"21",X"00",X"03",X"61",X"91",X"1C",X"19",X"18",X"00",X"03",X"51",X"01",X"14",
		X"19",X"0F",X"00",X"03",X"42",X"11",X"1E",X"13",X"17",X"00",X"03",X"35",X"67",X"0F",X"0A",X"0B",
		X"00",X"03",X"28",X"90",X"14",X"13",X"17",X"00",X"03",X"19",X"01",X"21",X"0F",X"1D",X"00",X"03",
		X"01",X"57",X"16",X"0F",X"19",X"00",X"02",X"92",X"30",X"0C",X"1F",X"24",X"00",X"02",X"87",X"77",
		X"14",X"14",X"15",X"00",X"02",X"79",X"87",X"1D",X"0B",X"15",X"00",X"02",X"69",X"59",X"0E",X"0F",
		X"0C",X"00",X"02",X"58",X"88",X"18",X"0A",X"10",X"00",X"02",X"46",X"75",X"14",X"1C",X"18",X"00",
		X"02",X"33",X"10",X"1A",X"10",X"24",X"00",X"02",X"29",X"17",X"15",X"10",X"16",X"00",X"02",X"25",
		X"52",X"0D",X"21",X"15",X"00",X"02",X"05",X"22",X"14",X"0B",X"18",X"00",X"01",X"76",X"35",X"17",
		X"1C",X"1D",X"00",X"01",X"65",X"35",X"15",X"0B",X"23",X"00",X"01",X"55",X"05",X"14",X"11",X"16",
		X"00",X"01",X"43",X"15",X"1C",X"0B",X"17",X"00",X"01",X"31",X"09",X"12",X"0F",X"0D",X"00",X"01",
		X"20",X"10",X"15",X"20",X"0E",X"00",X"01",X"17",X"55",X"0F",X"14",X"1D",X"00",X"01",X"05",X"02",
		X"20",X"0B",X"22",X"00",X"00",X"94",X"05",X"0E",X"1C",X"14",X"00",X"00",X"83",X"11",X"14",X"0B",
		X"23",X"00",X"00",X"70",X"01",X"0A",X"0A",X"0A",X"00",X"00",X"40",X"00",X"34",X"34",X"8E",X"3F",
		X"75",X"C6",X"07",X"BD",X"3B",X"16",X"35",X"B4",X"34",X"02",X"8D",X"05",X"B7",X"CD",X"6C",X"35",
		X"82",X"34",X"10",X"8E",X"CD",X"3E",X"4F",X"AB",X"84",X"30",X"01",X"8C",X"CD",X"6C",X"27",X"F9",
		X"8C",X"CD",X"74",X"26",X"F2",X"35",X"90",X"34",X"02",X"8D",X"04",X"A7",X"26",X"35",X"82",X"34",
		X"24",X"C6",X"0E",X"4F",X"C1",X"08",X"27",X"02",X"AB",X"A4",X"31",X"21",X"5A",X"26",X"F5",X"35",
		X"A4",X"86",X"32",X"34",X"02",X"10",X"8E",X"CD",X"74",X"8D",X"E4",X"A8",X"26",X"84",X"0F",X"27",
		X"0F",X"BD",X"40",X"91",X"7F",X"CD",X"00",X"7F",X"CD",X"01",X"6A",X"E4",X"27",X"12",X"20",X"E9",
		X"86",X"03",X"C6",X"04",X"8D",X"65",X"25",X"E9",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"D9",
		X"35",X"02",X"8E",X"3F",X"0C",X"10",X"8E",X"CF",X"A4",X"C6",X"2A",X"BD",X"3B",X"16",X"8D",X"91",
		X"B8",X"CD",X"6C",X"84",X"0F",X"27",X"02",X"8D",X"0F",X"10",X"8E",X"CD",X"3E",X"86",X"17",X"C6",
		X"04",X"8D",X"38",X"24",X"02",X"8D",X"01",X"39",X"8E",X"CD",X"3E",X"86",X"0A",X"BD",X"40",X"FA",
		X"8C",X"CD",X"66",X"25",X"F8",X"8E",X"CD",X"74",X"10",X"8E",X"CD",X"3E",X"86",X"06",X"BD",X"40",
		X"B1",X"10",X"8E",X"CD",X"66",X"8D",X"7A",X"8E",X"CD",X"7A",X"10",X"8E",X"CD",X"6C",X"86",X"08",
		X"8D",X"6F",X"BD",X"3F",X"88",X"10",X"8E",X"CD",X"74",X"20",X"46",X"34",X"16",X"C6",X"39",X"F7",
		X"CB",X"FF",X"1F",X"21",X"BD",X"40",X"F2",X"C1",X"0A",X"25",X"32",X"C1",X"24",X"22",X"2E",X"4A",
		X"26",X"F2",X"A6",X"61",X"BD",X"40",X"F2",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",X"40",
		X"F2",X"34",X"04",X"C4",X"0F",X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",X"22",
		X"0C",X"4A",X"26",X"EA",X"1C",X"FE",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"96",X"1A",X"01",X"20",
		X"F5",X"34",X"36",X"30",X"2E",X"8C",X"CF",X"A4",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",X"2E",
		X"30",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"EC",X"BD",X"3F",X"7C",X"BD",X"3F",X"A7",X"35",
		X"B6",X"34",X"36",X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"34",X"76",X"CC",X"00",
		X"00",X"1F",X"01",X"1F",X"02",X"CE",X"A0",X"00",X"86",X"39",X"36",X"34",X"36",X"34",X"36",X"34",
		X"36",X"34",X"36",X"34",X"36",X"34",X"B7",X"CB",X"FF",X"11",X"83",X"FF",X"EC",X"26",X"EB",X"35",
		X"F6",X"A6",X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",
		X"8D",X"EF",X"34",X"02",X"8D",X"EB",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",
		X"44",X"44",X"A7",X"81",X"35",X"82",X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",
		X"34",X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"0F",X"58",X"34",X"04",X"58",X"EB",X"E0",
		X"8E",X"CC",X"FC",X"3A",X"8D",X"CC",X"34",X"04",X"8D",X"C8",X"34",X"04",X"8D",X"C4",X"34",X"04",
		X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",X"89",X"00",
		X"19",X"30",X"1A",X"8D",X"B5",X"35",X"04",X"35",X"02",X"8D",X"BB",X"35",X"02",X"35",X"96",X"BD",
		X"F0",X"0F",X"86",X"0F",X"BD",X"4A",X"62",X"0F",X"D5",X"8E",X"11",X"70",X"86",X"F1",X"C6",X"22",
		X"10",X"8E",X"CD",X"3E",X"10",X"9C",X"EA",X"26",X"04",X"C6",X"55",X"20",X"07",X"10",X"9C",X"EE",
		X"26",X"02",X"C6",X"77",X"BD",X"4A",X"56",X"86",X"2B",X"BD",X"4A",X"50",X"30",X"89",X"03",X"00",
		X"86",X"15",X"97",X"DC",X"0A",X"DC",X"27",X"1B",X"1E",X"12",X"BD",X"3B",X"31",X"81",X"0A",X"2E",
		X"09",X"0D",X"D5",X"26",X"07",X"10",X"9F",X"D5",X"20",X"02",X"0F",X"D5",X"1E",X"12",X"BD",X"4A",
		X"50",X"20",X"E1",X"0D",X"D5",X"27",X"02",X"9E",X"D5",X"86",X"04",X"97",X"DC",X"10",X"8E",X"CD",
		X"6C",X"1E",X"12",X"BD",X"3B",X"31",X"1E",X"12",X"8A",X"F0",X"85",X"0F",X"26",X"02",X"8A",X"0F",
		X"BD",X"4A",X"56",X"0A",X"DC",X"1E",X"12",X"BD",X"3B",X"31",X"1E",X"12",X"BD",X"4A",X"56",X"0A",
		X"DC",X"26",X"F2",X"8E",X"13",X"80",X"C6",X"33",X"CE",X"4A",X"5F",X"DF",X"DF",X"CE",X"4A",X"59",
		X"86",X"0D",X"97",X"DC",X"86",X"02",X"97",X"E2",X"86",X"07",X"97",X"E1",X"86",X"0E",X"97",X"E7",
		X"8D",X"54",X"8E",X"3D",X"80",X"86",X"0D",X"97",X"DC",X"86",X"15",X"97",X"E2",X"8D",X"47",X"8E",
		X"67",X"80",X"86",X"0D",X"97",X"DC",X"86",X"28",X"97",X"E2",X"8D",X"3A",X"8E",X"13",X"36",X"10",
		X"8E",X"CF",X"A4",X"C6",X"11",X"CE",X"4A",X"56",X"DF",X"DF",X"CE",X"4A",X"50",X"86",X"03",X"97",
		X"DC",X"86",X"01",X"97",X"E2",X"86",X"0A",X"97",X"E1",X"86",X"15",X"97",X"E7",X"8D",X"17",X"8E",
		X"53",X"36",X"86",X"03",X"97",X"DC",X"86",X"04",X"97",X"E2",X"8D",X"0A",X"8E",X"F0",X"12",X"CC",
		X"40",X"00",X"BD",X"E0",X"09",X"39",X"9F",X"D9",X"34",X"04",X"C6",X"03",X"D7",X"E9",X"5C",X"D7",
		X"E6",X"E6",X"E4",X"10",X"9C",X"EA",X"27",X"05",X"10",X"9C",X"EC",X"26",X"02",X"C6",X"55",X"10",
		X"9C",X"EE",X"27",X"05",X"10",X"9C",X"F0",X"26",X"02",X"C6",X"77",X"96",X"E2",X"85",X"F0",X"26",
		X"02",X"8A",X"F0",X"AD",X"9F",X"A0",X"DF",X"86",X"2B",X"AD",X"C4",X"86",X"0A",X"AD",X"C4",X"1E",
		X"12",X"BD",X"3B",X"31",X"1E",X"12",X"AD",X"C4",X"0A",X"E9",X"26",X"F3",X"9F",X"D5",X"9E",X"D9",
		X"1E",X"01",X"D6",X"D6",X"9B",X"E7",X"1E",X"01",X"0F",X"DD",X"1E",X"12",X"BD",X"3B",X"31",X"1E",
		X"12",X"0D",X"DD",X"26",X"1A",X"34",X"02",X"86",X"04",X"91",X"E6",X"26",X"04",X"35",X"02",X"20",
		X"06",X"35",X"02",X"85",X"F0",X"26",X"08",X"8A",X"F0",X"85",X"0F",X"26",X"02",X"8A",X"0F",X"97",
		X"DD",X"03",X"DD",X"AD",X"9F",X"A0",X"DF",X"0A",X"E6",X"26",X"CF",X"9F",X"D5",X"9E",X"D9",X"1E",
		X"01",X"D6",X"D6",X"DB",X"E1",X"1E",X"01",X"96",X"E2",X"8B",X"01",X"19",X"97",X"E2",X"0A",X"DC",
		X"35",X"04",X"10",X"26",X"FF",X"62",X"39",X"34",X"12",X"9B",X"F2",X"19",X"24",X"02",X"86",X"99",
		X"97",X"F2",X"8E",X"CD",X"00",X"BD",X"40",X"FA",X"35",X"12",X"7E",X"5E",X"D8",X"34",X"16",X"C6",
		X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",X"C6",X"01",X"BD",X"41",X"10",
		X"58",X"8E",X"CC",X"06",X"3A",X"BD",X"40",X"F2",X"8D",X"61",X"96",X"F4",X"34",X"04",X"AB",X"E4",
		X"97",X"F4",X"96",X"F3",X"AB",X"E0",X"97",X"F3",X"8E",X"CC",X"12",X"BD",X"40",X"F2",X"8D",X"4B",
		X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",X"96",X"8E",X"CC",X"0E",X"BD",X"40",X"F2",X"8D",X"3B",
		X"8D",X"23",X"34",X"02",X"D7",X"F3",X"8E",X"CC",X"10",X"BD",X"40",X"F2",X"96",X"F4",X"8D",X"2B",
		X"8D",X"13",X"4D",X"27",X"04",X"0F",X"F3",X"0F",X"F4",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"41",
		X"16",X"8D",X"84",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",
		X"99",X"8B",X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",X"4F",X"C1",X"10",
		X"25",X"06",X"8B",X"0A",X"C0",X"10",X"20",X"F6",X"34",X"04",X"AB",X"E0",X"1F",X"89",X"35",X"82",
		X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",
		X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"10",X"8E",X"B0",X"00",X"8E",X"CC",X"16",X"BD",X"40",
		X"F2",X"8D",X"C8",X"E7",X"A4",X"C6",X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",X"5A",X"26",X"FB",
		X"8E",X"43",X"F6",X"AF",X"26",X"8E",X"20",X"80",X"AF",X"28",X"C6",X"0A",X"E7",X"22",X"6F",X"21",
		X"86",X"25",X"A7",X"23",X"86",X"3C",X"A7",X"24",X"86",X"77",X"A7",X"25",X"AD",X"B8",X"06",X"25",
		X"05",X"BD",X"44",X"B8",X"20",X"F6",X"C6",X"14",X"8E",X"CD",X"3E",X"31",X"2F",X"A6",X"A0",X"BD",
		X"40",X"FA",X"5A",X"26",X"F8",X"39",X"4F",X"E6",X"21",X"27",X"12",X"34",X"14",X"5A",X"CB",X"0F",
		X"E6",X"A5",X"58",X"BE",X"4A",X"68",X"AB",X"95",X"35",X"14",X"5A",X"26",X"EE",X"AE",X"28",X"30",
		X"8B",X"AF",X"2A",X"C6",X"0F",X"EB",X"21",X"A6",X"A5",X"BD",X"44",X"C1",X"E6",X"24",X"F7",X"C8",
		X"07",X"F6",X"C8",X"04",X"C4",X"07",X"26",X"08",X"E6",X"2E",X"27",X"74",X"6A",X"2E",X"20",X"70",
		X"8E",X"44",X"38",X"AF",X"26",X"1C",X"FE",X"39",X"34",X"04",X"E6",X"24",X"F7",X"C8",X"07",X"35",
		X"04",X"F1",X"C8",X"04",X"26",X"5A",X"54",X"26",X"13",X"E6",X"2E",X"27",X"02",X"6A",X"2E",X"8D",
		X"63",X"A1",X"22",X"26",X"04",X"A6",X"23",X"20",X"47",X"4A",X"20",X"44",X"54",X"26",X"13",X"E6",
		X"2E",X"27",X"02",X"6A",X"2E",X"8D",X"4D",X"A1",X"23",X"26",X"04",X"A6",X"22",X"20",X"31",X"4C",
		X"20",X"2E",X"E6",X"2E",X"27",X"04",X"6A",X"2E",X"20",X"26",X"C6",X"02",X"E7",X"2E",X"81",X"25",
		X"26",X"0E",X"6D",X"21",X"27",X"1A",X"8D",X"2C",X"6C",X"A4",X"6A",X"21",X"8D",X"40",X"20",X"0A",
		X"6C",X"21",X"8D",X"3A",X"6A",X"A4",X"26",X"08",X"1A",X"01",X"8E",X"43",X"F6",X"AF",X"26",X"39",
		X"8D",X"04",X"1C",X"FE",X"20",X"F4",X"C6",X"0F",X"EB",X"21",X"A7",X"A5",X"E6",X"25",X"AE",X"2A",
		X"BD",X"4A",X"50",X"39",X"C6",X"00",X"20",X"F6",X"34",X"06",X"86",X"04",X"BD",X"F0",X"09",X"35",
		X"86",X"34",X"06",X"E6",X"25",X"86",X"33",X"AE",X"2A",X"BD",X"4A",X"50",X"35",X"86",X"34",X"06",
		X"C6",X"00",X"20",X"F1",X"C6",X"66",X"D7",X"E9",X"C6",X"88",X"8D",X"04",X"C6",X"9A",X"20",X"20",
		X"34",X"36",X"8E",X"CC",X"88",X"BD",X"3B",X"31",X"1F",X"02",X"8E",X"CC",X"24",X"D6",X"E9",X"BD",
		X"3B",X"31",X"1E",X"12",X"BD",X"4A",X"50",X"1E",X"12",X"8C",X"CC",X"56",X"26",X"F1",X"35",X"B6",
		X"34",X"36",X"8E",X"CC",X"8A",X"BD",X"3B",X"31",X"1F",X"02",X"8E",X"CC",X"56",X"D6",X"E9",X"BD",
		X"3B",X"31",X"1E",X"12",X"BD",X"4A",X"50",X"1E",X"12",X"8C",X"CC",X"88",X"26",X"F1",X"35",X"B6",
		X"10",X"8E",X"B0",X"00",X"AF",X"28",X"CC",X"43",X"F6",X"ED",X"26",X"C6",X"19",X"E7",X"A4",X"C6",
		X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",X"5A",X"26",X"FB",X"E7",X"21",X"E7",X"22",X"6F",X"2F",
		X"86",X"32",X"A7",X"23",X"86",X"3C",X"A7",X"24",X"86",X"77",X"A7",X"25",X"AD",X"B8",X"06",X"25",
		X"05",X"BD",X"44",X"B8",X"20",X"F6",X"39",X"8E",X"25",X"60",X"8D",X"C4",X"C6",X"19",X"8E",X"CC",
		X"24",X"31",X"2F",X"A6",X"A0",X"BD",X"40",X"FA",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"88",
		X"BD",X"40",X"FA",X"C6",X"88",X"8D",X"30",X"86",X"34",X"C6",X"22",X"8E",X"48",X"6A",X"BD",X"4A",
		X"50",X"CE",X"45",X"B7",X"8E",X"CC",X"88",X"BD",X"40",X"F2",X"BD",X"46",X"14",X"D7",X"F7",X"0F",
		X"E9",X"C6",X"60",X"BD",X"44",X"E0",X"96",X"F7",X"8E",X"CC",X"88",X"BD",X"40",X"FA",X"86",X"22",
		X"97",X"E9",X"BD",X"44",X"E0",X"20",X"DD",X"86",X"51",X"8E",X"25",X"90",X"BD",X"4A",X"53",X"86",
		X"52",X"8E",X"25",X"A0",X"7E",X"4A",X"53",X"86",X"34",X"C6",X"00",X"8E",X"48",X"6A",X"BD",X"4A",
		X"50",X"8D",X"E4",X"8E",X"25",X"70",X"BD",X"45",X"20",X"C6",X"19",X"8E",X"CC",X"56",X"31",X"2F",
		X"A6",X"A0",X"BD",X"40",X"FA",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"8A",X"BD",X"40",X"FA",
		X"C6",X"88",X"8D",X"C3",X"86",X"34",X"C6",X"22",X"8E",X"48",X"7A",X"BD",X"4A",X"50",X"CE",X"46",
		X"13",X"8E",X"CC",X"8A",X"BD",X"40",X"F2",X"8D",X"1B",X"D7",X"F7",X"0F",X"E9",X"C6",X"70",X"BD",
		X"45",X"00",X"96",X"F7",X"8E",X"CC",X"8A",X"BD",X"40",X"FA",X"86",X"22",X"97",X"E9",X"BD",X"45",
		X"00",X"20",X"DE",X"39",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"04",X"32",X"62",X"6E",X"C4",X"B6",
		X"C8",X"04",X"84",X"03",X"BD",X"44",X"B8",X"B1",X"C8",X"04",X"26",X"E8",X"4D",X"27",X"E5",X"44",
		X"26",X"06",X"C1",X"18",X"27",X"DE",X"5A",X"39",X"44",X"26",X"D9",X"C1",X"40",X"27",X"D5",X"5C",
		X"39",X"A6",X"84",X"84",X"F0",X"27",X"07",X"CC",X"99",X"99",X"ED",X"81",X"ED",X"81",X"39",X"0F",
		X"F5",X"B6",X"CC",X"05",X"44",X"25",X"03",X"7E",X"5E",X"D3",X"8E",X"A0",X"4C",X"8D",X"E2",X"8E",
		X"A0",X"56",X"8D",X"DD",X"0D",X"60",X"27",X"5A",X"8E",X"A0",X"4C",X"10",X"8E",X"A0",X"56",X"BD",
		X"49",X"99",X"25",X"4E",X"1E",X"21",X"BD",X"49",X"5D",X"24",X"22",X"0C",X"F5",X"8E",X"48",X"E9",
		X"CC",X"42",X"00",X"BD",X"E0",X"09",X"86",X"10",X"A7",X"24",X"86",X"01",X"A7",X"A8",X"31",X"8E",
		X"A0",X"56",X"AF",X"A8",X"2D",X"8E",X"70",X"A0",X"AF",X"A8",X"2F",X"20",X"12",X"8E",X"A0",X"56",
		X"AF",X"C8",X"2D",X"8E",X"70",X"A0",X"AF",X"C8",X"2F",X"86",X"01",X"C6",X"42",X"8D",X"66",X"8E",
		X"A0",X"4C",X"AF",X"C8",X"2D",X"8E",X"20",X"A0",X"AF",X"C8",X"2F",X"4F",X"C6",X"41",X"8D",X"55",
		X"20",X"50",X"8E",X"A0",X"4C",X"BD",X"49",X"5D",X"24",X"21",X"0C",X"F5",X"8E",X"48",X"E9",X"CC",
		X"42",X"00",X"BD",X"E0",X"09",X"86",X"10",X"A7",X"24",X"4F",X"A7",X"A8",X"31",X"8E",X"A0",X"4C",
		X"AF",X"A8",X"2D",X"8E",X"20",X"A0",X"AF",X"A8",X"2F",X"20",X"11",X"8E",X"A0",X"4C",X"AF",X"C8",
		X"2D",X"8E",X"20",X"A0",X"AF",X"C8",X"2F",X"4F",X"C6",X"42",X"8D",X"19",X"0D",X"60",X"27",X"12",
		X"8E",X"A0",X"56",X"AF",X"C8",X"2D",X"8E",X"70",X"A0",X"AF",X"C8",X"2F",X"86",X"01",X"C6",X"41",
		X"8D",X"03",X"7E",X"3B",X"64",X"BD",X"49",X"63",X"24",X"23",X"0C",X"F5",X"34",X"02",X"8E",X"47",
		X"65",X"1F",X"98",X"5F",X"BD",X"E0",X"09",X"86",X"10",X"A7",X"24",X"35",X"02",X"A7",X"A8",X"31",
		X"AE",X"C8",X"2D",X"AF",X"A8",X"2D",X"AE",X"C8",X"2F",X"AF",X"A8",X"2F",X"39",X"BD",X"49",X"80",
		X"24",X"22",X"0C",X"F5",X"34",X"02",X"8E",X"47",X"65",X"1F",X"98",X"5F",X"BD",X"E0",X"09",X"86",
		X"08",X"A7",X"24",X"35",X"02",X"A7",X"A8",X"31",X"AE",X"C8",X"2D",X"AF",X"A8",X"2D",X"AE",X"C8",
		X"2F",X"AF",X"A8",X"2F",X"39",X"6F",X"C8",X"2C",X"E6",X"C8",X"31",X"26",X"0B",X"8E",X"0A",X"B0",
		X"C6",X"3C",X"34",X"04",X"C6",X"55",X"20",X"09",X"8E",X"58",X"B0",X"C6",X"34",X"34",X"04",X"C6",
		X"77",X"86",X"68",X"BD",X"4A",X"53",X"1F",X"98",X"31",X"47",X"C6",X"02",X"E7",X"2E",X"35",X"04",
		X"E7",X"24",X"8E",X"47",X"9D",X"AF",X"2C",X"AE",X"C8",X"2F",X"BD",X"49",X"D2",X"A6",X"42",X"81",
		X"42",X"27",X"21",X"ED",X"C8",X"32",X"AF",X"C8",X"34",X"10",X"AF",X"C8",X"36",X"86",X"01",X"BD",
		X"E0",X"37",X"AE",X"C4",X"A6",X"02",X"81",X"42",X"27",X"F3",X"EC",X"C8",X"32",X"AE",X"C8",X"34",
		X"10",X"AE",X"C8",X"36",X"BD",X"49",X"63",X"24",X"13",X"6D",X"C8",X"31",X"26",X"05",X"10",X"9F",
		X"EC",X"20",X"03",X"10",X"9F",X"F0",X"8E",X"CF",X"EA",X"BD",X"48",X"B8",X"BD",X"49",X"80",X"24",
		X"19",X"6D",X"C8",X"2C",X"27",X"1D",X"30",X"47",X"30",X"0F",X"10",X"8E",X"CD",X"66",X"C6",X"03",
		X"BD",X"3B",X"CF",X"BD",X"3F",X"88",X"86",X"05",X"8D",X"75",X"24",X"70",X"1F",X"12",X"BD",X"40",
		X"91",X"20",X"51",X"30",X"A9",X"32",X"9A",X"26",X"2C",X"8E",X"CF",X"96",X"BD",X"48",X"D3",X"31",
		X"26",X"AE",X"C8",X"2D",X"C6",X"04",X"BD",X"3B",X"CF",X"10",X"8E",X"CD",X"3E",X"6D",X"C8",X"31",
		X"26",X"05",X"10",X"9F",X"EA",X"20",X"03",X"10",X"9F",X"EE",X"30",X"47",X"30",X"0F",X"C6",X"14",
		X"BD",X"3B",X"CF",X"20",X"B1",X"BD",X"48",X"73",X"34",X"01",X"34",X"10",X"10",X"AC",X"E1",X"22",
		X"0F",X"8D",X"75",X"6D",X"C8",X"31",X"26",X"05",X"10",X"9F",X"EA",X"20",X"03",X"10",X"9F",X"EE",
		X"35",X"01",X"24",X"18",X"8E",X"A0",X"EA",X"31",X"47",X"AE",X"C8",X"2F",X"30",X"89",X"EA",X"F6",
		X"86",X"6A",X"E6",X"25",X"BD",X"4A",X"53",X"86",X"60",X"BD",X"E0",X"37",X"7E",X"E0",X"0F",X"34",
		X"26",X"20",X"0C",X"34",X"26",X"8E",X"CD",X"66",X"8D",X"24",X"86",X"04",X"25",X"01",X"4C",X"97",
		X"D5",X"8E",X"CD",X"74",X"8D",X"18",X"24",X"04",X"0A",X"D5",X"27",X"0E",X"30",X"0E",X"8C",X"CF",
		X"A4",X"25",X"F1",X"8E",X"CF",X"96",X"1C",X"FE",X"35",X"A6",X"1A",X"01",X"35",X"A6",X"34",X"10",
		X"31",X"47",X"31",X"2F",X"C6",X"03",X"BD",X"40",X"E1",X"A1",X"A0",X"26",X"07",X"5A",X"26",X"F6",
		X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",X"34",X"20",X"BD",X"48",X"D3",X"30",X"47",X"30",
		X"0F",X"C6",X"03",X"BD",X"3B",X"CF",X"AE",X"C8",X"2D",X"C6",X"04",X"BD",X"3B",X"CF",X"35",X"20",
		X"7E",X"3F",X"A7",X"34",X"30",X"1F",X"12",X"10",X"AC",X"62",X"27",X"0B",X"30",X"32",X"86",X"0E",
		X"BD",X"40",X"B1",X"31",X"32",X"20",X"F0",X"35",X"B0",X"6C",X"C8",X"2C",X"31",X"47",X"A6",X"C8",
		X"31",X"26",X"08",X"86",X"3C",X"A7",X"24",X"86",X"55",X"20",X"06",X"86",X"34",X"A7",X"24",X"86",
		X"77",X"1F",X"89",X"86",X"67",X"8E",X"29",X"5B",X"BD",X"4A",X"53",X"1F",X"98",X"8E",X"49",X"15",
		X"AF",X"2C",X"7E",X"49",X"C4",X"30",X"2F",X"10",X"8E",X"CD",X"3E",X"C6",X"14",X"BD",X"3B",X"CF",
		X"10",X"8E",X"CD",X"66",X"8E",X"CF",X"96",X"BD",X"48",X"D3",X"10",X"8E",X"CD",X"74",X"BD",X"3F",
		X"A7",X"AE",X"C8",X"2D",X"10",X"8E",X"CD",X"6C",X"C6",X"04",X"BD",X"3B",X"CF",X"8E",X"3F",X"75",
		X"10",X"8E",X"CD",X"66",X"C6",X"03",X"BD",X"3B",X"CF",X"BD",X"3F",X"88",X"8E",X"CD",X"3E",X"A6",
		X"C8",X"31",X"26",X"04",X"9F",X"EA",X"20",X"02",X"9F",X"EE",X"7E",X"47",X"68",X"10",X"8E",X"CD",
		X"6C",X"20",X"36",X"34",X"12",X"10",X"8E",X"CF",X"AA",X"AE",X"C8",X"2D",X"8D",X"2B",X"25",X"0C",
		X"31",X"2E",X"10",X"8C",X"CF",X"F8",X"25",X"F4",X"1C",X"FE",X"35",X"92",X"31",X"3A",X"35",X"92",
		X"34",X"12",X"10",X"8E",X"CD",X"6C",X"AE",X"C8",X"2D",X"8D",X"0E",X"25",X"EF",X"31",X"2E",X"10",
		X"8C",X"CF",X"96",X"25",X"F4",X"1C",X"FE",X"35",X"92",X"34",X"36",X"1E",X"12",X"C6",X"04",X"8D",
		X"17",X"C1",X"04",X"26",X"02",X"84",X"0F",X"A1",X"A0",X"22",X"05",X"25",X"07",X"5A",X"26",X"EF",
		X"1C",X"FE",X"35",X"B6",X"1A",X"01",X"35",X"B6",X"8C",X"C0",X"00",X"25",X"04",X"BD",X"40",X"E1",
		X"39",X"A6",X"80",X"39",X"8E",X"CC",X"16",X"BD",X"40",X"F2",X"BD",X"43",X"7B",X"8E",X"26",X"43",
		X"20",X"02",X"C6",X"03",X"A7",X"25",X"E7",X"A4",X"AF",X"28",X"C6",X"14",X"86",X"0A",X"30",X"2F",
		X"A7",X"80",X"5A",X"26",X"FB",X"8E",X"43",X"F6",X"AF",X"26",X"C6",X"0A",X"6F",X"21",X"E7",X"22",
		X"86",X"25",X"A7",X"23",X"AD",X"B8",X"06",X"25",X"15",X"10",X"AF",X"C8",X"36",X"ED",X"C8",X"32",
		X"86",X"03",X"BD",X"E0",X"37",X"10",X"AE",X"C8",X"36",X"EC",X"C8",X"32",X"20",X"E6",X"6E",X"B8",
		X"0C",X"4A",X"4F",X"55",X"53",X"54",X"2D",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",
		X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",
		X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"4A",X"7F",X"7E",X"4A",X"BF",X"7E",X"4A",X"F7",X"7E",X"4A",X"70",X"7E",X"4A",X"AD",X"7E",
		X"4A",X"E5",X"7E",X"4B",X"3A",X"7E",X"4B",X"2F",X"4B",X"5C",X"7E",X"4B",X"36",X"7E",X"4B",X"2B",
		X"34",X"67",X"10",X"8E",X"4B",X"C6",X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"11",X"35",X"E7",X"34",
		X"67",X"10",X"8E",X"4B",X"5C",X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"02",X"35",X"E7",X"BF",X"CA",
		X"04",X"48",X"10",X"AE",X"A6",X"EC",X"A1",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"10",X"BF",
		X"CA",X"02",X"C6",X"1A",X"F7",X"CA",X"00",X"88",X"04",X"5F",X"30",X"8B",X"39",X"34",X"67",X"10",
		X"8E",X"4B",X"C6",X"10",X"9F",X"D1",X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"14",X"35",X"E7",X"34",
		X"67",X"10",X"8E",X"4B",X"5C",X"10",X"9F",X"D1",X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"02",X"35",
		X"E7",X"CE",X"53",X"1F",X"33",X"C6",X"EE",X"C6",X"A6",X"C4",X"10",X"9E",X"D1",X"BD",X"4A",X"8E",
		X"6D",X"C0",X"2A",X"F4",X"39",X"34",X"67",X"10",X"8E",X"4B",X"C6",X"10",X"9F",X"D1",X"1A",X"FF",
		X"F7",X"CA",X"01",X"8D",X"14",X"35",X"E7",X"34",X"67",X"10",X"8E",X"4B",X"5C",X"10",X"9F",X"D1",
		X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"02",X"35",X"E7",X"97",X"D0",X"44",X"44",X"44",X"44",X"81",
		X"0A",X"2F",X"02",X"86",X"0A",X"10",X"9E",X"D1",X"BD",X"4A",X"8E",X"96",X"D0",X"84",X"0F",X"81",
		X"0A",X"2F",X"02",X"86",X"0A",X"10",X"9E",X"D1",X"7E",X"4A",X"8E",X"0C",X"F6",X"20",X"02",X"0F",
		X"F6",X"CE",X"4A",X"5C",X"20",X"09",X"0C",X"F6",X"20",X"02",X"0F",X"F6",X"CE",X"4A",X"53",X"10",
		X"8E",X"5D",X"7B",X"31",X"A6",X"10",X"AE",X"A6",X"AE",X"A1",X"E6",X"A0",X"0D",X"F6",X"27",X"01",
		X"5F",X"A6",X"A4",X"84",X"7F",X"AD",X"C4",X"6D",X"A0",X"2A",X"ED",X"39",X"4C",X"28",X"4C",X"3F",
		X"4C",X"56",X"4C",X"6D",X"4C",X"84",X"4C",X"9B",X"4C",X"B2",X"4C",X"C9",X"4C",X"E0",X"4C",X"F7",
		X"4D",X"0E",X"4D",X"25",X"4D",X"3C",X"4D",X"53",X"4D",X"6A",X"4D",X"81",X"4D",X"98",X"4D",X"AF",
		X"4D",X"C6",X"4D",X"DD",X"4D",X"ED",X"4E",X"04",X"4E",X"1B",X"4E",X"32",X"4E",X"50",X"4E",X"67",
		X"4E",X"7E",X"4E",X"95",X"4E",X"AC",X"4E",X"C3",X"4E",X"DA",X"4E",X"F1",X"4F",X"08",X"4F",X"1F",
		X"4F",X"3D",X"4F",X"54",X"4F",X"6B",X"4F",X"82",X"4F",X"99",X"4F",X"AA",X"4F",X"B8",X"4F",X"CF",
		X"4F",X"D8",X"4F",X"E8",X"4F",X"F8",X"4F",X"FC",X"50",X"05",X"50",X"0E",X"50",X"25",X"50",X"3C",
		X"50",X"42",X"50",X"52",X"50",X"6C",X"50",X"83",X"50",X"8F",X"50",X"9B",X"50",X"A7",X"50",X"B3",
		X"50",X"BF",X"50",X"CB",X"50",X"D7",X"50",X"E3",X"50",X"EF",X"50",X"FB",X"51",X"07",X"51",X"13",
		X"51",X"1F",X"51",X"2B",X"51",X"37",X"51",X"43",X"51",X"4F",X"51",X"5B",X"51",X"67",X"51",X"73",
		X"51",X"7F",X"51",X"8B",X"51",X"97",X"51",X"A8",X"50",X"83",X"51",X"B4",X"51",X"C0",X"51",X"CC",
		X"50",X"BF",X"51",X"D8",X"51",X"E4",X"51",X"F0",X"52",X"48",X"52",X"59",X"52",X"65",X"52",X"71",
		X"52",X"7D",X"52",X"89",X"52",X"93",X"52",X"9B",X"52",X"A7",X"52",X"AE",X"52",X"BA",X"52",X"C6",
		X"52",X"CA",X"52",X"D1",X"52",X"D8",X"52",X"F8",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",
		X"10",X"01",X"10",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",
		X"07",X"00",X"10",X"00",X"01",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"11",X"11",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"00",X"00",
		X"10",X"00",X"11",X"00",X"01",X"00",X"00",X"10",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"01",
		X"11",X"00",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"11",X"00",X"00",X"00",X"10",X"10",X"00",
		X"10",X"01",X"11",X"00",X"03",X"07",X"00",X"01",X"10",X"00",X"10",X"10",X"01",X"00",X"10",X"10",
		X"00",X"10",X"11",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"03",X"07",X"11",X"11",X"10",
		X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"10",X"01",
		X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"00",X"10",X"11",X"00",X"11",X"00",X"10",
		X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"10",X"00",
		X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",
		X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"10",X"00",
		X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"01",X"10",X"01",X"10",X"10",X"00",X"00",X"10",X"01",X"11",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",
		X"11",X"11",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"03",X"07",X"11",X"11",
		X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",
		X"11",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"11",X"10",X"00",X"10",
		X"01",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",
		X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"00",X"11",X"11",X"00",X"10",
		X"00",X"00",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",
		X"10",X"00",X"00",X"11",X"11",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"03",
		X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"01",X"10",
		X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",
		X"10",X"11",X"11",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"02",X"07",X"11",
		X"10",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"11",X"10",X"03",X"07",X"00",
		X"01",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"10",X"00",
		X"10",X"01",X"11",X"00",X"03",X"07",X"10",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"00",X"11",
		X"00",X"00",X"10",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"10",X"03",X"07",X"01",X"00",X"00",
		X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"10",X"11",
		X"11",X"10",X"04",X"07",X"01",X"10",X"11",X"00",X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",
		X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",X"10",X"00",X"00",X"10",X"01",X"00",X"01",X"00",
		X"03",X"07",X"10",X"00",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"01",X"10",X"10",X"00",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",
		X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"00",X"10",X"00",X"00",X"10",
		X"00",X"00",X"10",X"00",X"00",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",
		X"10",X"00",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"10",X"10",X"03",X"07",X"01",X"11",
		X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"11",X"11",X"00",X"10",X"10",X"00",X"10",X"01",X"00",
		X"10",X"00",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"11",X"00",X"10",
		X"10",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"11",
		X"00",X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"00",X"10",X"01",X"11",X"00",X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",
		X"10",X"00",X"10",X"10",X"00",X"10",X"01",X"01",X"00",X"01",X"01",X"00",X"00",X"10",X"00",X"04",
		X"07",X"01",X"00",X"01",X"00",X"10",X"00",X"00",X"10",X"10",X"00",X"00",X"10",X"10",X"01",X"00",
		X"10",X"10",X"01",X"00",X"10",X"10",X"01",X"00",X"10",X"01",X"10",X"11",X"00",X"03",X"07",X"10",
		X"00",X"10",X"10",X"00",X"10",X"01",X"01",X"00",X"00",X"10",X"00",X"01",X"01",X"00",X"10",X"00",
		X"10",X"10",X"00",X"10",X"03",X"07",X"01",X"00",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"01",
		X"01",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"03",X"07",X"01",X"11",X"10",
		X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"11",
		X"11",X"10",X"03",X"07",X"00",X"01",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"11",X"11",X"10",
		X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"00",X"03",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"11",X"11",X"10",X"03",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"01",X"11",X"00",X"10",X"00",X"10",
		X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",
		X"07",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"02",X"07",X"00",X"10",X"01",X"00",X"10",X"00",
		X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"02",X"07",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"01",X"02",X"10",X"10",X"01",X"07",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"03",X"07",
		X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"00",X"10",X"00",X"00",X"03",X"07",X"01",X"00",X"00",X"10",X"10",X"00",X"10",X"10",X"00",
		X"01",X"00",X"00",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"10",X"10",X"02",X"02",X"10",X"10",
		X"10",X"10",X"02",X"07",X"00",X"00",X"11",X"10",X"11",X"10",X"00",X"00",X"00",X"00",X"11",X"10",
		X"11",X"10",X"03",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"00",X"10",
		X"00",X"01",X"11",X"00",X"10",X"10",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"10",X"02",
		X"05",X"01",X"00",X"11",X"00",X"01",X"00",X"01",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",
		X"10",X"11",X"10",X"10",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"11",X"10",X"00",
		X"10",X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"02",
		X"05",X"11",X"10",X"10",X"00",X"11",X"10",X"00",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"10",
		X"00",X"11",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"01",
		X"00",X"01",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",X"02",
		X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"02",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",
		X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"11",X"10",X"02",
		X"05",X"11",X"10",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"10",X"02",X"05",X"11",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"00",X"10",
		X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"00",X"10",X"00",X"10",X"00",X"02",
		X"05",X"11",X"10",X"10",X"00",X"10",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"10",X"10",X"10",
		X"10",X"11",X"10",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",X"00",X"01",X"00",X"01",
		X"00",X"11",X"10",X"02",X"05",X"00",X"10",X"00",X"10",X"00",X"10",X"10",X"10",X"11",X"10",X"02",
		X"05",X"10",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"10",X"00",X"10",
		X"00",X"10",X"00",X"10",X"00",X"11",X"10",X"03",X"05",X"11",X"11",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"00",X"10",X"00",
		X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"00",X"10",X"02",X"05",X"11",X"10",
		X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"10",
		X"02",X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"00",X"20",X"4A",X"4F",X"55",
		X"53",X"54",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"20",
		X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",
		X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",
		X"43",X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",
		X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"03",X"05",X"10",X"00",X"10",X"10",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"01",
		X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"10",X"01",X"00",X"01",
		X"00",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"11",X"10",X"02",X"05",X"00",
		X"10",X"01",X"00",X"11",X"10",X"01",X"00",X"00",X"10",X"02",X"04",X"00",X"00",X"11",X"10",X"00",
		X"00",X"11",X"10",X"02",X"03",X"00",X"00",X"00",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",
		X"10",X"01",X"10",X"00",X"00",X"01",X"00",X"01",X"05",X"10",X"10",X"10",X"00",X"10",X"02",X"05",
		X"00",X"10",X"01",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"02",X"05",X"10",X"00",X"01",X"00",
		X"00",X"10",X"01",X"00",X"10",X"00",X"01",X"02",X"10",X"10",X"01",X"05",X"00",X"00",X"00",X"10",
		X"10",X"01",X"05",X"00",X"00",X"00",X"00",X"10",X"06",X"05",X"11",X"10",X"11",X"10",X"11",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"10",X"11",X"10",X"11",X"10",X"11",X"10",X"03",X"05",X"00",X"10",X"00",X"00",X"01",X"00",
		X"11",X"11",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"5A",X"6E",X"5A",X"8A",X"5A",X"FB",X"5B",
		X"0D",X"5B",X"18",X"5B",X"23",X"5A",X"9B",X"5A",X"B0",X"5A",X"B8",X"5A",X"C5",X"5A",X"E1",X"54",
		X"1F",X"54",X"2F",X"54",X"32",X"54",X"35",X"54",X"38",X"54",X"3A",X"54",X"50",X"54",X"5E",X"54",
		X"68",X"54",X"72",X"54",X"7D",X"54",X"8D",X"54",X"A2",X"54",X"B6",X"54",X"B8",X"54",X"BF",X"54",
		X"CD",X"54",X"E4",X"55",X"00",X"55",X"18",X"55",X"26",X"55",X"42",X"55",X"4D",X"55",X"54",X"55",
		X"5B",X"55",X"65",X"55",X"75",X"55",X"7E",X"55",X"89",X"55",X"94",X"55",X"A4",X"55",X"B4",X"55",
		X"BD",X"55",X"C7",X"55",X"CB",X"55",X"D5",X"55",X"E7",X"55",X"F6",X"56",X"07",X"56",X"17",X"56",
		X"23",X"56",X"2B",X"56",X"40",X"56",X"50",X"56",X"63",X"56",X"74",X"56",X"88",X"56",X"9F",X"56",
		X"AF",X"56",X"BE",X"56",X"D3",X"56",X"ED",X"56",X"FE",X"57",X"11",X"57",X"26",X"57",X"3A",X"57",
		X"57",X"57",X"7A",X"57",X"9A",X"57",X"AC",X"57",X"C5",X"57",X"DD",X"57",X"F5",X"58",X"0B",X"58",
		X"15",X"58",X"2D",X"58",X"43",X"58",X"61",X"58",X"88",X"58",X"8B",X"58",X"95",X"58",X"9B",X"58",
		X"B7",X"58",X"BF",X"58",X"D8",X"58",X"FA",X"59",X"15",X"59",X"1D",X"59",X"33",X"59",X"41",X"59",
		X"50",X"59",X"58",X"59",X"75",X"59",X"93",X"59",X"A3",X"59",X"B0",X"59",X"B9",X"59",X"D4",X"59",
		X"F6",X"5A",X"23",X"5A",X"28",X"5A",X"4F",X"5A",X"5D",X"5B",X"2D",X"5B",X"3D",X"5D",X"35",X"5D",
		X"43",X"5D",X"68",X"5D",X"2F",X"5D",X"22",X"5B",X"57",X"5B",X"59",X"5B",X"61",X"5B",X"69",X"5B",
		X"80",X"5B",X"93",X"5B",X"A1",X"5B",X"B1",X"5B",X"E6",X"5C",X"08",X"5C",X"11",X"5C",X"1C",X"5C",
		X"2C",X"5C",X"3E",X"5C",X"54",X"5C",X"62",X"5C",X"72",X"5C",X"83",X"5C",X"8A",X"5C",X"AC",X"5C",
		X"BC",X"5C",X"C9",X"5C",X"D5",X"5C",X"E7",X"5C",X"F0",X"5C",X"F2",X"5D",X"0D",X"5D",X"18",X"1E",
		X"12",X"23",X"0A",X"11",X"0B",X"17",X"0F",X"0A",X"13",X"1D",X"0A",X"19",X"20",X"0F",X"9C",X"02",
		X"05",X"80",X"05",X"00",X"80",X"07",X"05",X"80",X"01",X"AF",X"13",X"18",X"13",X"1E",X"13",X"0B",
		X"16",X"0A",X"1E",X"0F",X"1D",X"1E",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",X"8F",
		X"0B",X"16",X"16",X"0A",X"1D",X"23",X"1D",X"1E",X"0F",X"17",X"1D",X"0A",X"11",X"99",X"1C",X"0B",
		X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"1C",X"19",X"17",X"0A",X"0F",X"1C",X"1C",X"19",
		X"1C",X"8A",X"0B",X"16",X"16",X"0A",X"1C",X"19",X"17",X"1D",X"0A",X"19",X"95",X"1C",X"0B",X"17",
		X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",X"19",X"16",X"16",X"19",X"21",X"9D",X"1A",X"1C",X"0F",
		X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"0F",X"0A",X"1E",X"19",X"0A",X"0F",X"22",
		X"13",X"9E",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"1D",X"0A",X"0E",X"0F",
		X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",X"99",X"18",X"19",X"0A",X"0D",X"17",X"19",X"9D",X"0D",
		X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"10",X"1C",X"19",
		X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"17",X"1F",X"1D",X"1E",X"0A",X"0C",X"0F",X"0A",
		X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"1A",
		X"0A",X"1C",X"0B",X"1D",X"13",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"1E",X"0F",X"1D",X"9E",
		X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",X"0F",X"0A",X"1A",X"1C",X"19",X"1E",X"0F",X"0D",X"1E",
		X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"0D",X"19",X"16",X"19",X"1C",X"0A",X"1C",X"0B",
		X"17",X"0A",X"1E",X"0F",X"1D",X"9E",X"20",X"0F",X"1C",X"1E",X"13",X"0D",X"0B",X"16",X"0A",X"0C",
		X"0B",X"1C",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",X"0F",X"0A",X"0F",X"1C",X"1C",
		X"19",X"9C",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"1E",X"0F",X"1D",X"9E",X"0B",X"1F",X"1E",
		X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",X"1C",X"13",X"11",X"12",X"1E",
		X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",
		X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",X"10",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"0D",X"0F",
		X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",X"13",X"98",X"1D",X"16",X"0B",X"17",X"0A",X"1D",X"21",
		X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",
		X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",
		X"1E",X"0B",X"1C",X"9E",X"17",X"19",X"20",X"0F",X"0A",X"16",X"0F",X"10",X"9E",X"17",X"19",X"20",
		X"0F",X"0A",X"1C",X"13",X"11",X"12",X"9E",X"10",X"16",X"0B",X"9A",X"1D",X"19",X"1F",X"18",X"0E",
		X"0A",X"16",X"13",X"18",X"8F",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",X"18",X"11",
		X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",
		X"0A",X"0D",X"19",X"13",X"18",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1D",X"16",X"19",
		X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",
		X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1A",X"0B",X"13",X"0E",X"0A",X"0D",X"1C",X"0F",X"0E",
		X"13",X"1E",X"9D",X"10",X"1C",X"0F",X"0F",X"0A",X"17",X"0F",X"98",X"1E",X"19",X"1E",X"0B",X"16",
		X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"13",X"18",X"0A",X"17",X"13",X"18",X"1F",X"1E",X"0F",X"9D",
		X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"17",X"0F",X"18",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",
		X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1D",X"13",X"18",X"11",X"16",X"0F",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0E",X"1F",X"0B",X"16",X"0A",X"1A",X"16",
		X"0B",X"23",X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",
		X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",X"0B",X"11",X"0F",X"0A",
		X"1E",X"13",X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"11",
		X"0B",X"17",X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",X"1E",X"9D",X"0F",
		X"22",X"1E",X"1C",X"0B",X"0A",X"17",X"0B",X"18",X"0A",X"0F",X"20",X"0F",X"1C",X"A3",X"17",X"0F",
		X"18",X"0A",X"10",X"19",X"1C",X"0A",X"01",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"0A",X"11",
		X"0B",X"17",X"8F",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"19",
		X"0A",X"0E",X"0B",X"1E",X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",X"0F",X"8E",X"1A",X"1C",X"13",
		X"0D",X"13",X"18",X"11",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"0A",X"0A",
		X"0A",X"0A",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",
		X"9D",X"0A",X"0A",X"0A",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1D",X"16",X"19",X"1E",
		X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1F",X"18",
		X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",X"1C",
		X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",
		X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"0C",X"19",
		X"18",X"1F",X"1D",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"17",X"13",
		X"18",X"13",X"17",X"1F",X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"10",X"19",X"1C",X"0A",
		X"0B",X"18",X"23",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0E",X"13",X"10",X"10",X"13",X"0D",
		X"1F",X"16",X"1E",X"23",X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",X"16",X"0F",X"1E",X"1E",
		X"0F",X"1C",X"1D",X"0A",X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",
		X"1D",X"0D",X"19",X"1C",X"8F",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"0A",X"10",X"0B",X"0D",
		X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"9D",X"0D",X"16",X"0F",
		X"0B",X"1C",X"0A",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",
		X"19",X"1E",X"0B",X"16",X"9D",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",
		X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",
		X"0D",X"23",X"0D",X"16",X"8F",X"1D",X"0F",X"1E",X"0A",X"0B",X"1E",X"1E",X"1C",X"0B",X"0D",X"1E",
		X"0A",X"17",X"19",X"0E",X"0F",X"0A",X"17",X"0F",X"1D",X"1D",X"0B",X"11",X"8F",X"1D",X"0F",X"1E",
		X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"18",
		X"0B",X"17",X"8F",X"1F",X"1D",X"0F",X"0A",X"2C",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"01",
		X"0A",X"17",X"19",X"20",X"0F",X"2C",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",
		X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"02",X"0A",X"17",
		X"19",X"20",X"0F",X"2C",X"0A",X"1E",X"19",X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",X"0A",X"1E",
		X"12",X"0F",X"0A",X"20",X"0B",X"16",X"1F",X"8F",X"23",X"0F",X"9D",X"0B",X"0E",X"14",X"1F",X"1D",
		X"1E",X"17",X"0F",X"18",X"9E",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"1F",X"1D",X"0F",X"0A",X"2C",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"01",X"0A",X"10",X"16",X"0B",X"1A",X"2C",X"0A",X"1E",
		X"19",X"0A",X"0F",X"18",X"1E",X"0F",X"9C",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"10",
		X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"1D",X"0A",
		X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"8E",X"0C",X"23",X"0A",X"19",X"1A",X"0F",X"18",X"13",
		X"18",X"11",X"0A",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"19",X"1C",
		X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"9A",X"0B",X"18",X"0E",X"0A",X"1E",X"1F",
		X"1C",X"18",X"13",X"18",X"11",X"0A",X"11",X"0B",X"17",X"0F",X"0A",X"19",X"18",X"0A",X"0B",X"18",
		X"0E",X"0A",X"19",X"10",X"90",X"0A",X"0D",X"16",X"0F",X"0B",X"1C",X"0F",X"8E",X"12",X"13",X"11",
		X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",
		X"1D",X"0F",X"9E",X"0E",X"0B",X"13",X"16",X"23",X"0A",X"0C",X"1F",X"24",X"24",X"0B",X"1C",X"0E",
		X"9D",X"14",X"19",X"1F",X"1D",X"1E",X"0A",X"0D",X"12",X"0B",X"17",X"1A",X"13",X"19",X"18",X"9D",
		X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"1D",X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"1A",X"16",X"0B",
		X"23",X"0F",X"1C",X"0A",X"01",X"0A",X"17",X"19",X"20",X"0F",X"2C",X"0A",X"1E",X"19",X"0A",X"0D",
		X"0F",X"18",X"1E",X"0F",X"9C",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"13",X"18",X"0F",X"0A",
		X"0C",X"23",X"0A",X"1A",X"1C",X"0F",X"1D",X"1D",X"13",X"18",X"11",X"0A",X"0B",X"0E",X"20",X"0B",
		X"18",X"0D",X"8F",X"1A",X"1C",X"0F",X"1A",X"0B",X"1C",X"0F",X"0A",X"1E",X"19",X"0A",X"14",X"19",
		X"1F",X"1D",X"9E",X"0C",X"1F",X"24",X"24",X"0B",X"1C",X"0E",X"0A",X"0C",X"0B",X"13",X"1E",X"A9",
		X"1E",X"0F",X"0B",X"17",X"0A",X"21",X"0B",X"20",X"8F",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0B",
		X"21",X"0B",X"1C",X"0E",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"1E",X"0F",X"0B",X"17",X"0A",
		X"1A",X"16",X"0B",X"A3",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"0D",X"19",X"18",X"10",X"16",
		X"13",X"0D",X"1E",X"0A",X"27",X"0A",X"18",X"19",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0B",
		X"21",X"0B",X"1C",X"0E",X"0F",X"8E",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"0D",X"19",X"27",
		X"19",X"1A",X"0F",X"1C",X"0B",X"1E",X"13",X"19",X"18",X"0A",X"27",X"0A",X"0F",X"0B",X"0D",X"12",
		X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"03",X"00",X"00",X"00",X"0A",X"1A",X"19",X"13",
		X"18",X"1E",X"9D",X"21",X"0B",X"20",X"0F",X"8A",X"0C",X"0F",X"21",X"0B",X"1C",X"0F",X"0A",X"19",
		X"10",X"0A",X"1E",X"12",X"0F",X"0A",X"31",X"1F",X"18",X"0C",X"0F",X"0B",X"1E",X"0B",X"0C",X"16",
		X"0F",X"28",X"31",X"0A",X"1A",X"1E",X"0F",X"1C",X"19",X"0E",X"0B",X"0D",X"1E",X"23",X"96",X"11",
		X"16",X"0B",X"0E",X"13",X"0B",X"1E",X"19",X"1C",X"0A",X"21",X"0B",X"20",X"8F",X"03",X"00",X"00",
		X"00",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"0A",X"0C",X"19",X"1F",X"18",X"1E",X"A3",X"10",X"19",
		X"1C",X"0A",X"0E",X"13",X"1D",X"17",X"19",X"1F",X"18",X"1E",X"13",X"18",X"11",X"0A",X"10",X"13",
		X"1C",X"1D",X"1E",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"9C",X"18",X"19",X"0A",X"0C",X"19",X"1F",
		X"18",X"1E",X"23",X"0A",X"0B",X"21",X"0B",X"1C",X"0E",X"0F",X"8E",X"0D",X"19",X"16",X"16",X"0F",
		X"0D",X"1E",X"0F",X"0E",X"0A",X"03",X"00",X"00",X"00",X"0A",X"0C",X"19",X"1F",X"18",X"1E",X"A3",
		X"0F",X"11",X"11",X"0A",X"21",X"0B",X"20",X"8F",X"1D",X"1F",X"1C",X"20",X"13",X"20",X"0B",X"16",
		X"0A",X"21",X"0B",X"20",X"8F",X"0D",X"19",X"16",X"16",X"0F",X"0D",X"1E",X"0A",X"03",X"00",X"00",
		X"00",X"0A",X"1D",X"1F",X"1C",X"20",X"13",X"20",X"0B",X"16",X"0A",X"1A",X"19",X"13",X"18",X"1E",
		X"9D",X"18",X"19",X"0A",X"1D",X"1F",X"1C",X"20",X"13",X"20",X"0B",X"16",X"0A",X"1A",X"19",X"13",
		X"18",X"1E",X"1D",X"0A",X"0B",X"21",X"0B",X"1C",X"0E",X"0F",X"8E",X"0F",X"22",X"1E",X"1C",X"0B",
		X"0A",X"17",X"19",X"1F",X"18",X"1E",X"0A",X"0F",X"20",X"0F",X"1C",X"23",X"8A",X"2D",X"00",X"00",
		X"00",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"9D",X"12",X"19",X"17",X"0F",X"0A",X"19",X"10",X"0A",
		X"1E",X"12",X"8F",X"16",X"0B",X"20",X"0B",X"0A",X"1E",X"1C",X"19",X"16",X"96",X"1E",X"0F",X"17",
		X"1A",X"19",X"1C",X"0B",X"1C",X"23",X"0A",X"1D",X"0B",X"10",X"0F",X"1E",X"A3",X"1F",X"18",X"1E",
		X"13",X"16",X"0A",X"0B",X"0A",X"0D",X"19",X"18",X"1E",X"1C",X"19",X"16",X"0A",X"13",X"1D",X"0A",
		X"1A",X"1C",X"0F",X"1D",X"1D",X"0F",X"8E",X"03",X"AF",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",
		X"81",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"82",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1E",
		X"12",X"23",X"0A",X"18",X"0B",X"17",X"0F",X"0A",X"17",X"23",X"0A",X"16",X"19",X"1C",X"0E",X"A9",
		X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"13",X"18",X"13",X"1E",X"13",
		X"0B",X"16",X"9D",X"18",X"13",X"0D",X"0F",X"0A",X"14",X"19",X"1F",X"1D",X"1E",X"13",X"18",X"11",
		X"A9",X"17",X"0B",X"22",X"13",X"17",X"1F",X"17",X"0A",X"05",X"0A",X"0F",X"18",X"1E",X"1C",X"23",
		X"9D",X"1F",X"1D",X"0F",X"0A",X"27",X"17",X"19",X"20",X"0F",X"27",X"0A",X"1E",X"19",X"0A",X"1D",
		X"0F",X"16",X"0F",X"0D",X"1E",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",X"0A",X"0A",X"0A",X"0A",
		X"27",X"10",X"16",X"0B",X"1A",X"27",X"0A",X"1E",X"19",X"0A",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"2A",X"0D",X"2B",X"0A",X"01",X"09",X"08",X"02",X"0A",X"21",
		X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",
		X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",X"11",X"0B",X"17",X"0F",X"0A",X"19",X"20",X"0F",
		X"9C",X"0A",X"0A",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"21",X"0F",X"16",X"0D",
		X"19",X"17",X"0F",X"0A",X"1E",X"19",X"0A",X"14",X"19",X"1F",X"1D",X"9E",X"1E",X"19",X"0A",X"1D",
		X"1F",X"1C",X"20",X"13",X"20",X"0F",X"0A",X"0B",X"0A",X"14",X"19",X"1F",X"1D",X"9E",X"1E",X"12",
		X"0F",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"16",X"0B",X"18",X"0D",X"0F",X"0A",
		X"21",X"13",X"18",X"9D",X"13",X"18",X"0A",X"0B",X"0A",X"0D",X"19",X"16",X"16",X"13",X"1D",X"13",
		X"19",X"98",X"1A",X"13",X"0D",X"15",X"0A",X"1F",X"1A",X"0A",X"1E",X"12",X"0F",X"0A",X"0F",X"11",
		X"11",X"9D",X"0C",X"0F",X"10",X"19",X"1C",X"0F",X"0A",X"1E",X"12",X"0F",X"23",X"0A",X"12",X"0B",
		X"1E",X"0D",X"92",X"1E",X"19",X"0A",X"10",X"16",X"23",X"AD",X"1C",X"0F",X"1A",X"0F",X"0B",X"1E",
		X"0F",X"0E",X"16",X"23",X"0A",X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"1E",X"12",X"0F",X"0A",X"2C",
		X"10",X"16",X"0B",X"1A",X"2C",X"0A",X"0C",X"1F",X"1E",X"1E",X"19",X"98",X"17",X"0F",X"0F",X"1E",
		X"0A",X"1E",X"12",X"23",X"0A",X"0F",X"18",X"0F",X"17",X"13",X"0F",X"9D",X"0C",X"19",X"1F",X"18",
		X"0E",X"0F",X"1C",X"0A",X"2A",X"05",X"00",X"00",X"AB",X"12",X"1F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"2A",X"07",X"05",X"00",X"AB",X"1D",X"12",X"0B",X"0E",X"19",X"21",X"0A",X"16",X"19",X"1C",X"0E",
		X"0A",X"2A",X"01",X"05",X"00",X"00",X"AB",X"0A",X"1E",X"19",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",
		X"19",X"9C",X"13",X"18",X"1D",X"0F",X"1C",X"1E",X"0A",X"0B",X"0E",X"0E",X"13",X"1E",X"13",X"19",
		X"18",X"0B",X"16",X"0A",X"0D",X"19",X"13",X"18",X"1D",X"0A",X"10",X"19",X"9C",X"31",X"0E",X"1F",
		X"0B",X"16",X"0A",X"1A",X"16",X"0B",X"23",X"B1",X"1C",X"0F",X"0B",X"0E",X"23",X"0A",X"10",X"19",
		X"1C",X"8A",X"31",X"1D",X"13",X"18",X"11",X"16",X"0F",X"0A",X"1A",X"16",X"0B",X"23",X"B1",X"1A",
		X"1C",X"0F",X"1D",X"1D",X"8A",X"1E",X"12",X"13",X"1D",X"0A",X"13",X"1D",X"0A",X"14",X"19",X"1F",
		X"1D",X"1E",X"AE",X"0E",X"0F",X"1D",X"13",X"11",X"18",X"0F",X"0E",X"0A",X"0C",X"23",X"0A",X"21",
		X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",
		X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AE",X"0B",X"16",X"16",X"0A",X"1C",X"13",X"11",X"12",
		X"1E",X"1D",X"0A",X"1C",X"0F",X"1D",X"0F",X"1C",X"20",X"0F",X"8E",X"5D",X"B7",X"5D",X"C3",X"5D",
		X"CB",X"5D",X"D3",X"5D",X"D7",X"5D",X"E7",X"5D",X"EF",X"5D",X"F3",X"5D",X"F7",X"5D",X"FB",X"5E",
		X"0B",X"5E",X"1B",X"5E",X"2F",X"5E",X"33",X"5E",X"3B",X"5E",X"3F",X"5E",X"47",X"5E",X"57",X"5E",
		X"5B",X"5E",X"63",X"5E",X"6F",X"5E",X"77",X"5E",X"7B",X"5E",X"7F",X"5E",X"83",X"5E",X"93",X"5E",
		X"AB",X"5E",X"87",X"5E",X"B3",X"5E",X"8B",X"3E",X"50",X"99",X"09",X"36",X"90",X"33",X"0A",X"2E",
		X"A0",X"33",X"8B",X"2A",X"80",X"99",X"0D",X"30",X"80",X"99",X"8C",X"21",X"80",X"99",X"0E",X"37",
		X"80",X"99",X"8C",X"36",X"80",X"22",X"8F",X"36",X"80",X"22",X"0F",X"28",X"90",X"22",X"12",X"17",
		X"A0",X"99",X"10",X"17",X"A8",X"99",X"91",X"3A",X"80",X"33",X"13",X"24",X"B0",X"33",X"94",X"3A",
		X"20",X"88",X"95",X"2F",X"10",X"99",X"A3",X"2F",X"10",X"99",X"AF",X"23",X"D7",X"BB",X"42",X"5E",
		X"D7",X"BB",X"45",X"25",X"DF",X"44",X"43",X"34",X"E7",X"11",X"8B",X"28",X"16",X"BB",X"40",X"16",
		X"C0",X"33",X"42",X"6D",X"C0",X"33",X"46",X"20",X"D0",X"33",X"C7",X"30",X"80",X"22",X"45",X"4F",
		X"80",X"22",X"48",X"27",X"A0",X"22",X"3C",X"19",X"B0",X"22",X"4A",X"23",X"C0",X"22",X"CB",X"21",
		X"80",X"99",X"C9",X"24",X"60",X"33",X"23",X"59",X"60",X"33",X"CC",X"2A",X"40",X"88",X"CD",X"37",
		X"2A",X"11",X"4E",X"35",X"60",X"22",X"CF",X"28",X"16",X"BB",X"41",X"16",X"C0",X"33",X"42",X"6D",
		X"C0",X"33",X"46",X"20",X"D0",X"33",X"C7",X"34",X"20",X"22",X"EF",X"42",X"30",X"11",X"75",X"1B",
		X"40",X"11",X"F6",X"32",X"31",X"11",X"70",X"2E",X"41",X"11",X"71",X"38",X"51",X"11",X"F2",X"35",
		X"32",X"11",X"73",X"33",X"42",X"11",X"F4",X"34",X"33",X"11",X"F7",X"10",X"B6",X"44",X"F8",X"10",
		X"B6",X"DD",X"F9",X"10",X"B6",X"99",X"FA",X"11",X"46",X"11",X"DA",X"33",X"B0",X"11",X"5D",X"2A",
		X"B8",X"11",X"DE",X"24",X"57",X"11",X"62",X"36",X"57",X"55",X"63",X"5A",X"57",X"11",X"7B",X"49",
		X"77",X"11",X"7C",X"26",X"97",X"11",X"7D",X"3D",X"A7",X"77",X"FE",X"2E",X"77",X"11",X"7F",X"4D",
		X"77",X"77",X"FE",X"10",X"30",X"11",X"5F",X"10",X"40",X"11",X"60",X"10",X"50",X"11",X"6C",X"10",
		X"60",X"11",X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"62",X"7F",X"7E",X"62",X"4D",X"63",X"59",X"7E",X"63",X"2E",X"EF",X"24",X"7E",X"62",X"71",
		X"7E",X"63",X"36",X"7E",X"5E",X"EB",X"7E",X"63",X"3A",X"62",X"F1",X"86",X"7F",X"97",X"90",X"86",
		X"03",X"97",X"77",X"97",X"60",X"7E",X"63",X"E0",X"0F",X"8E",X"0F",X"8F",X"8E",X"AE",X"82",X"EC",
		X"84",X"84",X"80",X"C4",X"80",X"ED",X"81",X"8C",X"AF",X"E2",X"25",X"F3",X"86",X"01",X"BD",X"E0",
		X"37",X"8E",X"AF",X"E2",X"A6",X"84",X"84",X"20",X"A7",X"80",X"8C",X"B1",X"42",X"25",X"F5",X"CC",
		X"00",X"00",X"DD",X"97",X"ED",X"C8",X"18",X"ED",X"C8",X"1A",X"86",X"FF",X"97",X"6E",X"97",X"6F",
		X"97",X"70",X"BD",X"63",X"36",X"8E",X"5F",X"C5",X"AF",X"C8",X"2B",X"AE",X"C8",X"2B",X"30",X"05",
		X"AF",X"C8",X"2B",X"8C",X"60",X"10",X"10",X"24",X"03",X"21",X"A6",X"04",X"27",X"16",X"30",X"C8",
		X"18",X"A1",X"80",X"26",X"FC",X"6F",X"82",X"4D",X"2D",X"05",X"BD",X"4A",X"6A",X"20",X"05",X"84",
		X"7F",X"BD",X"4A",X"6D",X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"2B",X"A6",X"02",X"8D",X"41",
		X"86",X"08",X"BD",X"E0",X"37",X"AE",X"C8",X"2B",X"AD",X"94",X"AE",X"C8",X"2B",X"A6",X"03",X"A7",
		X"C8",X"2D",X"86",X"0A",X"A7",X"C8",X"33",X"A6",X"C8",X"18",X"8D",X"30",X"86",X"02",X"BD",X"E0",
		X"37",X"A6",X"C8",X"19",X"8D",X"26",X"86",X"02",X"BD",X"E0",X"37",X"A6",X"C8",X"1A",X"8D",X"1C",
		X"86",X"02",X"BD",X"E0",X"37",X"6A",X"C8",X"33",X"26",X"DD",X"6A",X"C8",X"2D",X"26",X"D3",X"20",
		X"8A",X"27",X"15",X"30",X"C8",X"18",X"6D",X"80",X"26",X"FC",X"A7",X"82",X"27",X"0A",X"2D",X"03",
		X"7E",X"4A",X"62",X"84",X"7F",X"7E",X"4A",X"65",X"39",X"39",X"5F",X"C9",X"11",X"02",X"00",X"60",
		X"10",X"12",X"09",X"00",X"60",X"74",X"13",X"07",X"12",X"60",X"DD",X"14",X"05",X"13",X"61",X"23",
		X"15",X"02",X"14",X"61",X"35",X"16",X"02",X"00",X"61",X"40",X"17",X"02",X"16",X"61",X"4B",X"18",
		X"01",X"17",X"5F",X"C9",X"00",X"01",X"15",X"5F",X"C9",X"00",X"05",X"18",X"5F",X"C9",X"9D",X"06",
		X"00",X"61",X"92",X"00",X"02",X"11",X"61",X"A7",X"1B",X"0A",X"9D",X"5F",X"C9",X"00",X"05",X"1B",
		X"CC",X"60",X"21",X"9E",X"75",X"ED",X"88",X"24",X"86",X"A0",X"A7",X"88",X"2D",X"A7",X"88",X"33",
		X"39",X"6A",X"C8",X"2D",X"2A",X"18",X"6C",X"C8",X"2D",X"EC",X"C8",X"11",X"10",X"83",X"FF",X"C0",
		X"2B",X"0C",X"A6",X"4B",X"81",X"78",X"22",X"12",X"CC",X"60",X"43",X"ED",X"C8",X"24",X"5F",X"4F",
		X"DD",X"32",X"39",X"A6",X"C8",X"11",X"2B",X"F6",X"20",X"E8",X"CC",X"60",X"5D",X"ED",X"C8",X"24",
		X"A6",X"C8",X"33",X"44",X"44",X"4C",X"A7",X"C8",X"2D",X"C6",X"01",X"20",X"E2",X"6A",X"C8",X"2D",
		X"26",X"F7",X"A6",X"C8",X"33",X"44",X"A7",X"C8",X"33",X"A7",X"C8",X"2D",X"CC",X"60",X"21",X"ED",
		X"C8",X"24",X"20",X"CA",X"8E",X"89",X"81",X"BD",X"60",X"A3",X"CC",X"7A",X"83",X"ED",X"A8",X"24",
		X"CC",X"01",X"23",X"ED",X"27",X"ED",X"A8",X"29",X"CC",X"00",X"81",X"ED",X"2A",X"E7",X"A8",X"27",
		X"E7",X"A8",X"28",X"E7",X"2F",X"CC",X"61",X"B9",X"9E",X"73",X"ED",X"88",X"24",X"86",X"60",X"A7",
		X"88",X"2D",X"39",X"34",X"10",X"DE",X"75",X"EE",X"C4",X"A6",X"42",X"81",X"20",X"26",X"F8",X"CC",
		X"8F",X"FF",X"8E",X"8E",X"C8",X"BD",X"E0",X"30",X"C6",X"07",X"6F",X"A5",X"5C",X"C1",X"36",X"25",
		X"F9",X"DE",X"2E",X"35",X"10",X"AF",X"2D",X"0C",X"A1",X"0C",X"AA",X"FC",X"00",X"1A",X"ED",X"A8",
		X"18",X"EC",X"98",X"0A",X"ED",X"A8",X"1A",X"86",X"04",X"A7",X"A8",X"33",X"39",X"CC",X"60",X"E6",
		X"9E",X"75",X"ED",X"88",X"24",X"39",X"EC",X"C8",X"20",X"27",X"0D",X"A6",X"C8",X"14",X"81",X"F8",
		X"27",X"15",X"CC",X"FF",X"00",X"DD",X"32",X"39",X"A6",X"C8",X"14",X"2E",X"05",X"CC",X"01",X"01",
		X"20",X"F3",X"CC",X"00",X"00",X"20",X"EE",X"CC",X"61",X"0D",X"ED",X"C8",X"24",X"A6",X"C8",X"14",
		X"2B",X"E0",X"CC",X"61",X"18",X"ED",X"C8",X"24",X"A6",X"C8",X"14",X"26",X"D5",X"A6",X"4F",X"2A",
		X"D1",X"20",X"DF",X"8E",X"74",X"DC",X"CC",X"F9",X"44",X"BD",X"4A",X"5C",X"8E",X"76",X"E3",X"CC",
		X"FA",X"44",X"7E",X"4A",X"5C",X"8E",X"89",X"81",X"BD",X"60",X"A3",X"CC",X"01",X"78",X"20",X"14",
		X"8E",X"89",X"B2",X"BD",X"60",X"A3",X"CC",X"00",X"F8",X"20",X"09",X"8E",X"89",X"E3",X"BD",X"60",
		X"A3",X"CC",X"00",X"80",X"ED",X"A8",X"2B",X"CC",X"00",X"08",X"ED",X"27",X"ED",X"A8",X"29",X"C6",
		X"D2",X"E7",X"2B",X"E7",X"A8",X"27",X"E7",X"A8",X"28",X"CC",X"61",X"70",X"ED",X"A8",X"24",X"39",
		X"EC",X"C8",X"2B",X"C3",X"FF",X"FF",X"ED",X"C8",X"2B",X"2F",X"0E",X"86",X"01",X"E6",X"C8",X"14",
		X"C1",X"02",X"26",X"01",X"4F",X"5F",X"DD",X"32",X"39",X"AE",X"4D",X"EC",X"02",X"ED",X"C8",X"24",
		X"20",X"F2",X"EE",X"C4",X"27",X"0E",X"A6",X"42",X"81",X"8F",X"26",X"F6",X"CC",X"EE",X"C2",X"ED",
		X"C8",X"24",X"20",X"EE",X"DE",X"2E",X"39",X"EE",X"C4",X"AE",X"C4",X"26",X"FA",X"CC",X"17",X"FF",
		X"8E",X"68",X"A5",X"BD",X"E0",X"30",X"DE",X"2E",X"39",X"A6",X"C8",X"2D",X"27",X"0E",X"6A",X"C8",
		X"2D",X"A6",X"C8",X"14",X"26",X"14",X"CC",X"01",X"00",X"DD",X"32",X"39",X"A6",X"C8",X"14",X"27",
		X"09",X"A6",X"4F",X"2B",X"05",X"CC",X"FF",X"00",X"20",X"EF",X"1F",X"31",X"AE",X"84",X"27",X"0A",
		X"A6",X"02",X"81",X"97",X"26",X"F6",X"A6",X"0F",X"A7",X"4F",X"CC",X"00",X"00",X"DD",X"32",X"39",
		X"86",X"80",X"97",X"B3",X"0F",X"90",X"86",X"08",X"BD",X"E0",X"37",X"8E",X"63",X"59",X"CC",X"48",
		X"00",X"BD",X"E0",X"09",X"BD",X"63",X"36",X"0F",X"8F",X"AE",X"9F",X"A0",X"0A",X"AE",X"84",X"27",
		X"1F",X"A6",X"02",X"2A",X"F8",X"81",X"97",X"27",X"F4",X"10",X"AE",X"0D",X"A6",X"02",X"10",X"AE",
		X"A4",X"10",X"AF",X"88",X"24",X"20",X"E6",X"8E",X"30",X"90",X"CC",X"00",X"11",X"7E",X"4A",X"53",
		X"86",X"0B",X"A7",X"4D",X"BD",X"62",X"27",X"86",X"08",X"BD",X"E0",X"37",X"6A",X"4D",X"26",X"F4",
		X"8E",X"A0",X"EA",X"6F",X"80",X"8C",X"A0",X"F2",X"25",X"F9",X"7E",X"3B",X"61",X"0F",X"B3",X"96",
		X"F5",X"27",X"08",X"8E",X"EF",X"21",X"BD",X"E0",X"2D",X"20",X"10",X"86",X"6D",X"A7",X"4D",X"BD",
		X"62",X"27",X"86",X"08",X"BD",X"E0",X"37",X"6A",X"4D",X"26",X"F4",X"CC",X"00",X"00",X"BD",X"E0",
		X"0C",X"8E",X"62",X"F1",X"BD",X"E0",X"15",X"86",X"04",X"BD",X"E0",X"37",X"BD",X"3B",X"2E",X"0F",
		X"90",X"86",X"31",X"A7",X"42",X"8E",X"63",X"59",X"CC",X"48",X"00",X"BD",X"E0",X"09",X"B6",X"CC",
		X"05",X"46",X"24",X"26",X"CC",X"03",X"84",X"ED",X"4D",X"6F",X"C8",X"10",X"8E",X"62",X"E9",X"BD",
		X"E0",X"15",X"BD",X"3B",X"43",X"BD",X"63",X"36",X"86",X"01",X"BD",X"E0",X"37",X"0C",X"11",X"EC",
		X"4D",X"27",X"07",X"C3",X"FF",X"FF",X"ED",X"4D",X"20",X"EE",X"BD",X"6B",X"A6",X"83",X"02",X"01",
		X"26",X"07",X"86",X"3C",X"A7",X"C8",X"10",X"20",X"DF",X"6A",X"C8",X"10",X"2E",X"DA",X"8E",X"62",
		X"DA",X"CC",X"49",X"00",X"BD",X"E0",X"09",X"7E",X"D0",X"00",X"86",X"05",X"BD",X"E0",X"37",X"BD",
		X"6B",X"A6",X"83",X"02",X"01",X"26",X"F3",X"20",X"82",X"00",X"07",X"C0",X"46",X"C0",X"3F",X"C0",
		X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"86",X"04",X"BD",X"E0",X"37",X"86",X"1E",X"A7",X"4D",X"BD",X"3B",X"2E",X"BE",X"E0",X"33",
		X"BD",X"E0",X"15",X"BD",X"63",X"36",X"86",X"19",X"D6",X"F2",X"5A",X"27",X"02",X"86",X"1A",X"BD",
		X"4A",X"62",X"86",X"3C",X"BD",X"E0",X"37",X"6A",X"4D",X"26",X"F7",X"7E",X"62",X"71",X"8E",X"EF",
		X"1B",X"BD",X"E0",X"2D",X"0C",X"B3",X"10",X"8E",X"12",X"00",X"CC",X"37",X"E2",X"8E",X"63",X"57",
		X"BD",X"87",X"93",X"CC",X"50",X"22",X"8E",X"38",X"E3",X"BD",X"4A",X"53",X"96",X"F2",X"85",X"F0",
		X"26",X"02",X"8A",X"F0",X"7E",X"4A",X"56",X"1F",X"09",X"CC",X"48",X"FF",X"BD",X"E0",X"0C",X"86",
		X"01",X"BD",X"E0",X"37",X"96",X"B3",X"2F",X"11",X"0F",X"B3",X"CC",X"00",X"00",X"BD",X"E0",X"0C",
		X"8E",X"63",X"01",X"CC",X"30",X"00",X"BD",X"E0",X"09",X"F6",X"C8",X"04",X"C4",X"30",X"27",X"DF",
		X"8E",X"CC",X"06",X"BD",X"3B",X"31",X"81",X"09",X"27",X"1E",X"96",X"F2",X"27",X"D1",X"81",X"02",
		X"24",X"04",X"C5",X"10",X"26",X"C9",X"C5",X"10",X"27",X"03",X"8B",X"99",X"19",X"8B",X"99",X"19",
		X"97",X"F2",X"8E",X"CD",X"00",X"BD",X"3B",X"3A",X"86",X"08",X"0F",X"60",X"C5",X"10",X"27",X"09",
		X"86",X"09",X"0C",X"60",X"C6",X"0A",X"BD",X"3B",X"2B",X"1F",X"89",X"BD",X"3B",X"2B",X"C6",X"0A",
		X"BD",X"3B",X"2B",X"8E",X"CC",X"02",X"BD",X"3B",X"34",X"BD",X"3B",X"55",X"D7",X"77",X"0F",X"90",
		X"CC",X"00",X"00",X"BD",X"E0",X"0C",X"86",X"30",X"A7",X"42",X"8E",X"EF",X"1E",X"BD",X"E0",X"2D",
		X"86",X"04",X"BD",X"E0",X"37",X"BD",X"3B",X"2E",X"BE",X"E0",X"33",X"BD",X"E0",X"15",X"CE",X"71",
		X"9B",X"AE",X"C1",X"EC",X"C1",X"80",X"30",X"88",X"5A",X"BD",X"4A",X"50",X"A6",X"C0",X"26",X"F5",
		X"DE",X"2E",X"8E",X"A0",X"4C",X"6F",X"80",X"8C",X"A0",X"60",X"25",X"F9",X"0F",X"36",X"0F",X"37",
		X"0F",X"AA",X"8E",X"CC",X"00",X"BD",X"3B",X"34",X"4F",X"58",X"49",X"58",X"49",X"58",X"49",X"58",
		X"49",X"DD",X"97",X"DD",X"54",X"DD",X"5E",X"8E",X"CC",X"14",X"BD",X"3B",X"31",X"6F",X"E2",X"81",
		X"03",X"23",X"08",X"6C",X"E4",X"81",X"06",X"23",X"02",X"6C",X"E4",X"8E",X"DE",X"11",X"10",X"8E",
		X"B1",X"AD",X"E6",X"E4",X"58",X"EC",X"85",X"ED",X"A4",X"86",X"02",X"A7",X"22",X"30",X"0E",X"31",
		X"23",X"8C",X"DF",X"99",X"25",X"EC",X"86",X"04",X"97",X"48",X"86",X"03",X"97",X"9F",X"86",X"01",
		X"97",X"A0",X"97",X"B0",X"86",X"5A",X"97",X"A7",X"0F",X"96",X"86",X"EA",X"97",X"9B",X"86",X"0D",
		X"97",X"3C",X"CC",X"00",X"00",X"DD",X"6E",X"DD",X"70",X"DD",X"73",X"DD",X"75",X"DD",X"38",X"DD",
		X"3A",X"0F",X"AF",X"0F",X"8E",X"0F",X"A1",X"8E",X"AE",X"82",X"EC",X"89",X"3A",X"B5",X"ED",X"81",
		X"8C",X"AF",X"E2",X"25",X"F5",X"86",X"01",X"BD",X"E0",X"37",X"8E",X"AF",X"E2",X"A6",X"89",X"3B",
		X"B6",X"8A",X"20",X"A7",X"80",X"8C",X"B1",X"42",X"25",X"F3",X"BD",X"E0",X"3A",X"86",X"01",X"BD",
		X"E0",X"37",X"10",X"8E",X"66",X"08",X"BD",X"65",X"EE",X"EC",X"A4",X"ED",X"84",X"10",X"8E",X"66",
		X"10",X"BD",X"65",X"EE",X"EC",X"A4",X"ED",X"84",X"96",X"90",X"2E",X"1F",X"CE",X"00",X"00",X"10",
		X"AE",X"C1",X"BD",X"65",X"EE",X"11",X"83",X"00",X"0E",X"25",X"F4",X"86",X"02",X"BD",X"E0",X"37",
		X"0A",X"90",X"8E",X"6B",X"C3",X"CC",X"11",X"FF",X"BD",X"E0",X"09",X"8E",X"83",X"7A",X"CC",X"20",
		X"FF",X"BD",X"E0",X"09",X"8E",X"8D",X"23",X"CC",X"09",X"00",X"BD",X"E0",X"09",X"FC",X"00",X"18",
		X"ED",X"A8",X"18",X"6F",X"2F",X"8E",X"00",X"64",X"AF",X"27",X"8E",X"88",X"8C",X"96",X"90",X"2E",
		X"03",X"8E",X"88",X"EE",X"AF",X"2D",X"96",X"77",X"BD",X"87",X"0E",X"96",X"60",X"27",X"2E",X"8E",
		X"8D",X"23",X"CC",X"09",X"00",X"BD",X"E0",X"09",X"FC",X"00",X"1C",X"ED",X"A8",X"18",X"C6",X"FF",
		X"E7",X"2F",X"8E",X"00",X"C8",X"AF",X"27",X"8E",X"88",X"BD",X"96",X"90",X"2E",X"03",X"8E",X"89",
		X"1F",X"AF",X"2D",X"96",X"77",X"BD",X"87",X"0E",X"86",X"08",X"BD",X"E0",X"37",X"8E",X"83",X"9F",
		X"CC",X"20",X"00",X"BD",X"E0",X"09",X"BE",X"E0",X"35",X"CC",X"68",X"FF",X"BD",X"E0",X"30",X"8E",
		X"EC",X"F8",X"CC",X"23",X"FF",X"BD",X"E0",X"09",X"8E",X"E7",X"85",X"CC",X"21",X"FF",X"BD",X"E0",
		X"09",X"CC",X"E7",X"1D",X"ED",X"2D",X"96",X"60",X"27",X"0E",X"8E",X"E7",X"85",X"CC",X"22",X"FF",
		X"BD",X"E0",X"09",X"CC",X"E7",X"51",X"ED",X"2D",X"96",X"90",X"10",X"2E",X"F9",X"6A",X"86",X"02",
		X"BD",X"E0",X"37",X"BD",X"6A",X"C7",X"8E",X"6B",X"20",X"CC",X"6F",X"00",X"BD",X"E0",X"09",X"86",
		X"FF",X"A7",X"42",X"6F",X"4D",X"6F",X"4F",X"0F",X"4B",X"86",X"02",X"BD",X"E0",X"37",X"96",X"4B",
		X"27",X"F7",X"EC",X"4E",X"8B",X"02",X"58",X"26",X"02",X"5C",X"4F",X"D5",X"4B",X"27",X"F5",X"ED",
		X"4E",X"D8",X"4B",X"D7",X"4B",X"10",X"AE",X"D8",X"0D",X"31",X"26",X"8D",X"21",X"E6",X"4F",X"2A",
		X"D8",X"86",X"01",X"BD",X"E0",X"37",X"10",X"BE",X"00",X"0E",X"31",X"2C",X"8D",X"10",X"86",X"01",
		X"BD",X"E0",X"37",X"10",X"BE",X"00",X"0E",X"31",X"A8",X"12",X"8D",X"02",X"20",X"BB",X"E6",X"27",
		X"C8",X"04",X"EB",X"25",X"BD",X"E0",X"1E",X"86",X"0A",X"A7",X"84",X"EC",X"24",X"ED",X"04",X"EC",
		X"22",X"ED",X"02",X"EC",X"26",X"ED",X"06",X"39",X"12",X"88",X"00",X"00",X"00",X"D3",X"1F",X"07",
		X"12",X"88",X"00",X"00",X"78",X"D3",X"1A",X"07",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",
		X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",
		X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"20",X"99",X"67",X"09",
		X"6A",X"C8",X"2F",X"26",X"2C",X"A6",X"C8",X"35",X"A7",X"C8",X"2F",X"6F",X"C8",X"2E",X"BD",X"80",
		X"D6",X"10",X"27",X"00",X"9F",X"A6",X"C8",X"35",X"81",X"0F",X"23",X"03",X"6A",X"C8",X"35",X"EC",
		X"07",X"ED",X"C8",X"2B",X"E6",X"0B",X"C1",X"D2",X"25",X"02",X"C6",X"D2",X"C0",X"05",X"BD",X"D7",
		X"BD",X"E6",X"C8",X"2E",X"27",X"7E",X"E1",X"4B",X"10",X"25",X"00",X"FD",X"C0",X"0F",X"E1",X"4B",
		X"10",X"22",X"01",X"1E",X"86",X"80",X"BD",X"D7",X"A8",X"8E",X"EF",X"7D",X"BD",X"E0",X"2D",X"CC",
		X"66",X"95",X"ED",X"C8",X"24",X"BD",X"D7",X"70",X"27",X"13",X"EC",X"C8",X"2B",X"A3",X"47",X"2B",
		X"07",X"83",X"00",X"0D",X"2A",X"14",X"20",X"05",X"C3",X"00",X"0D",X"2B",X"0D",X"CC",X"66",X"40",
		X"ED",X"C8",X"24",X"6F",X"C8",X"2E",X"5F",X"7E",X"67",X"55",X"A6",X"C8",X"17",X"81",X"18",X"26",
		X"05",X"86",X"0A",X"A7",X"C8",X"15",X"A6",X"4B",X"A1",X"C8",X"2E",X"27",X"22",X"25",X"10",X"A6",
		X"C8",X"11",X"2B",X"09",X"EC",X"C8",X"11",X"83",X"00",X"10",X"ED",X"C8",X"11",X"20",X"76",X"A6",
		X"C8",X"11",X"2E",X"71",X"EC",X"C8",X"11",X"C3",X"00",X"10",X"ED",X"C8",X"11",X"20",X"66",X"6F",
		X"C8",X"11",X"20",X"61",X"86",X"43",X"E6",X"4B",X"C1",X"65",X"25",X"08",X"86",X"7F",X"C1",X"A1",
		X"BD",X"D7",X"8C",X"12",X"A0",X"4B",X"27",X"24",X"2B",X"11",X"EC",X"C8",X"11",X"10",X"83",X"01",
		X"00",X"2C",X"23",X"C3",X"00",X"20",X"ED",X"C8",X"11",X"20",X"1B",X"EC",X"C8",X"11",X"10",X"83",
		X"FF",X"00",X"2F",X"12",X"83",X"00",X"20",X"ED",X"C8",X"11",X"20",X"0A",X"EC",X"C8",X"11",X"47",
		X"56",X"47",X"56",X"ED",X"C8",X"11",X"6D",X"C8",X"22",X"27",X"06",X"2B",X"0B",X"86",X"04",X"20",
		X"09",X"86",X"04",X"6D",X"C8",X"14",X"2A",X"02",X"86",X"FC",X"A7",X"C8",X"14",X"A7",X"4F",X"CC",
		X"00",X"00",X"DD",X"32",X"39",X"A6",X"4F",X"A7",X"C8",X"14",X"6D",X"C8",X"22",X"27",X"06",X"2B",
		X"0B",X"86",X"08",X"20",X"09",X"86",X"08",X"6D",X"C8",X"14",X"2A",X"02",X"86",X"F8",X"A7",X"C8",
		X"14",X"A7",X"4F",X"CC",X"00",X"00",X"DD",X"32",X"39",X"EC",X"C8",X"11",X"10",X"83",X"FF",X"40",
		X"2F",X"06",X"C3",X"FF",X"C0",X"ED",X"C8",X"11",X"CC",X"67",X"95",X"ED",X"C8",X"24",X"86",X"02",
		X"A7",X"C8",X"2D",X"20",X"A1",X"6A",X"C8",X"2D",X"2E",X"9C",X"CC",X"66",X"40",X"ED",X"C8",X"24",
		X"20",X"94",X"EC",X"C8",X"11",X"10",X"83",X"01",X"00",X"2C",X"DD",X"C3",X"00",X"10",X"ED",X"C8",
		X"11",X"20",X"D5",X"EC",X"47",X"10",X"83",X"FF",X"F9",X"2D",X"4D",X"10",X"83",X"01",X"21",X"2E",
		X"47",X"86",X"43",X"E6",X"4B",X"C1",X"65",X"25",X"08",X"86",X"7F",X"C1",X"A1",X"25",X"02",X"86",
		X"CE",X"A0",X"4B",X"27",X"26",X"2B",X"12",X"EC",X"C8",X"11",X"10",X"83",X"01",X"00",X"2C",X"06",
		X"C3",X"00",X"20",X"ED",X"C8",X"11",X"7E",X"67",X"55",X"EC",X"C8",X"11",X"10",X"83",X"FF",X"00",
		X"2F",X"06",X"83",X"00",X"20",X"ED",X"C8",X"11",X"7E",X"67",X"55",X"EC",X"C8",X"11",X"47",X"56",
		X"47",X"56",X"ED",X"C8",X"11",X"7E",X"67",X"55",X"BD",X"8E",X"8E",X"86",X"7F",X"A4",X"42",X"A7",
		X"42",X"86",X"3C",X"BD",X"E0",X"37",X"7E",X"E0",X"0F",X"C6",X"0C",X"E7",X"C8",X"17",X"BD",X"69",
		X"51",X"86",X"04",X"BD",X"E0",X"37",X"20",X"0C",X"63",X"4F",X"A6",X"C8",X"34",X"27",X"05",X"0A",
		X"AB",X"BD",X"D7",X"68",X"BD",X"8E",X"8E",X"C6",X"18",X"E7",X"C8",X"17",X"BD",X"69",X"51",X"86",
		X"04",X"BD",X"E0",X"37",X"BD",X"8E",X"8E",X"A6",X"C8",X"2D",X"84",X"FC",X"26",X"02",X"6F",X"4F",
		X"6A",X"C8",X"2D",X"2A",X"C4",X"86",X"03",X"A7",X"C8",X"12",X"FC",X"00",X"38",X"ED",X"C8",X"13",
		X"10",X"AE",X"C8",X"13",X"8D",X"2F",X"86",X"02",X"BD",X"E0",X"37",X"10",X"AE",X"C8",X"13",X"8D",
		X"24",X"10",X"AF",X"C8",X"13",X"86",X"06",X"BD",X"E0",X"37",X"6A",X"C8",X"12",X"26",X"E1",X"BD",
		X"8E",X"8E",X"CC",X"12",X"00",X"ED",X"84",X"86",X"02",X"BD",X"E0",X"37",X"CC",X"04",X"44",X"ED",
		X"C8",X"2E",X"7E",X"78",X"61",X"EC",X"47",X"46",X"56",X"1F",X"98",X"E6",X"4B",X"C0",X"0A",X"ED",
		X"C8",X"10",X"7E",X"82",X"09",X"6F",X"C8",X"34",X"A6",X"C8",X"34",X"C6",X"07",X"6F",X"C5",X"5C",
		X"C1",X"36",X"25",X"F9",X"A7",X"C8",X"34",X"86",X"02",X"A7",X"C8",X"14",X"8E",X"FF",X"F7",X"BD",
		X"E0",X"18",X"24",X"08",X"63",X"4F",X"60",X"C8",X"14",X"8E",X"01",X"23",X"AF",X"47",X"CC",X"00",
		X"00",X"DD",X"88",X"0F",X"8A",X"9E",X"73",X"27",X"0A",X"BD",X"D8",X"00",X"9E",X"75",X"27",X"03",
		X"BD",X"D8",X"00",X"8E",X"00",X"D1",X"96",X"8A",X"27",X"0A",X"8E",X"00",X"80",X"96",X"89",X"27",
		X"03",X"8E",X"00",X"3D",X"AF",X"4A",X"CC",X"66",X"40",X"ED",X"C8",X"24",X"8E",X"EF",X"78",X"BD",
		X"E0",X"2D",X"86",X"80",X"AA",X"42",X"A7",X"42",X"86",X"80",X"A7",X"C8",X"26",X"CC",X"8A",X"14",
		X"ED",X"4D",X"86",X"78",X"A7",X"C8",X"35",X"44",X"BD",X"D7",X"81",X"6F",X"C8",X"13",X"20",X"08",
		X"86",X"01",X"BD",X"E0",X"37",X"BD",X"D8",X"3D",X"6A",X"C8",X"15",X"2E",X"17",X"E6",X"C8",X"10",
		X"C0",X"02",X"2A",X"02",X"C6",X"06",X"E7",X"C8",X"10",X"8E",X"69",X"BF",X"EC",X"85",X"A7",X"C8",
		X"17",X"E7",X"C8",X"15",X"8E",X"69",X"CF",X"EC",X"C8",X"11",X"BD",X"D8",X"61",X"8D",X"02",X"20",
		X"CF",X"E6",X"C8",X"17",X"A6",X"4F",X"2A",X"02",X"CB",X"06",X"BE",X"00",X"34",X"3A",X"AF",X"C8",
		X"1C",X"E6",X"4B",X"C1",X"D2",X"25",X"0A",X"6F",X"C8",X"11",X"6F",X"C8",X"12",X"C6",X"D2",X"E7",
		X"4B",X"E7",X"C8",X"27",X"C0",X"0A",X"E7",X"C8",X"28",X"EC",X"47",X"C3",X"00",X"1B",X"ED",X"C8",
		X"29",X"BD",X"8E",X"83",X"96",X"AA",X"27",X"0E",X"96",X"AC",X"27",X"18",X"A6",X"C8",X"34",X"27",
		X"13",X"6F",X"C8",X"34",X"0A",X"AB",X"EC",X"C8",X"24",X"83",X"67",X"B3",X"24",X"06",X"CC",X"67",
		X"B3",X"ED",X"C8",X"24",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"AE",X"A2",X"AA",X"89",X"AE",
		X"AC",X"A4",X"A9",X"E8",X"3D",X"A4",X"A9",X"E8",X"3E",X"27",X"03",X"7E",X"DA",X"3E",X"39",X"00",
		X"08",X"0C",X"08",X"18",X"08",X"0C",X"08",X"FD",X"00",X"FE",X"80",X"FF",X"40",X"FF",X"A0",X"00",
		X"00",X"00",X"60",X"00",X"C0",X"01",X"80",X"03",X"00",X"5F",X"BD",X"6A",X"F3",X"BD",X"6A",X"93",
		X"ED",X"47",X"A6",X"C8",X"10",X"6A",X"C8",X"2D",X"2E",X"12",X"B6",X"B1",X"AE",X"A7",X"C8",X"2D",
		X"A6",X"C8",X"10",X"81",X"1E",X"27",X"10",X"8B",X"06",X"A7",X"C8",X"10",X"BD",X"6B",X"06",X"86",
		X"01",X"8E",X"69",X"DA",X"7E",X"E0",X"12",X"E6",X"2B",X"CB",X"03",X"E1",X"4B",X"27",X"1A",X"22",
		X"04",X"6A",X"4B",X"20",X"02",X"6C",X"4B",X"BD",X"6B",X"06",X"86",X"01",X"BD",X"E0",X"37",X"BD",
		X"6A",X"F3",X"BD",X"6A",X"93",X"ED",X"47",X"20",X"DE",X"8E",X"EF",X"83",X"BD",X"E0",X"2D",X"EC",
		X"42",X"4C",X"EE",X"C4",X"8E",X"D9",X"16",X"AF",X"C8",X"30",X"8E",X"6A",X"66",X"BD",X"E0",X"30",
		X"DE",X"2E",X"EC",X"47",X"ED",X"27",X"EC",X"4A",X"ED",X"2A",X"EC",X"C8",X"24",X"ED",X"A8",X"24",
		X"EF",X"A8",X"2B",X"CC",X"00",X"00",X"BD",X"D7",X"EA",X"86",X"02",X"BD",X"E0",X"37",X"BD",X"6A",
		X"93",X"20",X"F6",X"BD",X"6A",X"F3",X"10",X"9E",X"2C",X"BD",X"6A",X"9B",X"26",X"22",X"AE",X"C8",
		X"2B",X"ED",X"47",X"ED",X"07",X"EC",X"2A",X"CB",X"0A",X"ED",X"4A",X"ED",X"0A",X"86",X"24",X"A7",
		X"C8",X"10",X"BD",X"6B",X"06",X"8E",X"6A",X"63",X"86",X"01",X"7E",X"D7",X"C8",X"BD",X"6A",X"F3",
		X"7E",X"E0",X"0F",X"8D",X"03",X"26",X"42",X"39",X"10",X"AE",X"C4",X"10",X"AC",X"C8",X"24",X"26",
		X"23",X"A6",X"22",X"2A",X"1F",X"A6",X"A8",X"20",X"26",X"1A",X"A6",X"2B",X"81",X"C6",X"25",X"14",
		X"EC",X"27",X"C3",X"FF",X"FE",X"10",X"83",X"00",X"28",X"2F",X"06",X"10",X"83",X"00",X"F0",X"2D",
		X"03",X"1A",X"04",X"39",X"1C",X"FB",X"39",X"BE",X"6B",X"C1",X"4F",X"AB",X"82",X"8C",X"D0",X"00",
		X"26",X"F9",X"88",X"A1",X"27",X"02",X"0C",X"B2",X"39",X"A6",X"C8",X"10",X"8B",X"FA",X"A7",X"C8",
		X"10",X"2F",X"0B",X"BD",X"6B",X"06",X"86",X"05",X"8E",X"69",X"DA",X"7E",X"E0",X"12",X"0A",X"96",
		X"7E",X"E0",X"0F",X"10",X"AE",X"C8",X"1C",X"27",X"0C",X"6F",X"C8",X"1C",X"6F",X"C8",X"1D",X"BD",
		X"8E",X"9F",X"7E",X"D8",X"F4",X"39",X"A6",X"C8",X"10",X"80",X"06",X"2B",X"F8",X"10",X"BE",X"00",
		X"2A",X"31",X"A6",X"10",X"AF",X"C8",X"1C",X"BD",X"E0",X"24",X"BD",X"8E",X"70",X"7E",X"D8",X"F4",
		X"86",X"1E",X"BD",X"E0",X"37",X"CC",X"25",X"02",X"8D",X"66",X"26",X"F4",X"8D",X"62",X"27",X"FC",
		X"86",X"0F",X"BD",X"E0",X"37",X"CC",X"12",X"04",X"8D",X"56",X"26",X"E4",X"8D",X"52",X"27",X"FC",
		X"86",X"0F",X"BD",X"E0",X"37",X"CC",X"05",X"06",X"8D",X"46",X"26",X"E0",X"BD",X"3B",X"2E",X"1A",
		X"FF",X"CC",X"00",X"FF",X"FD",X"C0",X"00",X"CE",X"73",X"AB",X"8E",X"10",X"30",X"34",X"10",X"C6",
		X"11",X"A6",X"C0",X"88",X"9B",X"80",X"35",X"2B",X"10",X"27",X"05",X"BD",X"4A",X"50",X"20",X"F1",
		X"AE",X"E4",X"30",X"88",X"10",X"AF",X"E4",X"20",X"E8",X"8E",X"1B",X"E6",X"86",X"39",X"B7",X"CB",
		X"FF",X"8D",X"23",X"83",X"05",X"06",X"27",X"F1",X"30",X"1F",X"26",X"F0",X"6E",X"9F",X"FF",X"FE",
		X"ED",X"4D",X"EC",X"E1",X"ED",X"4F",X"86",X"01",X"BD",X"E0",X"37",X"8D",X"09",X"1F",X"01",X"EC",
		X"4D",X"AC",X"4D",X"6E",X"D8",X"0F",X"86",X"08",X"BA",X"C8",X"07",X"B7",X"C8",X"07",X"B6",X"C8",
		X"04",X"84",X"37",X"C6",X"F7",X"F4",X"C8",X"07",X"F7",X"C8",X"07",X"F6",X"C8",X"04",X"C4",X"07",
		X"39",X"90",X"00",X"0F",X"9E",X"CC",X"71",X"C8",X"ED",X"C8",X"13",X"CC",X"70",X"2F",X"ED",X"47",
		X"86",X"02",X"A7",X"C8",X"1C",X"86",X"20",X"BD",X"E0",X"37",X"20",X"5C",X"96",X"3C",X"27",X"02",
		X"0A",X"3C",X"8E",X"CC",X"14",X"BD",X"3B",X"31",X"A7",X"E2",X"8E",X"DE",X"11",X"10",X"8E",X"B1",
		X"AD",X"E6",X"22",X"27",X"04",X"6A",X"22",X"26",X"2A",X"E6",X"E4",X"CB",X"10",X"57",X"E6",X"85",
		X"25",X"04",X"54",X"54",X"54",X"54",X"C4",X"0F",X"E7",X"22",X"E6",X"0D",X"1D",X"2B",X"09",X"E3",
		X"A4",X"10",X"A3",X"06",X"2D",X"0B",X"20",X"07",X"E3",X"A4",X"10",X"A3",X"06",X"2E",X"02",X"EC",
		X"06",X"ED",X"A4",X"30",X"0E",X"31",X"23",X"8C",X"DF",X"99",X"25",X"C5",X"35",X"02",X"96",X"9B",
		X"81",X"E0",X"23",X"04",X"80",X"05",X"97",X"9B",X"96",X"9F",X"27",X"2C",X"0A",X"9F",X"26",X"66",
		X"BD",X"6E",X"01",X"CC",X"FF",X"E0",X"ED",X"A8",X"2B",X"86",X"01",X"A7",X"A8",X"14",X"86",X"01",
		X"A7",X"A8",X"2D",X"BD",X"6E",X"01",X"CC",X"01",X"3F",X"ED",X"A8",X"2B",X"86",X"07",X"A7",X"A8",
		X"14",X"86",X"FF",X"A7",X"A8",X"2D",X"20",X"3E",X"96",X"A0",X"27",X"3A",X"0A",X"A0",X"26",X"36",
		X"8E",X"86",X"D0",X"CC",X"69",X"FF",X"DE",X"0A",X"BD",X"E0",X"30",X"CC",X"00",X"EF",X"ED",X"2A",
		X"CC",X"00",X"14",X"ED",X"27",X"6F",X"A8",X"10",X"8E",X"86",X"D0",X"CC",X"69",X"FF",X"BD",X"E0",
		X"30",X"DE",X"2E",X"CC",X"00",X"EF",X"ED",X"2A",X"CC",X"01",X"06",X"ED",X"27",X"86",X"02",X"A7",
		X"A8",X"10",X"86",X"04",X"A7",X"24",X"0F",X"36",X"0F",X"37",X"0F",X"8F",X"86",X"FF",X"97",X"A2",
		X"86",X"01",X"97",X"B0",X"6F",X"C8",X"1F",X"6F",X"C8",X"23",X"6F",X"C8",X"27",X"6F",X"C8",X"2B",
		X"6F",X"C8",X"2F",X"6F",X"C8",X"33",X"96",X"9E",X"8B",X"01",X"19",X"97",X"9E",X"AD",X"D8",X"13",
		X"BD",X"D7",X"61",X"86",X"01",X"BD",X"E0",X"37",X"BD",X"6F",X"AC",X"CC",X"71",X"C8",X"ED",X"C8",
		X"13",X"AE",X"47",X"A6",X"03",X"30",X"04",X"8C",X"71",X"9B",X"25",X"03",X"8E",X"71",X"73",X"AF",
		X"47",X"A8",X"03",X"84",X"F0",X"27",X"1A",X"E6",X"03",X"8E",X"6F",X"CB",X"BD",X"6E",X"F0",X"8E",
		X"6F",X"D2",X"BD",X"6E",X"F0",X"8E",X"6F",X"D9",X"BD",X"6E",X"F0",X"8E",X"6F",X"E0",X"BD",X"6E",
		X"F0",X"AE",X"47",X"A6",X"03",X"85",X"01",X"27",X"06",X"A6",X"01",X"84",X"0F",X"97",X"8F",X"E6",
		X"03",X"C4",X"0E",X"8E",X"71",X"BC",X"AD",X"95",X"86",X"1E",X"BD",X"6E",X"64",X"BD",X"6E",X"53",
		X"BD",X"6E",X"C4",X"A6",X"D8",X"07",X"44",X"44",X"44",X"44",X"27",X"06",X"8E",X"89",X"81",X"BD",
		X"6E",X"17",X"A6",X"D8",X"07",X"84",X"0F",X"27",X"06",X"8E",X"89",X"B2",X"BD",X"6E",X"17",X"AE",
		X"47",X"A6",X"01",X"44",X"44",X"44",X"44",X"27",X"06",X"8E",X"89",X"E3",X"BD",X"6E",X"17",X"96",
		X"90",X"27",X"08",X"AE",X"47",X"A6",X"01",X"84",X"0F",X"97",X"8F",X"A6",X"C8",X"1C",X"27",X"03",
		X"6A",X"C8",X"1C",X"8E",X"6D",X"FE",X"A6",X"86",X"A7",X"C8",X"1B",X"4C",X"48",X"8E",X"6D",X"E2",
		X"EC",X"86",X"DD",X"AD",X"0F",X"AB",X"0F",X"AC",X"86",X"70",X"A7",X"4B",X"86",X"08",X"BD",X"E0",
		X"37",X"30",X"C4",X"96",X"AA",X"10",X"27",X"FE",X"43",X"96",X"AC",X"27",X"04",X"0A",X"AC",X"26",
		X"2D",X"DC",X"AD",X"83",X"00",X"01",X"2E",X"24",X"96",X"AB",X"81",X"02",X"22",X"20",X"8E",X"68",
		X"A8",X"CC",X"17",X"FF",X"BD",X"E0",X"09",X"0C",X"AB",X"86",X"FF",X"A7",X"A8",X"34",X"A6",X"C8",
		X"1B",X"27",X"03",X"6A",X"C8",X"1B",X"48",X"8E",X"6D",X"E2",X"EC",X"86",X"DD",X"AD",X"96",X"A1",
		X"27",X"BA",X"6A",X"4B",X"26",X"B6",X"96",X"90",X"27",X"AE",X"0C",X"8F",X"26",X"AA",X"0A",X"8F",
		X"20",X"A6",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",X"16",
		X"00",X"25",X"00",X"34",X"00",X"70",X"00",X"70",X"00",X"E1",X"01",X"51",X"01",X"C2",X"0A",X"0B",
		X"0C",X"DE",X"2C",X"8E",X"86",X"38",X"CC",X"6A",X"FF",X"BD",X"E0",X"30",X"DE",X"2E",X"CC",X"00",
		X"DF",X"ED",X"2A",X"6F",X"A8",X"10",X"39",X"A7",X"4B",X"EC",X"E1",X"ED",X"C8",X"11",X"AF",X"4D",
		X"86",X"3D",X"BD",X"E0",X"37",X"8E",X"8B",X"0E",X"CC",X"0F",X"FF",X"BD",X"E0",X"09",X"0C",X"A1",
		X"0C",X"AA",X"EC",X"4D",X"ED",X"2D",X"FC",X"00",X"1A",X"ED",X"A8",X"18",X"86",X"04",X"A7",X"A8",
		X"33",X"6F",X"A8",X"34",X"96",X"9F",X"27",X"04",X"86",X"02",X"97",X"B0",X"6A",X"4B",X"26",X"D0",
		X"6E",X"D8",X"11",X"AE",X"E1",X"AF",X"4F",X"8D",X"1A",X"96",X"90",X"27",X"04",X"AE",X"C4",X"26",
		X"F6",X"6E",X"D8",X"0F",X"AE",X"E1",X"AF",X"4F",X"A7",X"4B",X"8D",X"07",X"6A",X"4B",X"26",X"FA",
		X"6E",X"D8",X"0F",X"35",X"06",X"ED",X"C8",X"11",X"96",X"90",X"27",X"24",X"86",X"23",X"A7",X"C8",
		X"1E",X"A6",X"C8",X"1F",X"27",X"03",X"BD",X"6F",X"AC",X"86",X"01",X"BD",X"E0",X"37",X"A6",X"C8",
		X"1E",X"81",X"33",X"22",X"0B",X"31",X"C6",X"8B",X"04",X"A7",X"C8",X"1E",X"8D",X"1A",X"20",X"E9",
		X"6E",X"D8",X"11",X"31",X"C8",X"1F",X"31",X"24",X"6D",X"A4",X"26",X"FA",X"96",X"90",X"27",X"13",
		X"EC",X"84",X"ED",X"A4",X"EC",X"02",X"ED",X"22",X"A6",X"A4",X"27",X"07",X"E6",X"21",X"AE",X"22",
		X"7E",X"4A",X"53",X"39",X"A6",X"C8",X"1F",X"27",X"03",X"BD",X"6F",X"B4",X"31",X"C8",X"23",X"8D",
		X"12",X"31",X"C8",X"27",X"8D",X"0D",X"31",X"C8",X"2B",X"8D",X"08",X"31",X"C8",X"2F",X"8D",X"03",
		X"31",X"C8",X"33",X"A6",X"A4",X"27",X"08",X"6F",X"A4",X"5F",X"AE",X"22",X"7E",X"4A",X"53",X"39",
		X"34",X"16",X"A5",X"84",X"27",X"48",X"E5",X"84",X"27",X"46",X"10",X"AE",X"05",X"27",X"04",X"86",
		X"FF",X"A7",X"A4",X"A6",X"01",X"27",X"21",X"43",X"8E",X"AF",X"E2",X"10",X"8E",X"01",X"60",X"BD",
		X"6F",X"A1",X"AE",X"62",X"A6",X"02",X"43",X"94",X"4B",X"97",X"4B",X"A6",X"02",X"43",X"8E",X"AE",
		X"82",X"10",X"8E",X"01",X"60",X"BD",X"6F",X"A1",X"8E",X"EF",X"6A",X"BD",X"E0",X"2D",X"8E",X"81",
		X"A0",X"CC",X"27",X"FF",X"BD",X"E0",X"09",X"AE",X"62",X"EC",X"98",X"03",X"ED",X"2E",X"35",X"96",
		X"10",X"AE",X"05",X"27",X"02",X"6F",X"A4",X"A6",X"01",X"A7",X"E2",X"8E",X"AF",X"E2",X"10",X"8E",
		X"EB",X"98",X"A6",X"E4",X"43",X"A4",X"84",X"A7",X"84",X"A6",X"E4",X"A4",X"A0",X"AB",X"84",X"A7",
		X"80",X"8C",X"B1",X"42",X"25",X"EC",X"AE",X"63",X"A6",X"02",X"A7",X"E4",X"9A",X"4B",X"97",X"4B",
		X"8E",X"AE",X"82",X"10",X"8E",X"E9",X"37",X"A6",X"E4",X"43",X"A4",X"84",X"A7",X"84",X"A6",X"E4",
		X"A4",X"A0",X"AB",X"84",X"A7",X"80",X"8C",X"AF",X"E2",X"25",X"EC",X"A6",X"E0",X"35",X"16",X"ED",
		X"C8",X"15",X"EC",X"E1",X"ED",X"4F",X"86",X"01",X"BD",X"E0",X"37",X"EC",X"C8",X"15",X"6E",X"D8",
		X"0F",X"1F",X"89",X"E4",X"84",X"E7",X"80",X"31",X"3F",X"26",X"F6",X"39",X"CC",X"59",X"11",X"A7",
		X"C8",X"1F",X"20",X"06",X"CC",X"59",X"00",X"6F",X"C8",X"1F",X"8E",X"3A",X"60",X"BD",X"4A",X"53",
		X"96",X"9E",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"7E",X"4A",X"56",X"10",X"01",X"03",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"00",X"40",X"02",X"04",X"00",X"04",X"A0",X"6E",
		X"80",X"10",X"40",X"00",X"0C",X"00",X"00",X"53",X"11",X"2D",X"7D",X"54",X"11",X"33",X"9B",X"55",
		X"11",X"36",X"7D",X"56",X"11",X"1C",X"9B",X"57",X"11",X"1A",X"B6",X"58",X"11",X"0B",X"B6",X"FD",
		X"11",X"31",X"7D",X"FF",X"11",X"26",X"B6",X"FE",X"55",X"08",X"B6",X"FE",X"77",X"3F",X"B6",X"5B",
		X"11",X"30",X"7F",X"5C",X"11",X"2E",X"90",X"F5",X"11",X"1C",X"9B",X"F6",X"11",X"32",X"B6",X"FB",
		X"55",X"10",X"B6",X"FB",X"77",X"4F",X"B6",X"FC",X"11",X"38",X"7D",X"5A",X"11",X"11",X"78",X"40",
		X"01",X"00",X"00",X"30",X"01",X"00",X"02",X"40",X"01",X"00",X"04",X"60",X"02",X"00",X"00",X"33",
		X"01",X"00",X"06",X"60",X"01",X"00",X"08",X"33",X"03",X"00",X"41",X"24",X"02",X"00",X"75",X"06",
		X"01",X"01",X"7B",X"06",X"02",X"00",X"F7",X"80",X"03",X"00",X"08",X"35",X"03",X"00",X"01",X"26",
		X"02",X"00",X"85",X"07",X"03",X"01",X"FB",X"08",X"04",X"00",X"F7",X"06",X"02",X"00",X"08",X"05",
		X"1F",X"00",X"00",X"05",X"1F",X"00",X"04",X"05",X"1F",X"02",X"0A",X"04",X"2F",X"00",X"06",X"06",
		X"03",X"00",X"08",X"03",X"3F",X"00",X"31",X"02",X"4F",X"00",X"35",X"02",X"4F",X"02",X"BB",X"02",
		X"4F",X"00",X"B7",X"06",X"04",X"00",X"08",X"03",X"5F",X"00",X"F1",X"03",X"5F",X"00",X"F5",X"02",
		X"4F",X"02",X"FB",X"03",X"5F",X"00",X"F7",X"06",X"03",X"00",X"08",X"04",X"4F",X"00",X"01",X"02",
		X"6F",X"00",X"05",X"02",X"4F",X"02",X"4B",X"02",X"6F",X"00",X"47",X"08",X"05",X"00",X"08",X"02",
		X"6F",X"00",X"81",X"00",X"8F",X"00",X"85",X"00",X"6F",X"02",X"CB",X"00",X"8F",X"00",X"C7",X"08",
		X"05",X"00",X"08",X"03",X"7F",X"00",X"31",X"00",X"AF",X"00",X"B5",X"00",X"7F",X"03",X"BB",X"00",
		X"AF",X"00",X"F7",X"08",X"06",X"00",X"08",X"03",X"7F",X"00",X"01",X"00",X"AF",X"00",X"05",X"00",
		X"7F",X"03",X"0B",X"00",X"AF",X"00",X"87",X"08",X"06",X"00",X"08",X"03",X"7F",X"00",X"31",X"00",
		X"AF",X"00",X"B5",X"00",X"7F",X"03",X"BB",X"00",X"AF",X"00",X"F7",X"08",X"0F",X"00",X"08",X"03",
		X"7F",X"00",X"01",X"00",X"AF",X"00",X"05",X"00",X"7F",X"03",X"0B",X"00",X"AF",X"00",X"87",X"00",
		X"63",X"00",X"08",X"00",X"AF",X"00",X"31",X"00",X"AF",X"00",X"B5",X"00",X"7F",X"03",X"BB",X"00",
		X"AF",X"00",X"F7",X"00",X"64",X"00",X"08",X"00",X"AF",X"00",X"01",X"00",X"AF",X"00",X"05",X"00",
		X"7F",X"03",X"0B",X"00",X"AF",X"00",X"87",X"00",X"65",X"00",X"08",X"00",X"AF",X"00",X"31",X"00",
		X"AF",X"00",X"B5",X"00",X"7F",X"03",X"BB",X"00",X"AF",X"00",X"F7",X"00",X"6F",X"00",X"08",X"00",
		X"AF",X"00",X"01",X"00",X"AF",X"00",X"05",X"00",X"7F",X"03",X"0B",X"00",X"AF",X"00",X"87",X"00",
		X"86",X"00",X"08",X"00",X"AF",X"00",X"31",X"00",X"AF",X"00",X"B5",X"00",X"7F",X"03",X"BB",X"00",
		X"AF",X"00",X"F7",X"00",X"8F",X"00",X"08",X"00",X"AF",X"00",X"01",X"00",X"AF",X"00",X"05",X"00",
		X"7F",X"03",X"0B",X"00",X"AF",X"00",X"87",X"00",X"8F",X"00",X"08",X"10",X"F8",X"A0",X"11",X"87",
		X"A1",X"80",X"AB",X"79",X"7C",X"7C",X"79",X"81",X"7D",X"77",X"80",X"85",X"7C",X"85",X"87",X"74",
		X"76",X"73",X"72",X"79",X"87",X"77",X"80",X"79",X"72",X"87",X"A4",X"00",X"71",X"C8",X"71",X"C9",
		X"72",X"18",X"72",X"A1",X"72",X"F1",X"71",X"DF",X"39",X"8E",X"6F",X"E7",X"BD",X"6E",X"A3",X"86",
		X"0F",X"BD",X"6E",X"64",X"8E",X"6F",X"EB",X"BD",X"6E",X"A3",X"86",X"0F",X"7E",X"6D",X"2A",X"8E",
		X"70",X"2B",X"BD",X"6E",X"A3",X"86",X"1E",X"BD",X"6E",X"64",X"BD",X"6E",X"53",X"8E",X"72",X"00",
		X"CC",X"17",X"FF",X"BD",X"E0",X"09",X"AE",X"47",X"A6",X"02",X"A7",X"A8",X"2D",X"7E",X"6D",X"30",
		X"86",X"41",X"BD",X"E0",X"37",X"6A",X"C8",X"2D",X"2F",X"0B",X"8E",X"68",X"A5",X"CC",X"17",X"FF",
		X"BD",X"E0",X"09",X"20",X"EB",X"7E",X"68",X"A5",X"96",X"5C",X"27",X"48",X"96",X"52",X"27",X"44",
		X"CC",X"72",X"36",X"ED",X"C8",X"13",X"0F",X"A3",X"0F",X"A4",X"8E",X"6F",X"EF",X"BD",X"6E",X"A3",
		X"8E",X"6F",X"F3",X"7E",X"6E",X"A3",X"96",X"A3",X"9A",X"A4",X"27",X"05",X"8E",X"6F",X"F7",X"20",
		X"1B",X"96",X"52",X"27",X"08",X"8E",X"88",X"EE",X"86",X"30",X"BD",X"E6",X"A8",X"96",X"5C",X"27",
		X"08",X"8E",X"89",X"1F",X"86",X"30",X"BD",X"E6",X"A8",X"8E",X"6F",X"FB",X"BD",X"6E",X"A3",X"86",
		X"14",X"7E",X"6E",X"64",X"CC",X"72",X"74",X"ED",X"C8",X"13",X"0F",X"A5",X"0F",X"A6",X"8E",X"6F",
		X"FF",X"7E",X"6E",X"A3",X"8E",X"70",X"03",X"96",X"52",X"27",X"11",X"96",X"A5",X"26",X"DD",X"8E",
		X"88",X"EE",X"86",X"30",X"BD",X"E6",X"A8",X"8E",X"70",X"07",X"20",X"D0",X"96",X"5C",X"27",X"CC",
		X"96",X"A6",X"26",X"C8",X"8E",X"89",X"1F",X"86",X"30",X"BD",X"E6",X"A8",X"8E",X"70",X"0B",X"20",
		X"BB",X"96",X"52",X"27",X"2C",X"96",X"5C",X"27",X"28",X"CC",X"72",X"D2",X"ED",X"C8",X"13",X"86",
		X"FF",X"97",X"A3",X"97",X"A4",X"8E",X"70",X"0F",X"BD",X"6E",X"A3",X"86",X"0F",X"BD",X"6E",X"64",
		X"8E",X"70",X"13",X"BD",X"6E",X"A3",X"8E",X"70",X"17",X"BD",X"6E",X"A3",X"86",X"0F",X"7E",X"6D",
		X"2A",X"39",X"96",X"A3",X"2A",X"0C",X"8E",X"70",X"1F",X"96",X"A4",X"2A",X"08",X"8E",X"70",X"1B",
		X"20",X"03",X"8E",X"70",X"23",X"BD",X"6E",X"A3",X"0F",X"A3",X"0F",X"A4",X"86",X"14",X"7E",X"6E",
		X"64",X"8E",X"70",X"27",X"BD",X"6E",X"A3",X"86",X"1E",X"BD",X"6E",X"64",X"BD",X"6E",X"53",X"BD",
		X"6E",X"C4",X"AE",X"47",X"10",X"8E",X"89",X"E3",X"A6",X"84",X"26",X"04",X"A6",X"01",X"20",X"0C",
		X"10",X"8E",X"89",X"B2",X"85",X"0F",X"26",X"08",X"10",X"8E",X"89",X"81",X"44",X"44",X"44",X"44",
		X"84",X"0F",X"97",X"A2",X"10",X"AF",X"4D",X"F6",X"B1",X"BA",X"96",X"5C",X"27",X"05",X"96",X"52",
		X"27",X"01",X"54",X"E7",X"C8",X"1A",X"A6",X"01",X"84",X"0F",X"97",X"8F",X"8E",X"B1",X"42",X"6F",
		X"80",X"8C",X"B1",X"8D",X"25",X"F9",X"86",X"02",X"A7",X"C8",X"1D",X"86",X"06",X"A7",X"C8",X"19",
		X"10",X"8E",X"74",X"84",X"8E",X"B1",X"87",X"BD",X"E0",X"18",X"C6",X"0C",X"3D",X"E6",X"86",X"27",
		X"07",X"4A",X"2A",X"F9",X"86",X"05",X"20",X"F5",X"6C",X"86",X"31",X"A6",X"BD",X"E0",X"18",X"49",
		X"E6",X"A0",X"E0",X"3E",X"3D",X"AB",X"3E",X"8E",X"B1",X"42",X"6C",X"86",X"BD",X"74",X"17",X"6A",
		X"C8",X"19",X"26",X"CC",X"86",X"06",X"A7",X"C8",X"19",X"8E",X"B1",X"42",X"BD",X"E0",X"18",X"C6",
		X"8A",X"3D",X"E6",X"86",X"27",X"08",X"4C",X"81",X"45",X"25",X"F7",X"4F",X"20",X"F4",X"6C",X"86",
		X"BD",X"74",X"17",X"6A",X"C8",X"19",X"26",X"E1",X"7E",X"6D",X"5F",X"C8",X"DC",X"D3",X"C9",X"A4",
		X"D3",X"C9",X"A4",X"D2",X"D5",X"CF",X"C9",X"C8",X"F8",X"AE",X"D8",X"DF",X"C9",X"D3",X"DD",X"D6",
		X"DF",X"D8",X"A4",X"DA",X"C3",X"A4",X"CD",X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",
		X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",
		X"C4",X"D9",X"FB",X"A4",X"AD",X"A5",X"A6",X"AC",X"A4",X"CD",X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",
		X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",
		X"D9",X"F8",X"AE",X"DB",X"D0",X"D0",X"A4",X"CA",X"D3",X"DD",X"DC",X"C8",X"C9",X"A4",X"CA",X"DF",
		X"C9",X"DF",X"CA",X"CE",X"DF",X"D8",X"2E",X"34",X"02",X"0C",X"AA",X"8E",X"76",X"9F",X"CC",X"82",
		X"FF",X"BD",X"E0",X"09",X"35",X"02",X"8E",X"74",X"86",X"30",X"04",X"A1",X"84",X"24",X"FA",X"C6",
		X"08",X"E7",X"A8",X"35",X"3D",X"E3",X"02",X"ED",X"27",X"C3",X"00",X"06",X"ED",X"A8",X"29",X"E6",
		X"01",X"4F",X"ED",X"2A",X"E7",X"A8",X"27",X"C0",X"06",X"E7",X"A8",X"28",X"EC",X"4D",X"ED",X"2D",
		X"E6",X"C8",X"1A",X"E7",X"A8",X"2D",X"6A",X"C8",X"1D",X"2B",X"0B",X"BD",X"E0",X"18",X"3D",X"40",
		X"AB",X"A8",X"2D",X"A7",X"A8",X"2D",X"CC",X"00",X"00",X"ED",X"A8",X"1C",X"ED",X"A8",X"2B",X"6F",
		X"A8",X"34",X"86",X"04",X"A7",X"A8",X"33",X"EC",X"E1",X"ED",X"4F",X"86",X"01",X"BD",X"E0",X"37",
		X"6E",X"D8",X"0F",X"00",X"08",X"13",X"1A",X"26",X"2E",X"45",X"03",X"44",X"00",X"09",X"08",X"44",
		X"00",X"E5",X"13",X"50",X"00",X"16",X"1A",X"80",X"00",X"32",X"21",X"89",X"FF",X"39",X"26",X"89",
		X"FF",X"F9",X"2E",X"A2",X"FF",X"3A",X"45",X"D2",X"FE",X"C6",X"FF",X"44",X"FE",X"09",X"34",X"50",
		X"86",X"07",X"A7",X"C8",X"2D",X"CC",X"68",X"28",X"ED",X"C8",X"24",X"8E",X"EF",X"6D",X"BD",X"E0",
		X"2D",X"35",X"D0",X"34",X"50",X"8E",X"EF",X"97",X"BD",X"E0",X"2D",X"96",X"8E",X"A0",X"C8",X"34",
		X"97",X"8E",X"0A",X"A1",X"86",X"82",X"E6",X"43",X"8E",X"76",X"11",X"BD",X"E0",X"30",X"CC",X"00",
		X"00",X"ED",X"A8",X"2B",X"ED",X"A8",X"1C",X"ED",X"A8",X"27",X"EC",X"4A",X"C0",X"08",X"ED",X"2A",
		X"EC",X"47",X"C3",X"00",X"04",X"ED",X"27",X"6F",X"A8",X"35",X"EC",X"4D",X"10",X"83",X"89",X"E3",
		X"24",X"03",X"C3",X"00",X"31",X"ED",X"2D",X"EC",X"C8",X"11",X"ED",X"A8",X"11",X"A6",X"C8",X"14",
		X"A7",X"A8",X"14",X"6F",X"A8",X"22",X"6F",X"A8",X"23",X"6F",X"A8",X"16",X"6F",X"A8",X"10",X"A6",
		X"C8",X"33",X"A7",X"A8",X"33",X"6A",X"A8",X"33",X"26",X"09",X"1F",X"21",X"EE",X"E4",X"27",X"03",
		X"BD",X"75",X"3B",X"35",X"D0",X"BD",X"75",X"3B",X"7E",X"84",X"13",X"34",X"50",X"8E",X"EF",X"86",
		X"BD",X"E0",X"2D",X"10",X"AE",X"4D",X"A6",X"A8",X"2E",X"AE",X"E4",X"A7",X"88",X"2F",X"10",X"AE",
		X"A8",X"12",X"E6",X"A4",X"C1",X"04",X"24",X"01",X"5C",X"E7",X"A4",X"E7",X"88",X"2E",X"58",X"EB",
		X"A4",X"10",X"8E",X"75",X"A1",X"31",X"A5",X"A6",X"A4",X"AE",X"4D",X"AD",X"B8",X"01",X"10",X"AE",
		X"E4",X"6F",X"A8",X"33",X"A6",X"A8",X"35",X"26",X"08",X"63",X"A8",X"33",X"86",X"05",X"BD",X"E6",
		X"A8",X"0A",X"AA",X"AE",X"E4",X"10",X"AE",X"88",X"2B",X"27",X"08",X"0A",X"A1",X"CC",X"EE",X"C2",
		X"ED",X"A8",X"24",X"CC",X"77",X"AC",X"ED",X"05",X"86",X"04",X"A7",X"04",X"A6",X"02",X"84",X"7F",
		X"A7",X"02",X"35",X"D0",X"52",X"E6",X"B1",X"05",X"E6",X"A8",X"57",X"E6",X"B1",X"10",X"E6",X"A8",
		X"D6",X"48",X"1D",X"E3",X"C8",X"11",X"ED",X"C8",X"11",X"E3",X"4B",X"AB",X"C8",X"23",X"6F",X"C8",
		X"23",X"81",X"20",X"22",X"12",X"6C",X"C8",X"23",X"EC",X"C8",X"11",X"2A",X"07",X"43",X"50",X"82",
		X"FF",X"ED",X"C8",X"11",X"CC",X"20",X"00",X"ED",X"4B",X"A7",X"C8",X"27",X"80",X"06",X"A7",X"C8",
		X"28",X"A6",X"C8",X"14",X"8E",X"DC",X"D5",X"EC",X"86",X"EB",X"C8",X"16",X"E7",X"C8",X"16",X"89",
		X"00",X"1F",X"89",X"BD",X"DD",X"D2",X"10",X"83",X"01",X"20",X"2F",X"03",X"C3",X"FE",X"E4",X"10",
		X"83",X"00",X"04",X"2C",X"03",X"C3",X"01",X"1C",X"ED",X"47",X"C3",X"00",X"06",X"ED",X"C8",X"29",
		X"39",X"BD",X"78",X"E3",X"96",X"B0",X"BD",X"E0",X"37",X"BD",X"6A",X"F3",X"BD",X"75",X"B0",X"BD",
		X"77",X"9B",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"B0",X"02",X"AA",X"89",X"B0",X"00",X"A4",
		X"89",X"AF",X"F9",X"A4",X"A9",X"EA",X"97",X"84",X"7F",X"26",X"25",X"AE",X"47",X"10",X"AE",X"4A",
		X"A6",X"89",X"AE",X"A2",X"A4",X"89",X"AE",X"98",X"A4",X"A9",X"E8",X"3D",X"A4",X"A9",X"E8",X"44",
		X"27",X"03",X"BD",X"DA",X"3E",X"E6",X"4B",X"C1",X"E3",X"25",X"B6",X"0A",X"AA",X"7E",X"78",X"8A",
		X"A7",X"C8",X"35",X"BD",X"D9",X"C2",X"E7",X"C8",X"27",X"C0",X"06",X"E7",X"C8",X"28",X"A6",X"C8",
		X"14",X"27",X"08",X"2B",X"04",X"8B",X"FE",X"20",X"02",X"8B",X"02",X"A7",X"C8",X"14",X"EC",X"C8",
		X"11",X"2B",X"B8",X"47",X"56",X"47",X"56",X"43",X"50",X"82",X"FF",X"ED",X"C8",X"11",X"10",X"83",
		X"FF",X"E0",X"2D",X"A7",X"A6",X"C8",X"14",X"26",X"A2",X"B6",X"B1",X"B7",X"A7",X"C8",X"2D",X"BD",
		X"78",X"E3",X"86",X"0C",X"BD",X"E0",X"37",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"B0",X"02",
		X"AA",X"89",X"B0",X"00",X"A4",X"89",X"AF",X"F9",X"A4",X"A9",X"EA",X"98",X"84",X"7F",X"10",X"27",
		X"FF",X"4F",X"6A",X"C8",X"2D",X"26",X"D8",X"6C",X"C8",X"2D",X"96",X"A1",X"91",X"A2",X"24",X"CF",
		X"0C",X"A1",X"8E",X"EF",X"89",X"BD",X"E0",X"2D",X"86",X"0F",X"E6",X"43",X"8E",X"8E",X"AF",X"BD",
		X"E0",X"30",X"10",X"AF",X"C8",X"2B",X"EF",X"A8",X"2B",X"A6",X"C8",X"33",X"A7",X"A8",X"33",X"6F",
		X"A8",X"34",X"6F",X"2F",X"6F",X"A8",X"2E",X"86",X"08",X"A7",X"A8",X"14",X"CC",X"00",X"00",X"ED",
		X"A8",X"11",X"ED",X"A8",X"1A",X"6F",X"A8",X"22",X"6F",X"A8",X"16",X"6F",X"A8",X"10",X"FC",X"00",
		X"1A",X"ED",X"A8",X"18",X"EC",X"4D",X"ED",X"2D",X"CC",X"79",X"3C",X"ED",X"A8",X"24",X"EC",X"47",
		X"83",X"00",X"97",X"22",X"0A",X"63",X"2F",X"60",X"A8",X"14",X"CC",X"01",X"23",X"20",X"03",X"CC",
		X"FF",X"F7",X"ED",X"27",X"A6",X"4B",X"C6",X"A9",X"81",X"BB",X"22",X"08",X"C6",X"68",X"81",X"69",
		X"22",X"02",X"C6",X"45",X"4F",X"ED",X"2A",X"8E",X"79",X"24",X"AF",X"C8",X"2E",X"20",X"08",X"30",
		X"03",X"AF",X"C8",X"2E",X"BD",X"E0",X"37",X"BD",X"6A",X"F3",X"BD",X"E0",X"24",X"A6",X"D8",X"2E",
		X"BD",X"79",X"0E",X"AE",X"C8",X"2E",X"A6",X"4B",X"A7",X"C8",X"27",X"A0",X"01",X"A7",X"C8",X"28",
		X"A6",X"02",X"26",X"DB",X"86",X"07",X"BD",X"E0",X"37",X"BD",X"6A",X"F3",X"10",X"AE",X"4D",X"10",
		X"AE",X"B8",X"0A",X"31",X"A8",X"18",X"10",X"AF",X"C8",X"1C",X"BD",X"8E",X"89",X"86",X"08",X"BD",
		X"E0",X"37",X"10",X"AE",X"C8",X"1C",X"BD",X"8E",X"89",X"20",X"F2",X"AE",X"47",X"A6",X"89",X"AE",
		X"A2",X"AE",X"4A",X"A4",X"89",X"E8",X"42",X"9A",X"4B",X"97",X"4B",X"39",X"BD",X"6A",X"F3",X"BD",
		X"77",X"9B",X"96",X"90",X"2F",X"03",X"BD",X"78",X"B4",X"86",X"02",X"BD",X"E0",X"37",X"BD",X"78",
		X"8D",X"86",X"01",X"A7",X"C8",X"32",X"AE",X"9F",X"A0",X"0A",X"AE",X"84",X"27",X"4A",X"A6",X"02",
		X"81",X"03",X"26",X"F6",X"EC",X"4A",X"A3",X"0A",X"2A",X"04",X"43",X"50",X"82",X"FF",X"83",X"00",
		X"06",X"2C",X"E7",X"EC",X"47",X"A3",X"07",X"2A",X"04",X"43",X"50",X"82",X"FF",X"83",X"00",X"10",
		X"2C",X"D8",X"A6",X"88",X"2D",X"81",X"08",X"25",X"11",X"86",X"08",X"A7",X"88",X"2D",X"10",X"AE",
		X"84",X"E6",X"22",X"C1",X"04",X"26",X"03",X"A7",X"A8",X"2D",X"48",X"AB",X"88",X"32",X"A1",X"C8",
		X"32",X"25",X"B7",X"A7",X"C8",X"32",X"20",X"B2",X"86",X"03",X"A7",X"42",X"86",X"1E",X"A7",X"C8",
		X"2D",X"86",X"01",X"BD",X"E0",X"37",X"6A",X"C8",X"32",X"26",X"F6",X"A6",X"C8",X"33",X"27",X"2A",
		X"8E",X"78",X"5F",X"CC",X"04",X"FF",X"BD",X"E0",X"30",X"CC",X"02",X"22",X"ED",X"A8",X"2E",X"EC",
		X"47",X"ED",X"27",X"EC",X"4A",X"C0",X"06",X"ED",X"2A",X"EC",X"C8",X"20",X"C0",X"06",X"ED",X"A8",
		X"20",X"A6",X"C8",X"2D",X"A7",X"A8",X"2D",X"6F",X"A8",X"32",X"86",X"02",X"BD",X"E0",X"37",X"20",
		X"07",X"86",X"1E",X"A7",X"C8",X"2D",X"8D",X"25",X"AE",X"C8",X"20",X"EC",X"C8",X"2E",X"6A",X"C8",
		X"2D",X"27",X"0A",X"BD",X"4A",X"5C",X"86",X"02",X"BD",X"E0",X"37",X"20",X"EB",X"5F",X"BD",X"4A",
		X"5C",X"BD",X"77",X"9B",X"7E",X"E0",X"0F",X"BD",X"6A",X"F3",X"7E",X"E0",X"0F",X"EC",X"47",X"C4",
		X"FE",X"E7",X"48",X"46",X"56",X"1F",X"98",X"E6",X"4B",X"C0",X"05",X"C1",X"CE",X"23",X"02",X"C6",
		X"CE",X"81",X"88",X"23",X"02",X"86",X"88",X"ED",X"C8",X"20",X"E7",X"4B",X"1F",X"89",X"4F",X"58",
		X"49",X"ED",X"47",X"39",X"8E",X"78",X"D1",X"CC",X"02",X"FF",X"BD",X"E0",X"30",X"EC",X"47",X"ED",
		X"27",X"EC",X"4A",X"ED",X"2A",X"EC",X"C8",X"2E",X"ED",X"A8",X"2E",X"39",X"8D",X"E6",X"7E",X"78",
		X"61",X"86",X"44",X"BD",X"E0",X"37",X"6C",X"C8",X"2E",X"A6",X"C8",X"2E",X"81",X"04",X"23",X"EC",
		X"7E",X"E0",X"0F",X"BD",X"E0",X"24",X"A6",X"C8",X"14",X"2A",X"06",X"10",X"8E",X"79",X"1E",X"20",
		X"04",X"10",X"8E",X"79",X"21",X"EC",X"C8",X"11",X"2B",X"0D",X"83",X"00",X"80",X"2E",X"04",X"A6",
		X"A4",X"20",X"0B",X"A6",X"22",X"20",X"07",X"C3",X"00",X"80",X"2E",X"F3",X"A6",X"21",X"10",X"BE",
		X"00",X"28",X"31",X"A6",X"10",X"AF",X"C8",X"1C",X"BD",X"8E",X"70",X"7E",X"D8",X"F4",X"00",X"0C",
		X"06",X"00",X"06",X"0C",X"06",X"06",X"07",X"00",X"06",X"03",X"0C",X"06",X"07",X"00",X"06",X"43",
		X"12",X"06",X"07",X"18",X"0B",X"07",X"1E",X"0B",X"07",X"24",X"0B",X"00",X"10",X"AE",X"C8",X"2B",
		X"5F",X"A6",X"2B",X"A1",X"4B",X"27",X"38",X"25",X"21",X"E6",X"C8",X"11",X"C1",X"02",X"2C",X"1A",
		X"AE",X"47",X"A6",X"89",X"AE",X"B4",X"E6",X"C8",X"14",X"2A",X"04",X"A6",X"89",X"AE",X"90",X"AE",
		X"4A",X"5F",X"A4",X"89",X"E8",X"37",X"84",X"08",X"27",X"15",X"5F",X"A6",X"C8",X"11",X"81",X"FF",
		X"2D",X"0D",X"CC",X"7A",X"5E",X"ED",X"C8",X"24",X"86",X"04",X"A7",X"C8",X"2D",X"C6",X"01",X"34",
		X"04",X"EC",X"27",X"C3",X"FF",X"F4",X"A3",X"47",X"2A",X"52",X"C3",X"00",X"14",X"2B",X"3C",X"86",
		X"01",X"A7",X"C8",X"2E",X"AE",X"C8",X"20",X"27",X"12",X"A6",X"2B",X"E1",X"4B",X"22",X"25",X"A6",
		X"C8",X"14",X"27",X"6E",X"A6",X"C8",X"14",X"2B",X"3D",X"20",X"2A",X"A6",X"C8",X"14",X"2B",X"08",
		X"2E",X"0C",X"A6",X"4F",X"2B",X"1F",X"20",X"2E",X"81",X"FE",X"27",X"31",X"20",X"28",X"81",X"02",
		X"27",X"2B",X"20",X"11",X"A6",X"C8",X"14",X"2B",X"07",X"20",X"16",X"A6",X"C8",X"2E",X"26",X"23",
		X"A6",X"C8",X"14",X"2B",X"18",X"86",X"FF",X"35",X"04",X"DD",X"32",X"39",X"A6",X"C8",X"2E",X"26",
		X"12",X"A6",X"C8",X"14",X"2E",X"07",X"86",X"01",X"35",X"04",X"DD",X"32",X"39",X"4F",X"35",X"04",
		X"DD",X"32",X"39",X"EC",X"27",X"A3",X"47",X"2B",X"0B",X"10",X"83",X"00",X"97",X"2D",X"0E",X"83",
		X"01",X"2E",X"20",X"09",X"10",X"83",X"FF",X"69",X"2E",X"03",X"C3",X"01",X"2E",X"4D",X"2B",X"C0",
		X"20",X"CF",X"35",X"04",X"CC",X"7A",X"1F",X"ED",X"C8",X"24",X"86",X"06",X"A7",X"C8",X"2D",X"6A",
		X"C8",X"2D",X"27",X"0B",X"86",X"01",X"E6",X"4F",X"2A",X"01",X"40",X"5F",X"DD",X"32",X"39",X"0C",
		X"8E",X"6C",X"C8",X"34",X"8E",X"EF",X"8C",X"BD",X"E0",X"2D",X"AE",X"C8",X"2B",X"CC",X"78",X"87",
		X"ED",X"05",X"86",X"01",X"A7",X"04",X"A6",X"02",X"84",X"7F",X"A7",X"02",X"AE",X"4D",X"96",X"90",
		X"26",X"04",X"EC",X"84",X"20",X"02",X"EC",X"02",X"ED",X"C8",X"24",X"7E",X"8D",X"40",X"6A",X"C8",
		X"2D",X"27",X"06",X"CC",X"00",X"01",X"DD",X"32",X"39",X"CC",X"79",X"3C",X"ED",X"C8",X"24",X"CC",
		X"00",X"00",X"DD",X"32",X"39",X"BD",X"E0",X"18",X"49",X"C6",X"10",X"3D",X"8A",X"A0",X"1F",X"01",
		X"6C",X"84",X"39",X"96",X"8E",X"91",X"8F",X"25",X"4C",X"6A",X"C8",X"32",X"2E",X"0E",X"B6",X"B1",
		X"B4",X"A7",X"C8",X"32",X"9E",X"2C",X"A6",X"02",X"81",X"15",X"27",X"1A",X"86",X"45",X"E6",X"4B",
		X"C1",X"65",X"25",X"08",X"86",X"81",X"C1",X"A1",X"25",X"02",X"86",X"D0",X"5F",X"A0",X"4B",X"2A",
		X"0D",X"A6",X"C8",X"11",X"2B",X"08",X"CC",X"7A",X"CC",X"ED",X"C8",X"24",X"C6",X"01",X"6D",X"4F",
		X"2B",X"05",X"86",X"01",X"DD",X"32",X"39",X"86",X"FF",X"DD",X"32",X"39",X"CC",X"7A",X"83",X"ED",
		X"C8",X"24",X"5F",X"20",X"E9",X"0C",X"8E",X"6C",X"C8",X"34",X"AE",X"4D",X"AE",X"02",X"AF",X"C8",
		X"24",X"6E",X"84",X"4A",X"4F",X"55",X"53",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",
		X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",
		X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"6A",X"C8",X"32",X"2E",X"0E",
		X"B6",X"B1",X"B4",X"A7",X"C8",X"32",X"9E",X"2C",X"A6",X"02",X"81",X"15",X"27",X"3E",X"BD",X"80",
		X"D6",X"27",X"1C",X"EC",X"0A",X"A3",X"4A",X"10",X"2D",X"00",X"5B",X"10",X"B3",X"B1",X"BC",X"2D",
		X"0E",X"FC",X"B1",X"BF",X"ED",X"C8",X"2B",X"CC",X"7B",X"42",X"ED",X"C8",X"24",X"20",X"15",X"7E",
		X"7C",X"07",X"EC",X"C8",X"20",X"26",X"3C",X"EC",X"C8",X"11",X"2B",X"79",X"E3",X"C8",X"2B",X"2A",
		X"32",X"ED",X"C8",X"2B",X"EC",X"C8",X"11",X"B3",X"B1",X"C2",X"2B",X"69",X"CC",X"7B",X"66",X"ED",
		X"C8",X"24",X"86",X"02",X"20",X"58",X"EC",X"C8",X"11",X"2B",X"08",X"E3",X"C8",X"2B",X"2A",X"13",
		X"ED",X"C8",X"2B",X"C6",X"01",X"6A",X"C8",X"2D",X"2E",X"07",X"CC",X"7B",X"42",X"ED",X"C8",X"24",
		X"5F",X"20",X"43",X"7E",X"7B",X"0B",X"10",X"B3",X"B1",X"C5",X"2E",X"7B",X"AE",X"47",X"10",X"AE",
		X"4A",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"29",X"26",X"6C",X"FC",X"B1",X"C8",X"ED",X"C8",
		X"2B",X"20",X"12",X"EC",X"C8",X"11",X"2A",X"08",X"E3",X"C8",X"2B",X"2B",X"D6",X"ED",X"C8",X"2B",
		X"6A",X"C8",X"2D",X"2E",X"10",X"CC",X"7B",X"E1",X"ED",X"C8",X"24",X"B6",X"B1",X"CC",X"A7",X"C8",
		X"2D",X"C6",X"01",X"20",X"01",X"5F",X"A6",X"4B",X"81",X"D3",X"25",X"07",X"A6",X"C8",X"11",X"10",
		X"2A",X"00",X"AA",X"A6",X"4F",X"2B",X"05",X"86",X"01",X"DD",X"32",X"39",X"86",X"FF",X"DD",X"32",
		X"39",X"EC",X"C8",X"11",X"2A",X"08",X"E3",X"C8",X"2B",X"2B",X"98",X"ED",X"C8",X"2B",X"C6",X"01",
		X"6A",X"C8",X"2D",X"2E",X"0D",X"B6",X"B1",X"CF",X"A7",X"C8",X"2D",X"CC",X"7B",X"A3",X"ED",X"C8",
		X"24",X"5F",X"20",X"C2",X"7E",X"7B",X"0B",X"CC",X"7C",X"1E",X"ED",X"C8",X"24",X"EC",X"4A",X"ED",
		X"C8",X"2B",X"A6",X"88",X"14",X"A7",X"C8",X"2F",X"B6",X"B1",X"D2",X"A7",X"C8",X"2D",X"6A",X"C8",
		X"2D",X"2F",X"E1",X"E6",X"4B",X"C1",X"D3",X"25",X"17",X"BD",X"80",X"D6",X"27",X"1E",X"EC",X"07",
		X"C3",X"00",X"3F",X"10",X"A3",X"47",X"2D",X"14",X"C3",X"FF",X"82",X"10",X"A3",X"47",X"2E",X"0C",
		X"A6",X"C8",X"11",X"2B",X"17",X"E6",X"C8",X"2C",X"E1",X"4B",X"25",X"10",X"CC",X"7C",X"56",X"ED",
		X"C8",X"24",X"C6",X"01",X"20",X"07",X"CC",X"7C",X"1E",X"ED",X"C8",X"24",X"5F",X"A6",X"C8",X"2F",
		X"A1",X"C8",X"14",X"26",X"0A",X"6A",X"C8",X"2E",X"2B",X"05",X"6F",X"C8",X"2E",X"63",X"4F",X"7E",
		X"7B",X"D3",X"A6",X"4B",X"81",X"D3",X"25",X"18",X"A6",X"C8",X"11",X"2B",X"13",X"CC",X"7C",X"87",
		X"ED",X"C8",X"24",X"C6",X"01",X"20",X"E8",X"CC",X"7C",X"72",X"ED",X"C8",X"24",X"5F",X"20",X"DF",
		X"AE",X"4D",X"6E",X"98",X"02",X"6A",X"C8",X"32",X"2E",X"0E",X"B6",X"B1",X"B4",X"A7",X"C8",X"32",
		X"9E",X"2C",X"A6",X"02",X"81",X"15",X"27",X"3D",X"BD",X"80",X"D6",X"27",X"1B",X"EC",X"0A",X"A3",
		X"4A",X"10",X"2D",X"00",X"61",X"B3",X"B1",X"D4",X"2D",X"0E",X"FC",X"B1",X"D7",X"ED",X"C8",X"2B",
		X"CC",X"7C",X"F5",X"ED",X"C8",X"24",X"20",X"47",X"7E",X"7D",X"58",X"EC",X"C8",X"20",X"26",X"43",
		X"EC",X"C8",X"11",X"2B",X"3A",X"E3",X"C8",X"2B",X"2A",X"39",X"ED",X"C8",X"2B",X"EC",X"C8",X"11",
		X"B3",X"B1",X"DA",X"2B",X"2A",X"CC",X"7C",X"F5",X"ED",X"C8",X"24",X"86",X"02",X"A7",X"C8",X"2D",
		X"C6",X"01",X"7E",X"7D",X"BF",X"EC",X"C8",X"11",X"2B",X"08",X"E3",X"C8",X"2B",X"2A",X"14",X"ED",
		X"C8",X"2B",X"C6",X"01",X"6A",X"C8",X"2D",X"2E",X"07",X"CC",X"7C",X"CB",X"ED",X"C8",X"24",X"5F",
		X"7E",X"7D",X"BF",X"7E",X"7C",X"95",X"10",X"B3",X"B1",X"DD",X"2E",X"AC",X"AE",X"47",X"10",X"AE",
		X"4A",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"29",X"10",X"26",X"01",X"56",X"FC",X"B1",X"E0",
		X"ED",X"C8",X"2B",X"20",X"14",X"EC",X"C8",X"11",X"2A",X"08",X"E3",X"C8",X"2B",X"2B",X"D4",X"ED",
		X"C8",X"2B",X"C6",X"01",X"6A",X"C8",X"2D",X"2E",X"0D",X"B6",X"B1",X"E7",X"A7",X"C8",X"2D",X"CC",
		X"7E",X"47",X"ED",X"C8",X"24",X"5F",X"20",X"67",X"CC",X"7D",X"6F",X"ED",X"C8",X"24",X"EC",X"4A",
		X"ED",X"C8",X"2B",X"A6",X"88",X"14",X"A7",X"C8",X"2F",X"B6",X"B1",X"ED",X"A7",X"C8",X"2D",X"6A",
		X"C8",X"2D",X"10",X"2F",X"00",X"CE",X"A6",X"C8",X"11",X"10",X"2B",X"00",X"C3",X"E6",X"4B",X"C1",
		X"D3",X"25",X"17",X"BD",X"80",X"D6",X"27",X"1B",X"EC",X"07",X"C3",X"00",X"2D",X"10",X"A3",X"47",
		X"2D",X"11",X"C3",X"FF",X"A6",X"10",X"A3",X"47",X"2E",X"09",X"E6",X"C8",X"2C",X"E1",X"4B",X"10",
		X"25",X"00",X"9D",X"CC",X"7E",X"3A",X"ED",X"C8",X"24",X"C6",X"01",X"A6",X"C8",X"2F",X"A1",X"C8",
		X"14",X"26",X"1A",X"6A",X"C8",X"2E",X"2B",X"15",X"6F",X"C8",X"2E",X"63",X"4F",X"20",X"0E",X"A6",
		X"4B",X"81",X"D3",X"25",X"08",X"A6",X"C8",X"11",X"2B",X"03",X"7E",X"7C",X"7D",X"A6",X"C8",X"14",
		X"27",X"53",X"2A",X"22",X"34",X"04",X"EC",X"C8",X"11",X"58",X"49",X"58",X"49",X"58",X"49",X"35",
		X"04",X"10",X"AE",X"4A",X"AE",X"47",X"31",X"A6",X"A6",X"89",X"AE",X"83",X"A4",X"A9",X"E8",X"37",
		X"27",X"33",X"6F",X"4F",X"20",X"22",X"34",X"04",X"EC",X"C8",X"11",X"58",X"49",X"58",X"49",X"58",
		X"49",X"35",X"04",X"10",X"AE",X"4A",X"AE",X"47",X"31",X"A6",X"A6",X"89",X"AE",X"C1",X"A4",X"A9",
		X"E8",X"37",X"27",X"11",X"86",X"FF",X"A7",X"4F",X"CC",X"7E",X"7A",X"ED",X"C8",X"24",X"86",X"08",
		X"A7",X"C8",X"2D",X"C6",X"01",X"A6",X"C8",X"22",X"27",X"02",X"A7",X"4F",X"A6",X"4F",X"2B",X"05",
		X"86",X"01",X"DD",X"32",X"39",X"86",X"FF",X"DD",X"32",X"39",X"CC",X"7D",X"6F",X"ED",X"C8",X"24",
		X"5F",X"7E",X"7D",X"AB",X"7E",X"7C",X"95",X"EC",X"C8",X"11",X"2A",X"08",X"E3",X"C8",X"2B",X"2B",
		X"F3",X"ED",X"C8",X"2B",X"6A",X"C8",X"2D",X"2E",X"1D",X"6C",X"C8",X"2D",X"EC",X"C8",X"11",X"10",
		X"B3",X"B1",X"E9",X"2D",X"11",X"CC",X"7D",X"35",X"ED",X"C8",X"24",X"B6",X"B1",X"E4",X"A7",X"C8",
		X"2D",X"C6",X"01",X"7E",X"7D",X"BF",X"5F",X"7E",X"7D",X"BF",X"5F",X"6A",X"C8",X"2D",X"2E",X"A5",
		X"7E",X"7C",X"95",X"CC",X"7E",X"93",X"ED",X"C8",X"24",X"EC",X"4A",X"ED",X"C8",X"2B",X"86",X"15",
		X"A7",X"C8",X"2D",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"29",
		X"10",X"27",X"FE",X"89",X"6A",X"C8",X"2D",X"10",X"2F",X"FD",X"EA",X"EC",X"C8",X"11",X"C3",X"FF",
		X"C0",X"2B",X"18",X"E6",X"C8",X"2C",X"E1",X"4B",X"25",X"11",X"CC",X"7E",X"C5",X"ED",X"C8",X"24",
		X"C6",X"01",X"7E",X"7E",X"25",X"CC",X"7E",X"93",X"ED",X"C8",X"24",X"5F",X"7E",X"7E",X"25",X"6A",
		X"C8",X"32",X"2E",X"0E",X"B6",X"B1",X"B4",X"A7",X"C8",X"32",X"9E",X"2C",X"A6",X"02",X"81",X"15",
		X"27",X"41",X"BD",X"80",X"D6",X"10",X"27",X"00",X"B0",X"EC",X"0A",X"A3",X"4A",X"10",X"2D",X"00",
		X"1B",X"B3",X"B1",X"EF",X"2D",X"4B",X"CC",X"80",X"AF",X"ED",X"C8",X"24",X"5F",X"A6",X"4B",X"81",
		X"D3",X"25",X"06",X"A6",X"C8",X"14",X"2B",X"01",X"5C",X"7E",X"80",X"3F",X"10",X"B3",X"B1",X"F2",
		X"2E",X"2F",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"29",X"10",
		X"26",X"01",X"40",X"CC",X"7F",X"2D",X"ED",X"C8",X"24",X"5F",X"7E",X"80",X"3F",X"CC",X"7E",X"CF",
		X"ED",X"C8",X"24",X"EC",X"C8",X"11",X"10",X"B3",X"B1",X"F5",X"2D",X"ED",X"C6",X"01",X"7E",X"80",
		X"3F",X"CC",X"7F",X"58",X"ED",X"C8",X"24",X"E6",X"0B",X"E7",X"C8",X"2C",X"A6",X"88",X"14",X"A7",
		X"C8",X"2F",X"B6",X"B1",X"F9",X"A7",X"C8",X"2D",X"6A",X"C8",X"2D",X"10",X"2F",X"00",X"F8",X"E6",
		X"4B",X"C1",X"D3",X"25",X"05",X"A6",X"C8",X"11",X"2A",X"05",X"E1",X"C8",X"2C",X"23",X"10",X"CC",
		X"7F",X"79",X"ED",X"C8",X"24",X"C6",X"01",X"20",X"07",X"CC",X"7F",X"58",X"ED",X"C8",X"24",X"5F",
		X"A6",X"C8",X"2F",X"A1",X"C8",X"14",X"10",X"26",X"00",X"A5",X"6A",X"C8",X"2E",X"10",X"2B",X"00",
		X"9E",X"6F",X"C8",X"2E",X"63",X"4F",X"7E",X"80",X"2F",X"CC",X"7F",X"AA",X"ED",X"C8",X"24",X"E6",
		X"4B",X"E7",X"C8",X"2C",X"B6",X"B1",X"FC",X"A7",X"C8",X"2D",X"6A",X"C8",X"2D",X"10",X"2F",X"00",
		X"A6",X"A6",X"C8",X"11",X"10",X"2B",X"00",X"9B",X"E6",X"C8",X"2C",X"E1",X"4B",X"10",X"25",X"00",
		X"92",X"CC",X"80",X"4D",X"ED",X"C8",X"24",X"C6",X"01",X"A6",X"4B",X"81",X"D0",X"25",X"07",X"A6",
		X"C8",X"11",X"10",X"2A",X"FC",X"A7",X"A6",X"C8",X"14",X"27",X"54",X"2A",X"22",X"34",X"04",X"EC",
		X"C8",X"11",X"58",X"49",X"58",X"49",X"58",X"49",X"35",X"04",X"10",X"AE",X"4A",X"AE",X"47",X"31",
		X"A6",X"A6",X"89",X"AE",X"83",X"A4",X"A9",X"E8",X"37",X"27",X"34",X"6F",X"4F",X"20",X"22",X"34",
		X"04",X"EC",X"C8",X"11",X"58",X"49",X"58",X"49",X"58",X"49",X"35",X"04",X"10",X"AE",X"4A",X"AE",
		X"47",X"31",X"A6",X"A6",X"89",X"AE",X"C1",X"A4",X"A9",X"E8",X"37",X"27",X"12",X"86",X"FF",X"A7",
		X"4F",X"CC",X"80",X"5A",X"ED",X"C8",X"24",X"B6",X"B1",X"FF",X"A7",X"C8",X"2D",X"C6",X"01",X"A6",
		X"C8",X"22",X"27",X"02",X"A7",X"4F",X"A6",X"4F",X"2B",X"0E",X"86",X"01",X"DD",X"32",X"39",X"A6",
		X"C8",X"14",X"27",X"EB",X"4F",X"DD",X"32",X"39",X"86",X"FF",X"DD",X"32",X"39",X"CC",X"7F",X"AA",
		X"ED",X"C8",X"24",X"5F",X"7E",X"7F",X"C9",X"7E",X"7E",X"CF",X"5F",X"6A",X"C8",X"2D",X"2E",X"CF",
		X"7E",X"7E",X"CF",X"CC",X"80",X"73",X"ED",X"C8",X"24",X"E6",X"4B",X"E7",X"C8",X"2C",X"86",X"15",
		X"A7",X"C8",X"2D",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"AE",X"A2",X"A4",X"A9",X"E8",X"29",
		X"10",X"27",X"FE",X"9F",X"6A",X"C8",X"2D",X"10",X"2F",X"FE",X"44",X"EC",X"C8",X"11",X"C3",X"FF",
		X"C0",X"2B",X"18",X"E6",X"C8",X"2C",X"E1",X"4B",X"25",X"11",X"CC",X"80",X"A5",X"ED",X"C8",X"24",
		X"C6",X"01",X"7E",X"80",X"2F",X"CC",X"80",X"73",X"ED",X"C8",X"24",X"5F",X"7E",X"80",X"2F",X"CC",
		X"7E",X"CF",X"ED",X"C8",X"24",X"5F",X"A6",X"C8",X"14",X"10",X"27",X"FF",X"72",X"A6",X"C8",X"20",
		X"27",X"10",X"AE",X"47",X"A6",X"89",X"AE",X"A2",X"AE",X"4A",X"A4",X"89",X"E8",X"37",X"27",X"02",
		X"C6",X"01",X"4F",X"DD",X"32",X"39",X"9E",X"73",X"27",X"5C",X"96",X"A8",X"27",X"0A",X"9E",X"75",
		X"27",X"54",X"96",X"A9",X"27",X"4D",X"20",X"4E",X"10",X"9E",X"75",X"27",X"46",X"96",X"A9",X"26",
		X"42",X"E6",X"0B",X"E0",X"4B",X"25",X"01",X"50",X"E7",X"E2",X"EC",X"07",X"A3",X"47",X"25",X"05",
		X"43",X"53",X"C3",X"FF",X"FF",X"4D",X"26",X"06",X"E1",X"E4",X"22",X"02",X"E7",X"E4",X"E6",X"2B",
		X"E0",X"4B",X"25",X"01",X"50",X"E7",X"E2",X"EC",X"27",X"A3",X"47",X"25",X"05",X"43",X"53",X"C3",
		X"FF",X"FF",X"4D",X"26",X"06",X"E1",X"E4",X"22",X"02",X"E7",X"E4",X"E1",X"61",X"35",X"06",X"25",
		X"02",X"9E",X"75",X"1C",X"FB",X"39",X"1A",X"04",X"39",X"EC",X"47",X"10",X"83",X"00",X"04",X"2E",
		X"03",X"CC",X"00",X"04",X"10",X"83",X"01",X"20",X"2D",X"03",X"CC",X"01",X"20",X"ED",X"47",X"10",
		X"BE",X"00",X"2E",X"BD",X"8E",X"89",X"86",X"05",X"BD",X"E0",X"37",X"10",X"BE",X"00",X"2E",X"BD",
		X"8E",X"9F",X"10",X"BE",X"00",X"30",X"BD",X"8E",X"89",X"86",X"08",X"BD",X"E0",X"37",X"10",X"BE",
		X"00",X"30",X"BD",X"8E",X"9F",X"10",X"BE",X"00",X"32",X"BD",X"8E",X"89",X"86",X"0C",X"BD",X"E0",
		X"37",X"10",X"BE",X"00",X"32",X"BD",X"8E",X"9F",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"A9",X"E8",
		X"28",X"AA",X"A9",X"E8",X"2A",X"A4",X"89",X"AE",X"A2",X"9A",X"4B",X"97",X"4B",X"7E",X"E0",X"0F",
		X"86",X"05",X"A7",X"C8",X"10",X"10",X"AE",X"4E",X"BD",X"65",X"EE",X"86",X"0A",X"BD",X"E0",X"37",
		X"10",X"AE",X"4E",X"BD",X"65",X"EE",X"86",X"2A",X"A7",X"84",X"86",X"0A",X"BD",X"E0",X"37",X"6A",
		X"C8",X"10",X"26",X"E1",X"BD",X"82",X"40",X"86",X"02",X"BD",X"E0",X"37",X"10",X"8E",X"ED",X"19",
		X"86",X"05",X"A7",X"C8",X"12",X"AE",X"4E",X"BC",X"00",X"00",X"26",X"05",X"8E",X"F1",X"45",X"20",
		X"0C",X"BC",X"00",X"04",X"26",X"05",X"8E",X"31",X"51",X"20",X"02",X"AE",X"04",X"AF",X"C8",X"10",
		X"8D",X"17",X"10",X"AF",X"C8",X"13",X"86",X"08",X"BD",X"E0",X"37",X"10",X"AE",X"C8",X"13",X"6A",
		X"C8",X"12",X"26",X"D1",X"8D",X"3A",X"7E",X"E0",X"0F",X"AE",X"C8",X"10",X"A6",X"A0",X"27",X"2F",
		X"84",X"0F",X"C6",X"11",X"3D",X"A6",X"3F",X"84",X"F0",X"44",X"44",X"44",X"44",X"26",X"0A",X"AE",
		X"C8",X"10",X"30",X"01",X"AF",X"C8",X"10",X"20",X"E3",X"27",X"E1",X"81",X"01",X"26",X"02",X"C4",
		X"F0",X"E7",X"84",X"30",X"89",X"01",X"00",X"8C",X"98",X"00",X"22",X"D0",X"4A",X"20",X"EA",X"39",
		X"E6",X"27",X"C8",X"04",X"EB",X"25",X"BD",X"E0",X"1B",X"CC",X"12",X"00",X"ED",X"84",X"10",X"AE",
		X"4E",X"EC",X"22",X"ED",X"02",X"EC",X"24",X"ED",X"C8",X"10",X"ED",X"04",X"EC",X"26",X"C8",X"04",
		X"CB",X"0B",X"C8",X"04",X"ED",X"06",X"39",X"DC",X"73",X"26",X"07",X"DF",X"73",X"96",X"A7",X"97",
		X"A8",X"39",X"DF",X"75",X"96",X"A7",X"97",X"A9",X"39",X"0F",X"36",X"0C",X"A5",X"20",X"04",X"0F",
		X"37",X"0C",X"A6",X"C6",X"25",X"D7",X"AC",X"30",X"84",X"27",X"58",X"10",X"AE",X"0D",X"27",X"47",
		X"10",X"AE",X"A8",X"18",X"27",X"41",X"6C",X"A4",X"2E",X"49",X"27",X"04",X"6A",X"A4",X"20",X"43",
		X"0F",X"A3",X"0F",X"A4",X"86",X"80",X"A7",X"A4",X"AE",X"0D",X"34",X"10",X"86",X"30",X"BD",X"E6",
		X"A8",X"8E",X"78",X"61",X"CC",X"02",X"FF",X"BD",X"E0",X"30",X"EC",X"47",X"C3",X"00",X"06",X"ED",
		X"27",X"EC",X"4A",X"ED",X"2A",X"86",X"64",X"35",X"10",X"E6",X"88",X"2E",X"ED",X"A8",X"2E",X"8E",
		X"EF",X"80",X"BD",X"E0",X"2D",X"20",X"0C",X"96",X"90",X"2A",X"08",X"96",X"A0",X"27",X"04",X"86",
		X"02",X"97",X"B0",X"8E",X"81",X"39",X"CC",X"20",X"00",X"BD",X"E0",X"30",X"EC",X"47",X"ED",X"27",
		X"EC",X"4A",X"ED",X"2A",X"AE",X"4D",X"86",X"50",X"BD",X"E6",X"B1",X"BD",X"85",X"C1",X"8E",X"EF",
		X"B7",X"BD",X"E0",X"2D",X"11",X"93",X"73",X"26",X"08",X"DC",X"75",X"DD",X"73",X"96",X"A9",X"97",
		X"A8",X"CC",X"00",X"00",X"DD",X"75",X"AE",X"4D",X"AE",X"04",X"6A",X"06",X"26",X"19",X"96",X"90",
		X"2A",X"15",X"96",X"52",X"9A",X"5C",X"26",X"10",X"34",X"40",X"DE",X"0A",X"8E",X"61",X"F0",X"CC",
		X"34",X"00",X"BD",X"E0",X"30",X"35",X"40",X"39",X"8E",X"83",X"4B",X"CC",X"09",X"FF",X"BD",X"E0",
		X"30",X"86",X"16",X"A7",X"A8",X"2D",X"AE",X"4D",X"AF",X"2D",X"39",X"AE",X"4D",X"E6",X"88",X"2E",
		X"8D",X"16",X"86",X"08",X"BD",X"E0",X"37",X"96",X"90",X"27",X"05",X"6A",X"C8",X"2D",X"26",X"EB",
		X"AE",X"4D",X"5F",X"8D",X"03",X"7E",X"E0",X"0F",X"A6",X"88",X"30",X"8E",X"29",X"6C",X"BD",X"4A",
		X"53",X"30",X"89",X"03",X"00",X"86",X"6D",X"7E",X"4A",X"53",X"86",X"01",X"BD",X"E0",X"37",X"EE",
		X"C4",X"27",X"F7",X"A6",X"42",X"2A",X"F8",X"DF",X"93",X"30",X"C4",X"AE",X"84",X"27",X"F0",X"A6",
		X"02",X"2A",X"F8",X"A4",X"42",X"85",X"01",X"27",X"F2",X"8D",X"3D",X"24",X"EE",X"20",X"E0",X"86",
		X"01",X"BD",X"E0",X"37",X"96",X"A8",X"27",X"02",X"0A",X"A8",X"96",X"A9",X"27",X"02",X"0A",X"A9",
		X"EE",X"C4",X"27",X"EB",X"A6",X"42",X"81",X"89",X"26",X"F6",X"DF",X"93",X"30",X"C4",X"AE",X"84",
		X"27",X"DD",X"A6",X"02",X"2A",X"F8",X"8D",X"10",X"25",X"E6",X"AE",X"84",X"27",X"E2",X"A6",X"02",
		X"2A",X"F8",X"8D",X"04",X"24",X"F4",X"20",X"D8",X"9F",X"49",X"EC",X"47",X"A3",X"88",X"29",X"2E",
		X"34",X"EC",X"07",X"10",X"A3",X"C8",X"29",X"2E",X"2C",X"A3",X"47",X"DD",X"34",X"EC",X"88",X"27",
		X"E1",X"C8",X"27",X"22",X"20",X"A1",X"C8",X"28",X"25",X"1B",X"10",X"AE",X"98",X"1C",X"AE",X"D8",
		X"1C",X"E0",X"C8",X"28",X"58",X"58",X"2B",X"03",X"3A",X"20",X"03",X"50",X"31",X"A5",X"BD",X"DC",
		X"21",X"25",X"05",X"9E",X"49",X"1C",X"FE",X"39",X"9E",X"49",X"A6",X"42",X"A4",X"02",X"85",X"01",
		X"26",X"07",X"85",X"02",X"10",X"27",X"F1",X"0D",X"3F",X"85",X"04",X"26",X"5A",X"85",X"08",X"26",
		X"35",X"E6",X"C8",X"26",X"EB",X"4B",X"E0",X"0B",X"A6",X"88",X"17",X"81",X"0C",X"23",X"09",X"C0",
		X"08",X"2A",X"01",X"50",X"C1",X"03",X"20",X"07",X"C0",X"0A",X"2A",X"01",X"50",X"C1",X"02",X"22",
		X"15",X"A6",X"4F",X"A8",X"0F",X"2A",X"0F",X"DC",X"34",X"2A",X"07",X"A6",X"4F",X"2A",X"07",X"7E",
		X"85",X"0B",X"A6",X"4F",X"2A",X"F9",X"E6",X"C8",X"26",X"1D",X"ED",X"E3",X"E6",X"88",X"26",X"1D",
		X"A3",X"E1",X"E3",X"0A",X"A3",X"4A",X"27",X"05",X"2B",X"4C",X"7E",X"85",X"0B",X"8E",X"EF",X"CE",
		X"BD",X"E0",X"2D",X"9E",X"49",X"20",X"4A",X"8E",X"EF",X"9D",X"BD",X"E0",X"2D",X"9E",X"49",X"A6",
		X"42",X"81",X"97",X"27",X"0C",X"A6",X"02",X"81",X"97",X"27",X"12",X"BD",X"84",X"B7",X"7E",X"84",
		X"13",X"A6",X"02",X"81",X"97",X"27",X"F4",X"BD",X"85",X"D7",X"7E",X"84",X"13",X"1E",X"13",X"BD",
		X"85",X"D7",X"1E",X"13",X"7E",X"84",X"13",X"E6",X"0B",X"E0",X"4B",X"10",X"2A",X"00",X"60",X"10",
		X"27",X"00",X"76",X"7E",X"85",X"2D",X"9E",X"49",X"BD",X"84",X"E0",X"A6",X"02",X"81",X"97",X"27",
		X"05",X"BD",X"85",X"2D",X"20",X"07",X"1E",X"13",X"BD",X"85",X"D7",X"1E",X"13",X"1A",X"01",X"39",
		X"34",X"50",X"A6",X"42",X"84",X"7F",X"A7",X"42",X"CC",X"00",X"00",X"ED",X"C8",X"1A",X"10",X"AE",
		X"4D",X"CC",X"EE",X"C2",X"ED",X"C8",X"24",X"AD",X"B8",X"10",X"EE",X"62",X"10",X"AE",X"4D",X"A6",
		X"A8",X"2F",X"AE",X"E4",X"AE",X"0D",X"AD",X"B8",X"16",X"35",X"D0",X"9E",X"49",X"1E",X"13",X"BD",
		X"84",X"E0",X"1E",X"13",X"A6",X"42",X"81",X"97",X"27",X"8D",X"8D",X"03",X"7E",X"84",X"13",X"9E",
		X"49",X"1E",X"13",X"BD",X"85",X"99",X"1E",X"13",X"BD",X"85",X"AD",X"20",X"0C",X"9E",X"49",X"1E",
		X"13",X"BD",X"85",X"AD",X"1E",X"13",X"BD",X"85",X"99",X"9E",X"49",X"DC",X"34",X"27",X"58",X"2A",
		X"2C",X"A6",X"88",X"14",X"2F",X"06",X"40",X"8B",X"02",X"A7",X"88",X"14",X"40",X"8B",X"02",X"47",
		X"A7",X"C8",X"22",X"86",X"FF",X"A7",X"0F",X"A6",X"C8",X"14",X"2C",X"06",X"40",X"80",X"02",X"A7",
		X"C8",X"14",X"8B",X"02",X"40",X"47",X"A7",X"88",X"22",X"6F",X"4F",X"20",X"2A",X"A6",X"88",X"14",
		X"2C",X"06",X"40",X"80",X"02",X"A7",X"88",X"14",X"8B",X"02",X"40",X"47",X"A7",X"C8",X"22",X"6F",
		X"0F",X"A6",X"C8",X"14",X"2F",X"06",X"40",X"8B",X"02",X"A7",X"C8",X"14",X"40",X"8B",X"02",X"47",
		X"A7",X"88",X"22",X"86",X"FF",X"A7",X"4F",X"39",X"CE",X"86",X"FE",X"A7",X"88",X"23",X"EC",X"88",
		X"11",X"2F",X"09",X"43",X"50",X"82",X"FF",X"47",X"56",X"ED",X"88",X"11",X"39",X"86",X"02",X"A7",
		X"88",X"23",X"EC",X"88",X"11",X"2C",X"09",X"43",X"50",X"82",X"FF",X"47",X"56",X"ED",X"88",X"11",
		X"39",X"BE",X"86",X"36",X"CC",X"00",X"22",X"AB",X"80",X"5A",X"26",X"FB",X"81",X"32",X"27",X"06",
		X"AE",X"9F",X"A0",X"08",X"6C",X"01",X"39",X"4F",X"E6",X"88",X"27",X"E0",X"C8",X"27",X"82",X"00",
		X"EB",X"88",X"28",X"89",X"00",X"E0",X"C8",X"28",X"82",X"00",X"2A",X"09",X"8D",X"AB",X"86",X"FB",
		X"A7",X"88",X"23",X"20",X"07",X"8D",X"B6",X"86",X"05",X"A7",X"88",X"23",X"EC",X"07",X"A3",X"47",
		X"E3",X"88",X"29",X"A3",X"C8",X"29",X"2A",X"18",X"A6",X"88",X"14",X"2F",X"06",X"80",X"02",X"40",
		X"A7",X"88",X"14",X"A6",X"C8",X"14",X"40",X"48",X"A7",X"88",X"22",X"86",X"FF",X"A7",X"0F",X"39",
		X"A6",X"88",X"14",X"2C",X"06",X"40",X"80",X"02",X"A7",X"88",X"14",X"A6",X"C8",X"14",X"40",X"48",
		X"A7",X"88",X"22",X"6F",X"0F",X"39",X"F3",X"20",X"86",X"04",X"BD",X"E0",X"37",X"96",X"9D",X"81",
		X"DF",X"22",X"F5",X"86",X"01",X"BD",X"E0",X"37",X"AE",X"C8",X"2B",X"A6",X"89",X"B0",X"02",X"A8",
		X"89",X"EB",X"B8",X"84",X"20",X"A8",X"89",X"B0",X"02",X"A7",X"89",X"B0",X"02",X"84",X"20",X"26",
		X"43",X"E6",X"C8",X"2D",X"30",X"85",X"AF",X"C8",X"2B",X"E6",X"C8",X"14",X"30",X"85",X"8C",X"FF",
		X"F2",X"2D",X"D0",X"8C",X"01",X"28",X"2E",X"CB",X"AF",X"47",X"6C",X"C8",X"10",X"A6",X"C8",X"10",
		X"BD",X"86",X"EE",X"86",X"06",X"BD",X"E0",X"37",X"A6",X"C8",X"10",X"BD",X"86",X"F5",X"6C",X"C8",
		X"10",X"A6",X"C8",X"10",X"BD",X"86",X"EE",X"86",X"06",X"BD",X"E0",X"37",X"A6",X"C8",X"10",X"BD",
		X"86",X"F5",X"20",X"A4",X"6C",X"C8",X"10",X"A6",X"C8",X"10",X"BD",X"86",X"EE",X"86",X"06",X"BD",
		X"E0",X"37",X"A6",X"C8",X"10",X"BD",X"86",X"F5",X"A6",X"C8",X"10",X"84",X"03",X"26",X"E5",X"6C",
		X"4B",X"A6",X"4B",X"81",X"EF",X"25",X"DD",X"86",X"80",X"9A",X"4B",X"97",X"4B",X"7E",X"E0",X"0F",
		X"A6",X"C8",X"10",X"BD",X"86",X"F5",X"6C",X"C8",X"10",X"E6",X"4B",X"C1",X"DF",X"23",X"02",X"6A",
		X"4B",X"A6",X"C8",X"10",X"BD",X"86",X"EE",X"86",X"06",X"BD",X"E0",X"37",X"20",X"E2",X"34",X"02",
		X"BD",X"E0",X"24",X"20",X"05",X"34",X"02",X"BD",X"E0",X"21",X"35",X"02",X"10",X"BE",X"00",X"2C",
		X"84",X"03",X"48",X"31",X"A6",X"48",X"31",X"A6",X"BD",X"8E",X"70",X"7E",X"D8",X"F4",X"34",X"02",
		X"BD",X"87",X"19",X"6A",X"E4",X"26",X"F9",X"35",X"82",X"34",X"11",X"AE",X"04",X"27",X"2F",X"6C",
		X"05",X"6C",X"06",X"26",X"04",X"6A",X"05",X"6A",X"06",X"A6",X"05",X"81",X"05",X"22",X"1F",X"48",
		X"AB",X"05",X"80",X"03",X"5F",X"AE",X"61",X"E3",X"06",X"1A",X"F0",X"FD",X"CA",X"04",X"CC",X"07",
		X"03",X"FD",X"CA",X"06",X"EC",X"08",X"FD",X"CA",X"02",X"86",X"0A",X"B7",X"CA",X"00",X"35",X"91",
		X"34",X"10",X"AE",X"04",X"27",X"3B",X"A6",X"05",X"27",X"37",X"D6",X"90",X"2A",X"05",X"C6",X"07",
		X"BD",X"3B",X"2B",X"4A",X"A7",X"05",X"81",X"04",X"22",X"25",X"48",X"AB",X"05",X"5F",X"AE",X"E4",
		X"E3",X"06",X"34",X"01",X"1A",X"F0",X"FD",X"CA",X"04",X"CC",X"07",X"03",X"FD",X"CA",X"06",X"EC",
		X"08",X"FD",X"CA",X"02",X"CC",X"1A",X"EE",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"01",X"86",
		X"01",X"35",X"90",X"34",X"01",X"1A",X"F0",X"FD",X"CA",X"04",X"EC",X"81",X"88",X"04",X"C8",X"04",
		X"FD",X"CA",X"06",X"BF",X"CA",X"02",X"1F",X"20",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"81",
		X"34",X"10",X"DC",X"6E",X"DD",X"6A",X"DC",X"70",X"DD",X"6C",X"EE",X"9F",X"A0",X"0A",X"EE",X"C4",
		X"26",X"02",X"35",X"90",X"A6",X"42",X"2A",X"F6",X"81",X"82",X"26",X"05",X"EC",X"C8",X"2B",X"27",
		X"ED",X"E6",X"C8",X"14",X"10",X"AE",X"E4",X"AE",X"A1",X"EC",X"85",X"E3",X"47",X"10",X"83",X"FF",
		X"F6",X"2C",X"03",X"C3",X"01",X"2E",X"10",X"83",X"01",X"24",X"2F",X"03",X"C3",X"FE",X"D2",X"1F",
		X"01",X"A6",X"4B",X"81",X"58",X"22",X"08",X"96",X"6A",X"26",X"C3",X"8D",X"27",X"20",X"BF",X"81",
		X"91",X"22",X"12",X"31",X"27",X"96",X"6B",X"26",X"02",X"8D",X"19",X"96",X"6C",X"26",X"AF",X"31",
		X"27",X"8D",X"11",X"20",X"A9",X"81",X"AA",X"25",X"A5",X"96",X"6D",X"26",X"A1",X"31",X"A8",X"15",
		X"8D",X"02",X"20",X"9A",X"E6",X"A4",X"26",X"0A",X"AC",X"21",X"25",X"11",X"AC",X"23",X"22",X"0D",
		X"20",X"08",X"AC",X"21",X"22",X"04",X"AC",X"23",X"22",X"03",X"6C",X"B8",X"05",X"39",X"88",X"82",
		X"00",X"00",X"28",X"00",X"BA",X"A0",X"6A",X"00",X"00",X"9E",X"01",X"15",X"A0",X"6B",X"01",X"01",
		X"0D",X"00",X"60",X"A0",X"6C",X"00",X"00",X"36",X"00",X"C8",X"A0",X"6D",X"88",X"82",X"00",X"00",
		X"10",X"00",X"D2",X"A0",X"6A",X"01",X"00",X"86",X"00",X"24",X"A0",X"6B",X"01",X"00",X"DA",X"00",
		X"78",X"A0",X"6C",X"00",X"00",X"1E",X"00",X"E0",X"A0",X"6D",X"FF",X"C4",X"FF",X"E2",X"FF",X"F1",
		X"FF",X"F8",X"00",X"00",X"00",X"08",X"00",X"0F",X"00",X"1E",X"00",X"3C",X"61",X"DA",X"61",X"DA",
		X"A0",X"4C",X"39",X"D9",X"E8",X"0D",X"00",X"1E",X"8A",X"45",X"8A",X"AA",X"82",X"79",X"A0",X"36",
		X"82",X"67",X"E6",X"A8",X"A0",X"A3",X"8A",X"A6",X"EF",X"D3",X"EF",X"D6",X"EF",X"DF",X"EF",X"E2",
		X"EF",X"D9",X"EF",X"DC",X"EF",X"E5",X"00",X"00",X"EF",X"BA",X"55",X"20",X"65",X"61",X"DA",X"61",
		X"DA",X"A0",X"56",X"60",X"D9",X"E8",X"22",X"00",X"20",X"8A",X"4D",X"8A",X"AA",X"82",X"7F",X"A0",
		X"37",X"82",X"67",X"E6",X"A8",X"A0",X"A4",X"8A",X"A6",X"EF",X"D3",X"EF",X"D6",X"EF",X"DF",X"EF",
		X"E2",X"EF",X"D9",X"EF",X"DC",X"EF",X"E5",X"00",X"00",X"EF",X"C1",X"77",X"20",X"66",X"DD",X"B2",
		X"DD",X"B2",X"A0",X"4C",X"39",X"D9",X"E8",X"0D",X"00",X"1E",X"8A",X"45",X"8A",X"AA",X"82",X"79",
		X"A0",X"36",X"82",X"67",X"E6",X"A8",X"A0",X"A3",X"8A",X"A6",X"EF",X"D3",X"EF",X"D6",X"EF",X"DF",
		X"EF",X"E2",X"EF",X"D9",X"EF",X"DC",X"EF",X"E5",X"EF",X"C8",X"EF",X"BA",X"55",X"20",X"65",X"DD",
		X"B9",X"DD",X"B9",X"A0",X"56",X"60",X"D9",X"E8",X"22",X"00",X"20",X"8A",X"4D",X"8A",X"AA",X"82",
		X"7F",X"A0",X"37",X"82",X"67",X"E6",X"A8",X"A0",X"A4",X"8A",X"A6",X"EF",X"D3",X"EF",X"D6",X"EF",
		X"DF",X"EF",X"E2",X"EF",X"D9",X"EF",X"DC",X"EF",X"E5",X"EF",X"C8",X"EF",X"C1",X"77",X"20",X"66",
		X"EE",X"C2",X"EE",X"C2",X"00",X"00",X"00",X"00",X"E8",X"22",X"00",X"22",X"8A",X"55",X"8A",X"A7",
		X"74",X"C3",X"00",X"00",X"8A",X"7D",X"E6",X"B1",X"00",X"00",X"A0",X"B0",X"EF",X"A2",X"EF",X"A5",
		X"EF",X"AE",X"EF",X"B1",X"EF",X"A8",X"EF",X"AB",X"EF",X"B4",X"00",X"00",X"EF",X"92",X"11",X"10",
		X"6D",X"7A",X"83",X"7B",X"0B",X"00",X"00",X"00",X"00",X"E8",X"22",X"00",X"22",X"8A",X"55",X"8A",
		X"A7",X"74",X"C3",X"00",X"00",X"8A",X"7D",X"E6",X"B1",X"00",X"00",X"A0",X"B0",X"EF",X"A2",X"EF",
		X"A5",X"EF",X"AE",X"EF",X"B1",X"EF",X"A8",X"EF",X"AB",X"EF",X"B4",X"00",X"00",X"EF",X"92",X"11",
		X"05",X"6D",X"7A",X"83",X"7C",X"95",X"00",X"00",X"00",X"00",X"E8",X"22",X"00",X"24",X"8A",X"55",
		X"8A",X"A7",X"74",X"C3",X"00",X"00",X"8A",X"7D",X"E6",X"B1",X"00",X"00",X"A0",X"B0",X"EF",X"A2",
		X"EF",X"A5",X"EF",X"AE",X"EF",X"B1",X"EF",X"A8",X"EF",X"AB",X"EF",X"B4",X"00",X"00",X"EF",X"92",
		X"11",X"57",X"6D",X"7A",X"83",X"7E",X"CF",X"00",X"00",X"00",X"00",X"E8",X"22",X"00",X"26",X"8A",
		X"55",X"8A",X"A7",X"74",X"C3",X"00",X"00",X"8A",X"7D",X"E6",X"A8",X"00",X"00",X"A0",X"B0",X"EF",
		X"A2",X"EF",X"A5",X"EF",X"AE",X"EF",X"B1",X"EF",X"A8",X"EF",X"AB",X"EF",X"B4",X"00",X"00",X"EF",
		X"92",X"11",X"15",X"6D",X"7A",X"83",X"66",X"40",X"00",X"00",X"00",X"00",X"E8",X"22",X"00",X"00",
		X"8A",X"55",X"8A",X"A7",X"74",X"AE",X"00",X"00",X"8A",X"7D",X"E6",X"A8",X"00",X"00",X"A0",X"B0",
		X"EF",X"A2",X"EF",X"A5",X"EF",X"AE",X"EF",X"B1",X"00",X"00",X"00",X"00",X"EF",X"B4",X"00",X"00",
		X"EF",X"92",X"11",X"10",X"6D",X"55",X"55",X"11",X"55",X"55",X"DD",X"55",X"55",X"77",X"77",X"11",
		X"77",X"77",X"DD",X"77",X"77",X"11",X"11",X"DD",X"11",X"11",X"DD",X"11",X"11",X"00",X"10",X"00",
		X"71",X"00",X"50",X"A0",X"6E",X"00",X"12",X"00",X"E7",X"00",X"80",X"A0",X"6F",X"00",X"14",X"00",
		X"17",X"00",X"89",X"A0",X"70",X"00",X"16",X"00",X"7F",X"00",X"D2",X"A0",X"71",X"39",X"4A",X"4F",
		X"55",X"53",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"20",X"49",X"4E",X"43",X"2E",X"01",X"7E",X"E0",X"0F",X"AE",X"4D",X"BD",X"87",X"50",X"27",
		X"F6",X"96",X"38",X"A7",X"C8",X"16",X"0C",X"38",X"20",X"5B",X"D1",X"39",X"26",X"57",X"0F",X"88",
		X"0F",X"89",X"0F",X"8A",X"AE",X"9F",X"A0",X"0A",X"AE",X"84",X"27",X"12",X"A6",X"02",X"2A",X"F8",
		X"81",X"82",X"26",X"05",X"EC",X"88",X"2B",X"27",X"EF",X"BD",X"D8",X"00",X"20",X"EA",X"DC",X"6E",
		X"DD",X"6A",X"DC",X"70",X"DD",X"6C",X"96",X"8A",X"26",X"04",X"96",X"6D",X"27",X"67",X"96",X"89",
		X"26",X"08",X"96",X"6B",X"27",X"51",X"96",X"6C",X"27",X"54",X"96",X"88",X"26",X"04",X"96",X"6A",
		X"27",X"3E",X"8E",X"88",X"5C",X"96",X"3C",X"26",X"27",X"8E",X"88",X"3E",X"20",X"22",X"96",X"3A",
		X"A7",X"C8",X"16",X"0C",X"3A",X"86",X"01",X"BD",X"E0",X"37",X"E6",X"C8",X"16",X"A6",X"42",X"81",
		X"09",X"27",X"97",X"96",X"38",X"91",X"39",X"26",X"EC",X"D1",X"3B",X"26",X"E8",X"8E",X"88",X"3E",
		X"BD",X"87",X"B0",X"BD",X"E0",X"18",X"24",X"05",X"46",X"25",X"1A",X"20",X"11",X"46",X"25",X"07",
		X"8E",X"8A",X"5D",X"96",X"6A",X"27",X"31",X"8E",X"8A",X"65",X"96",X"6B",X"27",X"2A",X"8E",X"8A",
		X"6D",X"96",X"6C",X"27",X"23",X"8E",X"8A",X"75",X"96",X"6D",X"27",X"1C",X"8E",X"8A",X"5D",X"96",
		X"6A",X"27",X"15",X"8E",X"8A",X"65",X"96",X"6B",X"27",X"0E",X"8E",X"8A",X"6D",X"96",X"6C",X"27",
		X"07",X"8E",X"8A",X"75",X"96",X"6D",X"26",X"9D",X"6C",X"98",X"06",X"DE",X"2E",X"EC",X"02",X"ED",
		X"47",X"EC",X"04",X"ED",X"4A",X"AF",X"C8",X"20",X"AE",X"4D",X"AE",X"88",X"2C",X"A6",X"42",X"81",
		X"09",X"26",X"04",X"0C",X"39",X"20",X"02",X"0C",X"3B",X"BD",X"E0",X"2D",X"86",X"1E",X"A7",X"C8",
		X"10",X"10",X"AE",X"4D",X"EC",X"B8",X"0A",X"ED",X"C8",X"1A",X"86",X"0C",X"BD",X"8E",X"05",X"AE",
		X"C8",X"20",X"10",X"AE",X"94",X"BD",X"65",X"EE",X"A6",X"84",X"8A",X"10",X"10",X"AE",X"4D",X"E6",
		X"A8",X"2E",X"ED",X"84",X"A6",X"C8",X"10",X"81",X"14",X"2E",X"4C",X"BD",X"8E",X"4D",X"E6",X"C8",
		X"10",X"1F",X"98",X"43",X"47",X"84",X"0F",X"88",X"04",X"A7",X"07",X"1F",X"89",X"81",X"03",X"2F",
		X"02",X"C6",X"03",X"E7",X"1D",X"88",X"04",X"40",X"4C",X"4C",X"84",X"0F",X"1F",X"89",X"AB",X"05",
		X"EB",X"1B",X"A7",X"05",X"E7",X"1B",X"E6",X"07",X"C8",X"04",X"EB",X"05",X"E1",X"4B",X"23",X"09",
		X"E6",X"4B",X"5C",X"E0",X"05",X"C8",X"04",X"E7",X"07",X"10",X"AE",X"4D",X"E6",X"A8",X"2E",X"A6",
		X"84",X"8A",X"10",X"ED",X"84",X"ED",X"16",X"86",X"01",X"BD",X"E0",X"37",X"BD",X"8E",X"99",X"86",
		X"12",X"A7",X"84",X"EC",X"47",X"47",X"56",X"E7",X"04",X"86",X"0D",X"A7",X"06",X"6A",X"C8",X"10",
		X"10",X"26",X"FF",X"7B",X"AE",X"4D",X"EC",X"84",X"ED",X"C8",X"24",X"86",X"20",X"A7",X"C8",X"35",
		X"44",X"A7",X"C8",X"15",X"86",X"02",X"A7",X"C8",X"26",X"6F",X"C8",X"13",X"6F",X"C8",X"16",X"20",
		X"05",X"86",X"01",X"BD",X"E0",X"37",X"AD",X"D8",X"24",X"DC",X"32",X"26",X"6E",X"6A",X"C8",X"13",
		X"2E",X"0A",X"86",X"4B",X"A7",X"C8",X"13",X"64",X"C8",X"35",X"27",X"69",X"BD",X"8E",X"4D",X"AE",
		X"C8",X"20",X"10",X"AE",X"94",X"BD",X"65",X"EE",X"10",X"AE",X"4D",X"10",X"AE",X"2C",X"30",X"88",
		X"EC",X"E6",X"C8",X"26",X"8D",X"1F",X"5A",X"8D",X"1C",X"5A",X"8D",X"19",X"6A",X"C8",X"15",X"2E",
		X"09",X"6C",X"C8",X"26",X"A6",X"C8",X"35",X"A7",X"C8",X"15",X"A6",X"C8",X"35",X"44",X"26",X"B1",
		X"6C",X"C8",X"16",X"20",X"AC",X"34",X"04",X"C4",X"07",X"26",X"07",X"C6",X"02",X"E7",X"C8",X"26",
		X"E7",X"E4",X"E6",X"A5",X"6D",X"C8",X"16",X"27",X"08",X"C1",X"55",X"27",X"0A",X"C1",X"77",X"27",
		X"06",X"A6",X"84",X"8A",X"10",X"ED",X"84",X"30",X"0A",X"35",X"84",X"AE",X"4D",X"AE",X"88",X"2A",
		X"27",X"03",X"BD",X"E0",X"2D",X"BD",X"8E",X"8E",X"AE",X"C8",X"20",X"6A",X"98",X"06",X"10",X"AE",
		X"94",X"BD",X"65",X"EE",X"DE",X"2E",X"AE",X"4D",X"AD",X"98",X"14",X"8D",X"04",X"DC",X"32",X"20",
		X"5F",X"EC",X"98",X"0A",X"ED",X"C8",X"1A",X"CC",X"DC",X"E6",X"ED",X"C8",X"20",X"CC",X"00",X"00",
		X"ED",X"C8",X"11",X"6F",X"C8",X"14",X"6F",X"C8",X"16",X"6F",X"C8",X"10",X"6F",X"C8",X"13",X"6F",
		X"C8",X"15",X"6F",X"C8",X"22",X"6F",X"C8",X"23",X"86",X"80",X"AA",X"42",X"A7",X"42",X"86",X"0C",
		X"7E",X"8D",X"F6",X"CC",X"00",X"D2",X"ED",X"4A",X"86",X"3C",X"BD",X"E0",X"37",X"AE",X"4D",X"BD",
		X"87",X"50",X"DE",X"2E",X"AE",X"4D",X"AD",X"98",X"14",X"AE",X"4D",X"EC",X"84",X"ED",X"C8",X"24",
		X"8D",X"AF",X"BD",X"8E",X"4D",X"AE",X"4D",X"A6",X"98",X"1A",X"BD",X"E0",X"37",X"AD",X"D8",X"24",
		X"6D",X"C8",X"13",X"26",X"05",X"5D",X"10",X"26",X"01",X"4A",X"E7",X"C8",X"13",X"E6",X"4F",X"2A",
		X"01",X"40",X"E6",X"C8",X"15",X"27",X"05",X"6A",X"C8",X"15",X"26",X"23",X"AE",X"C8",X"20",X"8B",
		X"04",X"E6",X"86",X"27",X"1A",X"86",X"08",X"A7",X"C8",X"15",X"6F",X"C8",X"16",X"30",X"85",X"AF",
		X"C8",X"20",X"8C",X"DD",X"2C",X"26",X"08",X"AE",X"4D",X"AE",X"88",X"22",X"BD",X"E0",X"2D",X"6A",
		X"C8",X"16",X"2F",X"0B",X"E6",X"C8",X"22",X"27",X"AC",X"BD",X"8E",X"8E",X"5F",X"20",X"1F",X"BD",
		X"8E",X"8E",X"DC",X"32",X"AE",X"C8",X"20",X"A6",X"06",X"A7",X"C8",X"14",X"A6",X"80",X"A7",X"C8",
		X"16",X"AD",X"94",X"A7",X"C8",X"17",X"A6",X"4F",X"2A",X"04",X"60",X"C8",X"14",X"50",X"BD",X"DD",
		X"D2",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"89",X"B0",X"02",X"A4",X"A9",X"EA",X"98",X"84",X"7F",
		X"10",X"27",X"00",X"F4",X"A6",X"89",X"AE",X"A8",X"A4",X"A9",X"E8",X"37",X"27",X"11",X"9A",X"4B",
		X"97",X"4B",X"6F",X"4F",X"A6",X"C8",X"22",X"2A",X"01",X"40",X"8B",X"03",X"A7",X"C8",X"22",X"8D",
		X"08",X"8D",X"5A",X"7E",X"8D",X"45",X"A7",X"C8",X"17",X"E6",X"4B",X"E7",X"C8",X"27",X"C0",X"13",
		X"E7",X"C8",X"28",X"20",X"0F",X"A7",X"C8",X"17",X"E6",X"4B",X"C0",X"06",X"E7",X"C8",X"27",X"C0",
		X"0D",X"E7",X"C8",X"28",X"EC",X"47",X"C3",X"00",X"10",X"ED",X"C8",X"29",X"6F",X"C8",X"26",X"5F",
		X"A6",X"4F",X"2A",X"02",X"C6",X"06",X"EB",X"C8",X"17",X"AE",X"C8",X"18",X"3A",X"AF",X"C8",X"1C",
		X"AE",X"C8",X"1A",X"27",X"0A",X"C1",X"0C",X"25",X"0A",X"E0",X"C8",X"17",X"CB",X"0C",X"3A",X"AF",
		X"C8",X"1E",X"39",X"3A",X"AF",X"C8",X"1E",X"C6",X"02",X"E7",X"C8",X"26",X"39",X"DE",X"2E",X"10",
		X"AE",X"C8",X"1E",X"27",X"2E",X"BD",X"E0",X"2A",X"EC",X"22",X"9B",X"30",X"DB",X"31",X"ED",X"04",
		X"10",X"AE",X"24",X"EC",X"A1",X"ED",X"06",X"10",X"AF",X"02",X"30",X"0A",X"10",X"AE",X"C8",X"1C",
		X"EC",X"22",X"9B",X"30",X"DB",X"31",X"ED",X"04",X"10",X"AE",X"24",X"EC",X"A1",X"ED",X"06",X"10",
		X"AF",X"02",X"39",X"10",X"AE",X"C8",X"1C",X"27",X"F9",X"BD",X"E0",X"24",X"20",X"E2",X"10",X"AE",
		X"C8",X"1E",X"27",X"05",X"BD",X"E0",X"27",X"20",X"BF",X"10",X"AE",X"C8",X"1C",X"27",X"E3",X"BD",
		X"E0",X"21",X"20",X"CC",X"BD",X"8E",X"8E",X"CC",X"FF",X"80",X"ED",X"C8",X"11",X"6A",X"4B",X"6F",
		X"4C",X"6F",X"49",X"6F",X"C8",X"23",X"CC",X"00",X"00",X"ED",X"C8",X"20",X"CC",X"D8",X"58",X"ED",
		X"C8",X"30",X"6C",X"C8",X"15",X"7E",X"8F",X"6D",X"A6",X"C8",X"10",X"2A",X"08",X"AE",X"4D",X"AE",
		X"88",X"28",X"BD",X"E0",X"2D",X"6F",X"4C",X"6F",X"49",X"6F",X"C8",X"23",X"86",X"0A",X"A7",X"C8",
		X"15",X"CC",X"00",X"00",X"ED",X"C8",X"11",X"ED",X"C8",X"20",X"CC",X"D8",X"58",X"ED",X"C8",X"30",
		X"6F",X"C8",X"13",X"96",X"33",X"26",X"13",X"20",X"4A",X"BD",X"8E",X"4D",X"AE",X"4D",X"A6",X"98",
		X"1A",X"BD",X"E0",X"37",X"BD",X"D8",X"3D",X"5D",X"27",X"1B",X"5F",X"8E",X"DC",X"D5",X"AD",X"D8",
		X"30",X"A6",X"C8",X"15",X"2F",X"03",X"6A",X"C8",X"15",X"86",X"48",X"BD",X"8E",X"05",X"BD",X"D9",
		X"A3",X"26",X"D6",X"20",X"62",X"AE",X"4D",X"AE",X"88",X"1C",X"BD",X"E0",X"2D",X"6F",X"C8",X"13",
		X"20",X"11",X"BD",X"8E",X"4D",X"AE",X"4D",X"A6",X"98",X"1A",X"BD",X"E0",X"37",X"BD",X"D8",X"3D",
		X"5D",X"26",X"20",X"C6",X"04",X"8E",X"DC",X"D5",X"AD",X"D8",X"30",X"A6",X"C8",X"15",X"2F",X"07",
		X"6A",X"C8",X"15",X"86",X"48",X"20",X"02",X"86",X"60",X"BD",X"8E",X"05",X"BD",X"D9",X"A3",X"26",
		X"D1",X"20",X"24",X"BD",X"D8",X"13",X"5F",X"8E",X"DC",X"D5",X"AD",X"D8",X"30",X"AE",X"4D",X"AE",
		X"88",X"1E",X"BD",X"E0",X"2D",X"6F",X"C8",X"13",X"E6",X"C8",X"15",X"86",X"05",X"A7",X"C8",X"15",
		X"5D",X"2F",X"96",X"86",X"60",X"20",X"94",X"A6",X"C8",X"14",X"27",X"08",X"6F",X"4F",X"4D",X"2A",
		X"03",X"63",X"4F",X"40",X"8E",X"8F",X"B5",X"AE",X"86",X"AF",X"C8",X"20",X"6F",X"C8",X"16",X"6F",
		X"C8",X"15",X"86",X"01",X"A7",X"C8",X"13",X"CC",X"00",X"00",X"ED",X"C8",X"11",X"86",X"0C",X"A7",
		X"C8",X"17",X"7E",X"8D",X"EF",X"DC",X"E6",X"DC",X"ED",X"DC",X"F4",X"DC",X"FB",X"DD",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
