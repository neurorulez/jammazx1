library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bubbles_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bubbles_sound is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AA",X"0F",X"8E",X"00",X"7F",X"CE",X"04",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"00",
		X"C6",X"80",X"E7",X"02",X"86",X"37",X"A7",X"03",X"86",X"3C",X"A7",X"01",X"E7",X"02",X"CE",X"00",
		X"7F",X"6F",X"00",X"09",X"26",X"FB",X"86",X"3C",X"97",X"16",X"0E",X"20",X"FE",X"CE",X"F0",X"33",
		X"7E",X"F0",X"ED",X"10",X"FF",X"01",X"01",X"01",X"CE",X"F0",X"3E",X"7E",X"F0",X"ED",X"C0",X"FF",
		X"01",X"01",X"01",X"CE",X"A5",X"00",X"DF",X"16",X"CE",X"F0",X"5D",X"BD",X"F1",X"CF",X"CE",X"F0",
		X"8B",X"BD",X"F0",X"D8",X"BD",X"F1",X"73",X"CE",X"F0",X"90",X"7E",X"F0",X"ED",X"FE",X"34",X"02",
		X"16",X"60",X"D6",X"6E",X"FF",X"08",X"28",X"C8",X"2A",X"02",X"10",X"60",X"B6",X"3A",X"02",X"18",
		X"64",X"AC",X"64",X"FE",X"18",X"38",X"A1",X"38",X"02",X"14",X"68",X"90",X"34",X"02",X"12",X"60",
		X"7E",X"20",X"02",X"08",X"78",X"76",X"58",X"FF",X"18",X"22",X"00",X"C0",X"60",X"FC",X"01",X"01",
		X"FF",X"A0",X"FC",X"FF",X"08",X"18",X"F0",X"10",X"01",X"30",X"04",X"80",X"04",X"FE",X"30",X"CE",
		X"F0",X"95",X"8D",X"34",X"8D",X"14",X"8D",X"12",X"86",X"28",X"97",X"3D",X"73",X"00",X"25",X"8D",
		X"3E",X"73",X"00",X"25",X"86",X"1E",X"8D",X"0D",X"20",X"EA",X"86",X"30",X"97",X"3D",X"8D",X"2F",
		X"86",X"02",X"8D",X"01",X"39",X"16",X"CE",X"04",X"00",X"17",X"4A",X"26",X"FD",X"09",X"8C",X"00",
		X"00",X"26",X"F6",X"86",X"F0",X"97",X"21",X"39",X"A6",X"00",X"97",X"38",X"A6",X"01",X"97",X"21",
		X"A6",X"02",X"97",X"20",X"A6",X"03",X"97",X"25",X"A6",X"04",X"97",X"3D",X"39",X"8D",X"E9",X"8D",
		X"30",X"8D",X"58",X"96",X"3C",X"91",X"3D",X"26",X"F8",X"59",X"F7",X"04",X"00",X"8D",X"2D",X"8D",
		X"38",X"8D",X"5C",X"7D",X"00",X"21",X"27",X"E4",X"7D",X"00",X"22",X"26",X"E4",X"7D",X"00",X"25",
		X"27",X"DF",X"2B",X"05",X"7C",X"00",X"3D",X"20",X"D8",X"7A",X"00",X"3D",X"7A",X"00",X"3C",X"20",
		X"D0",X"7F",X"00",X"22",X"96",X"3D",X"97",X"3C",X"7F",X"00",X"3B",X"39",X"96",X"17",X"44",X"44",
		X"44",X"98",X"17",X"97",X"36",X"08",X"84",X"07",X"39",X"96",X"36",X"44",X"76",X"00",X"16",X"76",
		X"00",X"17",X"86",X"00",X"24",X"02",X"96",X"21",X"97",X"3B",X"39",X"96",X"3D",X"7A",X"00",X"3C",
		X"27",X"04",X"08",X"09",X"20",X"08",X"97",X"3C",X"D6",X"3B",X"54",X"7C",X"00",X"22",X"39",X"96",
		X"38",X"91",X"22",X"27",X"04",X"08",X"09",X"20",X"09",X"7F",X"00",X"22",X"96",X"21",X"90",X"20",
		X"97",X"21",X"39",X"7F",X"00",X"2F",X"7F",X"00",X"39",X"86",X"0E",X"97",X"30",X"7F",X"00",X"35",
		X"8D",X"9F",X"8D",X"A8",X"BD",X"F2",X"09",X"8D",X"B0",X"BD",X"F2",X"09",X"8D",X"BD",X"8D",X"79",
		X"8D",X"CD",X"8D",X"75",X"8D",X"0A",X"8D",X"71",X"8D",X"1D",X"8D",X"6D",X"8D",X"52",X"20",X"E2",
		X"96",X"34",X"7A",X"00",X"30",X"27",X"07",X"B6",X"00",X"21",X"26",X"0A",X"20",X"68",X"97",X"30",
		X"96",X"2F",X"9B",X"39",X"97",X"2F",X"39",X"96",X"2F",X"91",X"37",X"27",X"07",X"08",X"96",X"21",
		X"26",X"2A",X"20",X"29",X"7F",X"00",X"2F",X"7F",X"00",X"39",X"7F",X"00",X"35",X"DE",X"31",X"A6",
		X"00",X"97",X"2E",X"27",X"17",X"A6",X"01",X"97",X"33",X"A6",X"02",X"97",X"3A",X"A6",X"03",X"97",
		X"34",X"A6",X"04",X"97",X"37",X"86",X"05",X"BD",X"F5",X"74",X"DF",X"31",X"39",X"32",X"32",X"39",
		X"96",X"2E",X"27",X"06",X"91",X"21",X"26",X"04",X"20",X"03",X"08",X"09",X"39",X"7F",X"00",X"2E",
		X"96",X"33",X"97",X"2F",X"96",X"3A",X"97",X"39",X"39",X"96",X"35",X"9B",X"2F",X"97",X"35",X"2A",
		X"01",X"43",X"1B",X"B7",X"04",X"00",X"39",X"16",X"48",X"48",X"48",X"1B",X"CE",X"00",X"20",X"DF",
		X"1C",X"CE",X"F5",X"FD",X"BD",X"F5",X"74",X"C6",X"09",X"7E",X"F3",X"16",X"96",X"28",X"B7",X"04",
		X"00",X"DE",X"20",X"DF",X"29",X"DE",X"25",X"96",X"29",X"73",X"04",X"00",X"09",X"27",X"10",X"4A",
		X"26",X"FA",X"96",X"2A",X"73",X"04",X"00",X"09",X"27",X"05",X"4A",X"26",X"FA",X"20",X"E8",X"B6",
		X"04",X"00",X"2B",X"01",X"43",X"8B",X"00",X"B7",X"04",X"00",X"96",X"29",X"9B",X"22",X"97",X"29",
		X"96",X"2A",X"9B",X"23",X"97",X"2A",X"91",X"24",X"26",X"CB",X"96",X"27",X"27",X"06",X"9B",X"20",
		X"97",X"20",X"26",X"BD",X"39",X"86",X"01",X"20",X"0A",X"86",X"02",X"20",X"06",X"86",X"03",X"20",
		X"02",X"86",X"04",X"7F",X"00",X"20",X"97",X"1E",X"CE",X"FE",X"BA",X"A6",X"00",X"27",X"2D",X"7A",
		X"00",X"1E",X"27",X"06",X"4C",X"BD",X"F5",X"74",X"20",X"F1",X"08",X"DF",X"1C",X"BD",X"F5",X"74",
		X"DF",X"1A",X"DE",X"1C",X"A6",X"00",X"97",X"23",X"A6",X"01",X"EE",X"02",X"DF",X"21",X"8D",X"0F",
		X"DE",X"1C",X"08",X"08",X"08",X"08",X"DF",X"1C",X"9C",X"1A",X"26",X"E8",X"7E",X"F5",X"18",X"CE",
		X"00",X"24",X"81",X"00",X"27",X"15",X"81",X"03",X"27",X"09",X"C6",X"01",X"E7",X"00",X"08",X"80",
		X"02",X"20",X"EF",X"C6",X"91",X"E7",X"00",X"6F",X"01",X"08",X"08",X"C6",X"7E",X"E7",X"00",X"C6",
		X"F2",X"E7",X"01",X"C6",X"E9",X"E7",X"02",X"DE",X"21",X"4F",X"F6",X"00",X"1F",X"5C",X"D7",X"1F",
		X"D4",X"23",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",
		X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"48",X"48",X"48",X"48",X"48",X"B7",X"04",X"00",X"09",
		X"27",X"03",X"7E",X"00",X"24",X"39",X"36",X"A6",X"00",X"DF",X"1A",X"DE",X"1C",X"A7",X"00",X"08",
		X"DF",X"1C",X"DE",X"1A",X"08",X"5A",X"26",X"EF",X"32",X"39",X"CE",X"F6",X"57",X"DF",X"22",X"DE",
		X"22",X"A6",X"00",X"27",X"33",X"E6",X"01",X"C4",X"F0",X"D7",X"21",X"E6",X"01",X"08",X"08",X"DF",
		X"22",X"97",X"20",X"C4",X"0F",X"96",X"21",X"B7",X"04",X"00",X"96",X"20",X"CE",X"00",X"05",X"09",
		X"26",X"FD",X"4A",X"26",X"F7",X"7F",X"04",X"00",X"96",X"20",X"CE",X"00",X"05",X"09",X"26",X"FD",
		X"4A",X"26",X"F7",X"5A",X"26",X"DF",X"20",X"C7",X"39",X"7F",X"00",X"10",X"7F",X"00",X"11",X"39",
		X"96",X"10",X"8A",X"80",X"97",X"10",X"86",X"3C",X"97",X"11",X"39",X"86",X"04",X"BD",X"F3",X"90",
		X"96",X"11",X"48",X"48",X"43",X"BD",X"F4",X"4A",X"7C",X"00",X"24",X"BD",X"F4",X"4C",X"20",X"F8",
		X"16",X"58",X"1B",X"1B",X"1B",X"CE",X"F7",X"34",X"BD",X"F5",X"74",X"A6",X"00",X"16",X"84",X"0F",
		X"97",X"21",X"54",X"54",X"54",X"54",X"D7",X"20",X"A6",X"01",X"16",X"54",X"54",X"54",X"54",X"D7",
		X"22",X"84",X"0F",X"97",X"1E",X"DF",X"18",X"CE",X"F6",X"75",X"7A",X"00",X"1E",X"2B",X"08",X"A6",
		X"00",X"4C",X"BD",X"F5",X"74",X"20",X"F3",X"DF",X"25",X"BD",X"F4",X"86",X"DE",X"18",X"A6",X"02",
		X"97",X"27",X"BD",X"F4",X"98",X"DE",X"18",X"A6",X"03",X"97",X"23",X"A6",X"04",X"97",X"24",X"A6",
		X"05",X"16",X"A6",X"06",X"CE",X"FE",X"00",X"BD",X"F5",X"74",X"17",X"DF",X"28",X"7F",X"00",X"30",
		X"BD",X"F5",X"74",X"DF",X"2A",X"39",X"96",X"20",X"97",X"2F",X"DE",X"28",X"DF",X"1A",X"DE",X"1A",
		X"A6",X"00",X"9B",X"30",X"97",X"2E",X"9C",X"2A",X"27",X"26",X"D6",X"21",X"08",X"DF",X"1A",X"CE",
		X"00",X"31",X"96",X"2E",X"4A",X"26",X"FD",X"A6",X"00",X"B7",X"04",X"00",X"08",X"9C",X"2C",X"26",
		X"F1",X"5A",X"27",X"DA",X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"09",X"01",X"01",X"20",X"DF",
		X"96",X"22",X"8D",X"64",X"7A",X"00",X"2F",X"26",X"C1",X"96",X"13",X"9A",X"14",X"26",X"46",X"96",
		X"23",X"27",X"42",X"7A",X"00",X"24",X"27",X"3D",X"9B",X"30",X"97",X"30",X"DE",X"28",X"5F",X"96",
		X"30",X"7D",X"00",X"23",X"2B",X"06",X"AB",X"00",X"25",X"08",X"20",X"0B",X"AB",X"00",X"27",X"02",
		X"25",X"05",X"5D",X"27",X"08",X"20",X"0F",X"5D",X"26",X"03",X"DF",X"28",X"5C",X"08",X"9C",X"2A",
		X"26",X"DD",X"5D",X"26",X"01",X"39",X"DF",X"2A",X"96",X"22",X"27",X"06",X"8D",X"08",X"96",X"27",
		X"8D",X"16",X"7E",X"F3",X"F6",X"39",X"CE",X"00",X"31",X"DF",X"1C",X"DE",X"25",X"E6",X"00",X"08",
		X"BD",X"F3",X"16",X"DE",X"1C",X"DF",X"2C",X"39",X"4D",X"27",X"2B",X"DE",X"25",X"DF",X"1A",X"CE",
		X"00",X"31",X"97",X"1F",X"DF",X"1C",X"DE",X"1A",X"D6",X"1F",X"D7",X"1E",X"E6",X"01",X"54",X"54",
		X"54",X"54",X"08",X"DF",X"1A",X"DE",X"1C",X"A6",X"00",X"10",X"7A",X"00",X"1E",X"26",X"FA",X"A7",
		X"00",X"08",X"9C",X"2C",X"26",X"DE",X"39",X"8E",X"00",X"7F",X"7F",X"00",X"00",X"B6",X"04",X"02",
		X"C6",X"80",X"F7",X"04",X"02",X"7C",X"00",X"15",X"43",X"84",X"7F",X"36",X"84",X"5F",X"81",X"16",
		X"27",X"03",X"7F",X"00",X"13",X"81",X"18",X"27",X"03",X"7F",X"00",X"14",X"32",X"85",X"20",X"27",
		X"18",X"C6",X"7E",X"F1",X"EF",X"FD",X"26",X"05",X"BD",X"EF",X"FD",X"20",X"08",X"F1",X"DF",X"FD",
		X"26",X"07",X"BD",X"DF",X"FD",X"96",X"00",X"20",X"04",X"0E",X"F6",X"04",X"02",X"8D",X"20",X"7D",
		X"00",X"00",X"26",X"DD",X"0E",X"F6",X"04",X"02",X"96",X"10",X"9A",X"11",X"27",X"FE",X"4F",X"97",
		X"13",X"97",X"14",X"96",X"10",X"27",X"05",X"2B",X"03",X"7E",X"F3",X"69",X"7E",X"F3",X"7B",X"84",
		X"1F",X"26",X"01",X"39",X"4A",X"27",X"4C",X"81",X"0A",X"26",X"03",X"7E",X"F3",X"70",X"81",X"18",
		X"26",X"03",X"7E",X"F2",X"79",X"81",X"0F",X"22",X"0B",X"4A",X"BD",X"F3",X"90",X"7E",X"F3",X"F6",
		X"80",X"06",X"20",X"F5",X"81",X"16",X"27",X"F8",X"81",X"17",X"27",X"F4",X"81",X"18",X"22",X"0C",
		X"80",X"10",X"48",X"CE",X"FE",X"AE",X"8D",X"0C",X"EE",X"00",X"6E",X"00",X"80",X"18",X"BD",X"F2",
		X"17",X"7E",X"F2",X"2C",X"DF",X"1A",X"9B",X"1B",X"97",X"1B",X"96",X"1A",X"89",X"00",X"97",X"1A",
		X"DE",X"1A",X"39",X"CE",X"00",X"E0",X"86",X"20",X"8D",X"EA",X"09",X"26",X"FD",X"7F",X"04",X"00",
		X"5A",X"26",X"FD",X"73",X"04",X"00",X"DE",X"1A",X"8C",X"10",X"00",X"26",X"E9",X"39",X"0F",X"8E",
		X"00",X"7F",X"CE",X"FF",X"FF",X"5F",X"E9",X"00",X"09",X"8C",X"F0",X"00",X"26",X"F8",X"E1",X"00",
		X"27",X"01",X"3E",X"7F",X"04",X"02",X"CE",X"2E",X"E0",X"09",X"26",X"FD",X"BD",X"F3",X"2A",X"BD",
		X"F3",X"2A",X"BD",X"F3",X"2A",X"86",X"80",X"B7",X"04",X"02",X"86",X"01",X"BD",X"F3",X"90",X"BD",
		X"F3",X"F6",X"86",X"0B",X"BD",X"F3",X"90",X"BD",X"F3",X"F6",X"01",X"01",X"01",X"86",X"02",X"BD",
		X"F2",X"17",X"BD",X"F2",X"2C",X"F6",X"DF",X"FA",X"C1",X"7E",X"26",X"05",X"BD",X"DF",X"FA",X"20",
		X"AD",X"F6",X"EF",X"FA",X"C1",X"7E",X"26",X"A6",X"BD",X"EF",X"FA",X"20",X"A1",X"40",X"0F",X"00",
		X"99",X"09",X"02",X"00",X"F8",X"FF",X"F0",X"0F",X"02",X"21",X"26",X"02",X"80",X"00",X"FF",X"05",
		X"01",X"01",X"01",X"20",X"01",X"08",X"FF",X"FF",X"FF",X"01",X"01",X"0F",X"02",X"01",X"80",X"00",
		X"FF",X"01",X"20",X"01",X"23",X"00",X"03",X"20",X"00",X"FF",X"0E",X"E7",X"35",X"33",X"79",X"03",
		X"80",X"F2",X"FF",X"36",X"21",X"09",X"06",X"EF",X"03",X"C0",X"00",X"FF",X"20",X"11",X"07",X"07",
		X"04",X"00",X"D0",X"00",X"BB",X"01",X"08",X"00",X"47",X"01",X"01",X"22",X"00",X"DD",X"17",X"0B",
		X"0D",X"44",X"01",X"02",X"03",X"00",X"CC",X"01",X"FC",X"02",X"FC",X"03",X"F8",X"04",X"F8",X"06",
		X"F8",X"08",X"F4",X"0C",X"F4",X"10",X"F4",X"20",X"F2",X"40",X"F1",X"60",X"F1",X"80",X"F1",X"A0",
		X"F1",X"C0",X"F1",X"00",X"00",X"04",X"FF",X"FF",X"00",X"00",X"08",X"7F",X"D9",X"FF",X"D9",X"7F",
		X"24",X"00",X"24",X"08",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"08",X"00",X"40",X"80",
		X"00",X"FF",X"00",X"80",X"40",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",X"F5",X"D9",X"B0",X"7F",X"4E",
		X"24",X"09",X"00",X"09",X"24",X"4E",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"F4",X"00",X"E8",X"00",X"DC",X"00",X"E2",
		X"00",X"DC",X"00",X"E8",X"00",X"F4",X"00",X"00",X"10",X"59",X"7B",X"98",X"AC",X"B3",X"AC",X"98",
		X"7B",X"59",X"37",X"19",X"06",X"00",X"06",X"19",X"37",X"18",X"FF",X"FF",X"FF",X"BF",X"FF",X"FF",
		X"FF",X"7F",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"3F",X"FF",X"FF",
		X"FF",X"BF",X"30",X"83",X"78",X"69",X"5B",X"4E",X"42",X"37",X"2D",X"24",X"1C",X"15",X"0F",X"0A",
		X"06",X"03",X"01",X"00",X"01",X"03",X"06",X"0A",X"0F",X"15",X"1C",X"24",X"2D",X"37",X"42",X"4E",
		X"5B",X"69",X"78",X"88",X"99",X"AB",X"BE",X"D2",X"E7",X"FD",X"E7",X"D2",X"BE",X"AB",X"99",X"95",
		X"90",X"8C",X"88",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",X"F5",X"D9",X"B0",X"7F",X"4E",X"24",X"09",
		X"00",X"09",X"24",X"4E",X"52",X"37",X"00",X"00",X"00",X"10",X"54",X"73",X"26",X"03",X"00",X"00",
		X"10",X"95",X"11",X"41",X"03",X"ED",X"09",X"09",X"4B",X"14",X"0A",X"09",X"00",X"00",X"09",X"6A",
		X"F2",X"24",X"02",X"00",X"00",X"10",X"36",X"26",X"A0",X"00",X"00",X"00",X"16",X"54",X"57",X"31",
		X"00",X"00",X"00",X"20",X"85",X"46",X"41",X"02",X"0E",X"01",X"0E",X"27",X"51",X"36",X"00",X"00",
		X"00",X"0C",X"00",X"33",X"60",X"01",X"01",X"01",X"20",X"36",X"16",X"84",X"03",X"0E",X"01",X"0E",
		X"27",X"11",X"26",X"00",X"F0",X"05",X"08",X"A5",X"51",X"32",X"01",X"00",X"00",X"10",X"00",X"46",
		X"56",X"00",X"00",X"00",X"08",X"6A",X"14",X"27",X"01",X"FE",X"10",X"10",X"54",X"63",X"27",X"06",
		X"00",X"00",X"10",X"95",X"52",X"32",X"04",X"00",X"00",X"20",X"84",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"90",X"91",X"A2",X"3A",X"B4",X"5B",X"C6",X"7C",X"D8",X"9D",X"EA",X"BE",X"FC",X"DF",X"0E",
		X"01",X"01",X"02",X"02",X"04",X"88",X"40",X"08",X"08",X"40",X"88",X"01",X"01",X"02",X"02",X"03",
		X"04",X"05",X"06",X"07",X"08",X"09",X"0A",X"0C",X"08",X"80",X"10",X"78",X"18",X"70",X"20",X"60",
		X"28",X"58",X"30",X"50",X"40",X"48",X"01",X"02",X"02",X"03",X"03",X"03",X"06",X"06",X"06",X"06",
		X"0F",X"1F",X"36",X"55",X"74",X"91",X"A8",X"B9",X"CA",X"DB",X"EC",X"80",X"7C",X"78",X"74",X"70",
		X"74",X"78",X"7C",X"80",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"20",X"28",X"30",
		X"38",X"40",X"48",X"50",X"60",X"70",X"80",X"A0",X"B0",X"C0",X"20",X"10",X"0C",X"0A",X"08",X"07",
		X"06",X"05",X"04",X"01",X"02",X"04",X"08",X"09",X"0A",X"3F",X"4F",X"5F",X"6F",X"7F",X"68",X"58",
		X"48",X"38",X"28",X"18",X"1F",X"2F",X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",
		X"05",X"06",X"08",X"0A",X"0C",X"10",X"14",X"18",X"20",X"30",X"40",X"50",X"40",X"30",X"20",X"10",
		X"0C",X"0A",X"08",X"07",X"06",X"05",X"CC",X"BB",X"60",X"10",X"EE",X"AA",X"50",X"00",X"F0",X"43",
		X"F0",X"57",X"F3",X"69",X"F2",X"7D",X"F2",X"81",X"F2",X"79",X"2C",X"7C",X"12",X"0C",X"74",X"7C",
		X"1D",X"06",X"FC",X"7C",X"29",X"03",X"56",X"F8",X"04",X"0E",X"FF",X"00",X"04",X"01",X"01",X"7C",
		X"0D",X"0C",X"41",X"7C",X"12",X"06",X"74",X"7C",X"1D",X"03",X"79",X"7C",X"3F",X"08",X"F5",X"7C",
		X"30",X"06",X"14",X"7C",X"29",X"05",X"5B",X"18",X"F8",X"04",X"02",X"FF",X"00",X"23",X"06",X"01",
		X"F8",X"04",X"03",X"FF",X"00",X"23",X"02",X"AB",X"F8",X"04",X"07",X"FF",X"7C",X"29",X"15",X"5B",
		X"24",X"7C",X"23",X"10",X"5B",X"7C",X"14",X"08",X"74",X"3E",X"40",X"04",X"FF",X"3E",X"40",X"06",
		X"FF",X"7C",X"30",X"07",X"FF",X"7C",X"1D",X"10",X"F9",X"7C",X"0A",X"0C",X"41",X"3E",X"1E",X"08",
		X"7D",X"3E",X"1E",X"08",X"7D",X"18",X"3E",X"1E",X"06",X"7D",X"3E",X"1E",X"06",X"7D",X"3E",X"33",
		X"05",X"0A",X"3E",X"18",X"07",X"56",X"3E",X"1E",X"0D",X"0A",X"3E",X"33",X"0F",X"7D",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"F5",X"2F",X"7E",X"F5",X"74",X"F3",X"69",X"F4",X"C7",X"F0",X"01",X"F5",X"9E",X"F0",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
