-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "06CC8028B0802A880EA81A806A85AA0540B54085D4507C588BD4507E2C55532D";
    attribute INIT_01 of inst : label is "AAAAAAAAAAAAAAAAAAAAAABCA2AABA89AABA22C22AA2A82AAAAA9B328C8CAA20";
    attribute INIT_02 of inst : label is "70404E080E080E080E0809C101C101C10138203820382026AAAAAAAAAAAAAAAA";
    attribute INIT_03 of inst : label is "1CCE67FFFF00804FE7F820F820B143F8F8F0647C78E61CF639073820820A7040";
    attribute INIT_04 of inst : label is "A0E7207640EC81D903B287640EC81D22C8F23C8F23DDDDF00BBFF802FC78E3C7";
    attribute INIT_05 of inst : label is "8402C2108102BF5F9613F09439BDA99319804073D2239DA039D2239ED105A0E6";
    attribute INIT_06 of inst : label is "202AE00B08BF4680F6CCE383A826EF6B73B006E388B80CECDA97148B29712225";
    attribute INIT_07 of inst : label is "0000800000000CF555554F22212103C8884844433FFFF3F51517F28410FF0140";
    attribute INIT_08 of inst : label is "00E00000E0002488799ED83C0000000002087C078FB000000000020008A05400";
    attribute INIT_09 of inst : label is "295FDFC94FF3BAEBFF6DFFBAEBF9C94FF7F294FFFFF35F00000000012000030C";
    attribute INIT_0A of inst : label is "0010040000000000E2010ED0102CAFEFC2004090FC3FB1B18D000002F8CFFFFF";
    attribute INIT_0B of inst : label is "06003E0006CE00004001E3BFB78000000000087C3F60300000100001E001A100";
    attribute INIT_0C of inst : label is "BFFFFFFBDFFFDD7D77DB77DF5D7FFAF7FFFFF7EFFFFFB6FFF800000000100000";
    attribute INIT_0D of inst : label is "00000240000080064300617C47388BBFEBC0184238000007AFAC6BFFD6FFFD7F";
    attribute INIT_0E of inst : label is "4061801DE0001C0004913F3CFB06000000002F806FB0C0000009000BCEDC0030";
    attribute INIT_0F of inst : label is "FAFE97FD7EAFE773CFDFDB7DFDCF3FCEAFDFF52BFBFDFBEFFFD0000000000480";
    attribute INIT_10 of inst : label is "D2F8008424000000800000000E1C0503A202102A7F0C5084B41406C1F7FFEBF7";
    attribute INIT_11 of inst : label is "00000201019EC06F80000E00000107B3DFEE00000000024800CEFC3008000003";
    attribute INIT_12 of inst : label is "017FA67FEFFF7E7FFFE319FDFD55DFB5DF557F7F319FFFF9F9FFE7FE6BFD0000";
    attribute INIT_13 of inst : label is "00E80E33855FBF00388E2B1A0A069E4F4BA7A793D2C9E9F4F4B27A7D30000000";
    attribute INIT_14 of inst : label is "4D00292FC85D566502A9EC559365A884DDF5CA6736630A04C46CDA598C2819C1";
    attribute INIT_15 of inst : label is "B725E074D743369426F324A28539EE6BFF5232A54AE00D4FF39393500A4BF210";
    attribute INIT_16 of inst : label is "248AE99291E8E1C948F470F6A47A3872125D0C3113272FBDBE000F6010199398";
    attribute INIT_17 of inst : label is "53A7DBCA6035353535353525301A9A9A9A9A9A9F6E7B4DFF6FFFFFCFFFFF9FFC";
    attribute INIT_18 of inst : label is "FFFFAAAAFFEA74846A7494E929D253A4A7494E9A9D211A9D253A4A7494E929D2";
    attribute INIT_19 of inst : label is "FD145B8300000000871C00030002628C10A0029401DDDDDDFEAAABFFFEAA88AA";
    attribute INIT_1A of inst : label is "927D3A74000008000000048040618018700003800012401E1DDF800000000008";
    attribute INIT_1B of inst : label is "0820000000000001D74FA48A7FFFFFE633EE74E9FDF7FF7DD3A7DC633FFFFFF2";
    attribute INIT_1C of inst : label is "FF0000E000000040003FFD84800000FFD00001FB60000001F6C0000000000000";
    attribute INIT_1D of inst : label is "FDFD75DFDDEFFFE3FFF77BDFDD7F4FFFCAFFFA28ADBFF00000000000801B0C06";
    attribute INIT_1E of inst : label is "01F61B0003FE000018000F8000000000000000000100000006DFF8A2BFFE94FF";
    attribute INIT_1F of inst : label is "F3CBB7F59595BEFFFD0000000000400000600001B000E0000EF00001F6E00400";
    attribute INIT_20 of inst : label is "03F3F000000200000200001F7FFE9595BFACBB3DFFFEF7BF7BFF1FFBDFBDEFFF";
    attribute INIT_21 of inst : label is "041000301807C000070000001ECF7FB8000000000920033BF0C02000000F4BE0";
    attribute INIT_22 of inst : label is "99FFBFFDF9FFFF8C67F7F5577ED77D55FDFCC67FFFE7E7FF9FF9AFF400000080";
    attribute INIT_23 of inst : label is "2BA302C714D55464CAA8C9932AA3264EAA8C993AAA3264EFF7630000000005FE";
    attribute INIT_24 of inst : label is "491DD970F0B191316E0A0AAA32635464C58D5193167B9CB738EEE4923BB661E3";
    attribute INIT_25 of inst : label is "E72DCE3BB9248EED9879CEE8D0B5C535551932AA3264EAA8C993BFCC539C777B";
    attribute INIT_26 of inst : label is "4D7C20444194F3E71DDED247765C3C2C6444598282AA8C98D51931635464C59E";
    attribute INIT_27 of inst : label is "13FE046A5E0AE23480820335ED34711555555555565555D1726E4295559F0CC8";
    attribute INIT_28 of inst : label is "B6C82DB40A88B3152DBDA24742054678A23542338ACAB5446EEA054000001B9D";
    attribute INIT_29 of inst : label is "D8C1B04878C412322AAA288A2A22A28A2281551155511041415166E2D9144280";
    attribute INIT_2A of inst : label is "9554010AA4154555709489446EB0CEB44F47FFE44EE52803702E9AC04624EAC2";
    attribute INIT_2B of inst : label is "FFFA2012F4244141110181111110411B8AF0BC2ACA91BBBDB5FBD250A92AAB25";
    attribute INIT_2C of inst : label is "77DA54D1DDB5A913EABAAAB2AAA33FF82F7BFFF82F7BFFF87FF088C8A80A27A7";
    attribute INIT_2D of inst : label is "903505DF19A050281FFE7D03BB6B5377DA54D1DDB5A9A050281FFE7D03BB6B53";
    attribute INIT_2E of inst : label is "15C81FEEEEAEEFE6E23CFCCFD8DDD9DDE0061FCE383338E0990BBE33CFCF544E";
    attribute INIT_2F of inst : label is "0080FFFFFC3C03FC3C006E3F9F9800B0A5FC742EF7FF42EF8C807CDDDFC64E64";
    attribute INIT_30 of inst : label is "0D248361A70C249308201CF1E411C8238073C79047208E33407FFFFE1E01FE1E";
    attribute INIT_31 of inst : label is "CD44488166925D15555EC94921FFDFFF66C993264C993274E9933E12611A41A3";
    attribute INIT_32 of inst : label is "73248D26588B8445C8988B844638189485DDCB473FAECBFAECBFAECBFAECBFAE";
    attribute INIT_33 of inst : label is "FFB0473FADC3F3C9C23FCF23E2D6D3AA79B17D658444410242FF086186104043";
    attribute INIT_34 of inst : label is "C81D27920D527920DDD5355555557FD9CE7D45FDF11F9EE79FE398E3FE7CBFFB";
    attribute INIT_35 of inst : label is "7A5DE93E190975C0A1C0F1C2E1D5F1C341C0A1C00EC877C3D61727AE4F5DD11C";
    attribute INIT_36 of inst : label is "D555555AAEAAAAAAD5769DA56BBA6E99B6739F5169E7A5DE9E7A5DE9E7A5DE9E";
    attribute INIT_37 of inst : label is "557DBFF7DAABED5E4EA47AFEB654ECFE1F4927523D7F2A7637FB1650B2E59FBF";
    attribute INIT_38 of inst : label is "C0A1C00EC877C3D61727AE4F5DD11CC81D27920D527920DDD53FFDF554CF6F62";
    attribute INIT_39 of inst : label is "09C09E9013C82A06B8480CDAEF621D553D88A6B33EC5C0A1C0F1C2E1D5F1C341";
    attribute INIT_3A of inst : label is "1F411F401E9A1E911CBECA2376CE510DDF1A6CDC71C686F21E4BAA5CD6E04F48";
    attribute INIT_3B of inst : label is "E938AE90A65F61D4F1F1C3A707C62E155FFF1EAF9F411F401F411F401F411F40";
    attribute INIT_3C of inst : label is "51F0E9C54D5A5562AD27D6D249DFFFB95476780A7CBE5A011F350BB81117702A";
    attribute INIT_3D of inst : label is "4D728A8AC00022D5259D80002F35996A01C9494A4F200000000001D40B4B922B";
    attribute INIT_3E of inst : label is "9701764DBAE8AC000000000000000000000658096D527AB500000000BCDC4001";
    attribute INIT_3F of inst : label is "EF91800000000000176049DAC6A96B4014E747D23DC002ACCA9AE500093522A7";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "CEEBAB97BEEE11F8F2F4EBD3AF4ABF3DF957A5075D74CEF58E9D74C77AF75B66";
    attribute INIT_01 of inst : label is "555555555555555555555557F4C235D7C235F57F55F5555555556BAEEBAC47E3";
    attribute INIT_02 of inst : label is "F0C2C6185C105C105C1058C30BC30BC30B104170417041635555555555555555";
    attribute INIT_03 of inst : label is "1C0F9FCFE7FFFFFCFE7041B041E1D0846B1A02358D00B0AC3A0D1041041E30C2";
    attribute INIT_04 of inst : label is "C3A2D82DB05B60B6C16D86DB05B60B43D0B42D8B42F5F5F00BFC0F03FFC00200";
    attribute INIT_05 of inst : label is "1AFB0D6B5F647D85BEF9FD07066C976E526C9F77E4DBBE4DBBE4FBBF3A1FC3A3";
    attribute INIT_06 of inst : label is "39C5993E3E632BCE1E343F5E1CEDEFC0D5E72B2E407438D837CC739B81DDF396";
    attribute INIT_07 of inst : label is "180C4FE0C0678CF0000000000101028888C8C0033FFFF602222816C9990A75D9";
    attribute INIT_08 of inst : label is "0BB73DF7EF3F0994CFC3FCE4C6C36EE434D4C6DCE0FC87FC70DC84E63FFFFFE2";
    attribute INIT_09 of inst : label is "6B404019C8803AEA212510BAE84019C81006B500001722C861C60DCA50B72FBF";
    attribute INIT_0A of inst : label is "1B870139EE0F7FB901B7D823987FC6761786639C5054B1B18200000115D00001";
    attribute INIT_0B of inst : label is "CF508372FFFEC3F29B9738E0FC9F3CE1DC84D4C6E1FEFC87E3A6E5373B9FFFF7";
    attribute INIT_0C of inst : label is "FF02007DEE201D61084908585D44037B02007FFE3801FF910419C38DC7871C2D";
    attribute INIT_0D of inst : label is "737384E7F7FFDFC008C5F7C801097FCE709B848429F0A3FF272410881FC00FF1";
    attribute INIT_0E of inst : label is "A5F7E17727BEFDE7213281E78FDF80E30DB940DCF8FFF0DCB0D272D063F79FFC";
    attribute INIT_0F of inst : label is "3382D001C3A10073CC40094401CF2201B84005AE0B19F000012821871B872942";
    attribute INIT_10 of inst : label is "660E63FEFF0E20B84FE05C7F8C827F468010849FA3FE129414140110000093E6";
    attribute INIT_11 of inst : label is "71C370A073C3F0F8F2E37EB8729290F8723B90DC723394D1CFE386FDC39D3EE6";
    attribute INIT_12 of inst : label is "00884E8221706E440107390001DC21FC2177400073910041B82E0822E44280DC";
    attribute INIT_13 of inst : label is "FB004621DE05D01E11C4282A0A09C368E134729A394D1C368E1B4729A0000000";
    attribute INIT_14 of inst : label is "8F88FC804CBE6784B573A8AF8FEA7B3E02DBD58000A43ECA51F4680290FB30B7";
    attribute INIT_15 of inst : label is "097E0126B829A5CB5B265F56FB0C1FC001CD4FFFFFED6F8010D0C3E23F201336";
    attribute INIT_16 of inst : label is "47BFEE6F2D329837B28B44094B0CE604EC82E10BEBFCD00240A290FB9ECCC7BC";
    attribute INIT_17 of inst : label is "EC487D14991A4A4A4A4A4A5A5D8D2D2D2D2D2D23E0BEEA00C00001A000024005";
    attribute INIT_18 of inst : label is "AAAAFFFFFFBD89763D897B12F625EC4BD897B12F624D8F624EC49D893B127624";
    attribute INIT_19 of inst : label is "47FFFEF7CF0C2CF53FFF67BFFF78BFFB6B60C1EC01F5F5F5FFFFFEAAAAAA82AA";
    attribute INIT_1A of inst : label is "9A453A02000D03F9E39731381EF7DC3DDEBEFFAF9EA68F437668CF437660CF7E";
    attribute INIT_1B of inst : label is "D353FB7FDBE000000748A69A4000000E722074E8210D8841D3A440E720000006";
    attribute INIT_1C of inst : label is "812DB7EB812DB4A7BEE087E13801B9907730070FF720DB731FE0DB731B70DBF0";
    attribute INIT_1D of inst : label is "042175C01DE8100008077BC01D0840004E000EFBE240480030E380E1413FBF0F";
    attribute INIT_1E of inst : label is "531EFFCC6E2B6E187CDB98D86CDB98DC6EFF84A7F7FBFFC0012023EF80039C00";
    attribute INIT_1F of inst : label is "06DC301DBDBD800202801B6E30E21B7094FFDC27FCAFEDB723B6E6771FBFE637";
    attribute INIT_20 of inst : label is "8E1E1C3803053F8181FE000001013DBD80EDC36C000031A378400203D18C6000";
    attribute INIT_21 of inst : label is "E1A96E7B7E5C797FBF7C394E43E1C0EE4371C8CE53473F8E1BF70E60FB99D039";
    attribute INIT_22 of inst : label is "3A0885C1B910041CE400077087F085DD0001CE440106E0B8208B910A006C3906";
    attribute INIT_23 of inst : label is "2EE8B72FB9B803991A073236E81CC8FBA073236E81CC8F9C0C4A400000000221";
    attribute INIT_24 of inst : label is "B2600437C49734CBB2DD9D01CC8B0399172C0E644DE4D248C300092DC4486F99";
    attribute INIT_25 of inst : label is "359630C006CB71133BE6D99A65C92E5E00E64581CC8B96073226F22B2CE38884";
    attribute INIT_26 of inst : label is "4C16BD37BD7B0738E2236C98019DF1EEDD1EEFD77F40732340E646DD03991F38";
    attribute INIT_27 of inst : label is "4D54888028B1479A5AC897DAB75DA3C0000000000000008E22990FC0009C4B19";
    attribute INIT_28 of inst : label is "E2683BF5A88CF319B5D52A52415DCD320A80C17D2094240F3451400A952ABEE8";
    attribute INIT_29 of inst : label is "00043048F0C403922AAA2A0A2AA2E28820C155114455104141116FACCD1C2C58";
    attribute INIT_2A of inst : label is "80002940EA0000001080880F2EB08CF44B4D55544AA50803D03AB00B862648F0";
    attribute INIT_2B of inst : label is "AAAA2219F6E46C6C0004A10B0000009EABF428004E94AAB8FC515252B93BBC20";
    attribute INIT_2C of inst : label is "0821010A824202B6C0D003D40013D2948AA522948AA52294B1295E48C16225A6";
    attribute INIT_2D of inst : label is "7FFBAA8C149E8F47A49290B50484040821010A8242021E8F47A49290B5048404";
    attribute INIT_2E of inst : label is "A6A54BAAAAAAAB2FA2905000228190008A4E48064D001934005518290500ABF8";
    attribute INIT_2F of inst : label is "FE01FFFC003FFC003FFE7A920A03FF02004A21545EA215460A007A95572DF4CA";
    attribute INIT_30 of inst : label is "BAE9A6F77B9AEBA79EEA238EE14C8299288E3B85320A652900FFFE001FFE001F";
    attribute INIT_31 of inst : label is "282E9D29204649AEEEE4999A930000038F1E3C69D3E3C68D1E7CC774F67CD7C7";
    attribute INIT_32 of inst : label is "F4EDD664C5CAEAE57925CAFAE7AB25C0AF99B4CCF4BD2F03C0F4BD2F03C0F4BD";
    attribute INIT_33 of inst : label is "E372B4A96B1407E317889FFC300364FCFC640090C9899227A5FEFAAEAAE48F66";
    attribute INIT_34 of inst : label is "F0D529862952986294032ABEFFEEC5E718DE3E397721794ED01E63BA064CA072";
    attribute INIT_35 of inst : label is "472D1CA2C65925400D4009C13D5049C09D4049C06EA6743A8835626AC4D6C8D4";
    attribute INIT_36 of inst : label is "26666663333333331995B56FF6B75A1579C6378F9C347091CA472D1C347091CA";
    attribute INIT_37 of inst : label is "6254C0001B12A6441B10D4A89A061E5BBF000D886A54030F1AB1800400600000";
    attribute INIT_38 of inst : label is "4049C06EA6743A8835626AC4D6C8D4F0D52986295298629403200006244295B1";
    attribute INIT_39 of inst : label is "0940A63012F02101F222082B15B8803614E24B0A4B79400D4009C13D5049C09D";
    attribute INIT_3A of inst : label is "D6E1D6E1D5D7D508D46C5D6254A8EB09660244940A8B04BCD78AA1D43EA05318";
    attribute INIT_3B of inst : label is "E3406F8924961D6C1D7209682701AE035400962496E0D6E0D6E1D6E1D6E0D6E0";
    attribute INIT_3C of inst : label is "2260C0823C6812106B4119604E80003830B272067C627C03A62F8BC036178166";
    attribute INIT_3D of inst : label is "962444404000056901998001E4753A36014010940D40000000000760020CE05C";
    attribute INIT_3E of inst : label is "4001C0060260280000000000000000000000A8003424D04200000000A6020000";
    attribute INIT_3F of inst : label is "30820000000000005C000168CE10A20004C18D9940400495C12C4880002CC495";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "26726AFF0A6B7ACEC24E2938A462918C8C52311597FF8AF1AB17FE8D78D7FB7E";
    attribute INIT_01 of inst : label is "00000000000000000000000A039D60081D688228200200200A0009C92631EB3B";
    attribute INIT_02 of inst : label is "3041060826082608260820800480048004100090009000820000000000000000";
    attribute INIT_03 of inst : label is "F3399FFFFF3399C020182018201000DC0CBA02065D62B8060500100000003041";
    attribute INIT_04 of inst : label is "805248C49189231246248C491892310048521405017F55FF0ABF8FE3FFFFFFFF";
    attribute INIT_05 of inst : label is "1CE98E739C313C908F2D5CC7C89EC9939CCF264F713277132371323B98428053";
    attribute INIT_06 of inst : label is "8E59FE35359ACA6072EAC6E44E536EE583C82CBDB4B6BFAA4D59AD6B89F9CBD3";
    attribute INIT_07 of inst : label is "E7F3B00F3F982CF0000000000101028888C8C0033FFFF8133335F460CCE9788C";
    attribute INIT_08 of inst : label is "F62CCB2D12A4FF5B04B24A8305B2D8836FB305B05893449040B3479820804499";
    attribute INIT_09 of inst : label is "C6202037B80C4D342092104D340637B8080C6300000C8016593D8B37EE7CD964";
    attribute INIT_0A of inst : label is "167CFF6609F04024E2010EC014ACAFEFE23BDC64505444440500000003300000";
    attribute INIT_0B of inst : label is "32CF62CD9251024DF66C168090641080B06FBB0581259364817D9BEC1664812C";
    attribute INIT_0C of inst : label is "D1000016B4102080803F8020208205AD00001A34100061800420A27B027C139F";
    attribute INIT_0D of inst : label is "42C26FD80400B0166300617CC3388BBFEBC07FFFD950215088882C00018003A0";
    attribute INIT_0E of inst : label is "9B2C9EC41965A2541FEB608209126082CBE7F8B3209240B36CBECDBE5A426490";
    attribute INIT_0F of inst : label is "0D01480040D0188E38203F820238E030C820029404060C1000005964F604DFB9";
    attribute INIT_10 of inst : label is "2F89820584099F67300FB3802E140101F202100A7F05DEF7822222C008000418";
    attribute INIT_11 of inst : label is "4F02CF9CCCB24F204D82D1604DB66C9641226CB0412A6FBD325A05913E10A5D8";
    attribute INIT_12 of inst : label is "00081F8230C09980001DEE02026600DA00998080DEE0000666181823F04004B0";
    attribute INIT_13 of inst : label is "20C9C2020D1FBF04E67BC1155559627CB13E5A9F2D4F96B7CB5BE58DF0000000";
    attribute INIT_14 of inst : label is "A20D94D716000005C753B2783207863564E1A5A11B09326401858C2C24C998C1";
    attribute INIT_15 of inst : label is "5C19E1FFF52F6F9E7567B896C4B017E59F1941428529D2976B0B08836535C580";
    attribute INIT_16 of inst : label is "50156ED1D169B268C8B659346613689A3B09344BFF288882ECA2835FAD511512";
    attribute INIT_17 of inst : label is "B76DF9B6D3AB6B6B6B6B6B6B78DDBDBDBDBDBDB7429E7805E7FC0BFFF816FFF4";
    attribute INIT_18 of inst : label is "AAAAAAAAAA96EDA356EDADDB5BB6B76D6EDADDB5BB68DDBB6B76D6EDADDB5BB6";
    attribute INIT_19 of inst : label is "8410488904F3DB8BE082DC493447C20896AF3E9500AAAAAA0000000000002AAA";
    attribute INIT_1A of inst : label is "6D82C580004B0A209E0C0FE7792CB3CB11659459717DF8B2C444B8B244408891";
    attribute INIT_1B of inst : label is "B6EC02C01608000008B05B6D8000001BDC118B16020D80822C5823BDC000000B";
    attribute INIT_1C of inst : label is "00DB6D1600DB6D996580449FE00166083CC004092CF0B6CC1250B6CC16C0B64D";
    attribute INIT_1D of inst : label is "020082202210100408088420208030003D000DF7D04040082C9E009BBEC964F2";
    attribute INIT_1E of inst : label is "4C1269305832D9B44AB660B45AB660B058926DD804020010002027DF40037B00";
    attribute INIT_1F of inst : label is "0D34480A6A6A4100000096D9EA81F6CF5324B3D49365116CDA3D98441224982C";
    attribute INIT_20 of inst : label is "080810268284C0014200800080006A6A405344D200818C408400800420631004";
    attribute INIT_21 of inst : label is "9F76F996C9B026C9689026D9B2590089B2C104A9BEF4C9681644F8589760F626";
    attribute INIT_22 of inst : label is "7E08C30266000077B80809980368026602037B8000199860608FC100025B26C5";
    attribute INIT_23 of inst : label is "738AEF997C5EC67441C8CCCB8633A22E1C8CCC38633A20CF2573000000000020";
    attribute INIT_24 of inst : label is "69BECF23FA398577CDBE6F723336C674499B9199B6791C6279E766DA79DE47E4";
    attribute INIT_25 of inst : label is "6718DF7D99A4DF6691FD9CC2BBF6DFA7319D13723334CD8CE89B3CCE313CF3B3";
    attribute INIT_26 of inst : label is "EC171E3BDEE7476FBECCD34F3B48FCCE6179FA6FD39C8CCDB19D1266E46669DF";
    attribute INIT_27 of inst : label is "E401CCF1A1FD081AC808881F0000C40555555555565555FD005DEE9555FD7D5D";
    attribute INIT_28 of inst : label is "E172F90A282FCE5FCC33D7AFA0A5D03AA8A1C2810063C5D03114D00A952A40E2";
    attribute INIT_29 of inst : label is "84DB7DB937DB08188028A228A2A888AA89F4015451505554541558312E42AD22";
    attribute INIT_2A of inst : label is "E0023A8E01C1E8000D415410350B114FF2F6EEEFF32EDF881F71741FBEDDF5C7";
    attribute INIT_2B of inst : label is "7777FCE4F83F8383EEFA4EE4EEE51440DBFFEB407F6BAAA01D8F6DBDBABBBF57";
    attribute INIT_2C of inst : label is "46F64C5079EC98C8C02000280018110CA1CE450CA1CE450CCE19E07FDE1FF97B";
    attribute INIT_2D of inst : label is "F57A8C2340A010080B6D4D00F3D93146F64C5079EC98A010080B6D4D00F3D931";
    attribute INIT_2E of inst : label is "B86C3FAAAAAAA8D828148CC00BD5B8D50A340D801D0000740818468148CCFEDA";
    attribute INIT_2F of inst : label is "008100000000000000030284919CA5AAA5124461211C4611A0006A555D489974";
    attribute INIT_30 of inst : label is "4D24DBC9636D24D269201176042248448045D810892113C14080000000000000";
    attribute INIT_31 of inst : label is "6B365CFB6266C9505050CFC8A5029FF336EC9B336E8D3A24CC9B2692489A491B";
    attribute INIT_32 of inst : label is "F5A4ED2E26DB8B6DC9B6DB8B6E39B6F1B751424629AA6A9AA6AD2B4AD2B4A9AA";
    attribute INIT_33 of inst : label is "B89F5195CEF9C77844861DC5415C7F14E5B0B9E70DDCF907CED4E0C71C3E4E32";
    attribute INIT_34 of inst : label is "4C153B1B2553B1B2540D5AABEFBEBFFDEE7C48295DF9CE731635AD4AC5DBAC52";
    attribute INIT_35 of inst : label is "65899632E7DB2540014051C165DBD540B14151C02E0073CBA505808B01168514";
    attribute INIT_36 of inst : label is "C7878783C63C3C3C1E3F1FC54C19E5FBFF7B9F12162658996A65AD96B65AD963";
    attribute INIT_37 of inst : label is "6948F0500B4A471E59E6C294D0AE4C2B81400CF3614A57261053C91600E00F3F";
    attribute INIT_38 of inst : label is "4151C02E0073CBA505808B011685144C153B1B2553B1B2540D5C14069568A2B4";
    attribute INIT_39 of inst : label is "0140ECD802CC300AC60A0092F2B280D64ACA5E05C46D40014051C165DBD540B1";
    attribute INIT_3A of inst : label is "1DC01DC017CE17451CE38D21702269056838B854699500B31662B01558A0766C";
    attribute INIT_3B of inst : label is "E7242FF24254A15CD1F927E497268E2C1FFF57815DC11DC01DC11DC11DC11DC1";
    attribute INIT_3C of inst : label is "02802C234848D8A1ABCF55E7787FFFBAC0A07811743D7E01A91C8B2490164822";
    attribute INIT_3D of inst : label is "BC0A93D4000056E14A9B00034166734E001CA8CF68600000000003380565D10B";
    attribute INIT_3E of inst : label is "8E004320B32DA400000000000000000000018804D0BCC653000000000E4AE000";
    attribute INIT_3F of inst : label is "103D80000000000044302CA46C5845602EC80C722A8003279978150005A636C9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "67762BBF4A6E7D51DF4E3D38F4E3D18E8C7A31E52AC26854426AC26C2A5D5039";
    attribute INIT_01 of inst : label is "000000000000000000000002A88208A00208A82A80A8028000001DD86325F543";
    attribute INIT_02 of inst : label is "A000840014001400140010800280028002100050005000420000000000000000";
    attribute INIT_03 of inst : label is "10080733993F9FCFE7F00050000001CCC7782263BC2290441002182082002000";
    attribute INIT_04 of inst : label is "A002000400080010002004400080012040501405015555DFFAA00803E0400200";
    attribute INIT_05 of inst : label is "12F5894A5F3700DF4D7DEB4549BA52A54BAFF2279F9179F9139F913CF102A002";
    attribute INIT_06 of inst : label is "86193F1191B2CB6A1A72F0E2CE524069032AA5D249100008C9152D600966D1CB";
    attribute INIT_07 of inst : label is "EFF7600F7FB02CF0000000000101028888C8C0033FFFF8911115A468AD5F34AD";
    attribute INIT_08 of inst : label is "F2C5D1451429C997750C90BF788C4B3FA49F7897472705279F1704BBC820113F";
    attribute INIT_09 of inst : label is "000020042008082020481008200404200800000000000011867C71725E25CA29";
    attribute INIT_0A of inst : label is "E2E5F9AC1BE0806D8197D8730C5EC43617BEA1C8AC6B44448D00000000000000";
    attribute INIT_0B of inst : label is "747F1C5CA4917C9C92E5D13F27E9D73E97F69778BE48A7193D24B9A5D2E92045";
    attribute INIT_0C of inst : label is "000000021010000000000000000200840000000000000810002E82F97AE5E789";
    attribute INIT_0D of inst : label is "9C5CF6B0080000140841F7C8E3309FCA308B586698A022A22224688028000000";
    attribute INIT_0E of inst : label is "F9453E59FA28A285F932DEBAF264DF3C312F47174F249F1723135C91849AE927";
    attribute INIT_0F of inst : label is "20800000C18010082020000200208021980000020010200000004619F2F9C978";
    attribute INIT_10 of inst : label is "B473BC80A1F3FF2FE00F970028025FE68040003F81FF1212088886C000000040";
    attribute INIT_11 of inst : label is "9F7C5CFD5D0C9F4F5CBC512F9CDBE3219CCCE3179CC2E4D17484F8A672E648BB";
    attribute INIT_12 of inst : label is "0008040000000000000108020000000000000080108000000000000040400317";
    attribute INIT_13 of inst : label is "F3810A507E0CC11E89598B14444DEB5AF5AD78D6BC6B5E25AF12D78960000000";
    attribute INIT_14 of inst : label is "E24AC585168000032A99016A1D3BE37A50B9BB231214746829ADA60851D1B0B5";
    attribute INIT_15 of inst : label is "141BFE5046F2126205829A95561F046903BF424489496CC509E35882B16145A8";
    attribute INIT_16 of inst : label is "78C53FD99949A2ECCCA65176641368BB3A09B41403E22231822A10CD7BF54A24";
    attribute INIT_17 of inst : label is "162FCFCBC42965E165E165F16316F0B2F0B2F0BCBA325B0565420B7A8415D50C";
    attribute INIT_18 of inst : label is "00000000004BD78852C597AF0B165EBC2C597AF8B17316F5F162EBD7C58BAF5F";
    attribute INIT_19 of inst : label is "7904132A75F7C9A928204D525994A08610AF7A95000000000000000000000000";
    attribute INIT_1A of inst : label is "04020408003104AEBEE1E92F154517D16528A44A35269A8C59931A8C999F32AD";
    attribute INIT_1B of inst : label is "9A58060030080000208041040000000210100810020200802040202100000001";
    attribute INIT_1C of inst : label is "FFC92512FFC926FA28BF39392FFE2EE7B5DFF9F245E0925DE480925DE25F129E";
    attribute INIT_1D of inst : label is "00000020031810000800C620000010001000000000000007C33EFF3D7FD229F4";
    attribute INIT_1E of inst : label is "BDE592778BCC4BD05092EF104892EF178B24F6F00D0400100000000000002100";
    attribute INIT_1F of inst : label is "01000000000000000000624BE13D925F1F4917C527391625C4D4BB99E4C93FC5";
    attribute INIT_20 of inst : label is "F3EBE7CF02078041000080000000000000000010008000000000A00000000004";
    attribute INIT_21 of inst : label is "B92A4BA25297AE5228A7CE6B8C867F338C5E730B9345D213E299CB8722EE99CE";
    attribute INIT_22 of inst : label is "100000000000000420080000000000000200420000000000000101000188CA38";
    attribute INIT_23 of inst : label is "6576A4A9A52C64EEF089D9AD4237E6B50CDFDE54237E697BAD3D400000000020";
    attribute INIT_24 of inst : label is "CBBECD6FFD36FB425052B622766864EEF2E19BFBCBDD4E6E59E6779F7DDEDFF8";
    attribute INIT_25 of inst : label is "539B9679DDF5DF67B7FE997DA92A694B91BF3522766B74C9DDEDEEA7372CF33B";
    attribute INIT_26 of inst : label is "A82829021897E2CB3CEEFACF335BFD0DBED09414ADCCDFDE11BF34B844ECD2F7";
    attribute INIT_27 of inst : label is "037C00001C00E41137E0041037DF020AAAAAAAAAABAAAA3FAEE2EFEAAA2AE3A2";
    attribute INIT_28 of inst : label is "178000F002801941E18E05000080083400402841603C0A082C60000000002098";
    attribute INIT_29 of inst : label is "70000C01000004122A8228822A02420AA00154050400040505440020701EC300";
    attribute INIT_2A of inst : label is "1DDD83B0E11C0777781DC1C82AB00C111D1111011DC3C184100882C000000000";
    attribute INIT_2B of inst : label is "888888E4080982821109913111B05120C00E177B81C0111FE070870C03800070";
    attribute INIT_2C of inst : label is "3805898E020B1320D54555015544100310000003100000030006106234108E8C";
    attribute INIT_2D of inst : label is "E57AF220209F8FC7E00082BC0416263805898E020B131F8FC7E00082BC041626";
    attribute INIT_2E of inst : label is "4013FFBBBBFBB800201303FFD8C518A608627C8C3C1030F008E44041303EFE9E";
    attribute INIT_2F of inst : label is "FE7E000003C3FC03C3FC8300607F5A4D5A018B910000B91010006C377571007F";
    attribute INIT_30 of inst : label is "EB2EB8DCEE79E59E79EFE2080BEE17DC3F88202FB85F70013F000001E1FE01E1";
    attribute INIT_31 of inst : label is "4D224CDB43064944114551D88182B50B377C9D7275CDDF3778955CF3CFD75D7A";
    attribute INIT_32 of inst : label is "E7A4CF2F0C598E2CCDBC599E2E1BBC51E3DCCA4AA9AA6A9AA6ADAB6ADAB6AD2B";
    attribute INIT_33 of inst : label is "05C2F994C64972887D16CA58E0EFD7A651DD22F3FEEEFBD68D2A73CB2CBEEF35";
    attribute INIT_34 of inst : label is "C0142B0A0142B0A0158350000001554B5ADD5B050620A5A95125394A21B3220A";
    attribute INIT_35 of inst : label is "57895E2CC9D925C085C0D541E1563141214081C02EEC740A851587AF0F5F8214";
    attribute INIT_36 of inst : label is "3807F80C03C03FC0601E378FC819E5BB92D6B756CEB57AD5E357895E257895E2";
    attribute INIT_37 of inst : label is "505CD05C1A82E6165D00E0B880CC447318C00E80705C662200E3801400A000D4";
    attribute INIT_38 of inst : label is "4081C02EEC740A851587AF0F5F8214C0142B0A0142B0A015835417050465C7B0";
    attribute INIT_39 of inst : label is "05C0AC500BC0280AD818004257B618335ED868106F7DC085C0D541E156314121";
    attribute INIT_3A of inst : label is "14C014C015C61CC21471082151424105EC00101C28C182B0160AA8555AA05628";
    attribute INIT_3B of inst : label is "AF142B80085F01444160A56297A02E1057FF574F14C014C114C014C014C014C0";
    attribute INIT_3C of inst : label is "02C0202209C893806F48D3347800003900E178007CB47E012C0C091410122822";
    attribute INIT_3D of inst : label is "D018101200008420089500034F6432060090408408400000000007A00005810D";
    attribute INIT_3E of inst : label is "0000052082A132000000000000000000000280049046E4D200000000583C8000";
    attribute INIT_3F of inst : label is "945E000000000000405020246C10000024EA0E101200010091A0300004350482";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "5AFABEBEFBBA3E199235A8D6A35A8D6C6B51AD224AA3D084448AA2D0427FFA00";
    attribute INIT_01 of inst : label is "000000000000000000000000A2882008082088088008008008000BEAFEE8F866";
    attribute INIT_02 of inst : label is "669E6CF3CC51CCF3CCD3C98A399E799A79B14733CF334F260000000000000000";
    attribute INIT_03 of inst : label is "1FFFFCCE67CCE67FFFF3CF73CF227A49887A24C43D22116D4A6BB14734F2628E";
    attribute INIT_04 of inst : label is "CF76D96DB2DB65B6CB6D12DB2DB65BC4F17C5F17C5D55550FFFFFFFFE0400200";
    attribute INIT_05 of inst : label is "30901842132C40DA0A05598185681468C20C8E0D04703047070470683A7BCF77";
    attribute INIT_06 of inst : label is "89255953536C2C587F0DA2C21CC5604445B1A3092482AA223500E3184F42B900";
    attribute INIT_07 of inst : label is "EFF77FFF7FBFECF0000000000101028888C8C0033FFFFD53333194588B62AC8B";
    attribute INIT_08 of inst : label is "F205C104E021C9170C1000870090480724970090C8070400001706B8071F883B";
    attribute INIT_09 of inst : label is "108000000000000000480000000000000001080000020212087881725F25C821";
    attribute INIT_0A of inst : label is "02E5F92FFBFFFFECE2010ED2908C2FEFE2090CB4501444448D00000010800000";
    attribute INIT_0B of inst : label is "705F205C800E001C93E4320000E0300190E49700800087200324B92432E01E04";
    attribute INIT_0C of inst : label is "000000000000020208120800820000000000000000000000002182F106E407C9";
    attribute INIT_0D of inst : label is "0040E4BFFFFF1FF62300617C2021039FE7C033352150215222246C0000000000";
    attribute INIT_0E of inst : label is "B9043E4038209C043922E1860000E000412E48170000001724125C920806E000";
    attribute INIT_0F of inst : label is "00002002000000000000120000000000000008400000000000004821E201C97C";
    attribute INIT_10 of inst : label is "648380789803BF2F7FFF97FFEE140301D031086E7F14FFFDE888869000000000";
    attribute INIT_11 of inst : label is "1E005CBE5C101F00DC804E201C92E4020300E4100302E49170080080720180B8";
    attribute INIT_12 of inst : label is "0000000000000000000000000088204820220000000000000000000000000410";
    attribute INIT_13 of inst : label is "20D98E7389BFBF8C7EAC6B1444432935949ACA4D6526B2935949ACA4D0000000";
    attribute INIT_14 of inst : label is "8309C07265800002750033A7C20AC54930EA50A11998AC5920BF002662B17CC0";
    attribute INIT_15 of inst : label is "4857FFDB6FFECB37F141F61C11429644C4A5DD5AB52972925E9C80E2601C997A";
    attribute INIT_16 of inst : label is "4B750E25092406128490830942080084A904000AA8E88882402F50598E623D00";
    attribute INIT_17 of inst : label is "9325561255292DADA9292DADAA949496D6D494961A00D2A501554BA2AA966551";
    attribute INIT_18 of inst : label is "00000000001264AA5264B6ED6DDA9325264B6ED6DDAA949929325B76B6ED4992";
    attribute INIT_19 of inst : label is "00E380280DF7C9A9279E4D4000149E7AE31F7C63000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000800410A61BC1C292F950417C10520838835249A92455C9A928550A28D";
    attribute INIT_1B of inst : label is "925FFE7FF3F80000200000000000000000000000000500000000000000000000";
    attribute INIT_1C of inst : label is "01C924E201C924B82080C03920002E1865C0000005C0925C0000925C0240121C";
    attribute INIT_1D of inst : label is "000208000000000000000000020080000000000000000008043C00397DC021F0";
    attribute INIT_1E of inst : label is "1C00007008004B904092E0104892E0100800E4BFFCFFFFF00000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000000824BC203925F170017C40720E025C804B80000003804";
    attribute INIT_20 of inst : label is "0018000E0205FFC103FF80000000000000000000000042042040820102108000";
    attribute INIT_21 of inst : label is "B92A4B8242906E4027000E4F9008000390400C0B9245C0200201C80802E1920E";
    attribute INIT_22 of inst : label is "0000000000000000000002208120808800000000000000000000000002090A40";
    attribute INIT_23 of inst : label is "00708420210AAA1225542448D540112355424405450800389408400000000000";
    attribute INIT_24 of inst : label is "A0208807C00438421010A544000088000422200011C482494105494841540F82";
    attribute INIT_25 of inst : label is "209250415250104403E0821C290A4852AA008955091015542440E24124A082A4";
    attribute INIT_26 of inst : label is "0691EB8B1AD7002820A92828A281F2400E14852421554244A284000A88000071";
    attribute INIT_27 of inst : label is "E883FFFC00000AB000156ABFC820055000000000010000053040040000047100";
    attribute INIT_28 of inst : label is "FFFFFA0EFFFFE7FE1E7FF8FFFD6FD571550A14AB9FC0001563041AB56AD55587";
    attribute INIT_29 of inst : label is "F7DF71F6C7DFEAB5F775577555553DF55DF7BBFABBBFFBBABAAA9577FFFFFF6F";
    attribute INIT_2A of inst : label is "FFFC444F1EFFFFFF82223FD5610FD1AAA0AAAABAA0081E6ABF77F7DFBEFBFDF7";
    attribute INIT_2B of inst : label is "5555538DA2422424AAA22A8AAA0AAF55B441FFFFFE3FFFE7038FF8E347FC7F8F";
    attribute INIT_2C of inst : label is "FFF27671FDF4EC55EBBFAF47EAAABFFFEFFFFFFFEFFFFFFFFFFFAAD501255051";
    attribute INIT_2D of inst : label is "654E81DF55E070381FFF7FC3FBE9D9FFF27671FDF4ECE070381FFF7FC3FBE9D9";
    attribute INIT_2E of inst : label is "FFFFFFEEEEAEEFD56ABFFFC0309652C0097144D97D1365F40803BEABFFFCAA94";
    attribute INIT_2F of inst : label is "55D0AAAAAAAAAAAAAAA9567FFFF9FFF1FFFFF00EFFFF00EFAA8049FDDFFE20FF";
    attribute INIT_30 of inst : label is "249000A04124920100301CF1F011E023C073C7C047808EABE855555555555555";
    attribute INIT_31 of inst : label is "420A0042A8C400FAEBAE1892DA52E554D9B366C0000408102040A24820482089";
    attribute INIT_32 of inst : label is "84C91648215328A995B15338A8B7B1610B4514ACE51946519461184611846118";
    attribute INIT_33 of inst : label is "B3633955CF8156001B08583C219A4C96C0C498B68CCCF15629001CF3CF3C692E";
    attribute INIT_34 of inst : label is "9C4000000000000003C05FEBAABBBA021081166DD63329CA5C4C731B8DFBB8DB";
    attribute INIT_35 of inst : label is "2CA4B29280100000540004001408840084004400008107C000006420C8400E40";
    attribute INIT_36 of inst : label is "7FF8000FF9FFC0007FCEA3AAABABEBFB80842045A292CA4B292CA4B292CA4B29";
    attribute INIT_37 of inst : label is "2A874A5681543A400050050E0822131DB988002802871109883C822411408595";
    attribute INIT_38 of inst : label is "004400008107C000006420C8400E409C4000000000000003C05295A2A8001150";
    attribute INIT_39 of inst : label is "04000000081C05011024F22921D93C004764110F03B000540004001408840084";
    attribute INIT_3A of inst : label is "430743074018400E400054510408A284008684000358000740E8054022000000";
    attribute INIT_3B of inst : label is "0852807367231428041A900A4091202240000008430F43074307430743074307";
    attribute INIT_3C of inst : label is "2808C01125B6021000820800069FFF822404020000C00EE201B080D2A501A548";
    attribute INIT_3D of inst : label is "220344050000F189E3400000A802403101401451040000000000040806082850";
    attribute INIT_3E of inst : label is "4301F402195000000000000000000000000120000020030100000000F6F62000";
    attribute INIT_3F of inst : label is "39310000000000001F4001008004A6000A20A04D4C80021640440680000AD01C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "5EAFEABFFEEA3E909215A856A15A856C2B50AD5116B2C9A5AA36B2CCD2DDF172";
    attribute INIT_01 of inst : label is "000000000000000000000008208A80A80A888208208202200A000ABFAAA8FA42";
    attribute INIT_02 of inst : label is "628E6C73CC51CC73CC51CD8A398E798A39314731CF3147260000000000000000";
    attribute INIT_03 of inst : label is "FFFFFFFFFFF3F9F03813CF31C762F2F7BB8803DDC4C4112C5A69B1471476628E";
    attribute INIT_04 of inst : label is "4F66D12DA25B44B6896D12DA25B44B45D775DD775DD5555F0EA00802BFFFFFFF";
    attribute INIT_05 of inst : label is "B09048C232AC42FA68674B939211112256648E8B24745247452474593E3B4F67";
    attribute INIT_06 of inst : label is "012509D1D11A2A5A1882884B14E280BA7BA2B100000000000A8673902CA29B20";
    attribute INIT_07 of inst : label is "C7E2200C3F102CF0000000000101028888C8C0033FFFF1666222555EABAE24AB";
    attribute INIT_08 of inst : label is "E4E89A69168C924279BEDA3E7D3E93BE49227D279FB241B7DFA24113E8A05591";
    attribute INIT_09 of inst : label is "000000000000000000000000000000000000000000000047DF39FA248F48934C";
    attribute INIT_0A of inst : label is "F448F24401E000058197D810843EC53207814A8407805505AA80000000000000";
    attribute INIT_0B of inst : label is "268E7E8936D17EC92449E7BFB7CDE7BF27C9227D3F6D327DBE491249E44DA169";
    attribute INIT_0C of inst : label is "000000000000000000000000000000000000000000000000040F20727C49F3D2";
    attribute INIT_0D of inst : label is "DE9E49100000A0140C63FFC8A5085FCB308B02B1080FDC02A82D540000000000";
    attribute INIT_0E of inst : label is "12699C9DF34D22D1F2487F3CFB767FBEFA449FA26FB6DFA24FA48927DEDC4DB7";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000000000000000081F7CE4FC923D";
    attribute INIT_10 of inst : label is "C9F93E8525F91E46200F23002A435FA1804210BF81FE08400AA0B55000000000";
    attribute INIT_11 of inst : label is "CE7E891E89BECE6F893E914FC9244FB7DFEE4FA7DFE8492426DEFD3724F7ED13";
    attribute INIT_12 of inst : label is "00000000000000000000000000000000000000000000000000000000000087A7";
    attribute INIT_13 of inst : label is "F7800210FE08C51E47200AA5505A36ED1B768DBB46DDA36ED1B768DBB0000000";
    attribute INIT_14 of inst : label is "BA2AAB49C5800004302045B22A02C0488B44504534C6A55E9F0000531A95703D";
    attribute INIT_15 of inst : label is "A3D20000000000430910D31598AAA8BA358D40A142EB656982828E8AAAD27170";
    attribute INIT_16 of inst : label is "544B9E6D65B3CF36B2D9E59B592CF2CDA49679611664C4C5196F96894A6014D0";
    attribute INIT_17 of inst : label is "A5484F1D917ECA4A4A4A4ECEC8BF6765252525210404B29B03A537274A6C6E91";
    attribute INIT_18 of inst : label is "88888888889DBB22FDBB295252A4A5494A93B7676EC8BF6ECEDD94A9295252A4";
    attribute INIT_19 of inst : label is "7D145B8378E3930248A2981B6DC1228814AE3A9500AAAAAA888888888888AA88";
    attribute INIT_1A of inst : label is "00000002007A06CF1CFDE247A069A39A704D34536049303E9DDFB03EDDDFB830";
    attribute INIT_1B of inst : label is "2488008004080000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "FF924914FF9249134D3FFD924FFF44FFC89FFDFB68902489F6D02489F49FA4C9";
    attribute INIT_1D of inst : label is "00000000000000180000000000000000000000000000080FEF9CFF92389B4CE6";
    attribute INIT_1E of inst : label is "C9F6DB27D3EE91241A244FA412244FA7D3B64910010000100000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000080F491CBBF248E426DA391B24D17489EE913DDF6ED93E9";
    attribute INIT_20 of inst : label is "FBF3F7E480808000420080000000000000000000000000000000400000000000";
    attribute INIT_21 of inst : label is "124091349827C49B48B7E4913EDF7FB93E9F7FA124909B7BF4DC93DFB44F27E4";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000203D3E0FD";
    attribute INIT_23 of inst : label is "32D8E53B29D991C99923933AE48E4CCB9239332E58E5DE941A5AC00000000000";
    attribute INIT_24 of inst : label is "9641B62B07196C629914ECD9EDDEB3DBB97ACF6EF4A0D659A20C9B24832C560C";
    attribute INIT_25 of inst : label is "3596688326CB20DA15838EB6314C8A666CF6EF59EDDEBD67B772506B2CD1064D";
    attribute INIT_26 of inst : label is "EE972E59DEE31034419365906D8AC1865B1CA7653B367B7724F6665C91C99D28";
    attribute INIT_27 of inst : label is "EF7C1DFFDFCEEAB1FFE04AB1FE78055AAAAAAAAAAAAAAAEFEAFFAFEAAABEEAAA";
    attribute INIT_28 of inst : label is "73FFFBFEFFFEFFEFDCFFFEFFE128D57D02FDFAABD05D75D57F07D0E1C38755FF";
    attribute INIT_29 of inst : label is "F69A69F0A69F6ABFFFFFFFFFFFFFBFFFFDE7FFFFFFFFFFFFFFFC1574FFEE676F";
    attribute INIT_2A of inst : label is "A003005001802800D70000156ACC99AAAAAAAAAAAAABD56AB06F769F34FAA9A7";
    attribute INIT_2B of inst : label is "FFFFFA6DFB7FB7B7FFFFFFFFFFFFFF55EE6126C0612780109349449AE0000600";
    attribute INIT_2C of inst : label is "E6DB667FEDB6CC55F07FC177F00ABC0020C63C0020C63C007800AAFFFDBFFFFF";
    attribute INIT_2D of inst : label is "757AFFFF55BFDFEFFDB66D9FDB6D99E6DB667FEDB6CCFFDFEFFDB66D9FDB6D99";
    attribute INIT_2E of inst : label is "C0FFFF00000003D56ABE600FB18971517E644F7A4401E91090FFFEABE603AADB";
    attribute INIT_2F of inst : label is "00070000000000000001576FCC06A500A5BF37FFEFF37FFFAA806FC000003EFF";
    attribute INIT_30 of inst : label is "9249269348924924926031021800000000C40800000000AB0380000000000000";
    attribute INIT_31 of inst : label is "BACE2001E15249AAFEAEB0B2934DCE94D9B366CD9B3264D9B326612492249244";
    attribute INIT_32 of inst : label is "F4C996E591CA28E515A1CA28E4A5A1EC8E623D89C6F1BC6F1BC6F1BC6F1BC6F1";
    attribute INIT_33 of inst : label is "EB1302A96B828128192D849F339B68E824C74CB6C8889217295498A28A24892E";
    attribute INIT_34 of inst : label is "001500002150000217C00AABEFBEBFA318C012B8772D7B5EC29EE7B857DF8570";
    attribute INIT_35 of inst : label is "E8DBA373900925400140014001400140014001400A0050028005000A00140014";
    attribute INIT_36 of inst : label is "4000000FFE0000007FF47D1FC145541528C63004B36E8DBA36E8DBA36E8DBA36";
    attribute INIT_37 of inst : label is "001059B2400083CD0000002000000041F5E10000001000000086807403F2593A";
    attribute INIT_38 of inst : label is "4001400A0050028005000A00140014001500002150000217C0066C9000000410";
    attribute INIT_39 of inst : label is "054000000A8000001070F000041C3C0010700000083140014001400140014001";
    attribute INIT_3A of inst : label is "1407140714001400140000015000000540000054000002A0140A805402A00000";
    attribute INIT_3B of inst : label is "A000AA00005401400140010005002A0054001400140F14071407140714071407";
    attribute INIT_3C of inst : label is "8407120883FF200C101020088000002804045000500050E0000009008512010A";
    attribute INIT_3D of inst : label is "008020203FFFF803F0207FFD50880480FE220220909FFFFFFFFFFC03F0900480";
    attribute INIT_3E of inst : label is "20FFF890440241FFFFFFFFFFFFFFFFFFFFF807F202010008FFFFFFFFFFFF1FFE";
    attribute INIT_3F of inst : label is "7B77FFFFFFFFFFFFFF8F92011102109FC1501000803FF8402401007FF2400900";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "30444014504015C2CCC3130C4C3130C1862618C727962BB286079725D902A94B";
    attribute INIT_01 of inst : label is "AAAAAAAAAAAAAAAAAAAAAAA082AAA28AAAA2A28A2AA2A82AAAAAB1114444570B";
    attribute INIT_02 of inst : label is "638E4C73CC71CC73CC71C98E398E798E3931C731CF31C726AAAAAAAAAAAAAAAA";
    attribute INIT_03 of inst : label is "100E640201FFFFC020134F714762D37C9EB9124F5CE2516C5A7BB1C71C77638E";
    attribute INIT_04 of inst : label is "CF26D16DA2DB45B68B6D16DA2DB45BC5F57DDF17CDD555500AA00802A0400200";
    attribute INIT_05 of inst : label is "53C3394E583B804507B8BB6B6CFAE6CDA9966068B3030B3030B303059A39CF27";
    attribute INIT_06 of inst : label is "6C702C9595F981707A802930E35F62F9060D6E0000000000FD11A94948E0C586";
    attribute INIT_07 of inst : label is "EFF77FFF7FBFFCF0000000000101028888C8C0033FFFF7FDD99978708EF1B28E";
    attribute INIT_08 of inst : label is "F6EDDB6DF6EDDB777DBEDBBF7DBEDBBF6DB77DB7DFB77DB7DFB77DBBEFBFDDBB";
    attribute INIT_09 of inst : label is "000000000000000000000000000000000000000000000057DF7DFB76DF6DDB6D";
    attribute INIT_0A of inst : label is "F6EDFB6FFBFFFFEEE2000780000E77FFE01188840381FFAF5080000000000000";
    attribute INIT_0B of inst : label is "76DF7EDDB6DF7EDDB6EDF7BFB7EDF7BFB7EDB77DBF6DB77DBF6DBB6DF6EDBF6D";
    attribute INIT_0C of inst : label is "000000000000000000000000000000000000000000000000042FBEFB7EEDF7DB";
    attribute INIT_0D of inst : label is "DEDEEDBFFFFFBFFE2100707C000007DFF5E002394800600FFD7A840000000000";
    attribute INIT_0E of inst : label is "BB6DBEDDFB6DBEDDFB6EFFBEFB76FFBEFB6EDFB76FB6DFB76FB6DDB7DEDEEDB7";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000000000000000085F7DF6FDDB7D";
    attribute INIT_10 of inst : label is "EDFBBEFDBDFBBF6F7FFFB7FFF71C0201D00000247F969CE53FF5E83000000000";
    attribute INIT_11 of inst : label is "DF7EDDBEDDBEDF6FDDBEDF6FDDB6EFB7DFEEEFB7DFEEEDB776DEFDB776F7EDBB";
    attribute INIT_12 of inst : label is "00000000000000000000000000000000000000000000000000000000000087B7";
    attribute INIT_13 of inst : label is "20F802108BAFFF884E62144FFAFFC24FE127F093F849FC24FE127F0930000000";
    attribute INIT_14 of inst : label is "601897841700000495D168B800DB99A444140731128430740854570800C1CCC0";
    attribute INIT_15 of inst : label is "1058000000000049572258C44601F6F91E12374E9D60DEE46020380625E105D1";
    attribute INIT_16 of inst : label is "31D54F90914826C848A41164241208B21209045417B1919DAE1ACF6D296AB722";
    attribute INIT_17 of inst : label is "366D4C4FC017E7E7E7E7E3636009B1B1B1B1B1B5EA3629FF27FFFE5FFFFD9FFC";
    attribute INIT_18 of inst : label is "D7D7D7D7D7CFDF802FDF9FBF3F7E7EFCFDF8D9B1B36009B36366C6CD8D9B1B36";
    attribute INIT_19 of inst : label is "7DF7DBAB7DF7DBAB6FBEDD5B6DD5BEFAF7BF7EF781FFFFFFF5F5F5F5F5F5FFD7";
    attribute INIT_1A of inst : label is "00000002007B0EEFBEFDEB6FB56DB7DB756DB7DB756DBABEDDDFBABEDDDFBAB5";
    attribute INIT_1B of inst : label is "B6DFFEFFF7FC0000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "FFDB6DF6FFDB6DBB6DBFFDBB6FFF6EFFEDDFFDFB6DDFB6DDF6DFB6DDF6DFB6DD";
    attribute INIT_1D of inst : label is "00000000000000000000000000000000000000000000080FEFBEFFBB7DDB6DF6";
    attribute INIT_1E of inst : label is "DDF6DB77DBEEDBB7DBB6EFB7DBB6EFB7DBB6EDBFFDFFFFF80000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000080F6DBEFBFB6DF776DB7DDB76DF76DDEEDBBDDF6EDBBED";
    attribute INIT_20 of inst : label is "FBFBF7EEFEFDFFFF7FFFC0000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "BB6ADBB6DAB7EEDB6FB7EEDBBEDF7FBBBEDF7FBBB6DDDB7BF6DDDBDFB6EFB7EE";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000203DBEAFD";
    attribute INIT_23 of inst : label is "25061585AC6C6EF666DDECC51B77B3146DDECC51B77B334321A5000000000000";
    attribute INIT_24 of inst : label is "491CC9233196830AC2D616377B316EF66285BBD99A19296638E6649239964661";
    attribute INIT_25 of inst : label is "4A598E3999248E65919849418D632B0B1BBD99B77B3346DDECCD0C94B31C7332";
    attribute INIT_26 of inst : label is "11698B0C6B1B42C71CCC924732C8CC24A0C2B0B58D8DDECCD3BD11A34CE44286";
    attribute INIT_27 of inst : label is "EF7FEABDDFCEEAB1FFE06AB1FE78755000000000010000004000100000010440";
    attribute INIT_28 of inst : label is "7FFFFBFEFFFEFFEFDCFFFEFFE12BD57D02FDFAABD05D75D56F0413E7CF9F559F";
    attribute INIT_29 of inst : label is "F69A69F0A69F0ABFFFFFFFFFFFFFBFFFFDE7FFFFFFFFFFFFFFFC1574FFEFFF6F";
    attribute INIT_2A of inst : label is "FFFF7FFFFFBFFFFFDCFFFFD56ACC99AAAAAAAAAAAAABD50AB06F769F34FAA9A7";
    attribute INIT_2B of inst : label is "FFFFFBEDFB7FB7B7FFFFFFFFFFFFFF55B9FFFE3FFFFFFFFFFF7FFFFB9FFFFEFF";
    attribute INIT_2C of inst : label is "DFFFEEF7DFFFDD55CE0038440FEAB40000C60C0000C60C0018002AFFFDBFFFFF";
    attribute INIT_2D of inst : label is "FAA17FF055A7D3E9FFFFFFBFBFFFBBDFFFEEF7DFFFDCE7D3E9FFFFFFBFBFFFBB";
    attribute INIT_2E of inst : label is "FFFFFF00000000156ABE603FD874CECF9F1F17C99C8926700CFFE0ABE603FF6A";
    attribute INIT_2F of inst : label is "01800000000000000001564FCC06A5FFA53F37FFEFF37FF82A8039C0007FBEFF";
    attribute INIT_30 of inst : label is "4DB4D269374D36D34D38300000007000E0C0006001C002ABC000000000000000";
    attribute INIT_31 of inst : label is "4DA0C181630249550005E2E848FF9FFF66CD9B366CD9B366CD9B3E9A699A69B3";
    attribute INIT_32 of inst : label is "5BA44D872C0B9605C33C0B9606333C18E199E3673D2F4BD2F4BD2F4BD2F4BD2F";
    attribute INIT_33 of inst : label is "BD904F95CE49E2B84C578AC5E06E93B455B322EBA666498F84AAC24924926CBB";
    attribute INIT_34 of inst : label is "FF02FFFFD42FFFFD403FC554104015A94A4049E85D1FCE7387F5AD68FC488FD0";
    attribute INIT_35 of inst : label is "7F09FC3E4909243FF03FF03FF03FF03FF03FF03F81FC0FE07FC0FF81FF03FF03";
    attribute INIT_36 of inst : label is "C000000003FFFFFF80357D5FC55040516A5290127C27F09FC27F09FC27F09FC2";
    attribute INIT_37 of inst : label is "00181FF7C000C05F4000003000000060A04400000018000000C6093049A24FBF";
    attribute INIT_38 of inst : label is "8002803400A00D001A0034006800680068000002800000280007FDF000000600";
    attribute INIT_39 of inst : label is "02800000050000000808000006020000180800000C0680028002800280028002";
    attribute INIT_3A of inst : label is "680068006800680068000000A00000028000002800000140680D002801400000";
    attribute INIT_3B of inst : label is "4000340000680280068006001A005400A8006800E80068006800680068006800";
    attribute INIT_3C of inst : label is "000000000000000000000000000000500000A000A000A0000000A20001440003";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "EF1D800000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "044440145040178A8C80120048012001002400CAB30402A0951304015020056B";
    attribute INIT_01 of inst : label is "55555555555555555555555DFD555DF55555FD5FD5FD57D55555511144445E2A";
    attribute INIT_02 of inst : label is "628B6C536C516C536C516D8A2D8A6D8A2DB145B14DB145B75555555555555555";
    attribute INIT_03 of inst : label is "100E67FE01FF807FE0134DF145E3DBBD10A0028850E211EC7A6F3145145F628B";
    attribute INIT_04 of inst : label is "4DF6D1ADA35B46B68D6D1ADA35B46B47D5F5FD1F4FD555500AA00802A07F03F8";
    attribute INIT_05 of inst : label is "7A8A3DEB502202452234A50A045C0F5EB5144038A201CA2018A201851A2F4DF7";
    attribute INIT_06 of inst : label is "2860A816165B03431F7F570680023CA7C2602A0000000000A87C800E9AA08614";
    attribute INIT_07 of inst : label is "EFF77FFF7FBFECF0000000000101028888C8C0033FFFF3F55111204088FBA288";
    attribute INIT_08 of inst : label is "F6EDDB6DF6EDDB777DBEDBBF7DBEDBBF6DB77DB7DFB77DB7DFB77DBBEFBFDDBB";
    attribute INIT_09 of inst : label is "000000000000000000000000000000000000000000000017DF7DFB76DF6DDB6D";
    attribute INIT_0A of inst : label is "F6EDFB6FFBFFFFED81DFF8318C7EC5320FC73D28038000500080000000000000";
    attribute INIT_0B of inst : label is "76DF7EDDB6DF7EDDB6EDF7BFB7EDF7BFB7EDB77DBF6DB77DBF6DBB6DF6EDBF6D";
    attribute INIT_0C of inst : label is "000000000000000000000000000000000000000000000000002FBEFB7EEDF7DB";
    attribute INIT_0D of inst : label is "DEDEEDBFFFFFBFF40462FBE06318DFC330070E5A500060000280040000000000";
    attribute INIT_0E of inst : label is "BB6DBEDDFB6DBEDDFB6EFFBEFB76FFBEFB6EDFB76FB6DFB76FB6DDB7DEDEEDB7";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000000000000000005F7DF6FDDB7D";
    attribute INIT_10 of inst : label is "EDFBBEFDBDFBBF6F7FFFB7FFEA437FA100318C5F91FE2948400A001000000000";
    attribute INIT_11 of inst : label is "DF7EDDBEDDBEDF6FDDBEDF6FDDB6EFB7DFEEEFB7DFEEEDB776DEFDB776F7EDBB";
    attribute INIT_12 of inst : label is "00000000000000000000000000000000000000000000000000000000000007B7";
    attribute INIT_13 of inst : label is "FF808631EE0ACD1F1CF6B000050FA24FD127E893F449FA24FD127E8930000000";
    attribute INIT_14 of inst : label is "6808801E74000004F580FBB1D44A8FC1F6EEAA211F08204503BBFE3C20811039";
    attribute INIT_15 of inst : label is "785000000000004F5661D0C487D5E2A7DC03360C18411C1E7D5D5A0220079D10";
    attribute INIT_16 of inst : label is "31800D000100008000800240000001200000009FEAA0809FCE12AF7DAD555730";
    attribute INIT_17 of inst : label is "12255F6262213131313131313110989898989897BA6421FF77FFFE4FFFFE9FF8";
    attribute INIT_18 of inst : label is "802A802A806244C44244C48989131226244C48989131109131226244C4898913";
    attribute INIT_19 of inst : label is "7DF7DBAB7DF7DBAB6FBEDD5B6DD5BEFAF7BF7EF70000000000AA00AA00AA002A";
    attribute INIT_1A of inst : label is "00000000007B0EEFBEFDEB6FB56DB7DB756DB7DB756DBABEDDDFBABEDDDFBAB5";
    attribute INIT_1B of inst : label is "B6DFFEFFF7F80000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "FFDB6DF6FFDB6DBB6DBFFDBB6FFF6EFFEDDFFDFB6DDFB6DDF6DFB6DDF6DFB6DD";
    attribute INIT_1D of inst : label is "00000000000000000000000000000000000000000000000FEFBEFFBB7DDB6DF6";
    attribute INIT_1E of inst : label is "DDF6DB77DBEEDBB7DBB6EFB7DBB6EFB7DBB6EDBFFDFFFFF00000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000000F6DBEFBFB6DF776DB7DDB76DF76DDEEDBBDDF6EDBBED";
    attribute INIT_20 of inst : label is "FBFBF7EEFEFDFFFF7FFF80000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "BB6ADBB6DAB7EEDB6FB7EEDBBEDF7FBBBEDF7FBBB6DDDB7BF6DDDBDFB6EFB7EE";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000003DBEAFD";
    attribute INIT_23 of inst : label is "368E5517A8F008400E10801EB842007AE10801EB842005A283D6800000000000";
    attribute INIT_24 of inst : label is "00188B22239F472A8BD47804200708400F5C21002D14355430C4400031124445";
    attribute INIT_25 of inst : label is "0D550C3110000C459111CFA39D47EA3C021002842005AA1080168A1AAA186220";
    attribute INIT_26 of inst : label is "BAAFC79CEF3A01861888000622C888E7D1CEA3D5160108014A108AD52A522B45";
    attribute INIT_27 of inst : label is "0880000220310ABE001F8ABE0187855FFFFFFFFFFFFFFFFE9BAEFFFFFFEB8FFF";
    attribute INIT_28 of inst : label is "8000020080010010230001001DCC1572FD0204AB2FA28A1570F7DC18306055E0";
    attribute INIT_29 of inst : label is "0555550F5550EAB0000000000000200001140000000000000003D56700100048";
    attribute INIT_2A of inst : label is "0000800000400000200000157533555555555555554C1AEABF508550AA855554";
    attribute INIT_2B of inst : label is "00000209024024240000000000000055C0000100000000000080000400000100";
    attribute INIT_2C of inst : label is "749255582924AA55FFFFFF77FFEABBFFFF39F7FFFF39F7FFEFFFAAC001200000";
    attribute INIT_2D of inst : label is "4000000F55F83C1E09244960524955749255582924ABB83C1E09244960524955";
    attribute INIT_2E of inst : label is "000000FFFFFFFFD56AB19FFFCCC758C79E2A1BD09001424008001EAB19FF2A02";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFD57F033F95A005AC0C800100C8007AA807D3FFF802080";
    attribute INIT_30 of inst : label is "0490402015041241043FDFFFFFFFFFFFFF7FFFFFFFFFFEABFFFFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "4C804081C12249EAAAAFAAA001FFFFFD42850A142850A142850A3A08210820A1";
    attribute INIT_32 of inst : label is "228084A5680904048118090404111808C088AD0155354D5354D5354D5354D535";
    attribute INIT_33 of inst : label is "1F89479485C1E0AF809F8281A172BAA01680F2ACAEEEC105102A8EFBEFB078A1";
    attribute INIT_34 of inst : label is "006800000280000028000AAAAAAABFB0842381C0009E421087D08420F8000F80";
    attribute INIT_35 of inst : label is "7E89FA3C0B0926800280028002800280028002803400A00D001A003400680068";
    attribute INIT_36 of inst : label is "FFFFFFF0060000000014952572A24A112C2108E07A27E89FA27E89FA27E89FA2";
    attribute INIT_37 of inst : label is "FFC83FF7DFFE40325FFFFF90FFFFFF2091C00FFFFFC87FFFFE42001800C00FBF";
    attribute INIT_38 of inst : label is "3FF03F81FC0FE07FC0FF81FF03FF03FF02FFFFD42FFFFD403FCFFDF7FFFFF207";
    attribute INIT_39 of inst : label is "F43FFFFFE87FFFFFD9180FFFF20603FFC818FFFFE40C3FF03FF03FF03FF03FF0";
    attribute INIT_3A of inst : label is "03F803F803FF03FF03FFFFFD0FFFFFF43FFFFF43FFFFFA1F03E87F03FA1FFFFF";
    attribute INIT_3B of inst : label is "1FFF01FFFF43F43FF03FF0FFC0FF81FF03FF03FF43F003F803F803F803F803F8";
    attribute INIT_3C of inst : label is "7BF8EDF77C00DFF3EFEFDFF77FFFFF87FBF80FFC0FFC0F1FFFFE00FF7801FEF0";
    attribute INIT_3D of inst : label is "FF7FDFDFC00007FC0FDF8002AF77FB7F01DDFDDF6F600000000003FC0F6FFB7F";
    attribute INIT_3E of inst : label is "DF00076FBBFDBE0000000000000000000007F80DFDFEFFF7000000000000E001";
    attribute INIT_3F of inst : label is "EF2180000000000000706DFEEEFDEF603EAFEFFF7FC007BFDBFEFF800DBFF6FF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
