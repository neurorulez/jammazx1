library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"20",X"E3",X"7B",X"A5",X"CD",X"D0",X"0A",X"85",X"CC",X"85",X"CB",X"85",X"CE",X"A9",X"20",X"85",
		X"CD",X"20",X"59",X"69",X"2C",X"02",X"20",X"30",X"FB",X"20",X"A2",X"4B",X"46",X"75",X"90",X"FC",
		X"A5",X"76",X"29",X"01",X"0A",X"AA",X"49",X"02",X"A8",X"BD",X"99",X"77",X"8D",X"00",X"40",X"BD",
		X"9A",X"77",X"8D",X"01",X"40",X"B9",X"99",X"77",X"0A",X"85",X"03",X"B9",X"9A",X"77",X"2A",X"29",
		X"1F",X"09",X"40",X"85",X"04",X"8D",X"00",X"30",X"8D",X"00",X"34",X"E6",X"76",X"D0",X"30",X"E6",
		X"77",X"A6",X"20",X"B5",X"64",X"29",X"0F",X"85",X"10",X"55",X"64",X"4A",X"85",X"11",X"4A",X"4A",
		X"65",X"11",X"65",X"10",X"A6",X"1F",X"A4",X"77",X"C0",X"80",X"D0",X"08",X"D5",X"FA",X"D0",X"02",
		X"F6",X"FB",X"95",X"FA",X"18",X"75",X"FB",X"C9",X"10",X"90",X"02",X"A9",X"0F",X"85",X"D3",X"20",
		X"FF",X"7A",X"20",X"E1",X"4B",X"B0",X"42",X"20",X"D4",X"6F",X"20",X"6B",X"65",X"10",X"1E",X"20",
		X"9D",X"6C",X"B0",X"19",X"A5",X"74",X"D0",X"0F",X"20",X"59",X"66",X"20",X"97",X"64",X"20",X"10",
		X"68",X"20",X"9E",X"4A",X"20",X"22",X"63",X"20",X"DC",X"66",X"20",X"F7",X"60",X"20",X"7E",X"6A",
		X"20",X"F6",X"6E",X"A9",X"7F",X"AA",X"20",X"1F",X"7A",X"20",X"DA",X"79",X"AD",X"EC",X"02",X"F0",
		X"03",X"CE",X"EC",X"02",X"0D",X"E7",X"02",X"D0",X"03",X"4C",X"11",X"60",X"4C",X"14",X"60",X"B2",
		X"A5",X"42",X"25",X"43",X"30",X"03",X"4C",X"C7",X"7B",X"18",X"60",X"A5",X"8A",X"05",X"13",X"10",
		X"07",X"A5",X"76",X"29",X"20",X"F0",X"01",X"60",X"4C",X"59",X"71",X"A0",X"01",X"20",X"59",X"71",
		X"A4",X"1E",X"C8",X"98",X"4C",X"EB",X"79",X"46",X"71",X"A2",X"07",X"BD",X"19",X"02",X"F0",X"02",
		X"10",X"0A",X"CA",X"10",X"F6",X"24",X"71",X"30",X"02",X"86",X"72",X"60",X"A0",X"1A",X"E0",X"04",
		X"B0",X"07",X"88",X"8A",X"D0",X"03",X"88",X"30",X"E9",X"B9",X"00",X"02",X"F0",X"F8",X"30",X"F6",
		X"85",X"0C",X"B9",X"63",X"02",X"38",X"FD",X"7C",X"02",X"E9",X"03",X"C9",X"FA",X"90",X"E7",X"B9",
		X"84",X"02",X"FD",X"9D",X"02",X"E9",X"03",X"C9",X"FA",X"90",X"DB",X"B9",X"A5",X"02",X"38",X"FD",
		X"BE",X"02",X"85",X"09",X"B9",X"63",X"02",X"FD",X"7C",X"02",X"4A",X"66",X"09",X"0A",X"F0",X"0E",
		X"10",X"C4",X"49",X"FE",X"D0",X"C0",X"A5",X"09",X"49",X"FF",X"69",X"00",X"85",X"09",X"B9",X"C6",
		X"02",X"38",X"FD",X"DF",X"02",X"85",X"0A",X"B9",X"84",X"02",X"FD",X"9D",X"02",X"4A",X"66",X"0A",
		X"0A",X"F0",X"0E",X"10",X"A1",X"49",X"FE",X"D0",X"9D",X"A5",X"0A",X"49",X"FF",X"69",X"00",X"85",
		X"0A",X"A9",X"04",X"E0",X"01",X"F0",X"07",X"B0",X"08",X"20",X"D5",X"61",X"D0",X"03",X"20",X"DE",
		X"61",X"C0",X"19",X"B0",X"10",X"69",X"2A",X"46",X"0C",X"B0",X"14",X"69",X"1E",X"46",X"0C",X"B0",
		X"0E",X"69",X"3C",X"90",X"0A",X"F0",X"05",X"20",X"DE",X"61",X"D0",X"03",X"20",X"D5",X"61",X"C5",
		X"09",X"90",X"1F",X"C5",X"0A",X"90",X"1B",X"85",X"0C",X"4A",X"18",X"65",X"0C",X"6A",X"85",X"0C",
		X"A5",X"0A",X"65",X"09",X"6A",X"C5",X"0C",X"B0",X"09",X"8A",X"48",X"20",X"A1",X"62",X"68",X"AA",
		X"A0",X"00",X"4C",X"16",X"61",X"24",X"73",X"10",X"02",X"69",X"08",X"69",X"1C",X"60",X"69",X"1C",
		X"48",X"AD",X"1A",X"02",X"4A",X"68",X"B0",X"02",X"69",X"12",X"60",X"B9",X"00",X"02",X"29",X"07",
		X"85",X"09",X"AD",X"0A",X"2C",X"29",X"18",X"05",X"09",X"9D",X"00",X"02",X"B9",X"A5",X"02",X"9D",
		X"A5",X"02",X"B9",X"63",X"02",X"9D",X"63",X"02",X"B9",X"C6",X"02",X"9D",X"C6",X"02",X"B9",X"84",
		X"02",X"9D",X"84",X"02",X"B9",X"21",X"02",X"9D",X"21",X"02",X"B9",X"42",X"02",X"9D",X"42",X"02",
		X"60",X"A0",X"FF",X"24",X"12",X"30",X"2D",X"C8",X"C8",X"B1",X"10",X"45",X"0A",X"91",X"03",X"88",
		X"C9",X"F0",X"B0",X"17",X"B1",X"10",X"91",X"03",X"C8",X"C8",X"B1",X"10",X"91",X"03",X"C8",X"B1",
		X"10",X"45",X"09",X"91",X"03",X"CA",X"10",X"DF",X"4C",X"55",X"7A",X"B1",X"10",X"45",X"09",X"91",
		X"03",X"C8",X"D0",X"F1",X"C8",X"B1",X"10",X"85",X"14",X"C8",X"B1",X"10",X"C9",X"F0",X"B0",X"2C",
		X"C8",X"C8",X"51",X"10",X"29",X"0F",X"85",X"13",X"51",X"10",X"45",X"09",X"91",X"03",X"88",X"B1",
		X"10",X"48",X"A5",X"14",X"91",X"03",X"88",X"A5",X"13",X"45",X"0A",X"51",X"10",X"91",X"03",X"88",
		X"68",X"91",X"03",X"C8",X"C8",X"C8",X"CA",X"10",X"CB",X"4C",X"55",X"7A",X"45",X"14",X"29",X"07",
		X"48",X"51",X"10",X"45",X"0A",X"91",X"03",X"88",X"68",X"51",X"10",X"45",X"09",X"91",X"03",X"B0",
		X"E4",X"20",X"E7",X"74",X"B0",X"62",X"E0",X"01",X"D0",X"06",X"C0",X"19",X"D0",X"08",X"CA",X"C8",
		X"8A",X"D0",X"16",X"20",X"F8",X"62",X"A9",X"A0",X"9D",X"19",X"02",X"A9",X"00",X"9D",X"3A",X"02",
		X"9D",X"5B",X"02",X"C0",X"19",X"90",X"0D",X"B0",X"3F",X"A9",X"00",X"9D",X"19",X"02",X"C0",X"19",
		X"F0",X"21",X"B0",X"34",X"20",X"62",X"6F",X"B9",X"00",X"02",X"29",X"03",X"49",X"02",X"4A",X"6A",
		X"6A",X"09",X"3F",X"85",X"7F",X"A9",X"A0",X"99",X"00",X"02",X"A9",X"00",X"99",X"21",X"02",X"99",
		X"42",X"02",X"60",X"20",X"F8",X"62",X"D0",X"DF",X"8A",X"A6",X"1E",X"D6",X"6F",X"AA",X"A9",X"81",
		X"8D",X"EB",X"02",X"A9",X"05",X"85",X"DE",X"60",X"AD",X"E9",X"02",X"8D",X"E8",X"02",X"A5",X"22",
		X"F0",X"C5",X"AD",X"1A",X"02",X"4A",X"A9",X"00",X"B0",X"02",X"A9",X"20",X"20",X"44",X"6C",X"4C",
		X"D7",X"62",X"A5",X"76",X"29",X"03",X"F0",X"01",X"60",X"AD",X"1A",X"02",X"F0",X"0A",X"10",X"05",
		X"A0",X"17",X"4C",X"0D",X"77",X"4C",X"C5",X"63",X"20",X"FA",X"67",X"A5",X"22",X"F0",X"07",X"AD",
		X"19",X"02",X"F0",X"E4",X"30",X"E2",X"AD",X"EA",X"02",X"F0",X"03",X"CE",X"EA",X"02",X"CE",X"E8",
		X"02",X"D0",X"D5",X"A9",X"01",X"8D",X"E8",X"02",X"AE",X"E7",X"02",X"F0",X"CB",X"AD",X"EA",X"02",
		X"F0",X"05",X"EC",X"EE",X"02",X"B0",X"C1",X"AD",X"E9",X"02",X"38",X"E9",X"06",X"C9",X"20",X"90",
		X"03",X"8D",X"E9",X"02",X"AD",X"0A",X"2C",X"4A",X"6E",X"E0",X"02",X"4A",X"6E",X"E0",X"02",X"4A",
		X"6E",X"E0",X"02",X"69",X"04",X"C9",X"12",X"90",X"02",X"E9",X"10",X"8D",X"9E",X"02",X"AD",X"0A",
		X"2C",X"0A",X"A9",X"00",X"AA",X"A0",X"10",X"90",X"05",X"CA",X"A9",X"1F",X"A0",X"F0",X"8C",X"3B",
		X"02",X"8D",X"7D",X"02",X"8E",X"BF",X"02",X"A0",X"02",X"A5",X"D3",X"F0",X"0C",X"AD",X"EE",X"02",
		X"38",X"ED",X"E7",X"02",X"C9",X"04",X"90",X"01",X"88",X"8C",X"1A",X"02",X"B9",X"C2",X"63",X"A8",
		X"4C",X"16",X"77",X"17",X"37",X"A5",X"76",X"0A",X"D0",X"0C",X"AD",X"0A",X"2C",X"29",X"03",X"AA",
		X"BD",X"57",X"64",X"8D",X"5C",X"02",X"A5",X"22",X"F0",X"05",X"AD",X"EB",X"02",X"D0",X"05",X"CE",
		X"E8",X"02",X"F0",X"01",X"60",X"A9",X"0A",X"8D",X"E8",X"02",X"A0",X"19",X"A5",X"22",X"F0",X"0F",
		X"A2",X"AA",X"AD",X"1A",X"02",X"4A",X"B0",X"02",X"A2",X"40",X"EC",X"0A",X"2C",X"B0",X"03",X"20",
		X"5B",X"64",X"84",X"18",X"A2",X"1A",X"20",X"22",X"4A",X"20",X"E7",X"49",X"85",X"13",X"A5",X"0C",
		X"85",X"12",X"A5",X"18",X"18",X"69",X"21",X"A8",X"A2",X"3B",X"20",X"22",X"4A",X"20",X"E7",X"49",
		X"20",X"32",X"4A",X"85",X"7A",X"A5",X"18",X"C9",X"19",X"D0",X"17",X"A6",X"D3",X"E0",X"03",X"90",
		X"02",X"A2",X"03",X"AD",X"0A",X"2C",X"3D",X"4F",X"64",X"10",X"03",X"1D",X"53",X"64",X"65",X"7A",
		X"85",X"7A",X"A0",X"03",X"A9",X"01",X"85",X"0F",X"A6",X"18",X"85",X"18",X"4C",X"C8",X"64",X"9F",
		X"8F",X"8F",X"87",X"60",X"70",X"70",X"78",X"F0",X"00",X"00",X"10",X"88",X"B9",X"00",X"02",X"D0",
		X"07",X"88",X"10",X"F8",X"A0",X"19",X"38",X"60",X"30",X"F7",X"C9",X"40",X"90",X"0A",X"4A",X"4A",
		X"AA",X"BD",X"E8",X"02",X"10",X"EB",X"18",X"60",X"AD",X"7D",X"02",X"38",X"F9",X"63",X"02",X"10",
		X"02",X"49",X"FF",X"C9",X"08",X"B0",X"DA",X"AD",X"9E",X"02",X"38",X"F9",X"84",X"02",X"10",X"02",
		X"49",X"FF",X"C9",X"08",X"B0",X"CB",X"60",X"A2",X"00",X"A5",X"22",X"D0",X"03",X"86",X"FF",X"60",
		X"24",X"73",X"30",X"F9",X"24",X"FE",X"10",X"F5",X"AD",X"EB",X"02",X"D0",X"F0",X"E6",X"FF",X"A5",
		X"FF",X"C9",X"02",X"90",X"05",X"C9",X"0F",X"B0",X"E4",X"60",X"86",X"18",X"A9",X"03",X"85",X"0F",
		X"A2",X"19",X"A5",X"79",X"85",X"7A",X"A0",X"07",X"B9",X"19",X"02",X"F0",X"06",X"88",X"C4",X"0F",
		X"D0",X"F6",X"60",X"86",X"0E",X"A9",X"12",X"99",X"19",X"02",X"A5",X"7A",X"20",X"FE",X"70",X"A6",
		X"0E",X"C9",X"80",X"6A",X"85",X"0A",X"18",X"7D",X"21",X"02",X"30",X"08",X"C9",X"70",X"90",X"0A",
		X"A9",X"6F",X"D0",X"06",X"C9",X"91",X"B0",X"02",X"A9",X"91",X"99",X"3A",X"02",X"A5",X"7A",X"20",
		X"01",X"71",X"A6",X"0E",X"C9",X"80",X"6A",X"85",X"0D",X"18",X"7D",X"42",X"02",X"30",X"08",X"C9",
		X"70",X"90",X"0A",X"A9",X"6F",X"D0",X"06",X"C9",X"91",X"B0",X"02",X"A9",X"91",X"99",X"5B",X"02",
		X"A2",X"00",X"A5",X"0A",X"10",X"01",X"CA",X"86",X"09",X"A6",X"18",X"C9",X"80",X"6A",X"18",X"65",
		X"0A",X"18",X"7D",X"BE",X"02",X"99",X"BE",X"02",X"A5",X"09",X"7D",X"7C",X"02",X"99",X"7C",X"02",
		X"A2",X"00",X"A5",X"0D",X"10",X"01",X"CA",X"86",X"0C",X"A6",X"18",X"C9",X"80",X"6A",X"18",X"65",
		X"0D",X"18",X"7D",X"DF",X"02",X"99",X"DF",X"02",X"A5",X"0C",X"7D",X"9D",X"02",X"99",X"9D",X"02",
		X"A0",X"27",X"E0",X"01",X"90",X"02",X"A0",X"1F",X"4C",X"17",X"77",X"A5",X"42",X"25",X"43",X"10",
		X"0A",X"A5",X"22",X"D0",X"03",X"20",X"44",X"78",X"A9",X"FF",X"60",X"A5",X"21",X"4A",X"F0",X"18",
		X"A0",X"01",X"20",X"59",X"71",X"A0",X"02",X"A6",X"43",X"10",X"01",X"88",X"84",X"1E",X"A5",X"76",
		X"29",X"10",X"D0",X"04",X"98",X"20",X"EB",X"79",X"46",X"1E",X"20",X"95",X"6C",X"A0",X"02",X"20",
		X"59",X"71",X"A0",X"03",X"20",X"59",X"71",X"A0",X"04",X"20",X"59",X"71",X"A0",X"05",X"20",X"59",
		X"71",X"A9",X"20",X"85",X"01",X"A9",X"64",X"A2",X"39",X"20",X"1F",X"7A",X"A9",X"70",X"20",X"EA",
		X"7A",X"A6",X"1E",X"B4",X"42",X"84",X"0C",X"98",X"18",X"65",X"41",X"85",X"0D",X"20",X"C5",X"66",
		X"A4",X"0C",X"C8",X"20",X"C5",X"66",X"A4",X"0C",X"C8",X"C8",X"20",X"C5",X"66",X"0E",X"03",X"20",
		X"26",X"7B",X"A5",X"7B",X"29",X"1F",X"C9",X"07",X"D0",X"2E",X"E6",X"41",X"A5",X"41",X"C9",X"03",
		X"90",X"1A",X"A6",X"1E",X"A9",X"FF",X"95",X"42",X"A2",X"00",X"86",X"1E",X"86",X"41",X"A2",X"F0",
		X"86",X"77",X"A5",X"42",X"10",X"03",X"20",X"C7",X"7B",X"4C",X"95",X"6C",X"E6",X"0D",X"A6",X"0D",
		X"A9",X"F4",X"85",X"77",X"A9",X"0B",X"95",X"44",X"A5",X"77",X"D0",X"08",X"A9",X"FF",X"85",X"42",
		X"85",X"43",X"30",X"D4",X"A5",X"76",X"29",X"07",X"D0",X"2C",X"A6",X"0D",X"B4",X"44",X"2C",X"07",
		X"24",X"10",X"01",X"C8",X"2C",X"06",X"24",X"10",X"03",X"88",X"30",X"10",X"C0",X"0B",X"B0",X"0E",
		X"C0",X"01",X"F0",X"04",X"A0",X"00",X"F0",X"0C",X"A0",X"0B",X"D0",X"08",X"A0",X"24",X"C0",X"25",
		X"90",X"02",X"A0",X"00",X"94",X"44",X"A9",X"00",X"60",X"46",X"73",X"A5",X"22",X"F0",X"21",X"AD",
		X"19",X"02",X"30",X"1C",X"F0",X"1A",X"AD",X"EF",X"02",X"F0",X"15",X"0E",X"03",X"20",X"66",X"73",
		X"10",X"0E",X"A0",X"57",X"20",X"13",X"77",X"A5",X"76",X"29",X"03",X"D0",X"03",X"CE",X"EF",X"02",
		X"60",X"24",X"73",X"10",X"FB",X"AD",X"EF",X"02",X"29",X"F0",X"C9",X"60",X"B0",X"02",X"A9",X"60",
		X"48",X"A2",X"12",X"A9",X"50",X"86",X"10",X"85",X"11",X"A2",X"00",X"86",X"09",X"86",X"0A",X"86",
		X"12",X"20",X"21",X"62",X"A2",X"07",X"68",X"85",X"09",X"20",X"96",X"6E",X"A9",X"00",X"85",X"09",
		X"4C",X"96",X"6E",X"A9",X"06",X"8D",X"EE",X"02",X"A2",X"00",X"8A",X"9D",X"00",X"02",X"9D",X"00",
		X"03",X"E8",X"D0",X"F7",X"60",X"B9",X"44",X"00",X"0A",X"A8",X"D0",X"0D",X"A5",X"42",X"25",X"43",
		X"30",X"07",X"A2",X"B0",X"A9",X"56",X"4C",X"18",X"7A",X"4C",X"F8",X"79",X"A2",X"20",X"A9",X"00",
		X"85",X"19",X"BD",X"00",X"02",X"D0",X"04",X"CA",X"10",X"F8",X"60",X"10",X"63",X"20",X"B6",X"70",
		X"4A",X"4A",X"4A",X"4A",X"E0",X"19",X"D0",X"07",X"A5",X"76",X"29",X"01",X"4A",X"F0",X"01",X"38",
		X"7D",X"00",X"02",X"30",X"25",X"E0",X"19",X"F0",X"13",X"B0",X"17",X"CE",X"E7",X"02",X"D0",X"05",
		X"A0",X"7F",X"8C",X"EC",X"02",X"A9",X"00",X"9D",X"00",X"02",X"F0",X"CB",X"20",X"1B",X"6A",X"4C",
		X"15",X"67",X"AD",X"E9",X"02",X"8D",X"E8",X"02",X"D0",X"EB",X"9D",X"00",X"02",X"29",X"F0",X"18",
		X"69",X"10",X"E0",X"19",X"D0",X"02",X"A9",X"F0",X"A8",X"BD",X"A5",X"02",X"85",X"05",X"BD",X"63",
		X"02",X"85",X"06",X"BD",X"C6",X"02",X"85",X"07",X"BD",X"84",X"02",X"85",X"08",X"4C",X"E5",X"67",
		X"85",X"1B",X"06",X"1B",X"10",X"15",X"E0",X"19",X"B0",X"11",X"29",X"3C",X"4A",X"4A",X"A8",X"84",
		X"1C",X"B9",X"F8",X"02",X"85",X"1D",X"30",X"03",X"20",X"BE",X"48",X"A0",X"00",X"18",X"BD",X"21",
		X"02",X"10",X"01",X"88",X"7D",X"A5",X"02",X"9D",X"A5",X"02",X"85",X"05",X"98",X"7D",X"63",X"02",
		X"C9",X"20",X"90",X"2A",X"E0",X"1A",X"D0",X"06",X"20",X"EB",X"67",X"4C",X"E7",X"66",X"24",X"1B",
		X"10",X"1A",X"A4",X"1D",X"30",X"16",X"C0",X"04",X"B0",X"12",X"CE",X"E7",X"02",X"CE",X"FF",X"02",
		X"A4",X"1C",X"A9",X"00",X"9D",X"00",X"02",X"99",X"F8",X"02",X"F0",X"DF",X"29",X"1F",X"9D",X"63",
		X"02",X"29",X"7F",X"85",X"06",X"18",X"A0",X"00",X"BD",X"42",X"02",X"10",X"01",X"88",X"7D",X"C6",
		X"02",X"9D",X"C6",X"02",X"85",X"07",X"98",X"7D",X"84",X"02",X"C9",X"18",X"90",X"08",X"F0",X"04",
		X"A9",X"17",X"D0",X"02",X"A9",X"00",X"9D",X"84",X"02",X"85",X"08",X"BD",X"00",X"02",X"29",X"03",
		X"A8",X"B9",X"0C",X"68",X"A8",X"20",X"A8",X"6B",X"4C",X"E7",X"66",X"AD",X"E9",X"02",X"8D",X"E8",
		X"02",X"98",X"48",X"A0",X"17",X"20",X"0D",X"77",X"68",X"A8",X"A9",X"00",X"8D",X"1A",X"02",X"8D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
