-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_1N is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_1N is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_1N_0 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000037CEF4D74C31FFEFB9EB9E76D37DB",
		INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => x"D2BF7851D567979A7195052467C145E697B190517FC5F1FF5B2B5BCAF0564694",
		INIT_03 => x"9A991250425E2479969F15B679679A72925925EA662C675D92EC76BD3E5D2BB1",
		INIT_04 => x"5557263777774B67E2491767FFFF24911662481552595CB89B4952055555D510",
		INIT_05 => x"129CB5FC820209CDF2755D732720AD4F2556BC8CB49C85D40B943CE9B3A30955",
		INIT_06 => x"04107B9CB5C8041241C51049071625489A762D89AE995740169CB5FC82020BD0",
		INIT_07 => x"F2FD9156F0F55B73DCF73DCF749F9A55558A2F44104172268D65559800000000",
		INIT_08 => x"814555754BD2024B082691B60669142C2B52E54ACEFD029616C3E6839AF2BF2B",
		INIT_09 => x"3984641282825A8915635502528D08A0A8A6041226D49B50B58A8B5860B582E3",
		INIT_0A => x"849649088255542E084927508D28D08D2BD1241E4220955554C2453984641504",
		INIT_0B => x"E24176CDB76CDB505DB36DDB366D572495269651AA226A2E6A8D555555E482E0",
		INIT_0C => x"8DC3884CD5FC04048D83884CD5FC04048D43884CD5D555509191909549A59090",
		INIT_0D => x"05557915791579157915793D91103B7F37011155DB3C04048D83884CD5FC0404",
		INIT_0E => x"FCC4C484855555042F0825665224A467543895C3756289355555556E92D8E18E",
		INIT_0F => x"22DE10878B694260420209AE89E7807230927E827878E4A464276425AE8E6917",
		INIT_10 => x"00109A2190919095C15909D989549E69481078A25958B6858926C040406B7819",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"3131313131313131000000F020202020202020202020202000000088003E8355",
		INIT_15 => x"000000000000000000000000000000000000000000000000000000F131313131",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"7142209AAA8A49429AA6021202120A2BA461768AAA9116765446745547656220",
		INIT_1B => x"00000000000000000000F468A04802409AB246465021202120212064858A802B",
		INIT_1C => x"666666666099AAAAAAAAA999AAAAAA999998030499998881477722A666666665",
		INIT_1D => x"000000000000000F405163204666B0B999905622128BBBBBBBBBAA9655320904",
		INIT_1E => x"404191222122212221222042020845555202846402804666666666666666666A",
		INIT_1F => x"0000000F40805555550899999999999926023AA02040AAAAAAA224248AB220A8",
		INIT_20 => x"FDFDFDFDFDFDFDFDFDFAFCECECECECECECECECECE94444444000000000000000",
		INIT_21 => x"CCEBFDF0232132012120CDFAFCE0CCE9FDF0021003301211310DF8FCE0CCEBFD",
		INIT_22 => x"E9FDF0CDF8FCE0C460ECEBFDF0CDFAFCE0075676045575470CE9FDF0CDF8FCE0",
		INIT_23 => x"E6FCCCCD0FFCE688888444FDFDFDFDFDFDFDFDFDFDFAFCECECECECECECECECEC",
		INIT_24 => x"000000000000000000000000000B6FFCCCCD0FFFE6FCCCCF0FFEE6FCCCCE0FFD",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"576767640EEEEEEEEEEF567676764AF57647F5767648F57643F56767644CCCCE",
		INIT_27 => x"20020F576767643F50E53F70E72F60E61F70E70F60E63F70E72F60E61F40E40F",
		INIT_28 => x"0000F76767676767640F63F72F61F70F63F5767642F567676764BF56764C2020",
		INIT_29 => x"40C5767648F5767660C776764BF70C7EF60C6DF70C7CF60C6FF40C4E44444000",
		INIT_2A => x"567646F57640D57640D576444444F50C5DF70C7CF60C6FF70C7EF60C6DF57676",
		INIT_2B => x"767640C5767642F576488844F567640C567646F57640D57640D57644F567640C",
		INIT_2C => x"C567644AAAF567640E56764BF567640E56764888F5764BF5767640C5767641F5",
		INIT_2D => x"72F60E61F57676767676767640CCCCCCCCCC888F57640E57647F57648F567640",
		INIT_2E => x"F57648F50E53F70E72F60E61F70E70F60E63F70E72F60E61F70E70F60E63F70E",
		INIT_2F => x"7676767649F5766AF79F68F5676764FF57668F7BF6AF56492020200CCECEECEC",
		INIT_30 => x"7649F5767640C576764B000F5766AF79F68F56767676767647F7BF6AF57668F5",
		INIT_31 => x"2F60E61F57640F56767676406666666666666220F567640C567647F567640E56",
		INIT_32 => x"70E70F60E63F70E72F60E61F70E70F60E63F70E72F60E61F70E70F60E63F70E7",
		INIT_33 => x"F576767676418A88888A88888A88888A84F7676767640F57663F70E72F60E61F",
		INIT_34 => x"0E65F70C74F60C67F70E56767646F69F78F60C57F70C66F60C75F40C64F77F66",
		INIT_35 => x"40CCCCC8F5767676766AF69F78F60C57F70C76F60C65F40C74F67F76F7676764",
		INIT_36 => x"450000000CCCCCCCCCF576764BF5767640F5767649F5767642F576764BF57676",
		INIT_37 => x"0C7CF60C6FF40C4EF50C55F60C64F70C57640C77F60C66F40C45F567640C5676",
		INIT_38 => x"002020F567640C567646F50C56F60C65F70C57640C74F60C67F40C46F50C5DF7",
		INIT_39 => x"94C3595A3594E0D65A0D6510D650435959403595E3596E3595C3594575202313",
		INIT_3A => x"0000000000000000000000000000000000007164C3594A0D6590D6500D653235",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000E00",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1N_1 : RAMB16_S2
	generic map (
		INIT_00 => x"000000000000000000000000000000000001061841851860C20410C008104100",
		INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => x"0C3C92975E5DFA7BF7DE2081CD8001DFF013A421000CC30020FE200FA1196088",
		INIT_03 => x"709FC975C9CE7F18F334A211DF5E7BF9F5E7BC033C84EB10C63DC20C430060D7",
		INIT_04 => x"00CF1C8CCCCCF1FBD3C681FBEEEE3C680C6B8D0CD3C7BC5C7E04C2A377565D72",
		INIT_05 => x"88EC40FE46A30A4313CCD4190D28342528008434907480420F50B82011910956",
		INIT_06 => x"8C0C24EC40668F01C0403C0701071F084E08B08E410D580188EC405446A30901",
		INIT_07 => x"5B14CC005BD309AA6A9AA6A9539F4E5D690F060C0C304639A668090E22222220",
		INIT_08 => x"9B5E033F81A2873B0CA021D527081DA42B3720DA4631638CCEEAD38BCE53C53C",
		INIT_09 => x"071D1C35072385E50DE09B4BA0E20CE30CC300F30D8C36366343E6343A634310",
		INIT_0A => x"8CC430806256020D88C4E3CE2CD0CD0CC3C3220E241995803A53DB071D1C3B21",
		INIT_0B => x"F7D71F07C1F07CB407C1F07C1F90AB138D3CF1D0D237D033D24B775580DCE4D9",
		INIT_0C => x"01030C8C123C484401030C8C123C484401030C8C12200330707070734F3C7172",
		INIT_0D => x"01557FD56A9555554015403DD55C3F3BB741599199FC484401430C8C123C4844",
		INIT_0E => x"FC0000000200331C00081D03D03C1C1DCF3CFB42DCDBCF33775581079078000C",
		INIT_0F => x"6A10C8F4A8432BDBABE1AD278D2826D198E1F72B23285C5C5C5E1E1E0FEF890F",
		INIT_10 => x"002220307070707B50C7C7C7C734F3C74003FE83939A84290E4372DAEA49898E",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"7665544776655447000000F776655447766554477665544700000088006083D5",
		INIT_15 => x"000000000000000000000000000000000000000000000000000000F776655447",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"8144405444448B004422001000100B044441542424508805555645111005431A",
		INIT_1B => x"00000000000000000000F4444644400854180000100100010001094745440228",
		INIT_1C => x"4444444442554444444445554444445155522004555544404444303754444444",
		INIT_1D => x"000000000000000F00B140002444000155535460086444444444445455000104",
		INIT_1E => x"3129910001000100010000004080455550400046400004444444444444444446",
		INIT_1F => x"0000000F00885555552455555555555507408644001044444444300000454882",
		INIT_20 => x"B8888888888888888886FBB8888888888888888886233112220001123AAAAAAA",
		INIT_21 => x"C997FBB0300330010210D997FBB0C997FBB0031113101131320997FBB0C996FB",
		INIT_22 => x"95FBB0C995FBB0D770E994FBB0C994FBB0045774074645440994FBB0C994FBB0",
		INIT_23 => x"CBFCCCCC08FCCB13311331FAAAAAAAAAAAAAAAAAA995FAAAAAAAAAAAAAAAAAA9",
		INIT_24 => x"000000000000000000000000000788FCCCCD08FCCBFCCCCC08FCCBFCCCCC08FC",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"88888888E0123012303F8888888882F88885F888888DF8888AF8888888212232",
		INIT_27 => x"47756F88888888DF90F98F90F98F90F98F90F98F90F9BF90F9BF90F9BF90F9BF",
		INIT_28 => x"5674FA8888888888889F94F94F94F94F97F88888A7F88888888B2F88888E6576",
		INIT_29 => x"A0EA888885F88888A0EA888886F90E9AF90E9AF90E9AF90E99F90E9974567774",
		INIT_2A => x"88888BF88880D88880D888865454F90E9AF90E9AF90E99F90E99F90E99F88888",
		INIT_2B => x"888880D888888BF8888E5556F888880D88888AF88880D88880D88885F888880D",
		INIT_2C => x"D88888A674F888880E888885F888880E88888645F8888DF8888880D8888888F8",
		INIT_2D => x"9AF90F9AFA88888888888888AA5674567456747F88880F88885F8888DF888880",
		INIT_2E => x"F8888DF90F98F90F98F90F98F90F98F90F9BF90F9BF90F9BF90F9BF90F9AF90F",
		INIT_2F => x"88888888ACF888AFF9FF9FF888B888AF888AEF9DF9DF88AD98AB989746545464",
		INIT_30 => x"8884FB888880C88888B29AAF888AEF9EF9EF888B8888888885F9CF9CF888ADF8",
		INIT_31 => x"AF90F9AFA8880C88888888AAAB89AB89AB89AB88F888880D888889F888880E88",
		INIT_32 => x"90F99F90F98F90F98F90F98F90F98F90F9BF90F9BF90F9BF90F9BF90F9AF90F9",
		INIT_33 => x"FA8888888889A8B89AB98AB8A8B89AB98AFA888888880C888A9F90F99F90F99F",
		INIT_34 => x"0F94F90D94F90D97F90F888888A7F9BF9BF90E92F90E92F90E92F90E92F91F91",
		INIT_35 => x"8ABBBBBBF888888888AEF9EF9EF90E95F90E95F90E95F90E95F94F94FA888888",
		INIT_36 => x"89EFCEFCDAB89A89ABF88888B1FB888889F88888B0FB88888BF88888B2FB8888",
		INIT_37 => x"0E98F90E9BF90E9BF90D97F90D97F90E88880E96F90D96F90D96F888880D8888",
		INIT_38 => x"CFCEFDF888880D88888AF90D95F90D95F90E88880E95F90D94F90D94F90E98F9",
		INIT_39 => x"3843F3B43F381CFCE10FCE50FCE163F3B3B63F3A13F3A23F3903F3EFCEFDEFDE",
		INIT_3A => x"000000000000000000000000000000000000B3B8B3F3860FCE6CFCE20FCE083F",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000C00",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1N_2 : RAMB16_S2
	generic map (
		INIT_00 => x"000000000000000000000000000000000002092C928A24B2C928A2C820A2CB20",
		INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => x"A3E5D70D351454514D35064BCB8601145B30C501157A8E55A63EA2AFA00014E0",
		INIT_03 => x"D80DD4D3476837B5D36C5932C924514492451613760C32A0E974A9FA0B9296D2",
		INIT_04 => x"1A6F3C6EEEEE43F5234423F5CCCC34423EC7C02E6249544CC780CB29B99034D1",
		INIT_05 => x"4BD4620187233CD9B36660803C3CF08C306EC0F0FCC0C009AFBEB07A31DB3F90",
		INIT_06 => x"7843665462067813044BE24C112F332C07A9391C395E40004BD46A0287233C00",
		INIT_07 => x"E3B8C60EA3A33B4CD334CD3312F48766C0CD38F8074EEC70CC3060CDD951D951",
		INIT_08 => x"E4A0E9540C03332C8C33FCE1B33F120CF09B0A6CCB8123CBCB4B21DBCBE0EE0E",
		INIT_09 => x"8D3634DC23E3E820266028A7E8F38CB0CCB300CB12A44891A923189235A92321",
		INIT_0A => x"F804810CC390183E0F8004A08208A08208EE00118B32E406918B050D3634D504",
		INIT_0B => x"734D3F8FEBFAFE704FE3FAFEBF65AA22EE101048E833683368C1B9930630CBE2",
		INIT_0C => x"40C300000C7C400040C300000C7C400040C300000C4C69B2F2F0F0FB840410DB",
		INIT_0D => x"0AD55555555555555555403C804000000040CCCCCC7C400040C300000C7C4000",
		INIT_0E => x"FCCCCCCCCCC69B34AA283433C33C3436ACBCF7C9AAFCCD19B993383AC3ACA286",
		INIT_0F => x"3B07CBF1EC1F2FC72FCDBC7B3C70FD04C8F403331F1C3434343435343FEF0C67",
		INIT_10 => x"0000C332F2F0F0F7C12F2F0F0FB8404118231EC30F0EC1F0FC330BCBCB1C0E8C",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"7777777666666660000000F4444444477777777666666660000000AA00909024",
		INIT_15 => x"000000000000000000000000000000000000000000000000000000F444444447",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"1230433404140214240024041404304343412424340000004040404040440141",
		INIT_1B => x"00000000000000000000F3434111242334200424014041404140424110243101",
		INIT_1C => x"0440404040404040404040404040404040402413404051501040140104040404",
		INIT_1D => x"000000000000000F323041411000014040413424031404040404040404140010",
		INIT_1E => x"0011104040404040404042142422140404241241140300404040404040404043",
		INIT_1F => x"0000000F11110404040140404040404041243040410014040404010114114122",
		INIT_20 => x"15555555555555555110F115555555555555555110EFEDCDCFCDCDCDE0000000",
		INIT_21 => x"D550F550210000001000C550F550D550F550000110000131010550F550D550F1",
		INIT_22 => x"11F550D551F550C330C551F550D551F550011000000000110551F550D551F550",
		INIT_23 => x"30F3333301F330FEDDCFEEF115555555555555555111F1155555555555555551",
		INIT_24 => x"000000000000000000000000000001F3333301F330F3333301F330F3333301F3",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"222222220EDCFFEDCCEF2222222225F22221F2222221F22220F22222224CFEDC",
		INIT_27 => x"CFEDCF222222221F20C21F20C21F20C21F20C21F20C20F20C20F20C20F20C20F",
		INIT_28 => x"FEDDF22222222222221F25F25F25F25F24F2222224F2222222220F222220DDCC",
		INIT_29 => x"20C2222221F2222220C2222220F20C20F20C20F20C20F20C20F20C20FFEDCECC",
		INIT_2A => x"222220F22220C22220C22220FDFDF20C21F20C21F20C21F20C21F20C21F22222",
		INIT_2B => x"222220C2222220F22220ECEDF222220C222221F22220C22220C22221F222220C",
		INIT_2C => x"C222220DCFF222220C222221F222220C222220DFF22221F2222220C2222221F2",
		INIT_2D => x"20F20C20F22222222222222220FEDDCFEEDCFFCF22220C22221F22221F222220",
		INIT_2E => x"F22221F20C21F20C21F20C21F20C21F20C20F20C20F20C20F20C20F20C20F20C",
		INIT_2F => x"2222222221F22220F20F20F22222220F22220F20F20F2220CCFDDDCEEDDCFFEE",
		INIT_30 => x"2221F2222220D2222220DFDF22221F21F21F22222222222221F21F21F22221F2",
		INIT_31 => x"0F20C20F22220C2222222220DCCFEDDCFEEDCFFDF222220C222221F222220C22",
		INIT_32 => x"20C21F20C21F20C21F20C21F20C21F20C20F20C20F20C20F20C20F20C20F20C2",
		INIT_33 => x"F22222222220DDCCFEDDDFEECCFFEDCCCEF2222222220C22221F20C21F20C21F",
		INIT_34 => x"0C21F20D21F20D20F20C22222220F24F24F20C24F20C24F20C24F20C24F24F24",
		INIT_35 => x"24CFEDCFF22222222221F21F21F20C21F20C21F20C21F20C21F21F21F2222222",
		INIT_36 => x"20DCCEDDCFEEDCFEDFF2222221F2222225F2222221F2222224F2222220F22222",
		INIT_37 => x"0C21F20C20F20C20F20D20F20D20F20C22220C20F20D20F20D20F222220C2222",
		INIT_38 => x"CFFEDDF222220C222221F20D21F20D21F20C22220C21F20D21F20D21F20C21F2",
		INIT_39 => x"C1C03C0F03C0380F03C0F0340F00C03C3C0F03C0F03C0D03C0C03CEDDCFFEDDC",
		INIT_3A => x"0000000000000000000000000000000000000C31D03C03C0F07C0F07C0F00D03",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000F00",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1N_3 : RAMB16_S2
	generic map (
		INIT_00 => x"000000000000000000000000000000000001B4DF6D74DF5DB6D37DB6D36D74D3",
		INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => x"1BA659C71C1C7071C71C017E5EC0231C75EA3CC0002D3B004C344C0D0030824C",
		INIT_03 => x"34CB4071C0DF2D7CB07807E3071C71C071C71DF31D3A8E6C1B95C6E9B16DB857",
		INIT_04 => x"FFFF0F0CCCCCC1D131C3C1D133331C3C1D73428FF1C73424FC0028C3FFFF1C70",
		INIT_05 => x"28441000E00393C311CFF81E0208183A0FFDB8081CF800800DFC1E06E80293FF",
		INIT_06 => x"2C093444188C2E83C0E3BA0F030D3CA00C1736CE86CFFC0028441001E0039000",
		INIT_07 => x"491268E84949A2338CE338CEDA34E8FFFA020FEC4924DB3A3A8FFA0377773330",
		INIT_08 => x"1F4FFFDF83E003A00E8A30C303A33D7A4D34F4D3A07C036828423A03E8434434",
		INIT_09 => x"031C0C78030340220FD3D7C770D30E4A024000F03D8CF6305303053030430338",
		INIT_0A => x"2C0D2482E0FFFE0782C090890090890090CB020024B93FFFFC6003431C0C7300",
		INIT_0B => x"31C31D074DD374300741D374DD1C010A3F3C71D0D331D331D34FFFFFFF7C2479",
		INIT_0C => x"44030444403C444444030444403C444444030444403FFFF33330303FCF1C7030",
		INIT_0D => x"03C02A802A802A802A802ABC0444044444400000003C444444030444403C4444",
		INIT_0E => x"FC00020003FFFF0E80A00E01E01C0C0D4C3C73A9D4C0C7A3FFFFFE0520528A28",
		INIT_0F => x"05E003C81780070007001E07FE081C1340D01003A0A00C0C0C0C0C0E0C0F820F",
		INIT_10 => x"003A2003333030338033330303FCF1C78003C17380817818020042020281800E",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"0000000000000000000000F111111110000000000000000000000054007C43FF",
		INIT_15 => x"000000000000000000000000000000000000000000000000000000F111111110",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"1001010000001000000010000000000001000000001001000000000000000000",
		INIT_1B => x"00000000000000000000F0000000001000011000000000000000000000000201",
		INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => x"000000000000000F010000010000000000000000000000000000000000101112",
		INIT_1E => x"0100000000000000000000000000000000000000001010000000000000000000",
		INIT_1F => x"0000000F00000000000000000000000000000001001100000000000000000000",
		INIT_20 => x"00000000000000000000F0000000000000000000006555544777766540000000",
		INIT_21 => x"C000F000011111011110C000F000C000F000011111101101110000F000C000F0",
		INIT_22 => x"00F000C000F000C000C000F000C000F000011111011111110000F000C000F000",
		INIT_23 => x"00F0000000F00044444777F000000000000000000000F0000000000000000000",
		INIT_24 => x"0000000000000000000000000000A0F0000000F000F0000000F000F0000000F0",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"1111111107776666665F1111111110F11110F1111110F11110F1111111054444",
		INIT_27 => x"54444F111111110F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F",
		INIT_28 => x"6666F11111111111110F10F10F10F10F10F1111110F1111111110F1111105555",
		INIT_29 => x"10C1111110F1111110C1111110F10C10F10C10F10C10F10C10F10C1044444777",
		INIT_2A => x"111110F11110C11110C111106655F10C10F10C10F10C10F10C10F10C10F11111",
		INIT_2B => x"111110C1111110F111104477F111110C111110F11110C11110C11110F111110C",
		INIT_2C => x"C111110665F111110C111110F111110C11111054F11110F1111110C1111110F1",
		INIT_2D => x"10F10C10F111111111111111105555544444777F11110C11110F11110F111110",
		INIT_2E => x"F11110F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C",
		INIT_2F => x"1111111110F11110F10F10F11111110F11110F10F10F11105544444777776666",
		INIT_30 => x"1110F1111110C1111110655F11110F10F10F11111111111110F10F10F11110F1",
		INIT_31 => x"0F10C10F11110C11111111106665555544444777F111110C111110F111110C11",
		INIT_32 => x"10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C10F10C1",
		INIT_33 => x"F111111111107777666665555544444447F1111111110C11110F10C10F10C10F",
		INIT_34 => x"0C10F10C10F10C10F10C11111110F10F10F10C10F10C10F10C10F10C10F10F10",
		INIT_35 => x"10544447F11111111110F10F10F10C10F10C10F10C10F10C10F10F10F1111111",
		INIT_36 => x"105554444777776665F1111110F1111110F1111110F1111110F1111110F11111",
		INIT_37 => x"0C10F10C10F10C10F10C10F10C10F10C11110C10F10C10F10C10F111110C1111",
		INIT_38 => x"766666F111110C111110F10C10F10C10F10C11110C10F10C10F10C10F10C10F1",
		INIT_39 => x"3C63D3C63D3C14F4F10F4F1CF4F053D3D3C53D3C73D3C53D3C43D34444777777",
		INIT_3A => x"000000000000000000000000000000000000DF0C53D3C1CF4F18F4F18F4F053D",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000F00",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
