-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu1 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "8E55537FC8E55FFFFFFFFFFFFFFFFFFF4355F5C5FFFFFFFFFFFF510FF7EEF6C1";
    attribute INIT_01 of inst : label is "559D156E7B45555556EFDEB6CC2109B082C6CDBC2CA114D24BCC68CADD54234B";
    attribute INIT_02 of inst : label is "A52B10812AD4449744D3585134D5D2CFFC8A12F45066206C259D156E7B455555";
    attribute INIT_03 of inst : label is "A101101000001007C29D88652913A1CE10AA82EC1BA2B3B9A466495752FF0BB2";
    attribute INIT_04 of inst : label is "9090AD2B31304D6F834008B041A919C955C71220412023207BBB81EEEE0463BB";
    attribute INIT_05 of inst : label is "43C4C135BC84C4C119090FB05850F2E22C8185058FE22C81E1909A999C9C4C11";
    attribute INIT_06 of inst : label is "B20483EC16143CB88B20614163F88B2078782548AC4DF9504DD2C521F452055C";
    attribute INIT_07 of inst : label is "4C95375C0ACA52650D3244FB106A18132571D74513113C4EBE122C81C444CF08";
    attribute INIT_08 of inst : label is "AE806BC6175545D5055367237B95EEA50F35085346609D527509D05C5323BD83";
    attribute INIT_09 of inst : label is "0B030B030B030B021E1A16121E1A16127A7132363070D370AE1B3C9D55553550";
    attribute INIT_0A of inst : label is "4E242C2EB57C341811F9B7131313030303030082C6CACEC2C6CACEC2C6CACEF3";
    attribute INIT_0B of inst : label is "35DD05D068586F3416E0B08244BD8C952150554932F27FB7222E4512A245A309";
    attribute INIT_0C of inst : label is "E69556C553DA55055FF0A452FFD55752C9573B082E7A339E843DDDCC80C26797";
    attribute INIT_0D of inst : label is "3083E8227C7783A8934561A23268AFCB3C2672EFBEFBC9289624A62508B08382";
    attribute INIT_0E of inst : label is "B354294F2B9B69D049E47D374BD2C1208A5943FEBEFD5309B4918E4924496492";
    attribute INIT_0F of inst : label is "114B1041177BC381B914BD1FDEFD1FD555D4209557D555F7122041C48D245D52";
    attribute INIT_10 of inst : label is "9A98A9813BFC53626A62A6971757D79714D89A98A9BBFC4884040544FA811488";
    attribute INIT_11 of inst : label is "D41D41D41C4777714D89A989DDDC53626A624044C04C04C048971757D79714D8";
    attribute INIT_12 of inst : label is "3EBBB945D0763E97BBB98F838F50F6E7D094DAC5F62DF601F43C214D89A9899D";
    attribute INIT_13 of inst : label is "5F5553AAAAAAA70D55531131432C90BE43FB896459B2D59AC1C5565054173256";
    attribute INIT_14 of inst : label is "2391757D72E69C99518659018E7929A7E7E3FFD6D2FCA0089FCF24FFF0FFF955";
    attribute INIT_15 of inst : label is "452DF75F729BDCC96475F729FBDD4C96791D7B972508990239175EE1C9588998";
    attribute INIT_16 of inst : label is "9E400000000000000000FFFEE7B7C00000D81C0BE4BFFFF73DB419414BFE52D6";
    attribute INIT_17 of inst : label is "ADB7D9EE400000185858BD7BB92F5A588A3D888A0089011A6E24BC9941719C34";
    attribute INIT_18 of inst : label is "154BED5C64D924BF229072151692248104224890492371DBA2685C7ADB2CB6CB";
    attribute INIT_19 of inst : label is "DF5A235D955955176C5F42E34234CA725645C6A5E654754959A929798949D949";
    attribute INIT_1A of inst : label is "E63723532AAE251463BB888E01E3B6426F1BE59741164123525DF798DD955995";
    attribute INIT_1B of inst : label is "7EA04228D7082020B28256D8A0A35C8D982D5B5D55956156D561B17DA0A820B6";
    attribute INIT_1C of inst : label is "9449C65246426F1BE5977DE6DEE48A0BF48934D7DA04228D0565F4893694934D";
    attribute INIT_1D of inst : label is "1E9022AA4DF6D74DF58618D88DDA37E8D998B323A9444EA51316E93A948C1A7A";
    attribute INIT_1E of inst : label is "CB0450F3B58B8C94B0796E6B923822BE612C854410B8810612C8904F63C8F26C";
    attribute INIT_1F of inst : label is "22B2934BA509EA06FDCC2D509BC6F965DF79B4A35198D561CF0A5F493C2F43B5";
    attribute INIT_20 of inst : label is "6CB8D84163CD8B2696472A9755A65F7845D0B1349DD195715158F556D5150B68";
    attribute INIT_21 of inst : label is "C900D32E95FCEE4A42E9C953A4A18275DCE6514A49793587E695357B7AA2EE81";
    attribute INIT_22 of inst : label is "9C4992BB90D4992BE53E24A6EA4B16326D2049D19154A49CCB58992545275294";
    attribute INIT_23 of inst : label is "2BB90690154899715415355FAD6E7A5F584527452D3FF641114505B4264BB789";
    attribute INIT_24 of inst : label is "34894BC7EB053D43D73D63C44C171D075DADD562458556A576AC44530815FC69";
    attribute INIT_25 of inst : label is "3609919B46F5BE5414E42685C55134D22420464E4A63423509D45D4DD45D4D19";
    attribute INIT_26 of inst : label is "E92E22508902249574861408D350991B2352F3CC822955B16D0FCAA35555D185";
    attribute INIT_27 of inst : label is "A7587E6915056490AC5B5628DD151496436328DD0545259908BFCAC12255F93C";
    attribute INIT_28 of inst : label is "535585235A24626141561CF69CDAE712FE9D1FF29A4B770A6510163523579B76";
    attribute INIT_29 of inst : label is "7A87203A9C2CACB279470A08294D9C4663A50C0F199CBF2255079C8DE5415558";
    attribute INIT_2A of inst : label is "A7507E49870AD524BFC86E72B6DBF52367B85C5B59CDBF6B954BFF2A5CD66FD6";
    attribute INIT_2B of inst : label is "C5C738E89E7199FF22767254D5552356D65D24DA7D64296423609E65CE9561D9";
    attribute INIT_2C of inst : label is "E792FE26DB76D55E7DA7FE69550428D5973A61B6FD91C2820A53A71298E94303";
    attribute INIT_2D of inst : label is "2F4DE7C9E7A69CE7FF672EE7D427B954DE6D67B6E3ED823423774DBB5DBF6CDA";
    attribute INIT_2E of inst : label is "41EEBCB898CB8982250B0998BF53A739FF67CB89F62752DBF52367BB2F674276";
    attribute INIT_2F of inst : label is "66D67F727AEDFFE4AF72795379E76A595C4BBFE25E887E230BB9024202089625";
    attribute INIT_30 of inst : label is "04DAEBC8093912D2CE9D751BAF1342EBC8E7C39E4A43E7E9F27944249053CFCF";
    attribute INIT_31 of inst : label is "C252B8907358D4AB65485C672794941555E7D61E69098550428D8D0E245EEBCA";
    attribute INIT_32 of inst : label is "519549D6179A55EEEE792FEB5976FD3CDAD67FA59CB59FDAE712FE9D1FF29A4B";
    attribute INIT_33 of inst : label is "EA69B6D427E672369B6D7FD0A9C51B3E50B89634635895054562356D50FC5255";
    attribute INIT_34 of inst : label is "509EC8E150936612FB893236F9D5CC9A60B9AD4276723A69B6D88D424E7E6723";
    attribute INIT_35 of inst : label is "4E1E138DDDDDDDDD7923789089182255552F89F41FFD24C2FD378F8694D2FEE2";
    attribute INIT_36 of inst : label is "9160734B1433491C13C91A08E28608E28608E28608E28608E28401C1FFDCCC78";
    attribute INIT_37 of inst : label is "BA0B7456A956000BDA98B700C52980B7A6741567001155B9977622C888AA8AC4";
    attribute INIT_38 of inst : label is "000AC98BA563F0450009D8B3A6984522E3F000C1D222E3F0000000FB05675270";
    attribute INIT_39 of inst : label is "56700BA2984567000BC33A98B7452956840B732E02EA984595840B74560003E7";
    attribute INIT_3A of inst : label is "0452670B7A62918BA674526000AD947452E3F000C1D222E3F0000000F0BA6374";
    attribute INIT_3B of inst : label is "8B7BA9522E3F000C1D222E3F00000F00B333337456A95670000FBA222958BA67";
    attribute INIT_3C of inst : label is "57539A747344F3E88B63E88B6788048BA956700B3A95B3F6700A684A6567BA26";
    attribute INIT_3D of inst : label is "8A00654380B2D8ADB4F1C75915490A280D507E1C724495345E700000B95A68B7";
    attribute INIT_3E of inst : label is "63F0B79580452E3370B84BA2E4637000B7A9526700B7A918B7041152E370BA91";
    attribute INIT_3F of inst : label is "D089A766548AD8F9653E5C3F891A265478F91BE85447EC39CA850F50FB890075";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "427003FFC4255FFFFFFFFFFFFFFFFFFF0C55F400FFFFFFFFFFFFA3C1FA13F330";
    attribute INIT_01 of inst : label is "000044000010000009B84104E42112D8446BA48C64E612A30764DC42680023C7";
    attribute INIT_02 of inst : label is "83200210118CCC830C001C43000801CDFC4231F0000A10242000440000100000";
    attribute INIT_03 of inst : label is "E03030704000001082710C4884000024080F0F1E03CBD3073CC1CFB331D53070";
    attribute INIT_04 of inst : label is "79702B9EE0A0171B4A87347000478787330E2110003A3C50377740DDDD026EF1";
    attribute INIT_05 of inst : label is "0082805C7F76828057978F6C70F803D13840C74F81D13840F575747878782805";
    attribute INIT_06 of inst : label is "E540E3DB1C3E0CF44E5031D3E0744E503DDED3A2BB0B5F480B514D33F0010271";
    attribute INIT_07 of inst : label is "C667417D96926CF2031D8280000487B1D9C05F4D1E3C002DDDD13950C74F81C4";
    attribute INIT_08 of inst : label is "3DD61F4202325897E1D93DB2C4CD13136E1309C2C1D9CB652D5CB034558EF880";
    attribute INIT_09 of inst : label is "969E929A9E969A91D5D9DDD1D1D5D9DC8986828A890402D43D0AA235031B2D7C";
    attribute INIT_0A of inst : label is "2703BB3BCB4747D7170D88545C545C545C545C5155595D55595D51595D51554E";
    attribute INIT_0B of inst : label is "0CAA00600E0A0F9800E0C8C1CC7564F5DA30188731B58000953901F313029909";
    attribute INIT_0C of inst : label is "3C78CB803430C30CBD60FA81FFED8EA1C75D37A4B5F5DA7C782FF7F4ECC27C7B";
    attribute INIT_0D of inst : label is "10ABD231C2DF228C73009BF139F2FFE6B097D1EBAEBA832A3A8CA80D0788728A";
    attribute INIT_0E of inst : label is "16AD1A803866DEF1CF5A1B0047CB807842276297B100710A6B41278019801B41";
    attribute INIT_0F of inst : label is "0BD40008BD48F9904E9076B03403C029E76210AF9DCBE7422110004C48A285E1";
    attribute INIT_10 of inst : label is "4958549100CC52612561522161612161149849585480CEE22AAA268281CCBC4C";
    attribute INIT_11 of inst : label is "D915915914133331498495851DDC526125610570130130130421616121611498";
    attribute INIT_12 of inst : label is "00C44ECCA02200D4C44ECE0263D880D799D4F5C411841388123821498495840C";
    attribute INIT_13 of inst : label is "FFFFF9555F555406AE000100A2515B49E984CF5833ED1A71C4327920C802055A";
    attribute INIT_14 of inst : label is "B0F02763591E7E5FA705DF2701CF073ED85A942A01FE498E66EE3FAAA0AAAAFF";
    attribute INIT_15 of inst : label is "801EFA78D92EAEA47C278D92AC2D6A47C709F37D1D2A66AB0F027CDF4752A668";
    attribute INIT_16 of inst : label is "F1C00000000000000000DC7FFFE7C00000E71D8D586AABA0A8E90E8087FEA1AB";
    attribute INIT_17 of inst : label is "413B1F43DAEAA2A806C46F4CC55824C5C5B84C64A8E5B724D3187F61C5C734ED";
    attribute INIT_18 of inst : label is "33048071487EF07510AC9931C514DE48710DE48437D20C20CDC4410820800410";
    attribute INIT_19 of inst : label is "34CE32EC79F09F48D804C0F2D32C7E95C1C3CE9C5D34E007372757070727D717";
    attribute INIT_1A of inst : label is "AF2D32D1FB013CA16EF1D824B7BD2281F84E22BBF3320C1201E34DECBC79F00E";
    attribute INIT_1B of inst : label is "D471003CB8842A1098C69F063192E14B04E27C239F09F49F09FC601330142008";
    attribute INIT_1C of inst : label is "99116C8F9381F84E22BBD379B77EC8034DF3EC4D4710034B29FC4DF3EC4F3EC4";
    attribute INIT_1D of inst : label is "027450A9E75D75D7C30F04B04BE32F04B313B846C9A31B268DBF93EC991A4CAC";
    attribute INIT_1E of inst : label is "E600B6D5BFE6E4FEE01F77FDFF10033AE23A4C722A7E487223A48424A92A4298";
    attribute INIT_1F of inst : label is "909BE12E12075703842461207E1388AEF4DE6ED2EC7CB9F82E0BC4DD982DE9BF";
    attribute INIT_20 of inst : label is "5144C313A0375F100500AEF1271034CCC83563004A71C0B023086D550712013E";
    attribute INIT_21 of inst : label is "5F6821B1308077C5C18B65D97D4A5B6C3C57D78BDF28830E3C732DD6CC0B5162";
    attribute INIT_22 of inst : label is "35D4309DF25D43097C199C25F2C09D9BDB75D430F0F4BDF4E6FD4F53D750D2FE";
    attribute INIT_23 of inst : label is "BC5F00062285F308C90C2D775BB7CC34CCCC12841C157BE3B30421727BC06FE4";
    attribute INIT_24 of inst : label is "DE7F8E108601905904904906251A0A022B923552048E7722EB652803080AD4B5";
    attribute INIT_25 of inst : label is "6CAE70AE5388E30D2C1C1C44137300C130C409C1C1F2F32E071C41C81C01C437";
    attribute INIT_26 of inst : label is "7DBF10106FC93CE39E42AE14B6DAE70B32E106066B9E1EE023805713238E70AB";
    attribute INIT_27 of inst : label is "FE79CBE737DEFF73B808CE8F331C78F1CEE98F33871E3C73387543623337D502";
    attribute INIT_28 of inst : label is "E2074FBAD4747BD3881D324D32793A41DDE77FF1E8075F637D7C9D6C96E37DD1";
    attribute INIT_29 of inst : label is "F7CD199DF81472E7C74D9CBE2785FA45D1BF298905F47F13F3CF82CB42C83774";
    attribute INIT_2A of inst : label is "1D71E7C75D1FB2007FE42FCBEF7C9C1B9F5D71C0C31781E4E707FF1FD079F379";
    attribute INIT_2B of inst : label is "971C28DDF1D05F7F13EDDDEC8377BACC73E7BD73C73E07BC96D077E726F9C7AF";
    attribute INIT_2C of inst : label is "3A01DD3D785E0D76934C07D7975C24B39C9BD7DF27D3672F81E1BE92744FCA62";
    attribute INIT_2D of inst : label is "3AD30C1F1D5FF05D547D1DBDF8FF6F8D30C30C9E1827A12DB2C9E781C785E079";
    attribute INIT_2E of inst : label is "F7D14477FE477F83FCAEB5F8E7C97C17557C477F7F16DB789C1B9F5A9AD6D96D";
    attribute INIT_2F of inst : label is "7C30C5D5F617551C60111359F7D5F3C7A107155FE56695990F6F23E1A384F94D";
    attribute INIT_30 of inst : label is "980104442F9389BF45F5D74411E01104464DE9F58DC97C5F1113423EF9DBA64E";
    attribute INIT_31 of inst : label is "C1D8F4F1F07CB9B6D79275CDBD756C03778D1C73C70A5D75C2CB4B47BE710446";
    attribute INIT_32 of inst : label is "3A12C85D79F5EAB193A01DD0C35E03B97830C03C7E0C30793A41DDE77FF1E807";
    attribute INIT_33 of inst : label is "DFE7BEF81D53D5D27BEF7FC87FDE0F9FD2F4FB2C11CCF302C4972D90366133DE";
    attribute INIT_34 of inst : label is "E07557D5E075FA01D74F15D1545D45F9FAC7EF81D3D5D3E7BEF8CB81CDD53D5D";
    attribute INIT_35 of inst : label is "10104400FA50FA509FF1D4FAD70A93EAAA1F4FB40FC79A4294B16D4268C1D5D3";
    attribute INIT_36 of inst : label is "1010234E34E249289185171C30C31C30C31C30C31C30C31C30C1C040A99A9841";
    attribute INIT_37 of inst : label is "111001111111222141110015111111440001111122006533132003DEEEFCECA4";
    attribute INIT_38 of inst : label is "2221411000040111222141004400000404011515111515122222224000001112";
    attribute INIT_39 of inst : label is "1112211111111122214111110011111155244140240111115555100111222141";
    attribute INIT_3A of inst : label is "1111112555511110000111122214103004040115151115151222222241000001";
    attribute INIT_3B of inst : label is "1000000040401151511151512222241100000001111111122224111111410000";
    attribute INIT_3C of inst : label is "0011100112CC5950055510C1110020C111111221111104011221111001111111";
    attribute INIT_3D of inst : label is "1044A221226A6377783732262226A2233737626210CC00011112222255544033";
    attribute INIT_3E of inst : label is "1512555511115111121550040111122255111111225511110011111511121111";
    attribute INIT_3F of inst : label is "26222A2A22266763B36262552222222216522663B3B62216627B722611224401";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "932C600039393FFFFFFFFFFFFFFFFFFF0C93F312FFFFFFFFFFFF38DBF299F123";
    attribute INIT_01 of inst : label is "0000000000000000023228E3963C8DC4E327385230DC8291853004A30F183010";
    attribute INIT_02 of inst : label is "D4B82B82BB6AF803B80B8E9E02D0A0000393E332188069313000000000000000";
    attribute INIT_03 of inst : label is "40000CCCC4000004C368CEA8882A82282EB72F2BACC9E9892662495291409CA4";
    attribute INIT_04 of inst : label is "D4D031CF7BC00D0F5BDBA120424D4D4D69E3538C890FBEB4BDFDC2F7F7CA4515";
    attribute INIT_05 of inst : label is "80EF003400B5EF004D4D347A7E3DAB844D62A7E3DB844D62D8D8D4D0D4DEF004";
    attribute INIT_06 of inst : label is "31494D1E9F8F66E11314A9F8F6E11314B615461B7D50C05D10C0011E321388C3";
    attribute INIT_07 of inst : label is "DF0C084964685506037CEF2C04844677C30A12269E8F6A32C2C44C52A7E3DBD1";
    attribute INIT_08 of inst : label is "36F62A138ABA08AB134A35B06665999B24AB8CA403C483030CCC38BC89551180";
    attribute INIT_09 of inst : label is "232F2F2B272723202C282424202C2825A266EAEEE84E2433368E6268EB4C41B2";
    attribute INIT_0A of inst : label is "2B8BB3B0E0A022A2222B6C6460606C6C686864676F6B6767636F6F6B6767636F";
    attribute INIT_0B of inst : label is "648802D291015874A58ED8C37801A0D8089C620E54C0EEEE3091C84910C8354F";
    attribute INIT_0C of inst : label is "145253229CD34D35541DF621401626A2BB64CA5571D1C47472CBBBB3B3632493";
    attribute INIT_0D of inst : label is "58E6D338D43E20503B5A00806833357863136C514514D6B960DAE1D88AD8ABEE";
    attribute INIT_0E of inst : label is "A365B8D934030483CFFD88B9880922339344B67860AAB58C46232B6213623621";
    attribute INIT_0F of inst : label is "202404B501550A5264180151C41141820C0868C830210C0B538272F8C086210B";
    attribute INIT_10 of inst : label is "0000040808CC20000000123030303032080000000400CC88800808EF2C2E0041";
    attribute INIT_11 of inst : label is "C040040040033330800000008CCC200000002012012012012230303030320800";
    attribute INIT_12 of inst : label is "65E264A0822765D222645C241A881D2F06F2A0AA7466446A649230800000000C";
    attribute INIT_13 of inst : label is "000000000000005010A6644426BAC7EFCAA64F01941050C0A254C28E008B6B83";
    attribute INIT_14 of inst : label is "F0D184805E04C78D3231CD7231CD0F360E0C0000E0008C9F888C3C0005000000";
    attribute INIT_15 of inst : label is "6E1500401E1E94F9344401E1AE956F8345112DBDAD6F91734D184B6F6B96F917";
    attribute INIT_16 of inst : label is "924000000000000000007CF2FDDB800000CB908D247331188E441C514503A287";
    attribute INIT_17 of inst : label is "38E20D8340F3F0C9200408A26402800700907008D9F8888018045083534D6AD8";
    attribute INIT_18 of inst : label is "E20DA5B000FC280024CD700668E310019A71001884006EBEB11019A3BEBAE79E";
    attribute INIT_19 of inst : label is "400D804CD3063021322023A06A04A70FCFFFBCBCBEFBD42F1F5F1F1F5F0FCF0F";
    attribute INIT_1A of inst : label is "3204A06A9C42340245156D4549454603726C884200E2293A83C400C01CD30660";
    attribute INIT_1B of inst : label is "F878A37013A93224CCE3302338E044814274C38430630630E30AC88038DA38E3";
    attribute INIT_1C of inst : label is "162951954603726C88420030C501678E00CC12AF878A3301930600CC126CC12A";
    attribute INIT_1D of inst : label is "20D224C34D34D34D8D34401E0130044419540149214624851955065216258192";
    attribute INIT_1E of inst : label is "A8890532486828F2C8805004019E78E33530019B50AC019B53001896F5AD6B32";
    attribute INIT_1F of inst : label is "24F2CA44940DDB8B222A3880DC9B2210800C31504CD0130A248C600DA2332A48";
    attribute INIT_20 of inst : label is "FBC0D7B876BC0225AB788CD78C59800F8056EE0298D4C624506322405BA88F2C";
    attribute INIT_21 of inst : label is "8D9DACB05902F3636A10934A36C7C90582234D734D43CD3404194273153FFBF5";
    attribute INIT_22 of inst : label is "C36DC53CD536DC5235903542B41434A34C136D8D4D8734D15306D4B60DB60CDE";
    attribute INIT_23 of inst : label is "CC0D052DA8445485A364409F0C5015800F80AA6A1400037BE02998263354307D";
    attribute INIT_24 of inst : label is "3F8FAC99CC8851851851851A146248024C04C4066AE0C048184461258D214D44";
    attribute INIT_25 of inst : label is "41CC5ACC8B2ECAA754343501999E22D3BAE0834343604A040D60D6096096050F";
    attribute INIT_26 of inst : label is "3CF78A9ABF66341037AB61C4141CC5AD8043AE3C0BEDAC8890DAC34B9040DAD8";
    attribute INIT_27 of inst : label is "3CF3E2CB4F3D1C7BA22426DF9934D4926D95DF99CD351456B850172F3B990762";
    attribute INIT_28 of inst : label is "002B50BCE332BFD80CAD413CF4F5951282CF200ED7853E373CFE3C0F80C0F3E0";
    attribute INIT_29 of inst : label is "DB7CBCBCD2A2B6C249348C4C8D29F167DA349290E8D1C0A34D3402C1114D9B96";
    attribute INIT_2A of inst : label is "64D76259410D3DA8503AB4CB4CDE37AC0D8CD36BEF6F5BD6598500A7EAF0F9F0";
    attribute INIT_2B of inst : label is "8D36826C924E8D00A343435419B93CE5D74D34D34D359D3640C9D34D28D35D89";
    attribute INIT_2C of inst : label is "91200634D535669D0F3D51C70D36A81934A350378DCD231323CA3458D68F24A4";
    attribute INIT_2D of inst : label is "A04D35451704DB400237363586358D24D34D3535454D4B05A0534D575D5355D5";
    attribute INIT_2E of inst : label is "4DF8ECD8D1ED8D37358C88DAC63736D00036CD8D61A054D537AC0D86B0604604";
    attribute INIT_2F of inst : label is "BEFBDBF8D9AFC0BE9673DCEBD36BFAEB1985011340FB03ECDD8D632AC328D103";
    attribute INIT_30 of inst : label is "44138ECDCDDCF4C128D34D0E3BD0438ECF70BCD007E7BEEFB3DCD2BEFBFA0CAC";
    attribute INIT_31 of inst : label is "834DF8D378DC17304D74D35A24940449B99A34D145A834D36A41413334D38ECE";
    attribute INIT_32 of inst : label is "94054134D4516A99995214634D3554B0D4D355145134D4D5952142CD200ED785";
    attribute INIT_33 of inst : label is "23D841C0372360FD841CC00B8F3E8CA3D9D8D0042348D9D14173040892099364";
    attribute INIT_34 of inst : label is "40D383F340D375A1458DE0F40A32A8D634C5DC037360F35841C6810343F2360F";
    attribute INIT_35 of inst : label is "A000600A55550000001368D7C5AC6346AA298DA1200DE3EB8DC4B0AB06E14163";
    attribute INIT_36 of inst : label is "6909128908108204204A238E38E38E38E38E38E38E38E38E38E1A0E077555503";
    attribute INIT_37 of inst : label is "1111111111111111511111111111111111111111110099AB9BA8AA476655446A";
    attribute INIT_38 of inst : label is "1111511111111111111151111111111111111111111111111111115111111111";
    attribute INIT_39 of inst : label is "1111111111111111115111111111111111111111111111111111111111111151";
    attribute INIT_3A of inst : label is "1111111111111111111111111115110111111111111111111111111151111111";
    attribute INIT_3B of inst : label is "1111111111111111111111111111151111111111111111111115111111511111";
    attribute INIT_3C of inst : label is "1111111110441110011110411100104111111111111111111111111111111111";
    attribute INIT_3D of inst : label is "1100222222200220232202222222022222220020214411111111111111111100";
    attribute INIT_3E of inst : label is "1111111111111111111111111111111111111111111111111111111111111111";
    attribute INIT_3F of inst : label is "0222222222220202222020222222222222022202222202220222202202220011";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "E07FF2C03E0FFFFFFFFFFFFFFFFFFFFFC7FFF1E0FFFFFFFFFFFFF0C1FF11F0D0";
    attribute INIT_01 of inst : label is "00000000000000000FFD4514B1044200100B0205078041C30190C3907FFE02CC";
    attribute INIT_02 of inst : label is "1B500500504C2C032C05010B0140C06100E0B03104033A060000000000000000";
    attribute INIT_03 of inst : label is "0080008084200003E07521C00C07080805C00031700027071DC1C733306970C8";
    attribute INIT_04 of inst : label is "3030DF0D3240073702C3082000030303F3C30004004CF40C332230CC88800000";
    attribute INIT_05 of inst : label is "03C9001CC0D0C9000303C4DC0C0C02300410C0C0C1300410C0303030303C9000";
    attribute INIT_06 of inst : label is "10C031370303048C010C3030304C010C30000F0C34DBC3FCDBF00F0B31004070";
    attribute INIT_07 of inst : label is "CD0700F80000000F0F30C9040E00003301CC3EC3030300E353300430C0C0C100";
    attribute INIT_08 of inst : label is "3340382043FFC4FF00C21C13C47F114307734086C0CF4F2D3CB4F43C000003C3";
    attribute INIT_09 of inst : label is "1C18181818181819555555555551515058549414143106F0334230784FC76FF0";
    attribute INIT_0A of inst : label is "09431F1C9454D418181C9D9191919D9D9D9D9D9CD4D4D4D4D4D0D0D0D0D0D0DC";
    attribute INIT_0B of inst : label is "0FCC134000F0C8100C80C1C0EC1B087F063618C313534444C04050B40C430C80";
    attribute INIT_0C of inst : label is "1C7FFFD0F071C71F3680D180400D8F007DFD8DCFF35340D4D0741414D0101C7E";
    attribute INIT_0D of inst : label is "C43170B3431007007534C3485300303C2071D70C30C377537C1D4C1C2E42E514";
    attribute INIT_0E of inst : label is "190553C0E033C0B0C767C750F901D00CE0C3F0122003FC43F10C091C0C1C0100";
    attribute INIT_0F of inst : label is "00C08E330DC042304400180300340330C73334031CC0C733000010EC006183F5";
    attribute INIT_10 of inst : label is "0000040440CC2000000010300000000208000000040CCCCCCC8443C905140C23";
    attribute INIT_11 of inst : label is "C000000008033330800000000CCC200000000000000000000000000000020800";
    attribute INIT_12 of inst : label is "004447C3C03F007C4447CF0701C1CC3FC0307090C010D01CC01D00800000004C";
    attribute INIT_13 of inst : label is "555555555555543B1CCEEFFFF300000002C447030000DC3090D0723C300F00FF";
    attribute INIT_14 of inst : label is "F87FC3C3DF2CF7C7E702C7E702C7CB1C646400300040C00CF7371D5555555555";
    attribute INIT_15 of inst : label is "14070C30DFB437BE1FC30DFB04370BE1C7F0D8C5F70BFB0387FC36317DF0BFB0";
    attribute INIT_16 of inst : label is "71C00000000000000003F6FDAFFF000003FB0021300CCD10007007300101007D";
    attribute INIT_17 of inst : label is "452D8761D030F4FCF0C30FC4470330C0301C120C00CCCCF0D1C010F0F1C7795C";
    attribute INIT_18 of inst : label is "B00053F00C741010F83C100106181C0071C1C00607001C71C1C0061851451451";
    attribute INIT_19 of inst : label is "B2C013FC31C41C42FD02E0B3C13F90C0C0C71C0C0C71C003030303030303C303";
    attribute INIT_1A of inst : label is "3F3D13D240731C00000000F000000FC0FD4F60F2CBB01C0700CB2C3CFC31C40C";
    attribute INIT_1B of inst : label is "D0D4108CFC0E007800D01C803423CB4F0DC0720B1C41C81C41C4F40B040D0814";
    attribute INIT_1C of inst : label is "000003000FC0FD4F60F2CB0CF00C1C822C071DCD0D4108CF01C82C071D0C71DC";
    attribute INIT_1D of inst : label is "00303800C71C71C7871C0CF04F2D3CF4F0000300000F00003C000D0000000300";
    attribute INIT_1E of inst : label is "0740303E0F070874740300C03071C723F0DC00430EC400730DC006314C5314ED";
    attribute INIT_1F of inst : label is "3813773743034D43D40905303F53D83CB2C33C33F03CF1C8074082C01D03C20F";
    attribute INIT_20 of inst : label is "00000C303004020300F00C7F070032C2C0143B014C783FF3C0301FF03F438137";
    attribute INIT_21 of inst : label is "870C002000B031C0D1C340C21C00013CF031C302C72E471C1C7F6FF3C3400030";
    attribute INIT_22 of inst : label is "F0C0F2CC700C0F2E1C1C0CB310CB0C21CF00C0F4F4F02C7603C00F03C303C0B0";
    attribute INIT_23 of inst : label is "0C07134C53007C03CF3F6FFF0F00C032C2C0531006A691F0B01450C031CB3C00";
    attribute INIT_24 of inst : label is "1FC70750374003803403003C00EF3C13C7003F0E10C070130000FE0C420C6C0C";
    attribute INIT_25 of inst : label is "0C0CB63F63DCF73F0C0C0C0063FB0140514000C0C0F3D13F030C00C00C00C003";
    attribute INIT_26 of inst : label is "34200601C7031C0B1FD82C34F0C0CB6013F00004C2F4FFF40FC04D050B2C760B";
    attribute INIT_27 of inst : label is "1C71C1C7C71C1C753D03FF0C331C7071D5C30C33471C1C77501AA042053F4F00";
    attribute INIT_28 of inst : label is "C13F1C13D880B1C700FC701C707110006347700F43011E031C300E3D13F031C3";
    attribute INIT_29 of inst : label is "CD5D741C7077D471C71D80000B097006C21C1C1DBC74C071C71C004F00C0FFF1";
    attribute INIT_2A of inst : label is "1C71C1C73CF5F460103D85C17C741EF52CD471F5D71705C442010075F172D172";
    attribute INIT_2B of inst : label is "071CF03471DBC74071C0C0CC4FFFD3FC71C71C71C71C0B1C33C0B1C30871C707";
    attribute INIT_2C of inst : label is "1080631C701C3FF4C71C01C7C71D8CFF0C21CF1D0747600006C21C00B0970707";
    attribute INIT_2D of inst : label is "13C71C071D2C712D001DB31CB42CC7FC71C71C1C0007013C13C1C701C701C071";
    attribute INIT_2E of inst : label is "C3C006CC706CC7031C0C0C7072C11C4B401C6CC72C13D0701EF52CD113F3C23C";
    attribute INIT_2F of inst : label is "5D75C5D6CC17406FC0DBCBF5DB35D5D7C601A931F4FDD3F40CC7070777DC7CF0";
    attribute INIT_30 of inst : label is "0004006C0B4B40F00870C310010004006D2D0870C4F15C571BCBF06D74E1F707";
    attribute INIT_31 of inst : label is "A0C0DC70C03CF1D3C31C71DE1C7C0C0FFFDE1C71C7630C71D8CF8F031C34006F";
    attribute INIT_32 of inst : label is "F3CCC01C7071C0D1D1080631C71C001C7071C01C701C707110006347700F4301";
    attribute INIT_33 of inst : label is "31CB2C7C0D31D35CB2C7C013C70C0D21D0CC7E3F31CC7FCCC02D3F07307631FF";
    attribute INIT_34 of inst : label is "F0304DC0F031D0C04CC753574F1F0872DCCB47C0D1D351CB2C704FC0C0D31D35";
    attribute INIT_35 of inst : label is "4241000000000000C301FC7FCB6331F00004C7DB0007FD581658D4D871406331";
    attribute INIT_36 of inst : label is "3234218EDBEDBEDB6F822104104104104104104104104104104080601110000C";
    attribute INIT_37 of inst : label is "000000000000000020000000000000000000000000441010033120232111112C";
    attribute INIT_38 of inst : label is "0000200000000000000020000000000000000000000000000000003000000000";
    attribute INIT_39 of inst : label is "0000000000000000002000000000000000000000000000000000000000000020";
    attribute INIT_3A of inst : label is "0000000000000000000000000002000000000000000000000000000030000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000030000000000000000000002000000200000";
    attribute INIT_3C of inst : label is "0000000000000010001010001000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0044000000011001000010000000100000001101000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "1000000000001010000101000000000000100010000010001000010010004400";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
