-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "2826B20DE92534A788C494A5014A1294249FF1112E050083EF6135DFDEA33339";
    attribute INIT_01 of inst : label is "30CD14E1C7A43AEFB35F87A6E1107AFFF94D199CD9080987F8807108A3FDE000";
    attribute INIT_02 of inst : label is "31518E8E746A12C81895650943ED62CA2A0AA4012A25488AA60509A1548050C2";
    attribute INIT_03 of inst : label is "1555DD75D55714D34F17499A1E7D3B9DD4EE6753B9D365994D97F9C9EC099A2A";
    attribute INIT_04 of inst : label is "0C22E7A8001F188B89414787A2FA801100000000015DA5656565369B4D30D345";
    attribute INIT_05 of inst : label is "D67B249994A8F555555C550467F2AF1541F9FDFFD114662E62C444019F8BF150";
    attribute INIT_06 of inst : label is "9C4D6FB78F59D236B6A13822153B7CCE9ECCCACC91E50059608820180A2E051C";
    attribute INIT_07 of inst : label is "8088B5DE44E28200827BE6BA8E2048608010410AF742220273B9ACCBCD2CF022";
    attribute INIT_08 of inst : label is "44A90C97F297C762E0AA9B33AF90404C976AD769917BB4A8259F70828ABDDE70";
    attribute INIT_09 of inst : label is "9057C00AC2BE01A002B0AF80049A146981469D9DDD279F2FD7A45E49C9792F26";
    attribute INIT_0A of inst : label is "F37D16B159F2ED770984E3A441245A02FCC00000000030C20C30822ECFBFAAEA";
    attribute INIT_0B of inst : label is "33BC8CBDD5A6B7AE66FECF09D741DB3131EA32B7D7C9C77414D989A626B5AD6F";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE7EA4140A5B8ACCCBD5DB2AB67779D6C602034E97";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF4400000052707270B54A5FFFF6F6F74000000001402D5297FFFDBDBD9";
    attribute INIT_10 of inst : label is "2826B20DE92534A788C494A5014A1294249FF1112E050083EF6135DFDEA33339";
    attribute INIT_11 of inst : label is "30CD14E1C7A43AEFB35F87A6E1107AFFF94D199CD9080987F8807108A3FDE000";
    attribute INIT_12 of inst : label is "31518E8E746A12C81895650943ED62CA2A0AA4012A25488AA60509A1548050C2";
    attribute INIT_13 of inst : label is "1555DD75D55714D34F17499A1E7D3B9DD4EE6753B9D365994D97F9C9EC099A2A";
    attribute INIT_14 of inst : label is "0C22E7A8001F188B89414787A2FA801100000000015DA5656565369B4D30D345";
    attribute INIT_15 of inst : label is "D67B249994A8F555555C550467F2AF1541F9FDFFD114662E62C444019F8BF150";
    attribute INIT_16 of inst : label is "9C4D6FB78F59D236B6A13822153B7CCE9ECCCACC91E50059608820180A2E051C";
    attribute INIT_17 of inst : label is "8088B5DE44E28200827BE6BA8E2048608010410AF742220273B9ACCBCD2CF022";
    attribute INIT_18 of inst : label is "44A90C97F297C762E0AA9B33AF90404C976AD769917BB4A8259F70828ABDDE70";
    attribute INIT_19 of inst : label is "9057C00AC2BE01A002B0AF80049A146981469D9DDD279F2FD7A45E49C9792F26";
    attribute INIT_1A of inst : label is "F37D16B159F2ED770984E3A441245A02FCC00000000030C20C30822ECFBFAAEA";
    attribute INIT_1B of inst : label is "33BC8CBDD5A6B7AE66FECF09D741DB3131EA32B7D7C9C77414D989A626B5AD6F";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE7EA4140A5B8ACCCBD5DB2AB67779D6C602034E97";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF4400000052707270B54A5FFFF6F6F74000000001402D5297FFFDBDBD9";
    attribute INIT_20 of inst : label is "2826B20DE92534A788C494A5014A1294249FF1112E050083EF6135DFDEA33339";
    attribute INIT_21 of inst : label is "30CD14E1C7A43AEFB35F87A6E1107AFFF94D199CD9080987F8807108A3FDE000";
    attribute INIT_22 of inst : label is "31518E8E746A12C81895650943ED62CA2A0AA4012A25488AA60509A1548050C2";
    attribute INIT_23 of inst : label is "1555DD75D55714D34F17499A1E7D3B9DD4EE6753B9D365994D97F9C9EC099A2A";
    attribute INIT_24 of inst : label is "0C22E7A8001F188B89414787A2FA801100000000015DA5656565369B4D30D345";
    attribute INIT_25 of inst : label is "D67B249994A8F555555C550467F2AF1541F9FDFFD114662E62C444019F8BF150";
    attribute INIT_26 of inst : label is "9C4D6FB78F59D236B6A13822153B7CCE9ECCCACC91E50059608820180A2E051C";
    attribute INIT_27 of inst : label is "8088B5DE44E28200827BE6BA8E2048608010410AF742220273B9ACCBCD2CF022";
    attribute INIT_28 of inst : label is "44A90C97F297C762E0AA9B33AF90404C976AD769917BB4A8259F70828ABDDE70";
    attribute INIT_29 of inst : label is "9057C00AC2BE01A002B0AF80049A146981469D9DDD279F2FD7A45E49C9792F26";
    attribute INIT_2A of inst : label is "F37D16B159F2ED770984E3A441245A02FCC00000000030C20C30822ECFBFAAEA";
    attribute INIT_2B of inst : label is "33BC8CBDD5A6B7AE66FECF09D741DB3131EA32B7D7C9C77414D989A626B5AD6F";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE7EA4140A5B8ACCCBD5DB2AB67779D6C602034E97";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF4400000052707270B54A5FFFF6F6F74000000001402D5297FFFDBDBD9";
    attribute INIT_30 of inst : label is "2826B20DE92534A788C494A5014A1294249FF1112E050083EF6135DFDEA33339";
    attribute INIT_31 of inst : label is "30CD14E1C7A43AEFB35F87A6E1107AFFF94D199CD9080987F8807108A3FDE000";
    attribute INIT_32 of inst : label is "31518E8E746A12C81895650943ED62CA2A0AA4012A25488AA60509A1548050C2";
    attribute INIT_33 of inst : label is "1555DD75D55714D34F17499A1E7D3B9DD4EE6753B9D365994D97F9C9EC099A2A";
    attribute INIT_34 of inst : label is "0C22E7A8001F188B89414787A2FA801100000000015DA5656565369B4D30D345";
    attribute INIT_35 of inst : label is "D67B249994A8F555555C550467F2AF1541F9FDFFD114662E62C444019F8BF150";
    attribute INIT_36 of inst : label is "9C4D6FB78F59D236B6A13822153B7CCE9ECCCACC91E50059608820180A2E051C";
    attribute INIT_37 of inst : label is "8088B5DE44E28200827BE6BA8E2048608010410AF742220273B9ACCBCD2CF022";
    attribute INIT_38 of inst : label is "44A90C97F297C762E0AA9B33AF90404C976AD769917BB4A8259F70828ABDDE70";
    attribute INIT_39 of inst : label is "9057C00AC2BE01A002B0AF80049A146981469D9DDD279F2FD7A45E49C9792F26";
    attribute INIT_3A of inst : label is "F37D16B159F2ED770984E3A441245A02FCC00000000030C20C30822ECFBFAAEA";
    attribute INIT_3B of inst : label is "33BC8CBDD5A6B7AE66FECF09D741DB3131EA32B7D7C9C77414D989A626B5AD6F";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE7EA4140A5B8ACCCBD5DB2AB67779D6C602034E97";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF4400000052707270B54A5FFFF6F6F74000000001402D5297FFFDBDBD9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "65D823424048190D41F927EFAFDF4FBE80401329F2162C07AC289E7E7E6623B3";
    attribute INIT_01 of inst : label is "EF7F328019641505A9A9513A6DB6318080DF8BD11B1D6BE0A82A9299B404D6DB";
    attribute INIT_02 of inst : label is "46227111889366FCDF7ADAFEF62095BFD6A7539F3F71B5FB486FAA77FEC7FECA";
    attribute INIT_03 of inst : label is "BBEF36D36DB4D3EFBCF0E3144532403A2908E9A403E04DE28133FA19F3C908C4";
    attribute INIT_04 of inst : label is "021D185000008274664450781D054449C000008B001008A0A0A0080802BEEBAE";
    attribute INIT_05 of inst : label is "915249466E025999999E502A184D57940A061201E14209D19D5051EA60741441";
    attribute INIT_06 of inst : label is "A9193A457EBC2D17776CAC26C04C82D5211BBB2B178A5503C92249B37372B7D2";
    attribute INIT_07 of inst : label is "FDEF533815F20822085FCB3DDA0240240800000BFE367C053AFB0E6B0E759471";
    attribute INIT_08 of inst : label is "870E11E0351E4C9685667F1D3EEB772404B54CE25AB6700025AD9DFDEF53389D";
    attribute INIT_09 of inst : label is "7087C0BB447E2FE02CD11F80053C1C5BE1C4B02FFE42AB4865DA108210420047";
    attribute INIT_0A of inst : label is "4043BA8AEF062599DEEF77F2A80A8891FEDE000000000000041040011A141051";
    attribute INIT_0B of inst : label is "CC53318FFECFC9F39D8536CDF289E8CE5D1FC5F86D4D21872FA6F6D9CB2D6B57";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC55CF30CEC21CB9BB37326EEDCCD55EA2464485BE";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF41000000572277026CDC00FFF000090000000000155B372ABFFC00002";
    attribute INIT_10 of inst : label is "65D823424048190D41F927EFAFDF4FBE80401329F2162C07AC289E7E7E6623B3";
    attribute INIT_11 of inst : label is "EF7F328019641505A9A9513A6DB6318080DF8BD11B1D6BE0A82A9299B404D6DB";
    attribute INIT_12 of inst : label is "46227111889366FCDF7ADAFEF62095BFD6A7539F3F71B5FB486FAA77FEC7FECA";
    attribute INIT_13 of inst : label is "BBEF36D36DB4D3EFBCF0E3144532403A2908E9A403E04DE28133FA19F3C908C4";
    attribute INIT_14 of inst : label is "021D185000008274664450781D054449C000008B001008A0A0A0080802BEEBAE";
    attribute INIT_15 of inst : label is "915249466E025999999E502A184D57940A061201E14209D19D5051EA60741441";
    attribute INIT_16 of inst : label is "A9193A457EBC2D17776CAC26C04C82D5211BBB2B178A5503C92249B37372B7D2";
    attribute INIT_17 of inst : label is "FDEF533815F20822085FCB3DDA0240240800000BFE367C053AFB0E6B0E759471";
    attribute INIT_18 of inst : label is "870E11E0351E4C9685667F1D3EEB772404B54CE25AB6700025AD9DFDEF53389D";
    attribute INIT_19 of inst : label is "7087C0BB447E2FE02CD11F80053C1C5BE1C4B02FFE42AB4865DA108210420047";
    attribute INIT_1A of inst : label is "4043BA8AEF062599DEEF77F2A80A8891FEDE000000000000041040011A141051";
    attribute INIT_1B of inst : label is "CC53318FFECFC9F39D8536CDF289E8CE5D1FC5F86D4D21872FA6F6D9CB2D6B57";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC55CF30CEC21CB9BB37326EEDCCD55EA2464485BE";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF41000000572277026CDC00FFF000090000000000155B372ABFFC00002";
    attribute INIT_20 of inst : label is "65D823424048190D41F927EFAFDF4FBE80401329F2162C07AC289E7E7E6623B3";
    attribute INIT_21 of inst : label is "EF7F328019641505A9A9513A6DB6318080DF8BD11B1D6BE0A82A9299B404D6DB";
    attribute INIT_22 of inst : label is "46227111889366FCDF7ADAFEF62095BFD6A7539F3F71B5FB486FAA77FEC7FECA";
    attribute INIT_23 of inst : label is "BBEF36D36DB4D3EFBCF0E3144532403A2908E9A403E04DE28133FA19F3C908C4";
    attribute INIT_24 of inst : label is "021D185000008274664450781D054449C000008B001008A0A0A0080802BEEBAE";
    attribute INIT_25 of inst : label is "915249466E025999999E502A184D57940A061201E14209D19D5051EA60741441";
    attribute INIT_26 of inst : label is "A9193A457EBC2D17776CAC26C04C82D5211BBB2B178A5503C92249B37372B7D2";
    attribute INIT_27 of inst : label is "FDEF533815F20822085FCB3DDA0240240800000BFE367C053AFB0E6B0E759471";
    attribute INIT_28 of inst : label is "870E11E0351E4C9685667F1D3EEB772404B54CE25AB6700025AD9DFDEF53389D";
    attribute INIT_29 of inst : label is "7087C0BB447E2FE02CD11F80053C1C5BE1C4B02FFE42AB4865DA108210420047";
    attribute INIT_2A of inst : label is "4043BA8AEF062599DEEF77F2A80A8891FEDE000000000000041040011A141051";
    attribute INIT_2B of inst : label is "CC53318FFECFC9F39D8536CDF289E8CE5D1FC5F86D4D21872FA6F6D9CB2D6B57";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC55CF30CEC21CB9BB37326EEDCCD55EA2464485BE";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF41000000572277026CDC00FFF000090000000000155B372ABFFC00002";
    attribute INIT_30 of inst : label is "65D823424048190D41F927EFAFDF4FBE80401329F2162C07AC289E7E7E6623B3";
    attribute INIT_31 of inst : label is "EF7F328019641505A9A9513A6DB6318080DF8BD11B1D6BE0A82A9299B404D6DB";
    attribute INIT_32 of inst : label is "46227111889366FCDF7ADAFEF62095BFD6A7539F3F71B5FB486FAA77FEC7FECA";
    attribute INIT_33 of inst : label is "BBEF36D36DB4D3EFBCF0E3144532403A2908E9A403E04DE28133FA19F3C908C4";
    attribute INIT_34 of inst : label is "021D185000008274664450781D054449C000008B001008A0A0A0080802BEEBAE";
    attribute INIT_35 of inst : label is "915249466E025999999E502A184D57940A061201E14209D19D5051EA60741441";
    attribute INIT_36 of inst : label is "A9193A457EBC2D17776CAC26C04C82D5211BBB2B178A5503C92249B37372B7D2";
    attribute INIT_37 of inst : label is "FDEF533815F20822085FCB3DDA0240240800000BFE367C053AFB0E6B0E759471";
    attribute INIT_38 of inst : label is "870E11E0351E4C9685667F1D3EEB772404B54CE25AB6700025AD9DFDEF53389D";
    attribute INIT_39 of inst : label is "7087C0BB447E2FE02CD11F80053C1C5BE1C4B02FFE42AB4865DA108210420047";
    attribute INIT_3A of inst : label is "4043BA8AEF062599DEEF77F2A80A8891FEDE000000000000041040011A141051";
    attribute INIT_3B of inst : label is "CC53318FFECFC9F39D8536CDF289E8CE5D1FC5F86D4D21872FA6F6D9CB2D6B57";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC55CF30CEC21CB9BB37326EEDCCD55EA2464485BE";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF41000000572277026CDC00FFF000090000000000155B372ABFFC00002";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "AC6C9B0B6A1152384EF2458DC31B9637206FE10252F489532F0C2A2E2E77895A";
    attribute INIT_01 of inst : label is "AE6C338E313D4041194D7F3E6DB936000F7FEFE2429152F897008088B0293B6D";
    attribute INIT_02 of inst : label is "63331D98ECCF199172982C30314719ABDAF44618AA4529CB18E7860F7C1F7C42";
    attribute INIT_03 of inst : label is "259659659659651451451441004B6CBF8DB2FF36EBBACDBCEB33FB59C7290866";
    attribute INIT_04 of inst : label is "3162E7A800004D8B98C44007E2FAF265A000001BA0462969696950A944249249";
    attribute INIT_05 of inst : label is "0D292DCCEB38BE1E1E1F96D16FBAAFE5B5FBEFFFFD69362EEA8F5A159F8BFC62";
    attribute INIT_06 of inst : label is "92154067CB9E9C07474CA967C71B0D8DB65E6BCC4F3395CA5B66DBBD9B9AF659";
    attribute INIT_07 of inst : label is "0C8E712C95F6C300C34FC7B9F08801000155155BFB167809D28080A20A4F1E3A";
    attribute INIT_08 of inst : label is "970E11E1B69CED9A8664FF9DBEE632209611E0B208F259002D3FDB4CCE782C93";
    attribute INIT_09 of inst : label is "2009C02D000E0A4009501380016C0014C000442445C1B569A3DC0E83D07A0F47";
    attribute INIT_0A of inst : label is "194EB083AF9775309C0C75F220AA42C5FEC144444444451555551574E1C3C74C";
    attribute INIT_0B of inst : label is "2B58AD2D8A8F21AD6E860F5F8705C229751B8D2CC39F87462CD14B873E39CE77";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC134F3A84E93F6EEEDDDDBBBB7750348266661C1E";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFBFFFFF0031134664ECCF00FF0FFFF01555555555513B33C03FC3FFFFC";
    attribute INIT_10 of inst : label is "AC6C9B0B6A1152384EF2458DC31B9637206FE10252F489532F0C2A2E2E77895A";
    attribute INIT_11 of inst : label is "AE6C338E313D4041194D7F3E6DB936000F7FEFE2429152F897008088B0293B6D";
    attribute INIT_12 of inst : label is "63331D98ECCF199172982C30314719ABDAF44618AA4529CB18E7860F7C1F7C42";
    attribute INIT_13 of inst : label is "259659659659651451451441004B6CBF8DB2FF36EBBACDBCEB33FB59C7290866";
    attribute INIT_14 of inst : label is "3162E7A800004D8B98C44007E2FAF265A000001BA0462969696950A944249249";
    attribute INIT_15 of inst : label is "0D292DCCEB38BE1E1E1F96D16FBAAFE5B5FBEFFFFD69362EEA8F5A159F8BFC62";
    attribute INIT_16 of inst : label is "92154067CB9E9C07474CA967C71B0D8DB65E6BCC4F3395CA5B66DBBD9B9AF659";
    attribute INIT_17 of inst : label is "0C8E712C95F6C300C34FC7B9F08801000155155BFB167809D28080A20A4F1E3A";
    attribute INIT_18 of inst : label is "970E11E1B69CED9A8664FF9DBEE632209611E0B208F259002D3FDB4CCE782C93";
    attribute INIT_19 of inst : label is "2009C02D000E0A4009501380016C0014C000442445C1B569A3DC0E83D07A0F47";
    attribute INIT_1A of inst : label is "194EB083AF9775309C0C75F220AA42C5FEC144444444451555551574E1C3C74C";
    attribute INIT_1B of inst : label is "2B58AD2D8A8F21AD6E860F5F8705C229751B8D2CC39F87462CD14B873E39CE77";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC134F3A84E93F6EEEDDDDBBBB7750348266661C1E";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFBFFFFF0031134664ECCF00FF0FFFF01555555555513B33C03FC3FFFFC";
    attribute INIT_20 of inst : label is "AC6C9B0B6A1152384EF2458DC31B9637206FE10252F489532F0C2A2E2E77895A";
    attribute INIT_21 of inst : label is "AE6C338E313D4041194D7F3E6DB936000F7FEFE2429152F897008088B0293B6D";
    attribute INIT_22 of inst : label is "63331D98ECCF199172982C30314719ABDAF44618AA4529CB18E7860F7C1F7C42";
    attribute INIT_23 of inst : label is "259659659659651451451441004B6CBF8DB2FF36EBBACDBCEB33FB59C7290866";
    attribute INIT_24 of inst : label is "3162E7A800004D8B98C44007E2FAF265A000001BA0462969696950A944249249";
    attribute INIT_25 of inst : label is "0D292DCCEB38BE1E1E1F96D16FBAAFE5B5FBEFFFFD69362EEA8F5A159F8BFC62";
    attribute INIT_26 of inst : label is "92154067CB9E9C07474CA967C71B0D8DB65E6BCC4F3395CA5B66DBBD9B9AF659";
    attribute INIT_27 of inst : label is "0C8E712C95F6C300C34FC7B9F08801000155155BFB167809D28080A20A4F1E3A";
    attribute INIT_28 of inst : label is "970E11E1B69CED9A8664FF9DBEE632209611E0B208F259002D3FDB4CCE782C93";
    attribute INIT_29 of inst : label is "2009C02D000E0A4009501380016C0014C000442445C1B569A3DC0E83D07A0F47";
    attribute INIT_2A of inst : label is "194EB083AF9775309C0C75F220AA42C5FEC144444444451555551574E1C3C74C";
    attribute INIT_2B of inst : label is "2B58AD2D8A8F21AD6E860F5F8705C229751B8D2CC39F87462CD14B873E39CE77";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC134F3A84E93F6EEEDDDDBBBB7750348266661C1E";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFBFFFFF0031134664ECCF00FF0FFFF01555555555513B33C03FC3FFFFC";
    attribute INIT_30 of inst : label is "AC6C9B0B6A1152384EF2458DC31B9637206FE10252F489532F0C2A2E2E77895A";
    attribute INIT_31 of inst : label is "AE6C338E313D4041194D7F3E6DB936000F7FEFE2429152F897008088B0293B6D";
    attribute INIT_32 of inst : label is "63331D98ECCF199172982C30314719ABDAF44618AA4529CB18E7860F7C1F7C42";
    attribute INIT_33 of inst : label is "259659659659651451451441004B6CBF8DB2FF36EBBACDBCEB33FB59C7290866";
    attribute INIT_34 of inst : label is "3162E7A800004D8B98C44007E2FAF265A000001BA0462969696950A944249249";
    attribute INIT_35 of inst : label is "0D292DCCEB38BE1E1E1F96D16FBAAFE5B5FBEFFFFD69362EEA8F5A159F8BFC62";
    attribute INIT_36 of inst : label is "92154067CB9E9C07474CA967C71B0D8DB65E6BCC4F3395CA5B66DBBD9B9AF659";
    attribute INIT_37 of inst : label is "0C8E712C95F6C300C34FC7B9F08801000155155BFB167809D28080A20A4F1E3A";
    attribute INIT_38 of inst : label is "970E11E1B69CED9A8664FF9DBEE632209611E0B208F259002D3FDB4CCE782C93";
    attribute INIT_39 of inst : label is "2009C02D000E0A4009501380016C0014C000442445C1B569A3DC0E83D07A0F47";
    attribute INIT_3A of inst : label is "194EB083AF9775309C0C75F220AA42C5FEC144444444451555551574E1C3C74C";
    attribute INIT_3B of inst : label is "2B58AD2D8A8F21AD6E860F5F8705C229751B8D2CC39F87462CD14B873E39CE77";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC134F3A84E93F6EEEDDDDBBBB7750348266661C1E";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFBFFFFF0031134664ECCF00FF0FFFF01555555555513B33C03FC3FFFFC";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "AD6DDD4B2A11523F8E2A45DEEBBDC77BA065011A44EB8957020448C8C9D6580A";
    attribute INIT_01 of inst : label is "1FC82DCE53AC1404044138AA829F3E7FFBA0E47301D033A0822A5081542FBB6D";
    attribute INIT_02 of inst : label is "3111888C446D515028EF2434B455B960DC37EB0D8AE421F5ECB4EB2A4A9A4A8A";
    attribute INIT_03 of inst : label is "40000000000000000000000003F97A93C5EA4E17A933443CDD1083C817C50A22";
    attribute INIT_04 of inst : label is "C095185000003054650D280015053973CAA220190144A949494918A854410410";
    attribute INIT_05 of inst : label is "97292CEED71B601FE01F6A80B7F557DAA00DFDFFF680C1D33505A000607402DC";
    attribute INIT_06 of inst : label is "00C44066F1EE9E18C8C61419E37B0DC8BE4E75E5C133C74E77DDF73F91EDE28B";
    attribute INIT_07 of inst : label is "5C77A8403E100000000BDE44D80000000020C302FD35BC101488A882A8EBA8C1";
    attribute INIT_08 of inst : label is "3A54A84FA7282D591E4470A8F0BAABBADBD68102CB40807D4352E31C37A040AB";
    attribute INIT_09 of inst : label is "30C040E186423A603A7180800340000420004CA2222534691A1F29652CE59C99";
    attribute INIT_0A of inst : label is "B068999339F273B2114A9436606E02DDFDC05444545469969A65C6B0E9D3C30D";
    attribute INIT_0B of inst : label is "ED5FB53DD3C565B5AE96AF6DE7C8FFEF671FE93E8F6DE6AEB71F7B3DEC98C63C";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE326478E76F124CCEDDD93BB277773F8355FFEDB5";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFAA63630077577777E23F00FFF9F9F9155555555114388FC03FFE7E7E4";
    attribute INIT_10 of inst : label is "AD6DDD4B2A11523F8E2A45DEEBBDC77BA065011A44EB8957020448C8C9D6580A";
    attribute INIT_11 of inst : label is "1FC82DCE53AC1404044138AA829F3E7FFBA0E47301D033A0822A5081542FBB6D";
    attribute INIT_12 of inst : label is "3111888C446D515028EF2434B455B960DC37EB0D8AE421F5ECB4EB2A4A9A4A8A";
    attribute INIT_13 of inst : label is "40000000000000000000000003F97A93C5EA4E17A933443CDD1083C817C50A22";
    attribute INIT_14 of inst : label is "C095185000003054650D280015053973CAA220190144A949494918A854410410";
    attribute INIT_15 of inst : label is "97292CEED71B601FE01F6A80B7F557DAA00DFDFFF680C1D33505A000607402DC";
    attribute INIT_16 of inst : label is "00C44066F1EE9E18C8C61419E37B0DC8BE4E75E5C133C74E77DDF73F91EDE28B";
    attribute INIT_17 of inst : label is "5C77A8403E100000000BDE44D80000000020C302FD35BC101488A882A8EBA8C1";
    attribute INIT_18 of inst : label is "3A54A84FA7282D591E4470A8F0BAABBADBD68102CB40807D4352E31C37A040AB";
    attribute INIT_19 of inst : label is "30C040E186423A603A7180800340000420004CA2222534691A1F29652CE59C99";
    attribute INIT_1A of inst : label is "B068999339F273B2114A9436606E02DDFDC05444545469969A65C6B0E9D3C30D";
    attribute INIT_1B of inst : label is "ED5FB53DD3C565B5AE96AF6DE7C8FFEF671FE93E8F6DE6AEB71F7B3DEC98C63C";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE326478E76F124CCEDDD93BB277773F8355FFEDB5";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFAA63630077577777E23F00FFF9F9F9155555555114388FC03FFE7E7E4";
    attribute INIT_20 of inst : label is "AD6DDD4B2A11523F8E2A45DEEBBDC77BA065011A44EB8957020448C8C9D6580A";
    attribute INIT_21 of inst : label is "1FC82DCE53AC1404044138AA829F3E7FFBA0E47301D033A0822A5081542FBB6D";
    attribute INIT_22 of inst : label is "3111888C446D515028EF2434B455B960DC37EB0D8AE421F5ECB4EB2A4A9A4A8A";
    attribute INIT_23 of inst : label is "40000000000000000000000003F97A93C5EA4E17A933443CDD1083C817C50A22";
    attribute INIT_24 of inst : label is "C095185000003054650D280015053973CAA220190144A949494918A854410410";
    attribute INIT_25 of inst : label is "97292CEED71B601FE01F6A80B7F557DAA00DFDFFF680C1D33505A000607402DC";
    attribute INIT_26 of inst : label is "00C44066F1EE9E18C8C61419E37B0DC8BE4E75E5C133C74E77DDF73F91EDE28B";
    attribute INIT_27 of inst : label is "5C77A8403E100000000BDE44D80000000020C302FD35BC101488A882A8EBA8C1";
    attribute INIT_28 of inst : label is "3A54A84FA7282D591E4470A8F0BAABBADBD68102CB40807D4352E31C37A040AB";
    attribute INIT_29 of inst : label is "30C040E186423A603A7180800340000420004CA2222534691A1F29652CE59C99";
    attribute INIT_2A of inst : label is "B068999339F273B2114A9436606E02DDFDC05444545469969A65C6B0E9D3C30D";
    attribute INIT_2B of inst : label is "ED5FB53DD3C565B5AE96AF6DE7C8FFEF671FE93E8F6DE6AEB71F7B3DEC98C63C";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE326478E76F124CCEDDD93BB277773F8355FFEDB5";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFAA63630077577777E23F00FFF9F9F9155555555114388FC03FFE7E7E4";
    attribute INIT_30 of inst : label is "AD6DDD4B2A11523F8E2A45DEEBBDC77BA065011A44EB8957020448C8C9D6580A";
    attribute INIT_31 of inst : label is "1FC82DCE53AC1404044138AA829F3E7FFBA0E47301D033A0822A5081542FBB6D";
    attribute INIT_32 of inst : label is "3111888C446D515028EF2434B455B960DC37EB0D8AE421F5ECB4EB2A4A9A4A8A";
    attribute INIT_33 of inst : label is "40000000000000000000000003F97A93C5EA4E17A933443CDD1083C817C50A22";
    attribute INIT_34 of inst : label is "C095185000003054650D280015053973CAA220190144A949494918A854410410";
    attribute INIT_35 of inst : label is "97292CEED71B601FE01F6A80B7F557DAA00DFDFFF680C1D33505A000607402DC";
    attribute INIT_36 of inst : label is "00C44066F1EE9E18C8C61419E37B0DC8BE4E75E5C133C74E77DDF73F91EDE28B";
    attribute INIT_37 of inst : label is "5C77A8403E100000000BDE44D80000000020C302FD35BC101488A882A8EBA8C1";
    attribute INIT_38 of inst : label is "3A54A84FA7282D591E4470A8F0BAABBADBD68102CB40807D4352E31C37A040AB";
    attribute INIT_39 of inst : label is "30C040E186423A603A7180800340000420004CA2222534691A1F29652CE59C99";
    attribute INIT_3A of inst : label is "B068999339F273B2114A9436606E02DDFDC05444545469969A65C6B0E9D3C30D";
    attribute INIT_3B of inst : label is "ED5FB53DD3C565B5AE96AF6DE7C8FFEF671FE93E8F6DE6AEB71F7B3DEC98C63C";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFE326478E76F124CCEDDD93BB277773F8355FFEDB5";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFAA63630077577777E23F00FFF9F9F9155555555114388FC03FFE7E7E4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "4909206050AA0C4065208AC2748C6B09CB855AAEC3E200A24D53C02C2D444D83";
    attribute INIT_01 of inst : label is "7912293020DA85AC12A111AF80C2B0404C608C443216AA3054003A95052E8596";
    attribute INIT_02 of inst : label is "63335DDAEEC8D002406209A524568DE406C118B3D26AA990504924049224922F";
    attribute INIT_03 of inst : label is "00000000000000000000000001813AB304E2CC13AB354C36D43003D816050866";
    attribute INIT_04 of inst : label is "844AE7A80001032B93F208004AFA9CFCAAA0A099AA81420202024D0283000000";
    attribute INIT_05 of inst : label is "08AB6DA8C0341FE0001E222C584AAF888A161201E8A40E2DDAF2280B9F8BFDAA";
    attribute INIT_06 of inst : label is "3BC4801C1830680CDCC8469786890391BD580123688855A59B26C96250C2E186";
    attribute INIT_07 of inst : label is "39234C220018000000202894E044090C128A28A009841020000A0A05F7945104";
    attribute INIT_08 of inst : label is "AD7AA9A96128094F094761B49A088880204514882298442090008D7963452205";
    attribute INIT_09 of inst : label is "37C0BFC1BE05F06FF26F917FFA45D3A45D3A422F761DB56D800380320600C812";
    attribute INIT_0A of inst : label is "B2AE810BA0D14220D6295D4910F94A9DFEE0555455545915D35115B0E1C3D34D";
    attribute INIT_0B of inst : label is "002000864A40C0C00202010471296400102CCCC0400431188B0000800239CE70";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC856CAAE6029113122624CCC0888211015F5CD840";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF11BF37FF02222222E01055FFF1F1F95555555554157804157FFC7C7C5";
    attribute INIT_10 of inst : label is "4909206050AA0C4065208AC2748C6B09CB855AAEC3E200A24D53C02C2D444D83";
    attribute INIT_11 of inst : label is "7912293020DA85AC12A111AF80C2B0404C608C443216AA3054003A95052E8596";
    attribute INIT_12 of inst : label is "63335DDAEEC8D002406209A524568DE406C118B3D26AA990504924049224922F";
    attribute INIT_13 of inst : label is "00000000000000000000000001813AB304E2CC13AB354C36D43003D816050866";
    attribute INIT_14 of inst : label is "844AE7A80001032B93F208004AFA9CFCAAA0A099AA81420202024D0283000000";
    attribute INIT_15 of inst : label is "08AB6DA8C0341FE0001E222C584AAF888A161201E8A40E2DDAF2280B9F8BFDAA";
    attribute INIT_16 of inst : label is "3BC4801C1830680CDCC8469786890391BD580123688855A59B26C96250C2E186";
    attribute INIT_17 of inst : label is "39234C220018000000202894E044090C128A28A009841020000A0A05F7945104";
    attribute INIT_18 of inst : label is "AD7AA9A96128094F094761B49A088880204514882298442090008D7963452205";
    attribute INIT_19 of inst : label is "37C0BFC1BE05F06FF26F917FFA45D3A45D3A422F761DB56D800380320600C812";
    attribute INIT_1A of inst : label is "B2AE810BA0D14220D6295D4910F94A9DFEE0555455545915D35115B0E1C3D34D";
    attribute INIT_1B of inst : label is "002000864A40C0C00202010471296400102CCCC0400431188B0000800239CE70";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC856CAAE6029113122624CCC0888211015F5CD840";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF11BF37FF02222222E01055FFF1F1F95555555554157804157FFC7C7C5";
    attribute INIT_20 of inst : label is "4909206050AA0C4065208AC2748C6B09CB855AAEC3E200A24D53C02C2D444D83";
    attribute INIT_21 of inst : label is "7912293020DA85AC12A111AF80C2B0404C608C443216AA3054003A95052E8596";
    attribute INIT_22 of inst : label is "63335DDAEEC8D002406209A524568DE406C118B3D26AA990504924049224922F";
    attribute INIT_23 of inst : label is "00000000000000000000000001813AB304E2CC13AB354C36D43003D816050866";
    attribute INIT_24 of inst : label is "844AE7A80001032B93F208004AFA9CFCAAA0A099AA81420202024D0283000000";
    attribute INIT_25 of inst : label is "08AB6DA8C0341FE0001E222C584AAF888A161201E8A40E2DDAF2280B9F8BFDAA";
    attribute INIT_26 of inst : label is "3BC4801C1830680CDCC8469786890391BD580123688855A59B26C96250C2E186";
    attribute INIT_27 of inst : label is "39234C220018000000202894E044090C128A28A009841020000A0A05F7945104";
    attribute INIT_28 of inst : label is "AD7AA9A96128094F094761B49A088880204514882298442090008D7963452205";
    attribute INIT_29 of inst : label is "37C0BFC1BE05F06FF26F917FFA45D3A45D3A422F761DB56D800380320600C812";
    attribute INIT_2A of inst : label is "B2AE810BA0D14220D6295D4910F94A9DFEE0555455545915D35115B0E1C3D34D";
    attribute INIT_2B of inst : label is "002000864A40C0C00202010471296400102CCCC0400431188B0000800239CE70";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC856CAAE6029113122624CCC0888211015F5CD840";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF11BF37FF02222222E01055FFF1F1F95555555554157804157FFC7C7C5";
    attribute INIT_30 of inst : label is "4909206050AA0C4065208AC2748C6B09CB855AAEC3E200A24D53C02C2D444D83";
    attribute INIT_31 of inst : label is "7912293020DA85AC12A111AF80C2B0404C608C443216AA3054003A95052E8596";
    attribute INIT_32 of inst : label is "63335DDAEEC8D002406209A524568DE406C118B3D26AA990504924049224922F";
    attribute INIT_33 of inst : label is "00000000000000000000000001813AB304E2CC13AB354C36D43003D816050866";
    attribute INIT_34 of inst : label is "844AE7A80001032B93F208004AFA9CFCAAA0A099AA81420202024D0283000000";
    attribute INIT_35 of inst : label is "08AB6DA8C0341FE0001E222C584AAF888A161201E8A40E2DDAF2280B9F8BFDAA";
    attribute INIT_36 of inst : label is "3BC4801C1830680CDCC8469786890391BD580123688855A59B26C96250C2E186";
    attribute INIT_37 of inst : label is "39234C220018000000202894E044090C128A28A009841020000A0A05F7945104";
    attribute INIT_38 of inst : label is "AD7AA9A96128094F094761B49A088880204514882298442090008D7963452205";
    attribute INIT_39 of inst : label is "37C0BFC1BE05F06FF26F917FFA45D3A45D3A422F761DB56D800380320600C812";
    attribute INIT_3A of inst : label is "B2AE810BA0D14220D6295D4910F94A9DFEE0555455545915D35115B0E1C3D34D";
    attribute INIT_3B of inst : label is "002000864A40C0C00202010471296400102CCCC0400431188B0000800239CE70";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC856CAAE6029113122624CCC0888211015F5CD840";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF11BF37FF02222222E01055FFF1F1F95555555554157804157FFC7C7C5";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "D9090660584F09E55A2112D765A6C94CE01E93394A0C2BE47B0035D151660B4B";
    attribute INIT_01 of inst : label is "4B36B8AEACE6900547ACBDFF8B8271BFB0E09C4CCB3B0770BCD5328164D84C96";
    attribute INIT_02 of inst : label is "6222599A888AD2821032412524CA45A26E5B39871868A132D61A65A1A621A608";
    attribute INIT_03 of inst : label is "000000000000000000000000000369822DAE08B6B8202026808002000A5D0866";
    attribute INIT_04 of inst : label is "0B2518500000CC946828807FA5051F2A000AA0902AC0636363630381C0000000";
    attribute INIT_05 of inst : label is "4972643900B60000001EA0D367BD57A835F9EFFFE28B31D66520A3F460740822";
    attribute INIT_06 of inst : label is "FE2B01A5BF7B6B2E7E6B42ABB6CD938C0081912B58CA5591C9224962D6C2ADB6";
    attribute INIT_07 of inst : label is "2B290880504A0000000429A76D404804828A28A90D04D6400022288EFBEFBEFB";
    attribute INIT_08 of inst : label is "70E1CD19016BCD6D235561A293580009004C0201261100AA1404052B29008045";
    attribute INIT_09 of inst : label is "00000040C0001000102000000042001020010404CC12AB420413102204408824";
    attribute INIT_0A of inst : label is "C0B10C2242C088CC522967A99DE996ADFDC1232323331450031050C408101041";
    attribute INIT_0B of inst : label is "4201080774605AE8432B41B76D8B60420A6456E930B72CD881021048416D7B50";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFD428125DE111400020400088000269125D5D4B94C";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF4100880000000000E01F11FF0909091555555555403807C47FC242424";
    attribute INIT_10 of inst : label is "D9090660584F09E55A2112D765A6C94CE01E93394A0C2BE47B0035D151660B4B";
    attribute INIT_11 of inst : label is "4B36B8AEACE6900547ACBDFF8B8271BFB0E09C4CCB3B0770BCD5328164D84C96";
    attribute INIT_12 of inst : label is "6222599A888AD2821032412524CA45A26E5B39871868A132D61A65A1A621A608";
    attribute INIT_13 of inst : label is "000000000000000000000000000369822DAE08B6B8202026808002000A5D0866";
    attribute INIT_14 of inst : label is "0B2518500000CC946828807FA5051F2A000AA0902AC0636363630381C0000000";
    attribute INIT_15 of inst : label is "4972643900B60000001EA0D367BD57A835F9EFFFE28B31D66520A3F460740822";
    attribute INIT_16 of inst : label is "FE2B01A5BF7B6B2E7E6B42ABB6CD938C0081912B58CA5591C9224962D6C2ADB6";
    attribute INIT_17 of inst : label is "2B290880504A0000000429A76D404804828A28A90D04D6400022288EFBEFBEFB";
    attribute INIT_18 of inst : label is "70E1CD19016BCD6D235561A293580009004C0201261100AA1404052B29008045";
    attribute INIT_19 of inst : label is "00000040C0001000102000000042001020010404CC12AB420413102204408824";
    attribute INIT_1A of inst : label is "C0B10C2242C088CC522967A99DE996ADFDC1232323331450031050C408101041";
    attribute INIT_1B of inst : label is "4201080774605AE8432B41B76D8B60420A6456E930B72CD881021048416D7B50";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFD428125DE111400020400088000269125D5D4B94C";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF4100880000000000E01F11FF0909091555555555403807C47FC242424";
    attribute INIT_20 of inst : label is "D9090660584F09E55A2112D765A6C94CE01E93394A0C2BE47B0035D151660B4B";
    attribute INIT_21 of inst : label is "4B36B8AEACE6900547ACBDFF8B8271BFB0E09C4CCB3B0770BCD5328164D84C96";
    attribute INIT_22 of inst : label is "6222599A888AD2821032412524CA45A26E5B39871868A132D61A65A1A621A608";
    attribute INIT_23 of inst : label is "000000000000000000000000000369822DAE08B6B8202026808002000A5D0866";
    attribute INIT_24 of inst : label is "0B2518500000CC946828807FA5051F2A000AA0902AC0636363630381C0000000";
    attribute INIT_25 of inst : label is "4972643900B60000001EA0D367BD57A835F9EFFFE28B31D66520A3F460740822";
    attribute INIT_26 of inst : label is "FE2B01A5BF7B6B2E7E6B42ABB6CD938C0081912B58CA5591C9224962D6C2ADB6";
    attribute INIT_27 of inst : label is "2B290880504A0000000429A76D404804828A28A90D04D6400022288EFBEFBEFB";
    attribute INIT_28 of inst : label is "70E1CD19016BCD6D235561A293580009004C0201261100AA1404052B29008045";
    attribute INIT_29 of inst : label is "00000040C0001000102000000042001020010404CC12AB420413102204408824";
    attribute INIT_2A of inst : label is "C0B10C2242C088CC522967A99DE996ADFDC1232323331450031050C408101041";
    attribute INIT_2B of inst : label is "4201080774605AE8432B41B76D8B60420A6456E930B72CD881021048416D7B50";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFD428125DE111400020400088000269125D5D4B94C";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF4100880000000000E01F11FF0909091555555555403807C47FC242424";
    attribute INIT_30 of inst : label is "D9090660584F09E55A2112D765A6C94CE01E93394A0C2BE47B0035D151660B4B";
    attribute INIT_31 of inst : label is "4B36B8AEACE6900547ACBDFF8B8271BFB0E09C4CCB3B0770BCD5328164D84C96";
    attribute INIT_32 of inst : label is "6222599A888AD2821032412524CA45A26E5B39871868A132D61A65A1A621A608";
    attribute INIT_33 of inst : label is "000000000000000000000000000369822DAE08B6B8202026808002000A5D0866";
    attribute INIT_34 of inst : label is "0B2518500000CC946828807FA5051F2A000AA0902AC0636363630381C0000000";
    attribute INIT_35 of inst : label is "4972643900B60000001EA0D367BD57A835F9EFFFE28B31D66520A3F460740822";
    attribute INIT_36 of inst : label is "FE2B01A5BF7B6B2E7E6B42ABB6CD938C0081912B58CA5591C9224962D6C2ADB6";
    attribute INIT_37 of inst : label is "2B290880504A0000000429A76D404804828A28A90D04D6400022288EFBEFBEFB";
    attribute INIT_38 of inst : label is "70E1CD19016BCD6D235561A293580009004C0201261100AA1404052B29008045";
    attribute INIT_39 of inst : label is "00000040C0001000102000000042001020010404CC12AB420413102204408824";
    attribute INIT_3A of inst : label is "C0B10C2242C088CC522967A99DE996ADFDC1232323331450031050C408101041";
    attribute INIT_3B of inst : label is "4201080774605AE8432B41B76D8B60420A6456E930B72CD881021048416D7B50";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFD428125DE111400020400088000269125D5D4B94C";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF4100880000000000E01F11FF0909091555555555403807C47FC242424";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "0425910928D11A2548224D0C9A193432234FF8D84E0190B1C7642BEDEDE23939";
    attribute INIT_01 of inst : label is "0EC80CC1D3055551040D57181C993C008E40C866410341600214781413FB3B69";
    attribute INIT_02 of inst : label is "39998CCC666D9BDB7BC96CB0B375B084DB36EB5D436E0DEDAD72CB172CB72CE5";
    attribute INIT_03 of inst : label is "000000000000000000000000025B6A93CDAA4F36A93644B8C810934847050B33";
    attribute INIT_04 of inst : label is "B09AE7A80000306B862888001AFACA80000008020B46A1C1C1C11A8946000000";
    attribute INIT_05 of inst : label is "272B6DCC9F592000001E82009FF7FFA08007FDFFE8A0C7799F8228019FDFE088";
    attribute INIT_06 of inst : label is "FF446347CB94840404041176CB320C79B64E65D4C133886A2599652D811F0209";
    attribute INIT_07 of inst : label is "849463358057FFFFFFB425D410110020014514590B020880007FFFFEFBEFBEFB";
    attribute INIT_08 of inst : label is "264CC8CCF400C553440471595860000DB731ACD698C66B2AAC96F084946B35B0";
    attribute INIT_09 of inst : label is "3FF1FFF1FF8FFC7FFC7FE3FFFF8FF3F8FF3F8D044531B56397595A6B4D69AD0B";
    attribute INIT_0A of inst : label is "903E8813AA5040232994C11660960000FCC0031121201841C70400CC183030C3";
    attribute INIT_0B of inst : label is "630D8C789A05270C641CDE01827093633013330FD781C3680C9B19AC66FBCE74";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3F4508422BD4911326224CC488BA5FC044CE0E2B";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF5400AA0000000000E01FFAFF090909C000000000003807FEBFC242427";
    attribute INIT_10 of inst : label is "0425910928D11A2548224D0C9A193432234FF8D84E0190B1C7642BEDEDE23939";
    attribute INIT_11 of inst : label is "0EC80CC1D3055551040D57181C993C008E40C866410341600214781413FB3B69";
    attribute INIT_12 of inst : label is "39998CCC666D9BDB7BC96CB0B375B084DB36EB5D436E0DEDAD72CB172CB72CE5";
    attribute INIT_13 of inst : label is "000000000000000000000000025B6A93CDAA4F36A93644B8C810934847050B33";
    attribute INIT_14 of inst : label is "B09AE7A80000306B862888001AFACA80000008020B46A1C1C1C11A8946000000";
    attribute INIT_15 of inst : label is "272B6DCC9F592000001E82009FF7FFA08007FDFFE8A0C7799F8228019FDFE088";
    attribute INIT_16 of inst : label is "FF446347CB94840404041176CB320C79B64E65D4C133886A2599652D811F0209";
    attribute INIT_17 of inst : label is "849463358057FFFFFFB425D410110020014514590B020880007FFFFEFBEFBEFB";
    attribute INIT_18 of inst : label is "264CC8CCF400C553440471595860000DB731ACD698C66B2AAC96F084946B35B0";
    attribute INIT_19 of inst : label is "3FF1FFF1FF8FFC7FFC7FE3FFFF8FF3F8FF3F8D044531B56397595A6B4D69AD0B";
    attribute INIT_1A of inst : label is "903E8813AA5040232994C11660960000FCC0031121201841C70400CC183030C3";
    attribute INIT_1B of inst : label is "630D8C789A05270C641CDE01827093633013330FD781C3680C9B19AC66FBCE74";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3F4508422BD4911326224CC488BA5FC044CE0E2B";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF5400AA0000000000E01FFAFF090909C000000000003807FEBFC242427";
    attribute INIT_20 of inst : label is "0425910928D11A2548224D0C9A193432234FF8D84E0190B1C7642BEDEDE23939";
    attribute INIT_21 of inst : label is "0EC80CC1D3055551040D57181C993C008E40C866410341600214781413FB3B69";
    attribute INIT_22 of inst : label is "39998CCC666D9BDB7BC96CB0B375B084DB36EB5D436E0DEDAD72CB172CB72CE5";
    attribute INIT_23 of inst : label is "000000000000000000000000025B6A93CDAA4F36A93644B8C810934847050B33";
    attribute INIT_24 of inst : label is "B09AE7A80000306B862888001AFACA80000008020B46A1C1C1C11A8946000000";
    attribute INIT_25 of inst : label is "272B6DCC9F592000001E82009FF7FFA08007FDFFE8A0C7799F8228019FDFE088";
    attribute INIT_26 of inst : label is "FF446347CB94840404041176CB320C79B64E65D4C133886A2599652D811F0209";
    attribute INIT_27 of inst : label is "849463358057FFFFFFB425D410110020014514590B020880007FFFFEFBEFBEFB";
    attribute INIT_28 of inst : label is "264CC8CCF400C553440471595860000DB731ACD698C66B2AAC96F084946B35B0";
    attribute INIT_29 of inst : label is "3FF1FFF1FF8FFC7FFC7FE3FFFF8FF3F8FF3F8D044531B56397595A6B4D69AD0B";
    attribute INIT_2A of inst : label is "903E8813AA5040232994C11660960000FCC0031121201841C70400CC183030C3";
    attribute INIT_2B of inst : label is "630D8C789A05270C641CDE01827093633013330FD781C3680C9B19AC66FBCE74";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3F4508422BD4911326224CC488BA5FC044CE0E2B";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF5400AA0000000000E01FFAFF090909C000000000003807FEBFC242427";
    attribute INIT_30 of inst : label is "0425910928D11A2548224D0C9A193432234FF8D84E0190B1C7642BEDEDE23939";
    attribute INIT_31 of inst : label is "0EC80CC1D3055551040D57181C993C008E40C866410341600214781413FB3B69";
    attribute INIT_32 of inst : label is "39998CCC666D9BDB7BC96CB0B375B084DB36EB5D436E0DEDAD72CB172CB72CE5";
    attribute INIT_33 of inst : label is "000000000000000000000000025B6A93CDAA4F36A93644B8C810934847050B33";
    attribute INIT_34 of inst : label is "B09AE7A80000306B862888001AFACA80000008020B46A1C1C1C11A8946000000";
    attribute INIT_35 of inst : label is "272B6DCC9F592000001E82009FF7FFA08007FDFFE8A0C7799F8228019FDFE088";
    attribute INIT_36 of inst : label is "FF446347CB94840404041176CB320C79B64E65D4C133886A2599652D811F0209";
    attribute INIT_37 of inst : label is "849463358057FFFFFFB425D410110020014514590B020880007FFFFEFBEFBEFB";
    attribute INIT_38 of inst : label is "264CC8CCF400C553440471595860000DB731ACD698C66B2AAC96F084946B35B0";
    attribute INIT_39 of inst : label is "3FF1FFF1FF8FFC7FFC7FE3FFFF8FF3F8FF3F8D044531B56397595A6B4D69AD0B";
    attribute INIT_3A of inst : label is "903E8813AA5040232994C11660960000FCC0031121201841C70400CC183030C3";
    attribute INIT_3B of inst : label is "630D8C789A05270C641CDE01827093633013330FD781C3680C9B19AC66FBCE74";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF3F4508422BD4911326224CC488BA5FC044CE0E2B";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF5400AA0000000000E01FFAFF090909C000000000003807FEBFC242427";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "8065D22B3803086558000085410A8215602FF1580E05500ACB2221C7C69138A9";
    attribute INIT_01 of inst : label is "188016E1C22695FDAABD06109904BA00811F2391411343400141701223FDE924";
    attribute INIT_02 of inst : label is "3111888C446E1B5B6B516DA1A154A84D01808050094405062142081420942084";
    attribute INIT_03 of inst : label is "00000000000000000000000003D9288944A2251288920314490F694794090A22";
    attribute INIT_04 of inst : label is "04600800000103803800000060002000000000002BC2E36363630381C0000000";
    attribute INIT_05 of inst : label is "272924889D65E000001EA22C684AAFA88A1A1201EA8C0CAEEAAAA20A212A0028";
    attribute INIT_06 of inst : label is "4555E00E81084001818046B40CA9046C95422D5AC0128C2865996504828D8414";
    attribute INIT_07 of inst : label is "00182914805ADB66DB3425F100000000029A69AD014041000020000000000000";
    attribute INIT_08 of inst : label is "14284884E820A24A02044E70584000049360A452B05229001496E000182914A0";
    attribute INIT_09 of inst : label is "37C9FFE1BE4FF86FF87F93FFFF0FC3E4DC3F4D000131142396515A6B4D69AD2E";
    attribute INIT_0A of inst : label is "101C0011021150220100906440A40204FCC01A01B0A01061041E794408101001";
    attribute INIT_0B of inst : label is "632D8CB11002162C6018D810004113631020322756904170087B18AC62908423";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF2201888421D6D557AEAB5DD6AAA1FA00CC4410E9";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFF00FF550000000000E01F50FF0909094000000000003807D43FC242425";
    attribute INIT_10 of inst : label is "8065D22B3803086558000085410A8215602FF1580E05500ACB2221C7C69138A9";
    attribute INIT_11 of inst : label is "188016E1C22695FDAABD06109904BA00811F2391411343400141701223FDE924";
    attribute INIT_12 of inst : label is "3111888C446E1B5B6B516DA1A154A84D01808050094405062142081420942084";
    attribute INIT_13 of inst : label is "00000000000000000000000003D9288944A2251288920314490F694794090A22";
    attribute INIT_14 of inst : label is "04600800000103803800000060002000000000002BC2E36363630381C0000000";
    attribute INIT_15 of inst : label is "272924889D65E000001EA22C684AAFA88A1A1201EA8C0CAEEAAAA20A212A0028";
    attribute INIT_16 of inst : label is "4555E00E81084001818046B40CA9046C95422D5AC0128C2865996504828D8414";
    attribute INIT_17 of inst : label is "00182914805ADB66DB3425F100000000029A69AD014041000020000000000000";
    attribute INIT_18 of inst : label is "14284884E820A24A02044E70584000049360A452B05229001496E000182914A0";
    attribute INIT_19 of inst : label is "37C9FFE1BE4FF86FF87F93FFFF0FC3E4DC3F4D000131142396515A6B4D69AD2E";
    attribute INIT_1A of inst : label is "101C0011021150220100906440A40204FCC01A01B0A01061041E794408101001";
    attribute INIT_1B of inst : label is "632D8CB11002162C6018D810004113631020322756904170087B18AC62908423";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF2201888421D6D557AEAB5DD6AAA1FA00CC4410E9";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFF00FF550000000000E01F50FF0909094000000000003807D43FC242425";
    attribute INIT_20 of inst : label is "8065D22B3803086558000085410A8215602FF1580E05500ACB2221C7C69138A9";
    attribute INIT_21 of inst : label is "188016E1C22695FDAABD06109904BA00811F2391411343400141701223FDE924";
    attribute INIT_22 of inst : label is "3111888C446E1B5B6B516DA1A154A84D01808050094405062142081420942084";
    attribute INIT_23 of inst : label is "00000000000000000000000003D9288944A2251288920314490F694794090A22";
    attribute INIT_24 of inst : label is "04600800000103803800000060002000000000002BC2E36363630381C0000000";
    attribute INIT_25 of inst : label is "272924889D65E000001EA22C684AAFA88A1A1201EA8C0CAEEAAAA20A212A0028";
    attribute INIT_26 of inst : label is "4555E00E81084001818046B40CA9046C95422D5AC0128C2865996504828D8414";
    attribute INIT_27 of inst : label is "00182914805ADB66DB3425F100000000029A69AD014041000020000000000000";
    attribute INIT_28 of inst : label is "14284884E820A24A02044E70584000049360A452B05229001496E000182914A0";
    attribute INIT_29 of inst : label is "37C9FFE1BE4FF86FF87F93FFFF0FC3E4DC3F4D000131142396515A6B4D69AD2E";
    attribute INIT_2A of inst : label is "101C0011021150220100906440A40204FCC01A01B0A01061041E794408101001";
    attribute INIT_2B of inst : label is "632D8CB11002162C6018D810004113631020322756904170087B18AC62908423";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF2201888421D6D557AEAB5DD6AAA1FA00CC4410E9";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF00FF550000000000E01F50FF0909094000000000003807D43FC242425";
    attribute INIT_30 of inst : label is "8065D22B3803086558000085410A8215602FF1580E05500ACB2221C7C69138A9";
    attribute INIT_31 of inst : label is "188016E1C22695FDAABD06109904BA00811F2391411343400141701223FDE924";
    attribute INIT_32 of inst : label is "3111888C446E1B5B6B516DA1A154A84D01808050094405062142081420942084";
    attribute INIT_33 of inst : label is "00000000000000000000000003D9288944A2251288920314490F694794090A22";
    attribute INIT_34 of inst : label is "04600800000103803800000060002000000000002BC2E36363630381C0000000";
    attribute INIT_35 of inst : label is "272924889D65E000001EA22C684AAFA88A1A1201EA8C0CAEEAAAA20A212A0028";
    attribute INIT_36 of inst : label is "4555E00E81084001818046B40CA9046C95422D5AC0128C2865996504828D8414";
    attribute INIT_37 of inst : label is "00182914805ADB66DB3425F100000000029A69AD014041000020000000000000";
    attribute INIT_38 of inst : label is "14284884E820A24A02044E70584000049360A452B05229001496E000182914A0";
    attribute INIT_39 of inst : label is "37C9FFE1BE4FF86FF87F93FFFF0FC3E4DC3F4D000131142396515A6B4D69AD2E";
    attribute INIT_3A of inst : label is "101C0011021150220100906440A40204FCC01A01B0A01061041E794408101001";
    attribute INIT_3B of inst : label is "632D8CB11002162C6018D810004113631020322756904170087B18AC62908423";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF2201888421D6D557AEAB5DD6AAA1FA00CC4410E9";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFF00FF550000000000E01F50FF0909094000000000003807D43FC242425";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
