-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_8N is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_8N is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_8N_0 : RAMB16_S2
	generic map (
		INIT_00 => x"0226064062606662206202226226062600000000000000000000000000000000",
		INIT_01 => x"2A41FFFF84D8FFFF0000FA05000057FF8901F90B0850FE9B86C8FFFFB921FFFF",
		INIT_02 => x"6662266266266662206242226226062626B9A420000C1C6E02C6702018006FF9",
		INIT_03 => x"FFFFFFFFFFFFFFFFFFFF0000FFF00000FFFF55F7FFFF7D1D0200FFFF322FFD88",
		INIT_04 => x"3FFF0FFFFFFFFFFF03F3BEEFFFFFC000FFFF5555FFFF5555FFFFFFFFFFF0FFF0",
		INIT_05 => x"FFFFFFFFFFFFFFFFFFFF0000FFFF0000FFF3BFF3FFFDFFF0FFC0FFE80FF0AFEC",
		INIT_06 => x"FFC3FFC3FFCFFFCFFFC3FFFFFFCFFF00FFFF000054000000FFFF0000FFFF0000",
		INIT_07 => x"FFFF0000FFFF057FFFC3FFC3FFC3FFC3FFC3FFFFFFC3FFFFFFFF0000FFFF0000",
		INIT_08 => x"FFFFDDDFFFFF7F000FC30FC3FFC3FFC30FC3FFFFFFC3FFFF0FFF0000FFFF0000",
		INIT_09 => x"C00001C04083080BE0C94258CE8B2040FFFF0000FFFF0000FFFF0000FFFF0000",
		INIT_0A => x"600208000040A0005A1844286828008800000081000081234000008410030003",
		INIT_0B => x"008012040410000230A0200852100000040001C00040002000010300C00002C1",
		INIT_0C => x"7000C882040211002420000084680400FFFF73D1FFE414106000010080046000",
		INIT_0D => x"424200080004008180801020C1820000FFFFF0DDFFFFF1CE4028006000200040",
		INIT_0E => x"18A40408100842324002000040C80000FFFF3F1FFFFF3D3C012008406A010600",
		INIT_0F => x"44080000400260000424080041810800FFFFA519FFFFC4051300000000000408",
		INIT_10 => x"66622662662666622062422262260626FFFF7007FFFF874A912600200842A012",
		INIT_11 => x"E26CFFFFBAE0FFFFB2B8FFFF62C9FFFF20622222622606262626266062606662",
		INIT_12 => x"000026EF00007F80B002FFFF0009FFFFB2B8FFFF62D9FFFFE221FFFFBAE2FFFF",
		INIT_13 => x"FFFDFFFDFFFDFFFD0000000000000000000000000000000000002FFF0000E200",
		INIT_14 => x"FFFFEABFFFFFFFFEABD5FFFF7EAFFFFF00000000000000000000000000000000",
		INIT_15 => x"04840484848084800484000084800480F000F00000000000F000F00000000000",
		INIT_16 => x"3FF53FF5555555553FF53FF555555555EBEBEBEBEBEBEBEBEBEBEBEBEBC0EBC0",
		INIT_17 => x"3FEB3FEAFEE3AAA0FFFFFFFFFF00FF00FFFFFFFF332C00005555AAAA5550AAA0",
		INIT_18 => x"FF0300AB0303AAAA0303AEAF03030000003003030003030305550AAA5555AAAA",
		INIT_19 => x"3B7B00007B787B78C30CC30C30C330C3C30CC30C30C330C3FF00FF0300300303",
		INIT_1A => x"0300000003000000030300007B787B78000000007B787B783B7B3B7B7B787B78",
		INIT_1B => x"FFFFFFFFFFFDFF20FFFFDF74FFFF775D00008E270000FFD00000000000000000",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FF00F00000000000AA80FD0000000000FFFFDFDFFFFFF7F7FFA8FFF400002D40",
		INIT_21 => x"07402AC157FD7D000007011FD5FFC005FD150B0755E0EE0021152F00FC000000",
		INIT_22 => x"7FF700047FF71B54FFD400002AA8055015145740000F00BF0000BE0002AA3FFF",
		INIT_23 => x"001F0000F4F00000800056A8F000000002400000000000005FD03C0000000030",
		INIT_24 => x"0000080000051FC0FF77BFFCEC530000FFFDFFFD555E07D4FFFF0015FA805557",
		INIT_25 => x"8FFF00FDFFFF015000000080454000000000000000280000AA00FFFFFFFFFFDD",
		INIT_26 => x"0000000100957FFF000A000020000E15500E02A0A0079BFF0003FF0077F7070F",
		INIT_27 => x"665C59BF7FF8FF422AAA03FFAAAAEAA000180000AA0A00010000000000180000",
		INIT_28 => x"0002008A020097D4000A5155AAA8800075C501E70DEAF9172D40681ED7FF8000",
		INIT_29 => x"06003FF8BDFF0000007E082803FF02A0BFBDDFBF8000EFBE5BDDEE204D540000",
		INIT_2A => x"0FD57DA2F82FA0AABBEF7F7B6EE7FC59A7F76AA0B79400000000000000000000",
		INIT_2B => x"057B7FD56AA8E9FFA8AE9AAAB8AAA6AABA2E1790AA000000AA80FFF3003001C5",
		INIT_2C => x"AA6AE8005BA900005578000000000000000000000000000000AAFFFF8022FFFF",
		INIT_2D => x"0AA500540A000A8002A900004A80000002C0D9990000E8F051FB7F5F7EE05749",
		INIT_2E => x"DFAAAAEFE9AA805400000000050000000020BF7E0802DF7BABBE2601B26A40AA",
		INIT_2F => x"7F7F2DD5EF3E6657000000005EFF00077FB9AEAA0002A1AA00020000BA8E000B",
		INIT_30 => x"0F00F00000000000400000000000000075DEFFFF5508FFEA5F81002AB59FFFCA",
		INIT_31 => x"FFFF0030CC0C0AAC0010FFF103C00000F3C003C00000000001C0D70000000000",
		INIT_32 => x"00FF0013FFFFFFFF00030003F4FFF3FFD55F03FEC00C0C0C000F000F0C0C0C0C",
		INIT_33 => x"0FDAFFFC8FF03FC0D0000000354017D7000000000F5003FF00000000003F000C",
		INIT_34 => x"FFF3ABFFFFF0F03C540005553C0C7C0CF300FFF803FF03F07FFF0FFFFD80503F",
		INIT_35 => x"3FF8000FE03FD000FFFFAFFFFFFFFFFF00000000000A000323FF7B3F0303EFEF",
		INIT_36 => x"AA070000F555025F02FFFFFFFFFFFFFFFFF5FFCC555530C3870D80077FD787DB",
		INIT_37 => x"FFFFAFAAFFFFAAAA0000015500005550071F57FFFFF4FFF5E1FFBFFF3FF6FFFF",
		INIT_38 => x"FD033C33CC00C7F83C33FC3CC03EC03F0FC003002AA00FC00000000003000000",
		INIT_39 => x"D030CEFE3FFAFF3F03FFFFFFFFFFFFFAC3FF43FFF3F3F0302FFFFFFDFC300000",
		INIT_3A => x"00000000F814000700000000007F0000FFFFFFFFFFFFFFFEFFFFFFFFF800E000",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE40F00030000D557EFDB00000000C3BEC17D",
		INIT_3C => x"FFFFFFFDFFFF76EEBFFF07FFFFFFFFFFFFFFFFFFFFFFFFFDFFFF47FFFFFFFFFF",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFF06FFFFFFFFFF05FF0000FFFF0011",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF77FFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8N_1 : RAMB16_S2
	generic map (
		INIT_00 => x"0226062222202220266622024624626600000000000000000000000000000000",
		INIT_01 => x"B88BFFFFFA0BFFFF0000D5FA00000005D205FFBF1819FFFF0382FFFFF23FFFFF",
		INIT_02 => x"2262624626262666066662024624626604D487C001F9406E29813C02E4007F44",
		INIT_03 => x"FFFFFFFFFFFFFFFFFFFF2222FFF02220FFFFA040FFFF00008B2BFFFFFBF44A22",
		INIT_04 => x"3FFF0FFFFFFFFFFF03F357FFFFFFE222FFFFAAAAFFFFAAAAFFFFFFFFFFF0FFF0",
		INIT_05 => x"FFFFFFFFFFFFFFFFFFFF2222FFFF2AAAFFF3FFF1F7FF5FF0FFC0355C0F107DD5",
		INIT_06 => x"FFC3FFC3FFCFFFCFFFC3DDDDFFCFDF77F540000000000000FFFF2222FFFF2222",
		INIT_07 => x"FFFF0000FFFF0000FFC3FFC3FFC3FFC3FFC3DDDDFFC3DDDDDFFF0000FFFF0000",
		INIT_08 => x"FFFF0000FFFF01000FC30FC3FFC3FFC30FC3DDDDFFC3DDDD0054000057FF0000",
		INIT_09 => x"55414070505F00230008400428870011FFFF0000FFFF0000FFFF0000FFFF000A",
		INIT_0A => x"471022184505AE26E028000801A2009080100420402201030404000100810043",
		INIT_0B => x"D173A22A14461A09400400002410010001012070000410002004204070100830",
		INIT_0C => x"04160000149198001142010118010001FFFF0C74FEE412082400108200000600",
		INIT_0D => x"04149046931004111820000002004000FFFF1D04FFFF1419200010018000A200",
		INIT_0E => x"11801080591102088040008423000000FFFF49C1FFFF9C010410204041A21048",
		INIT_0F => x"04000042044000244202008000100004FFFF0800FFFF04049016001004018010",
		INIT_10 => x"22626246262626660626620246246266FFFF0020FFFF09008148604092410080",
		INIT_11 => x"FFEFFFFFFFFBF73CFFFEFFFFFBFFFFFF26662202462462662266662226222622",
		INIT_12 => x"0000012400005800F318FFFFA39FFFFFFFFEFFFFFBFFFFFFFECBFFFFFFFFFFFF",
		INIT_13 => x"F22CF22CF22CF22C000000000000000000000000000000000000677F00005C00",
		INIT_14 => x"7FFFFAAFFFFFEBAB557FFFFF57AAFFFF00000000000000000000000000000000",
		INIT_15 => x"08480848484048400048000048400040FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_16 => x"3FF53FF5555555553FF53FF555555555FFFFFFFFFFFFFFFFFFFFFFFFFFC0FFC0",
		INIT_17 => x"3FEB3FEAFEF7AAA0FFFFFFFFFF00FF00FFFFFFFF73DC0000AAAA0000AAA00000",
		INIT_18 => x"FF0200FF0202FFFF0202FFFF0203000002020202020302030AAA0000AAAA0000",
		INIT_19 => x"07B70000B7B407B4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF02FF0202020202",
		INIT_1A => x"ABAA0000ABAA0000ABAB0003B7B4B7B400030003B7B4B7B437B737B7B7B4B7B4",
		INIT_1B => x"FFFFFFFFE5D8FFC0FFFF0000FFFF000000005FFF0000FD000000000000000000",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFF",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FC00700000000000FFC0F40000000000FFFF0802FFFF4004FFF9B7900000D000",
		INIT_21 => x"A400EFC35554F0000003AA83001F000AE0A82FE000102000459956C0A8000000",
		INIT_22 => x"FDF75DD6FFA70001FFF0000000010000FEA8EA00002F00548000FF000FFF3FFF",
		INIT_23 => x"000300004000000000000000CC2B0000040000000000000083C0FC0A4A208202",
		INIT_24 => x"00BA03E088000740FFF4FFF7B6DFF800FFFAFFFF8ABFEFFA05550008FFF807FF",
		INIT_25 => x"93FD00F4FF55000010000014000A2800800000000050000040FFFFFFFFFFFF35",
		INIT_26 => x"0012000B1192FFFFFFC5A088D08007FA03BF0BC0FEA037FF0E05FF00BBFF0291",
		INIT_27 => x"46587105FFF4FD013AAA00D4AAFF140000040000683700000000000000010000",
		INIT_28 => x"08002D55002000027ABD0300479F05E0C0005F6F0015A2000010C9870404F800",
		INIT_29 => x"E9E33F97D015AA0002BF815FEB5FC01569ABBE6AF800F8AE77B7ED407B400000",
		INIT_2A => x"0000CF7E546AAFBBEFA36AEEE6EFB9FBAEA2AA00B80000000000000000000000",
		INIT_2B => x"AA06F7AF017FDF7C2AAEAE8A2AAAEAA3AFA30000800000004220001F201FA840",
		INIT_2C => x"F82600001A4A000054055000000000000000000000000000004F3EFFF2FEFFFF",
		INIT_2D => x"0000454500A25415000800002800000062709F9D0000E7F0FEFFF7F7FB7AFEFD",
		INIT_2E => x"AE97F7BAFAD5A82A00000000005000018908EFFB625AFFEFF2054040FE7E2D40",
		INIT_2F => x"95F7037D5157F5DE0000000006590000D5A24AAEA9EEAAA3000000002A3A0000",
		INIT_30 => x"FA00F000000000000000000000000000C4827A11CBFE1054FBBA08061F76B555",
		INIT_31 => x"5FFF0030FC0C0FF1000CFF4000000000007003C00000000003804D0000000000",
		INIT_32 => x"01BF0007FFFFFFFF00030003F3FFF17F4FFF005FD60C0C0C000F000F0C0C0C0C",
		INIT_33 => x"FDBCFFF427703FC00000000000FF0D710000000000FF01FF00000000003F000C",
		INIT_34 => x"FFFA0000FAF938BC000005553E2C7E2CF30AF5D7A955ABF087FF0FFFFFC0801F",
		INIT_35 => x"0FFE00033E0D4000FFFFFFFFFFFFFFFF000A02AAABFFAAAB7CFF3FBFFFFFFFFF",
		INIT_36 => x"FFFF0000FFFF030F0C3F5D7FC30FD75FFF6FFFCEFFFFB0EB787EF800B0EB78BF",
		INIT_37 => x"FFFFFFFFFFFFFFFF0000000000000000C00003DF0000FDF0FE1F00FFFF6FFFC0",
		INIT_38 => x"F4333C33CC00CFD014137FF4C03C802B030000003FF007400000000003000000",
		INIT_39 => x"CFFFCFFFFFF7FFBF5BEB0000EBFF000003FF03FFF033F030FFFF1540FC300000",
		INIT_3A => x"00000000FF8200000000000000070000FFFFFFFFFFFFFFFFFFFFFFF6F8004800",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFFF7FFDF000F002500003FFFC14000000000C014C000",
		INIT_3C => x"FFFFFFFBFFF7EFEF1FFF046DFFFF7DFFFFFFFFFFFFFFF740FFFF045BFFFFFFFF",
		INIT_3D => x"FFFFD647FFFFFFFFFFFFFFFFFFFFD6FF7FFF07FFFFF7FFFF011D0000DFFF0000",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C98FFFF9DFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"0000000000000000FFFFFFFFDDDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8N_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0224262224220226262626266062666600000000000000000000000000000000",
		INIT_01 => x"FFEBFFFFBF9FFFFF0000028000007524C0D3FFFF34C2FFFF67D07FFFFAFFFFFF",
		INIT_02 => x"66626062662666222626622660626666010900758810025012400A081A00BE00",
		INIT_03 => x"FFFFFFFFFFFFFFFFFFFF3333FFF03330FFFF0000FFFF0000FFFFFF78FFD417FC",
		INIT_04 => x"0DFF0FF7FFFFFFFF0AA35555FFFFF333FFFF0000FFFF0000FFFFFFFFFFF0FFF0",
		INIT_05 => x"FFFFFFFFFFFFFFFFFFFF3333FFFF15557FF3FFF0EFFF0FF0EAA055542AA85554",
		INIT_06 => x"FFC3FFC3FFCFFFCFFFC3EEEEFFCFEF330000000000000000FFFF3333FFFF3333",
		INIT_07 => x"4FFF0000FFFF0000FFC3FFC3FFC3FFC3FFC3EEEEFFC3EEEE3FFF0000FF540000",
		INIT_08 => x"FFFF0000FFFF00000FC30FC3FFC3FFC30FC3EEEEFFC3EEEE00000000017F0000",
		INIT_09 => x"9C00855880834107840030920C830446FFFF0000FFFF0000FFFF0000FFFF0000",
		INIT_0A => x"022004000010006005298202122202008188D5450002955744C5454756451455",
		INIT_0B => x"00060000000400000401220000810120800454DD0200E565000044520C00501D",
		INIT_0C => x"0080008A000002022000100001120404FFFF0000DF4220158A6841442A8A5171",
		INIT_0D => x"940A00C0044011080020008004002040FFFF8140FFFF0040A82A1125488A0496",
		INIT_0E => x"48044000409652000010000002060000FFFF0010FFFF210182294514A4A61045",
		INIT_0F => x"04200000100404001000000800820000FFFD9124FDFF4A490A021411B20A2511",
		INIT_10 => x"666240426626662226266A2660626E66DFFF1040FFFF02088324010488628904",
		INIT_11 => x"FFFFDFD5FFFFC044FFFFFFFFFFFFFFF62626A626606266668A26262626622AA6",
		INIT_12 => x"00BE0000E0000000FFCFFFFFBFEFFFFFFFFFFFFFFFFFFFFFFFFFFFDCFFFFDC7F",
		INIT_13 => x"FABCFABCFABCFABC000000000000000000000000000000000000447600006000",
		INIT_14 => x"DAADFFAAED5DAFEAFFFFFFFFFFFFFFFF00000154000001540000000000000000",
		INIT_15 => x"04840484848084800004000084800000F000F00000000000F000F00000000000",
		INIT_16 => x"3FF51FF5555555553FF53FF555555555EBEBEBEBEBEBEBEBEBEBEBEBEBC0EBC0",
		INIT_17 => x"3FFB1FEAFEE1AAA0FFFF7FFFFF00FF00FFFFFFFF5104A0000000555500005550",
		INIT_18 => x"FF0300FF0303FFFF0303FFF00303000003030303030303030000055500005555",
		INIT_19 => x"007B00007B780078C30CC30C30C330C3C30CC30C30C330C3FF03FF0303030303",
		INIT_1A => x"0000000000000000000000007B787B78000000007B787B783B7B3B7B7B787B78",
		INIT_1B => x"FFFFFFFFFC80FFD0FFFF0000FFFF00000000BFFF002DD0000000000000000000",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF7FFFFFFFFFFFF",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"F400000000000000FFC0D00000000000FFFF0000FFFF00027FFE4103A8000000",
		INIT_21 => x"0001FFC357D04000880FFFFD0000007CFFF037FB0000F80024B8FFC000000000",
		INIT_22 => x"5F97B22A55BF20B8FFFC00002000000AFFFD5400003F0000F000FFC00FFF3FFF",
		INIT_23 => x"4000000000000000000300000ED00000000000000000000047F8FFFF8084DFFB",
		INIT_24 => x"005F001CFFC080005E65FD0B2DFFFC00FFFF4745FFFFD7150000000003FF001F",
		INIT_25 => x"41F200D0400000001E000000054000000000000000000000BBFFFFFFFFFFF500",
		INIT_26 => x"006603FF9BBAFFFF01708AAC00FA46540045FFF05550FFFF0A0055000FFF001E",
		INIT_27 => x"9ADF6000FFF005511EAA007FAAAA554000000000200100000000000000000000",
		INIT_28 => x"001040000000021401010382000088FE1FA8014008AA0000000099630000FF86",
		INIT_29 => x"D7FD13D040005700002FB800FFB8E8007FFB577DDBA0EF7BDD55B400F0000000",
		INIT_2A => x"0022D5DBAA00D6DEFABFFEFD9AEABF6EA2EAA400800000000000002100000820",
		INIT_2B => x"8A155F7B50A857FBABCA2ABEAAA2A82AA9FE0000000000008FBA0000F2AB05E0",
		INIT_2C => x"1FFFAA29FEFB0000A80A0000800000000000000000000000000580FBFBFFFD74",
		INIT_2D => x"002A5128A000AA00007F0000000000002470FFFF0000BFEABEA2EF7FDBA9BDEF",
		INIT_2E => x"ACAA7FFFFF4280AA000000000155000199B3FFFF639AFFFF00202AB80010AAA6",
		INIT_2F => x"754F005D7FBD5BDD0000000001B80000A8AB02A9AAA9AA8A000000000E2A0000",
		INIT_30 => x"F7F0C000000000000000000000000000B9B155FB7427EBAEF593BFADC46BDF5E",
		INIT_31 => x"0F0F00300C2C0FF0000FFC000000000000B803C000000000AAF08F0000000000",
		INIT_32 => x"D57F0003FFFF5CFF00030003F3FFF00F03FF000F000C0C0C000F000F0C0C0C0C",
		INIT_33 => x"DBFCFFD0BBB03FC0000000000AFF0FF00000000002FF00FF00000000001D002E",
		INIT_34 => x"FC0FFFFFAFAC3FFC055505557FFC7FFCF3AFF0C30C00FFF003FF2FFFFFC0C80F",
		INIT_35 => x"01FF00008F400000FFFF5555FFFF5555FFFF037FFFFF03030CFE1555EEEE5555",
		INIT_36 => x"000000020002EBAF0C3F0C3FC30FC30FFF00FFE100005F540787FE20FFFF07FF",
		INIT_37 => x"FFFF5555F50F5555AAAA0000ABFF0000C38A03CF28B0FCF0FFE1FE57F6FFF57F",
		INIT_38 => x"78333C33CC00C12CBC393FF3C03CC03F030000003FF003000000000001000000",
		INIT_39 => x"CEEEC555EFF055550EBE02A9BC0F7E178155C00050300030FFFF00F3FC10CC00",
		INIT_3A => x"00000000FFFF003F0000000000000000FFFFFFFFFFFFFFD5FFFFFDC0D02A0C00",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFFF10F30F0005000000001FFCC00000000000C228C33C",
		INIT_3C => x"FFFFFFFFFFFEFEFF27FF0000FFFF0527FFFFF764FFFF4000FFFF0004FFFF6D7F",
		INIT_3D => x"FFFF7D7FFFFFFFFFFFFFFFFEFFFFFEED0DFF22FFFF66FFFF0000000017FF0000",
		INIT_3E => x"FFFFFFFFFFFFFFFFEF77FFFF7F7CFFFFFFFFEFFBFFFFFBBBFFFFFFFFFFFFFFFF",
		INIT_3F => x"0000000000000000FFFFFFFFB7FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8N_3 : RAMB16_S2
	generic map (
		INIT_00 => x"0266066260064626266606646666666200000000000000000000000000000000",
		INIT_01 => x"FFFF7666FFFF7776000050280000246BC1A277F7791367E7FFFB677FFFFF767E",
		INIT_02 => x"666622266266206626660264666666620250004334004000C004081B03C2C560",
		INIT_03 => x"FFFFFFFFFFFFFFFFA06800001A000000FFFF0000FFFF0000FFFF6666FFE03216",
		INIT_04 => x"0FBF03F3FFFFFFFFEFFA000006810000FFFF0000FFFF0000FFFFFFFFFFF0FFF0",
		INIT_05 => x"FFFFFFFFFFFFFFFF06810000A0680000FFF3FFF0FFF00FF01FFD0000FFFD0000",
		INIT_06 => x"FFC3FFC3FFCFFFCFFAAFFFFFFA86FFF5000000000000000081A00000681A0000",
		INIT_07 => x"00570000FFFF0000FFC3FFC3FFC3FFC3FAAFFFFFFAAFFFFF07F5000040000000",
		INIT_08 => x"FFFF0000FFFF00030FC30FC3FFC3FFC32AAFFFFFFAAFFFFF0000000000000000",
		INIT_09 => x"A7B28007248B20034100200803020228FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0",
		INIT_0A => x"002EC41268220116012000206214080800800010004008038010200060038013",
		INIT_0B => x"9282110B9A08045900008008891208084308420700000A023446004847518007",
		INIT_0C => x"020244000882001A401242A000101008FFF90080F05000200006220000020406",
		INIT_0D => x"2700902020E100000000420000202002FFFF2049F7FF00829A20100010100018",
		INIT_0E => x"C2212010200080181000810008000A01FFFF8084FFFE8120440080188108010A",
		INIT_0F => x"84204080106014060000080040002008BFDC112292F3020A9208504002120509",
		INIT_10 => x"6666FAEF6266ABFE2666FFFF6666FFFF2D7C81407BD762120201080808800109",
		INIT_11 => x"FFFF9981FFFF0000FFFFFFFFFFFFFFF62666FFFE6666FEFA3266EFEE6206FEFE",
		INIT_12 => x"27FF0000FE400000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9987FFFF0124",
		INIT_13 => x"55545554555455540000000000000000000000000000000000A2000000000000",
		INIT_14 => x"FEF5FFFF55FFFFFFFFFFFFFFFFFFFFFF000055FE0000BD520000000000000000",
		INIT_15 => x"08480848484048400000000048400000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_16 => x"3FF50055555555553FF53FF555555555FFFFFFFFFFFFFFFFFFFFFFFFFFC0FFC0",
		INIT_17 => x"3FEA01EAAAA0AAA0FFFF07FFFF00FF00FFFFFFFF0000FFA05555AAAA5550AAA0",
		INIT_18 => x"FC000055000055550000555000000000020202020203020305550AAA5555AAAA",
		INIT_19 => x"00070000B7B40004FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF02FF0202020202",
		INIT_1A => x"000000000000000000030003B7B4B7B40003BFBFB7B4B7B437B737B7B7B4B7B4",
		INIT_1B => x"FFFFFFFFFFD0FFD0FFFF0000FFFF00000000DD458BF400000000BBBB0000BBBB",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"F000000000000000FF00C00000000000FFFFEFFFFFFFFEFFFFFD555440F90000",
		INIT_21 => x"0001FF6D5F400000FFBFFFD002AB000157E5FFB040000000F4D5FF0000000000",
		INIT_22 => x"401004000FBD155757FEABFEEB8A000FFFF00000003F0000F800FFC00FFFFFFF",
		INIT_23 => x"0000000000000000300100000400000000000000000000000F5DFFFF75FFFFFF",
		INIT_24 => x"0000EEFAE840BEAB2FF0FFEF0005FFFAFFFF02AAFFFFAA80000001FF007FF3E1",
		INIT_25 => x"00DB004AA800800003000000000000000015000056AA0000FFFFFD05FFFF5FFF",
		INIT_26 => x"AFFFFFFFFFFFFFFF0010FFFF0F65FFFF2F400A7C008E3FFF3F82000B3FFFEFA9",
		INIT_27 => x"1BAF8000FFD000000EAA003FAAFDF54000000000000C00000000000000000000",
		INIT_28 => x"00000000000800000080ABFF0000D55568D5A0A27D05AA0A00006B600000FFE0",
		INIT_29 => x"7E1000600000A12A00076DD8577F006A8BDEE757AAFBDB6D17BF000000000000",
		INIT_2A => x"0000BF7615C2B7ED656D6A6B777EA2E6AAB800000000000000008086000039A2",
		INIT_2B => x"D6BC77F6AA00FDFBAA1BAAFAAAAE6AAA2E30400000000000FF550A00FFFE0004",
		INIT_2C => x"015500A0000002800BC00000000000000000000000000000AEEA0007A555F400",
		INIT_2D => x"A800540005552AA0000000000000000061CDFFFF5EAAFFA8EF7D9EA6F7BFB7EB",
		INIT_2E => x"BAEE0000802A00000000000000AA0000B74EFFFFCD9EFFFF80A802AA0000A800",
		INIT_2F => x"DF9E0005EADFF6F70000000000290000A9AA01BE2AFAAA2E0000000000B80000",
		INIT_30 => x"F000C00000000000000000000000000008A089070020D857300F3401FA2008AA",
		INIT_31 => x"0FAF0030AC0E03C0AA0FF08000000000028403C000000000FF040F0000000000",
		INIT_32 => x"000F0003FFFFACFF00003FFF33FFC00F03FD000F0C0C0C0C000F000F0C0C0C0C",
		INIT_33 => x"BFFCFD002A803FC0000000003FFF0FF0000000000FFF003F00000000000C000C",
		INIT_34 => x"57FFFFF5FFFC3FFC0555A7557FFC7FFCF85FFAEBAC00FFF00BFFFFFFFFEACF83",
		INIT_35 => x"007F0000E10000007FFF0000FFFF0000FFFF033FFFFF0303A6FF0001CFCF1111",
		INIT_36 => x"0000002F002FFFFFFFFFAEBFFFFFEBAFFF88FFFF2082EABF0078FF867FFD00FF",
		INIT_37 => x"DFD4000000010000FFFF0000FFFF0000EAAA03EFAAAAFEF07FFE5FA32FFFFABF",
		INIT_38 => x"3C333C33CC00C03CFC3C0FC3C03E4017030000001FC003000000000000000000",
		INIT_39 => x"CCFC4444FFFA4000BFFFC000FFF50156C2AAC2A8A2B053F0FFFFAAF3D000CC00",
		INIT_3A => x"00000000007F00150000000000000000FFFFFFFFFFF7FFC3FFFFF400FFFF0C00",
		INIT_3B => x"FFFFFFFFFFFFFFFFFFFFD000FC00FFFF000000000FF4C33C00000002C33CC3BE",
		INIT_3C => x"FFFFFFFFFF76FFFF1FFF0000FFFF0001FFFF7400FFFF0000FFFF0000FFFF0001",
		INIT_3D => x"FFFFD7FFFFFFFFFFFFFFFFFBFFFFFEFB023F2FFFFFFEFFFF0000000005BF0000",
		INIT_3E => x"FFFFFFFFFFFFFFFFEF7EFFFFFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
