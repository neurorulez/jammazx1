library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"03",X"86",X"41",X"B5",X"33",X"85",X"37",X"0A",X"0A",X"85",X"8B",X"A2",X"4E",X"A9",X"06",X"A0",
		X"03",X"24",X"4E",X"70",X"04",X"A9",X"42",X"A0",X"0F",X"84",X"3E",X"20",X"76",X"68",X"A6",X"4F",
		X"86",X"3D",X"20",X"E4",X"7E",X"A5",X"27",X"85",X"2B",X"A5",X"28",X"85",X"2C",X"A6",X"37",X"BD",
		X"54",X"6C",X"85",X"8B",X"A2",X"47",X"A9",X"00",X"24",X"4E",X"70",X"04",X"A2",X"4E",X"A9",X"7E",
		X"20",X"76",X"68",X"20",X"A4",X"7E",X"A5",X"86",X"29",X"10",X"D0",X"0A",X"A0",X"03",X"B1",X"2B",
		X"29",X"0F",X"91",X"2B",X"10",X"1A",X"A9",X"65",X"A0",X"07",X"20",X"C9",X"7E",X"A6",X"37",X"BD",
		X"45",X"6C",X"0A",X"69",X"A4",X"A8",X"A9",X"57",X"20",X"C9",X"7E",X"A9",X"18",X"20",X"4F",X"7A",
		X"A6",X"41",X"CA",X"10",X"8C",X"60",X"18",X"65",X"8B",X"A8",X"8A",X"69",X"00",X"60",X"20",X"2D",
		X"7F",X"A2",X"00",X"A9",X"16",X"20",X"34",X"7A",X"A2",X"1C",X"A9",X"00",X"20",X"34",X"7A",X"A2",
		X"20",X"20",X"32",X"7A",X"A9",X"AD",X"20",X"57",X"7B",X"A9",X"17",X"4C",X"4F",X"7A",X"A5",X"90",
		X"F0",X"0F",X"C6",X"90",X"A2",X"08",X"20",X"32",X"7A",X"A9",X"95",X"20",X"57",X"7B",X"4C",X"29",
		X"7A",X"A8",X"A2",X"04",X"A9",X"02",X"24",X"97",X"10",X"0E",X"A5",X"AE",X"D0",X"11",X"A5",X"86",
		X"29",X"10",X"D0",X"0B",X"A9",X"01",X"A0",X"10",X"84",X"37",X"20",X"34",X"7A",X"A4",X"37",X"98",
		X"AA",X"A9",X"2F",X"4C",X"53",X"79",X"A5",X"90",X"F0",X"16",X"C6",X"90",X"A2",X"10",X"A9",X"06",
		X"20",X"34",X"7A",X"A2",X"08",X"20",X"32",X"7A",X"A9",X"95",X"20",X"57",X"7B",X"20",X"29",X"7A",
		X"A2",X"18",X"20",X"32",X"7A",X"A9",X"92",X"20",X"57",X"7B",X"A9",X"15",X"20",X"4F",X"7A",X"A5",
		X"62",X"29",X"0F",X"D0",X"20",X"A2",X"14",X"A9",X"07",X"24",X"62",X"50",X"0B",X"A9",X"08",X"20",
		X"34",X"7A",X"A2",X"2C",X"A9",X"0D",X"D0",X"07",X"20",X"34",X"7A",X"A2",X"28",X"A9",X"09",X"18",
		X"65",X"91",X"4C",X"34",X"7A",X"A2",X"24",X"A9",X"11",X"D0",X"F4",X"AB",X"69",X"79",X"69",X"84",
		X"69",X"8F",X"69",X"9F",X"69",X"DD",X"69",X"E6",X"69",X"04",X"6A",X"13",X"6A",X"22",X"6A",X"3A",
		X"6A",X"4E",X"6A",X"65",X"6A",X"74",X"6A",X"88",X"6A",X"9C",X"6A",X"B7",X"6A",X"CC",X"6A",X"D5",
		X"6A",X"F2",X"6A",X"1A",X"6B",X"C2",X"69",X"B5",X"69",X"93",X"69",X"E5",X"69",X"C9",X"69",X"CC",
		X"69",X"CF",X"69",X"D2",X"69",X"FF",X"64",X"03",X"65",X"D5",X"69",X"D9",X"69",X"00",X"18",X"06",
		X"36",X"3C",X"3C",X"12",X"00",X"BA",X"3C",X"00",X"66",X"2C",X"32",X"42",X"00",X"32",X"30",X"00",
		X"20",X"3E",X"1E",X"AC",X"32",X"3E",X"3C",X"00",X"32",X"20",X"00",X"20",X"3E",X"1E",X"AC",X"2C",
		X"32",X"3A",X"BC",X"00",X"20",X"3E",X"1E",X"2C",X"00",X"3E",X"30",X"26",X"3C",X"3A",X"80",X"26",
		X"30",X"3A",X"1E",X"38",X"3C",X"00",X"1A",X"32",X"26",X"30",X"BA",X"34",X"3E",X"3A",X"24",X"00",
		X"3A",X"3C",X"16",X"38",X"BC",X"3A",X"1E",X"2C",X"1E",X"1A",X"3C",X"00",X"32",X"34",X"3C",X"26",
		X"32",X"B0",X"00",X"34",X"32",X"26",X"30",X"3C",X"BA",X"0A",X"0C",X"82",X"0E",X"02",X"82",X"10",
		X"0C",X"82",X"14",X"02",X"82",X"04",X"0C",X"0C",X"82",X"04",X"12",X"02",X"82",X"34",X"1E",X"38",
		X"00",X"1A",X"32",X"26",X"B0",X"C4",X"16",X"3E",X"44",X"26",X"2C",X"26",X"16",X"38",X"46",X"00",
		X"20",X"3E",X"1E",X"2C",X"00",X"3C",X"16",X"30",X"2A",X"3A",X"00",X"1C",X"1E",X"3A",X"3C",X"38",
		X"32",X"46",X"1E",X"9C",X"1A",X"32",X"30",X"22",X"38",X"16",X"3C",X"3E",X"2C",X"16",X"3C",X"26",
		X"32",X"30",X"BA",X"46",X"32",X"3E",X"00",X"2C",X"16",X"30",X"1C",X"1E",X"1C",X"00",X"24",X"16",
		X"38",X"9C",X"3C",X"24",X"16",X"3C",X"00",X"42",X"16",X"3A",X"00",X"16",X"00",X"22",X"38",X"1E",
		X"16",X"3C",X"00",X"2C",X"16",X"30",X"1C",X"26",X"30",X"A2",X"3C",X"24",X"1E",X"00",X"1E",X"16",
		X"22",X"2C",X"1E",X"00",X"24",X"16",X"3A",X"00",X"2C",X"16",X"30",X"1C",X"1E",X"9C",X"3C",X"24",
		X"1E",X"00",X"1A",X"32",X"2C",X"3E",X"2E",X"18",X"26",X"16",X"00",X"24",X"16",X"3A",X"00",X"2C",
		X"16",X"30",X"1C",X"1E",X"9C",X"46",X"32",X"3E",X"00",X"24",X"16",X"40",X"1E",X"00",X"2C",X"16",
		X"30",X"1C",X"1E",X"9C",X"2C",X"26",X"20",X"1E",X"00",X"3A",X"3E",X"34",X"34",X"32",X"38",X"3C",
		X"00",X"26",X"3A",X"00",X"22",X"32",X"30",X"9E",X"46",X"32",X"3E",X"38",X"00",X"3C",X"38",X"26",
		X"34",X"00",X"26",X"3A",X"00",X"32",X"30",X"1E",X"00",X"42",X"16",X"C6",X"46",X"32",X"3E",X"00",
		X"16",X"38",X"1E",X"00",X"24",X"32",X"34",X"1E",X"2C",X"1E",X"3A",X"3A",X"2C",X"46",X"00",X"2E",
		X"16",X"38",X"32",X"32",X"30",X"1E",X"9C",X"1A",X"32",X"2E",X"2E",X"3E",X"30",X"26",X"1A",X"16",
		X"3C",X"26",X"32",X"30",X"00",X"3A",X"46",X"3A",X"3C",X"1E",X"2E",X"00",X"1C",X"1E",X"3A",X"3C",
		X"38",X"32",X"46",X"1E",X"9C",X"46",X"32",X"3E",X"00",X"1A",X"38",X"1E",X"16",X"3C",X"1E",X"1C",
		X"00",X"16",X"00",X"3C",X"42",X"32",X"00",X"2E",X"26",X"2C",X"1E",X"00",X"1A",X"38",X"16",X"3C",
		X"1E",X"B8",X"46",X"32",X"3E",X"00",X"28",X"3E",X"3A",X"3C",X"00",X"1C",X"1E",X"3A",X"3C",X"38",
		X"32",X"46",X"1E",X"1C",X"00",X"16",X"00",X"04",X"02",X"02",X"00",X"2E",X"1E",X"22",X"16",X"18",
		X"3E",X"1A",X"2A",X"00",X"2C",X"16",X"30",X"1C",X"1E",X"B8",X"3C",X"24",X"1E",X"38",X"1E",X"00",
		X"42",X"1E",X"38",X"1E",X"00",X"30",X"32",X"00",X"3A",X"3E",X"38",X"40",X"26",X"40",X"32",X"38",
		X"BA",X"1C",X"A5",X"02",X"4A",X"4A",X"4A",X"AA",X"BD",X"F2",X"76",X"85",X"46",X"0A",X"85",X"47",
		X"A6",X"01",X"BD",X"F6",X"76",X"85",X"0B",X"A5",X"02",X"29",X"0F",X"C9",X"09",X"90",X"04",X"49",
		X"0F",X"69",X"00",X"85",X"37",X"49",X"07",X"69",X"01",X"29",X"0F",X"AA",X"BD",X"E9",X"76",X"A4",
		X"0B",X"20",X"EF",X"70",X"85",X"58",X"A6",X"37",X"BD",X"E9",X"76",X"20",X"EF",X"70",X"85",X"59",
		X"60",X"A9",X"DA",X"A4",X"0B",X"30",X"08",X"A6",X"23",X"E0",X"02",X"D0",X"02",X"A9",X"90",X"20",
		X"EF",X"70",X"AA",X"A0",X"00",X"84",X"37",X"A0",X"07",X"20",X"C6",X"79",X"A8",X"4C",X"61",X"64",
		X"A5",X"5D",X"29",X"0F",X"F0",X"49",X"F8",X"A5",X"9E",X"38",X"E5",X"A2",X"AA",X"A5",X"9F",X"E5",
		X"A3",X"A8",X"A5",X"A0",X"E9",X"00",X"D8",X"90",X"36",X"F0",X"04",X"A2",X"99",X"A0",X"99",X"8A",
		X"D0",X"03",X"98",X"F0",X"2A",X"98",X"A4",X"AD",X"84",X"3A",X"A4",X"AE",X"84",X"3B",X"A0",X"00",
		X"84",X"A2",X"84",X"A3",X"20",X"63",X"64",X"A5",X"A2",X"A6",X"A3",X"24",X"97",X"30",X"04",X"A5",
		X"3A",X"A6",X"3B",X"85",X"95",X"86",X"96",X"05",X"96",X"F0",X"04",X"A9",X"7F",X"85",X"90",X"60",
		X"A5",X"0F",X"18",X"65",X"51",X"85",X"37",X"A5",X"10",X"65",X"4F",X"29",X"0F",X"A8",X"A2",X"03",
		X"86",X"41",X"B5",X"33",X"85",X"3A",X"0A",X"0A",X"AA",X"38",X"A5",X"37",X"FD",X"44",X"4E",X"85",
		X"38",X"98",X"FD",X"45",X"4E",X"90",X"12",X"D0",X"10",X"A6",X"3A",X"BD",X"54",X"6C",X"4A",X"4A",
		X"4A",X"AA",X"BD",X"63",X"6C",X"C5",X"38",X"B0",X"09",X"A6",X"41",X"CA",X"10",X"D2",X"A9",X"01",
		X"D0",X"05",X"A6",X"3A",X"BD",X"45",X"6C",X"A8",X"85",X"8E",X"20",X"76",X"75",X"88",X"D0",X"FA",
		X"F8",X"86",X"92",X"84",X"93",X"98",X"18",X"65",X"92",X"90",X"02",X"E6",X"93",X"C6",X"8E",X"D0",
		X"F5",X"85",X"92",X"D8",X"60",X"02",X"02",X"02",X"02",X"03",X"03",X"04",X"04",X"04",X"04",X"05",
		X"05",X"05",X"05",X"05",X"00",X"08",X"10",X"10",X"18",X"10",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"FF",X"80",X"40",X"20",X"68",X"A2",X"02",X"86",X"37",X"A9",X"00",X"85",X"5D",
		X"85",X"4D",X"85",X"49",X"B5",X"55",X"30",X"28",X"B5",X"5F",X"85",X"48",X"B5",X"5E",X"24",X"4E",
		X"70",X"0A",X"0A",X"26",X"48",X"26",X"49",X"0A",X"26",X"48",X"26",X"49",X"B5",X"5A",X"85",X"4C",
		X"B5",X"08",X"48",X"B5",X"07",X"AA",X"68",X"20",X"00",X"6D",X"A6",X"37",X"95",X"08",X"94",X"07",
		X"A9",X"00",X"85",X"49",X"8A",X"F0",X"02",X"A5",X"63",X"85",X"48",X"A9",X"80",X"85",X"4C",X"B4",
		X"5A",X"B5",X"5F",X"48",X"B5",X"5E",X"AA",X"68",X"20",X"FE",X"6C",X"A5",X"37",X"4A",X"AA",X"B5",
		X"58",X"85",X"48",X"B5",X"46",X"85",X"4C",X"A5",X"23",X"C9",X"02",X"D0",X"0C",X"A5",X"48",X"4A",
		X"18",X"65",X"48",X"85",X"48",X"90",X"02",X"E6",X"49",X"20",X"04",X"6D",X"48",X"8A",X"A6",X"37",
		X"95",X"5A",X"94",X"5E",X"68",X"95",X"5F",X"CA",X"CA",X"30",X"03",X"4C",X"6A",X"6C",X"60",X"86",
		X"4A",X"06",X"4A",X"2A",X"26",X"4A",X"2A",X"A8",X"A5",X"4A",X"2A",X"29",X"03",X"60",X"84",X"4D",
		X"85",X"4B",X"86",X"4A",X"A5",X"4C",X"45",X"4D",X"10",X"34",X"38",X"A5",X"4A",X"E5",X"48",X"A8",
		X"A5",X"4B",X"E5",X"49",X"90",X"16",X"D0",X"0D",X"C0",X"00",X"D0",X"09",X"85",X"4A",X"85",X"4B",
		X"85",X"4D",X"AA",X"A8",X"60",X"A6",X"4D",X"84",X"4A",X"85",X"4B",X"60",X"49",X"FF",X"AA",X"98",
		X"49",X"FF",X"A8",X"C8",X"D0",X"01",X"E8",X"8A",X"A6",X"4C",X"86",X"4D",X"90",X"E9",X"18",X"A5",
		X"4A",X"65",X"48",X"A8",X"A5",X"4B",X"65",X"49",X"90",X"DB",X"A9",X"FF",X"A8",X"B0",X"D6",X"20",
		X"84",X"66",X"A9",X"6B",X"85",X"69",X"A2",X"00",X"86",X"6A",X"A5",X"86",X"4A",X"B0",X"11",X"86",
		X"81",X"CA",X"86",X"79",X"86",X"7A",X"86",X"7D",X"86",X"7E",X"A0",X"07",X"A2",X"77",X"D0",X"11",
		X"A9",X"C0",X"85",X"81",X"CA",X"86",X"7B",X"86",X"7C",X"86",X"7F",X"86",X"80",X"A0",X"87",X"A2",
		X"77",X"20",X"B8",X"6F",X"A5",X"1D",X"18",X"65",X"51",X"A8",X"A5",X"1E",X"29",X"03",X"69",X"00",
		X"AA",X"98",X"38",X"E9",X"30",X"A8",X"8A",X"E9",X"00",X"B0",X"03",X"A0",X"00",X"98",X"24",X"4E",
		X"70",X"02",X"A0",X"00",X"84",X"38",X"85",X"39",X"18",X"65",X"4F",X"24",X"4E",X"70",X"08",X"29",
		X"0F",X"A0",X"E2",X"A2",X"51",X"D0",X"10",X"29",X"03",X"85",X"3A",X"A0",X"BC",X"A2",X"4B",X"24",
		X"38",X"10",X"04",X"A0",X"CE",X"A2",X"4B",X"86",X"2C",X"84",X"2B",X"0A",X"0A",X"A8",X"B1",X"2B",
		X"38",X"E5",X"53",X"85",X"1B",X"C8",X"B1",X"2B",X"29",X"0F",X"E5",X"54",X"85",X"1C",X"C8",X"B1",
		X"2B",X"38",X"E5",X"51",X"85",X"19",X"C8",X"B1",X"2B",X"29",X"03",X"E9",X"00",X"18",X"65",X"39",
		X"85",X"1A",X"A5",X"39",X"AA",X"0A",X"18",X"24",X"38",X"10",X"24",X"A5",X"3A",X"0A",X"A8",X"B9",
		X"07",X"78",X"85",X"2B",X"B9",X"08",X"78",X"85",X"2C",X"A0",X"00",X"E8",X"8A",X"0A",X"65",X"2D",
		X"91",X"69",X"A5",X"2E",X"69",X"00",X"C8",X"91",X"69",X"E6",X"69",X"E6",X"69",X"D0",X"0A",X"65",
		X"2D",X"85",X"2B",X"A5",X"2E",X"69",X"00",X"85",X"2C",X"A0",X"00",X"B1",X"2B",X"C8",X"AA",X"B1",
		X"2B",X"C8",X"C9",X"A0",X"90",X"3D",X"C9",X"D0",X"90",X"16",X"F0",X"03",X"4C",X"85",X"6F",X"C6",
		X"69",X"A0",X"00",X"B1",X"69",X"85",X"2C",X"C6",X"69",X"B1",X"69",X"85",X"2B",X"4C",X"2B",X"6E",
		X"85",X"37",X"98",X"18",X"65",X"2B",X"A0",X"00",X"91",X"69",X"86",X"2B",X"E6",X"69",X"A5",X"2C",
		X"69",X"00",X"91",X"69",X"E6",X"69",X"A5",X"37",X"29",X"0F",X"09",X"20",X"06",X"2B",X"2A",X"85",
		X"2C",X"D0",X"B6",X"86",X"3F",X"AA",X"B1",X"2B",X"85",X"3D",X"C8",X"B1",X"2B",X"C8",X"84",X"39",
		X"29",X"03",X"A8",X"8A",X"29",X"03",X"85",X"40",X"8A",X"6A",X"6A",X"6A",X"6A",X"85",X"4C",X"29",
		X"0F",X"85",X"41",X"A9",X"09",X"38",X"E5",X"41",X"AA",X"98",X"4A",X"66",X"3D",X"46",X"40",X"66",
		X"3F",X"CA",X"D0",X"F6",X"85",X"3E",X"A5",X"19",X"85",X"15",X"18",X"65",X"3D",X"85",X"19",X"A5",
		X"1A",X"85",X"16",X"65",X"3E",X"85",X"1A",X"24",X"4C",X"10",X"12",X"A5",X"3F",X"49",X"FF",X"AA",
		X"A5",X"40",X"49",X"FF",X"A8",X"E8",X"86",X"3F",X"D0",X"01",X"C8",X"84",X"40",X"A5",X"1B",X"85",
		X"17",X"18",X"65",X"3F",X"85",X"1B",X"A5",X"1C",X"85",X"18",X"65",X"40",X"85",X"1C",X"A5",X"1A",
		X"10",X"03",X"4C",X"80",X"6F",X"24",X"81",X"30",X"3F",X"A5",X"19",X"C5",X"1D",X"A5",X"1A",X"E5",
		X"1E",X"90",X"06",X"A9",X"80",X"85",X"81",X"B0",X"28",X"A5",X"1F",X"C5",X"1B",X"A5",X"20",X"E5",
		X"1C",X"90",X"7D",X"A9",X"80",X"85",X"81",X"A5",X"17",X"C5",X"1F",X"A5",X"18",X"30",X"12",X"E5",
		X"20",X"90",X"0E",X"20",X"6E",X"70",X"85",X"7A",X"84",X"79",X"8A",X"10",X"04",X"A9",X"8F",X"85",
		X"5D",X"A0",X"47",X"A2",X"77",X"20",X"B8",X"6F",X"A5",X"81",X"29",X"0F",X"D0",X"27",X"A5",X"19",
		X"C5",X"1D",X"A5",X"1A",X"E5",X"1E",X"90",X"48",X"20",X"22",X"70",X"24",X"81",X"70",X"07",X"85",
		X"7E",X"84",X"7D",X"4C",X"7F",X"6F",X"85",X"80",X"84",X"7F",X"A2",X"CF",X"86",X"81",X"A0",X"C7",
		X"A2",X"77",X"20",X"B8",X"6F",X"A5",X"1D",X"18",X"69",X"30",X"AA",X"A5",X"1E",X"69",X"00",X"E4",
		X"19",X"E5",X"1A",X"90",X"1A",X"A5",X"1B",X"C5",X"1F",X"A5",X"1C",X"30",X"13",X"E5",X"20",X"90",
		X"0F",X"20",X"6E",X"70",X"85",X"7C",X"84",X"7B",X"8A",X"30",X"04",X"A9",X"8F",X"85",X"5D",X"60",
		X"A4",X"39",X"4C",X"2B",X"6E",X"84",X"39",X"85",X"37",X"29",X"03",X"85",X"3F",X"A5",X"37",X"29",
		X"08",X"4A",X"85",X"38",X"8A",X"29",X"08",X"05",X"38",X"4A",X"4A",X"86",X"38",X"A8",X"8A",X"29",
		X"03",X"0A",X"06",X"3F",X"88",X"10",X"FA",X"85",X"3D",X"A5",X"37",X"4A",X"4A",X"6A",X"6A",X"85",
		X"4C",X"A9",X"00",X"85",X"40",X"4C",X"A4",X"6E",X"86",X"32",X"84",X"31",X"24",X"4E",X"70",X"26",
		X"A5",X"02",X"0A",X"A8",X"A2",X"00",X"B1",X"31",X"10",X"01",X"CA",X"18",X"65",X"0F",X"85",X"1D",
		X"8A",X"65",X"10",X"85",X"1E",X"C8",X"A2",X"00",X"B1",X"31",X"10",X"01",X"CA",X"18",X"65",X"0D",
		X"A8",X"8A",X"65",X"0E",X"D0",X"0C",X"A5",X"0F",X"85",X"1D",X"A5",X"10",X"85",X"1E",X"A4",X"0D",
		X"A5",X"0E",X"29",X"0F",X"85",X"20",X"84",X"1F",X"60",X"A5",X"19",X"38",X"E5",X"15",X"85",X"3D");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
