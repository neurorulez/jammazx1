-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "00005555000055550000555500005555000055550000555500005555616C2008";
    attribute INIT_01 of inst : label is "0CC00CC00C0C1D1D0FE11EF40E4A1B1E0FC31FD60F690FC30FC3163400005555";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFEFCDCCC3FBF3337FEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF0000000000000000FFFFFFFF3FE42AA8FFFFFFFF00000000";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5555000000000000";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_06 of inst : label is "123020081DD42A282BA92A280F78022031342A2813362AAA30302A2A0FC32028";
    attribute INIT_07 of inst : label is "1C8C03233234C8C03234C8C01C8C032310140000102000801F9728281E9C2A28";
    attribute INIT_08 of inst : label is "0DD1222A1DD408801D1C2A2A0FC328A80CC022281FD62AA80FC30A8200000000";
    attribute INIT_09 of inst : label is "0FC32A283FDF0A823FFF0A820C0C2A2A3CE40AA203032A2830302A2A1FD70A82";
    attribute INIT_0A of inst : label is "3FD70A820FD720000FC32A28303020201D942A280FD30AA20FC3282A0FC30880";
    attribute INIT_0B of inst : label is "80000000DAA2A222DA8A8000E40B1694302C080032342AAA1B1E20203A3C0A82";
    attribute INIT_0C of inst : label is "C4C0FCFC232B3337FFFFFFFF13333FFF4C4C0C0C313130305555000000000000";
    attribute INIT_0D of inst : label is "0000D8DC232333374103FFF34000FD3C13137EDFC8C0DCCCDDF9F7FBDDF9F7FF";
    attribute INIT_0E of inst : label is "C8C8CCC477F6303CFFFFFFFF2C8C480C1004FFFF3238302174ACDCCC1A3D3337";
    attribute INIT_0F of inst : label is "09110008406028081C0C01010CC0700008008EFF000040009FDD3C0C00003727";
    attribute INIT_10 of inst : label is "FFFFFFFF333303234900000102030233000D01015CCC404006200001300C4000";
    attribute INIT_11 of inst : label is "00000001FFFFFFFFC140380C0303E03C08008FCE0000C888301C3333DECCC8C0";
    attribute INIT_12 of inst : label is "DCCCC8C0FFFFFFFF33B703230020FFB2C080CC800061400000000000340CCCCC";
    attribute INIT_13 of inst : label is "000000004CC40880FFFFFFFF0020B3F2C8C03C0B0143702C340CCCCC00002223";
    attribute INIT_14 of inst : label is "CCC42339ECC800000303000001030203C040F3CFC888D7572CCC08C004043F7C";
    attribute INIT_15 of inst : label is "C040F3CFC888D757030300000103330FC3520888CCC800000303000021233331";
    attribute INIT_16 of inst : label is "D3F0ECCC0000F9F8000000000001000200000000EAABDFD60303000001030203";
    attribute INIT_17 of inst : label is "00000000000000000000000000000000CFF3BFFF0000362FFBF7CFCB0000EFFB";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000004880000000000000000FC0000000000";
    attribute INIT_19 of inst : label is "4C4C0C0C313130304C4C0C0C00000C0C31313030000030300C0C000030308880";
    attribute INIT_1A of inst : label is "0C0C0000C0800000C0C0000002030000FFFF0000FFFF00000203FC0000000000";
    attribute INIT_1B of inst : label is "1FD62AA84C4C0C0C000000000000000000000C0C35B930300000FC303030FC00";
    attribute INIT_1C of inst : label is "FFFF000055550000CCC800004440300C233300000111300CDCCCFCFC33373F3F";
    attribute INIT_1D of inst : label is "C000D555C000D555C000D555C000D555FFFFFFFFFFFFFFFFD4C4A8A8300C300C";
    attribute INIT_1E of inst : label is "00000000000000004C4C2C2C3131383800000000080020280C0C0C0C30303030";
    attribute INIT_1F of inst : label is "0003555700035557000355570003555700035557C000D5550C0C0C0C3030FC30";
    attribute INIT_20 of inst : label is "0D482F781332333D000000000000313C363C2223010383B34000C000C080F138";
    attribute INIT_21 of inst : label is "03300223333BEB882CC0F02C333EC000EB88003003230000E080B0E0F3320000";
    attribute INIT_22 of inst : label is "00133C1C0EC7EB8860203CCCCCC4C0003C3C3B3004400C0C0CC5000000003C1C";
    attribute INIT_23 of inst : label is "ECEC0000FFFFEB88000014044444C0003C3C3B3004400C0C333B022201030000";
    attribute INIT_24 of inst : label is "0040084024040791010202122090102400000000001400008880000000000000";
    attribute INIT_25 of inst : label is "00C0142401111119012020101004044402000000000000000040008400400000";
    attribute INIT_26 of inst : label is "0040084024040791010202122090102400220000000000000000000048400000";
    attribute INIT_27 of inst : label is "00C0142401111119012020101004044421100000000000000040000008408000";
    attribute INIT_28 of inst : label is "CCC4C1F1C040FBBF3B3844440000ECEC333F01011317EB88CCC4C1F1C040FBBF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "3FBF3F7F02330203E270C9F0CC80C0803CDC3C6C0E0B02033EBC353CE8B80000";
    attribute INIT_2B of inst : label is "0323011302330000FEFCFDFCCC80C0803FBF3F7F2E2B0203DCCCFCCCE0B0C080";
    attribute INIT_2C of inst : label is "0303000003033313FFFD2331C4C4FCEC0303031300000313FFFDDCCC0000FCEC";
    attribute INIT_2D of inst : label is "0CC100040000080A5777240C0000FEFC0CC100040000080A533706620000FCEC";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "B3B5333BBDBCCC00180CD88C4000CC00B3B5333BBDBC03CC3C9CC8884000C202";
    attribute INIT_31 of inst : label is "FBFFFFFF333341ACEFFCFFFCCCC041AC23BFFFFF7FF700A8C8ECFFFCFDF400A8";
    attribute INIT_32 of inst : label is "30243227000100335ECEECCC3E7E0033363C2223000180835ECEECCC3E7E33C0";
    attribute INIT_33 of inst : label is "3BFFFFFF331341ACEFFCFFFC4CC041AC23BFFFFF7DF700A8C8ECFFFCFD7400A8";
    attribute INIT_34 of inst : label is "033001013C0C011100C06040089040000F3301013C0C00084070604008901404";
    attribute INIT_35 of inst : label is "091101013C0C1028C0E06040089014040D0101013C0C0004C0F0604008902808";
    attribute INIT_36 of inst : label is "0F3301013C0C101440706040089028080D0101013C0C0008C0F0604008901404";
    attribute INIT_37 of inst : label is "0303000100002028C0C06018000000000B3301013C0C10284060604008901404";
    attribute INIT_38 of inst : label is "0303280900000000C0C0400000003C0C0303140500002028C0C0501400002808";
    attribute INIT_39 of inst : label is "2B0B00010000303CC4C44000000000001313000100000000E0E8400000003C0C";
    attribute INIT_3A of inst : label is "033001013C0C011100C06040089040000F3301013C0C00084070604408901404";
    attribute INIT_3B of inst : label is "091101013C0C1028C0E06040089014040D0101013C0C0004C0F0604008902808";
    attribute INIT_3C of inst : label is "0F3301013C0C101440706040089028080D0101013C0C0008C0F0604008901404";
    attribute INIT_3D of inst : label is "0303000100002028C0C06018000000000B3301013C0C10284060604008901404";
    attribute INIT_3E of inst : label is "0303280900000000C0C0400000003C0C0303140500002028C0C0501400002808";
    attribute INIT_3F of inst : label is "2B0B00010000303CC4C44000000000001313000100000000E0E8400000003C0C";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "AAAA0000AAAA0000AAAA0000AAAA0000AAAA0000AAAA0000AAAA00001CD00FBC";
    attribute INIT_01 of inst : label is "15552EE815152E2C14540FC311140CC015542FE910141FD715142B2BAAAA0000";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFFFFCCCCFFFF33337F7DE7DBFFF3FFFFDFFBFFFFFFFFFFFF";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF0000000000000000FFFFFFFF10042BFCFFFFFFFF382C0000";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000AAAA0000FFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_06 of inst : label is "2FEB300C262C0FC32EE8074333342BBA2B3A07432F692C6C3034303025380F86";
    attribute INIT_07 of inst : label is "C4C0313803132C4C03132C4CC4C0313800000000010204082F6903122D6823E3";
    attribute INIT_08 of inst : label is "262E0F872EEA0CC02E2E0C0C2DF80FD2272D0D852FE90FC3253C2FEB00000000";
    attribute INIT_09 of inst : label is "2F690FC30FC72FF30FD72FC30C0C0C0C0FD23DF8030307433A3A30300FC30FC3";
    attribute INIT_0A of inst : label is "0FC32FFF0FC33A3C0FC30FC33A3A30302D7807432FE93DF82F692FF22FE92EE8";
    attribute INIT_0B of inst : label is "000040000000C2220000C8882968D807333000082BBB2C4C0F0F30300FD72F7D";
    attribute INIT_0C of inst : label is "4000DCCC3FBF13335555FFFF0001373F0C0C8C8C303032320000AAAA0000FFFF";
    attribute INIT_0D of inst : label is "0000C0403FBF13330000C7F30000D8C400002737FCECCCC40000F7BF0000F7BF";
    attribute INIT_0E of inst : label is "BC6CC4C03B7AFABEFFFFFFFF00000C4C0000355C00003130DEB84CCC3EA73331";
    attribute INIT_0F of inst : label is "06220630809080800000280C0000002044C444C100000000ADECBEAF00000103";
    attribute INIT_10 of inst : label is "C573FFFF1BF3333B84C082C2313000100312222A84C0A8880110000404100820";
    attribute INIT_11 of inst : label is "00000000C57BFFFF0000CEC63131100244C444C10000544400002221CFD7ECCC";
    attribute INIT_12 of inst : label is "CFE4ECCCCD53FFFFD7F3333B131143110C4C0400031283920000000000000888";
    attribute INIT_13 of inst : label is "000000000000CCCCED53FFFF131143114C4C8004000093B30000488800001115";
    attribute INIT_14 of inst : label is "C040BC9C377E80000000000203330303AAA8FFFFFFFE00003CEC0CC800003D1C";
    attribute INIT_15 of inst : label is "AAA8FFFFFFFE0000030B0002000013070001FEFC7EFEC08023330000301C0333";
    attribute INIT_16 of inst : label is "E3F0F6FC0000DCCC0000000000020003BCEC0000FDDCC0410000000203330303";
    attribute INIT_17 of inst : label is "000000000000000000000000000000002FCFDFF700001333DFF3FC6F0000FFFF";
    attribute INIT_18 of inst : label is "04040000000040400101000000004440FC000000000001010000084544400000";
    attribute INIT_19 of inst : label is "0C0C8C8C303032320C0C8C8C0000CCCC70703232000033330C0C444030300000";
    attribute INIT_1A of inst : label is "0C0C4040ECC84040ECC80101233B4440FFFF0101FFFF4440233B084500000000";
    attribute INIT_1B of inst : label is "2FE90FC30C0C8C8C00000000000000000000CCCCFC30323200003B7730300845";
    attribute INIT_1C of inst : label is "000000000000AAAA340C000000009C8C301C000000003236C4C0FCFC03133F3F";
    attribute INIT_1D of inst : label is "EAAAC000EAAAC000EAAAC000EAAAC000FFFFFFFFFFFFFFFFE8E8C0C0300C300C";
    attribute INIT_1E of inst : label is "02224440022244400C0C8C8C38383232246C1111A84400000C0CCCCC30303333";
    attribute INIT_1F of inst : label is "AAAB0003AAAB0003AAAB0003AAAB0003AAAB0003EAAAC0000C0CCCCC30303B77";
    attribute INIT_20 of inst : label is "F2A41114010193B00000000000001C0C1333BDFD00006DCB800040004040D000";
    attribute INIT_21 of inst : label is "00102333333F1331F040323C333F4800133102030333000070C0F270F3330000";
    attribute INIT_22 of inst : label is "23291CCC01711331380CFCCC4040C8803E3C0CC000003C0C0040000000001CCC";
    attribute INIT_23 of inst : label is "7FFFEAAA1454DBB988808000000040003E3C0CC000003C0C1404002300002333";
    attribute INIT_24 of inst : label is "C04000C01222C00002010201440401200000300800000000CCC0000000000000";
    attribute INIT_25 of inst : label is "0C003000000004800300A84400001020010000000000000000000C4000008080";
    attribute INIT_26 of inst : label is "C04000C01222C000020102014404012003100000000000000000000044C00000";
    attribute INIT_27 of inst : label is "0C003000000004800300A84400001020102000000000000000000000040C4840";
    attribute INIT_28 of inst : label is "C0C2C0803C4CFFFFFCDC00000000C04013337FFF00001333C0C2C0803C4CFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "3FFF33370130233BF330C4C00000CCC00CCC33371D1423393FFCDCCC00002008";
    attribute INIT_2B of inst : label is "3333031300000002FFFCDCCC0C40ECC83FFF33370000233BCCCCDCCC1474ECC8";
    attribute INIT_2C of inst : label is "01010002000003034EC6BCDC0000FFFE3323000100000303FCDC44400000FFFE";
    attribute INIT_2D of inst : label is "0220000000000003393000000000F3320220000000000003030300000000F77E";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "3F7A777F989C6E6AA4F0C4C00000E4603F7A777F989C2F6FCCC4FFFE00006339";
    attribute INIT_31 of inst : label is "FFFF7FD70313360EFFFC7DF4C0409C0CFBFFFDFF03132A5EEFFCFF7CC040A85C";
    attribute INIT_32 of inst : label is "0F1A03130000091BADFCFDDD3626A9B91333BFFF00006CC9ADFCFDDD3626F9F8";
    attribute INIT_33 of inst : label is "3FFF7FF70313360EFFFCFDF4C0409C0CFBFFFFFF03132A5EEFFCFFFCC040A85C";
    attribute INIT_34 of inst : label is "033200080404032180C0100004404880033300080404033F808010000440CCC4";
    attribute INIT_35 of inst : label is "0622000804040732C0D010000440C4C40232000804041332C0C0100004408888";
    attribute INIT_36 of inst : label is "03330008040413328080100004408888023200080404033FC0C010000440CCC4";
    attribute INIT_37 of inst : label is "2B0B00000000323EC0C0000000009C8C0733000804040732809010000440C4C4";
    attribute INIT_38 of inst : label is "0303000000003236E0E8000000009C8C0303000000003236C0C0000000009C8C";
    attribute INIT_39 of inst : label is "030300000000323EC0C002020000A888030380800000222AC0C000000000BC8C";
    attribute INIT_3A of inst : label is "033200080404032180C0100004404880033300080404033F808010000440CCC4";
    attribute INIT_3B of inst : label is "0622000804040732C0D010000440C4C40232000804041332C0C0100004408888";
    attribute INIT_3C of inst : label is "03330008040413328080100004408888023200080404033FC0C010000440CCC4";
    attribute INIT_3D of inst : label is "2B0B00000000323EC0C0000000009C8C0733000804040732809010000440C4C4";
    attribute INIT_3E of inst : label is "0303000000003236E0E8000000009C8C0303000000003236C0C0000000009C8C";
    attribute INIT_3F of inst : label is "030300000000323EC0C002020000A888030380800000222AC0C000000000BC8C";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "3333333303030303FFFFFFFFFCFCFCFCCCCCCCCCC0C0C0C0000000002418241C";
    attribute INIT_01 of inst : label is "1DD50CC01D1D0C0C1EF40FE11B1E0E4A1FD60FC31A3C1FD71F9603213F3F3F3F";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFFFD40407FFF0101CBE3755DFFFB1004FFFB1004FFFF1004";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF0000000000005555FFFFFFFF8552C003FFFFFFFFAFFA3FFC";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000005555";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_06 of inst : label is "0761300C0C842F692EE82F691B3C033021302F6907632EEE30343A3A0F92252C";
    attribute INIT_07 of inst : label is "4CC8133223318CC423318CC44CC8133200000000012004800FC329380FC82B69";
    attribute INIT_08 of inst : label is "0C84272F0CC00CC00C0C2E2E0FD22DF80D85272D0FC32FE90F960FC300000000";
    attribute INIT_09 of inst : label is "0FC32F692FCF0FD32FFF0FC30C0C2E2E2DF01FF203032F6930303A3A0FC30FC3";
    attribute INIT_0A of inst : label is "2FC30FD70FC330140FC32F69303030300DD02F690FC31FF20FC32D7A0FC30CC0";
    attribute INIT_0B of inst : label is "800040008AA2E2228A8AC000A14A52853138080023312EEE0F0F30302F7D0FD7";
    attribute INIT_0C of inst : label is "C080FCEC373F0000FFFFFFFF02233FBF00000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000C8C8373700000002EFF30000F86C02022F9FDCC4000088A8F7BF88A8F7BF";
    attribute INIT_0E of inst : label is "9CCC000000C04000A00A00000000C080382C500500000203FCFC40403F3F0101";
    attribute INIT_0F of inst : label is "3F3F340CFCFC3C4C2E8F171FC040F4C44E47CEEB000000000300000100002323";
    attribute INIT_10 of inst : label is "00000000004000000C4000405FDE5676222B0003C000C0C023330227FBF4D040";
    attribute INIT_11 of inst : label is "000000000000000080006C4C5FDFF4644E47CECB0000DCCCC880FFFF03110000";
    attribute INIT_12 of inst : label is "010000000000000044C00000D1B1EBB3B7F59D9501300110888088800223BFFF";
    attribute INIT_13 of inst : label is "CCC43FFFF55DB13800000000D1B1E3B3FFF5391F000231390223FFFF00003337";
    attribute INIT_14 of inst : label is "C8C0363CBDDC00003FBFFFFF3A2E333F8000F7DFDDDC82023CCF0CC0333B3F3F";
    attribute INIT_15 of inst : label is "8000F7DFDDDC8202FFFFC73F23230FF38203DCDCDCDC4000FFFFCCCC0C8A3FBD";
    attribute INIT_16 of inst : label is "04040000733D0000FCDCCCC4377F3FBF14440000BFBECAC33FBFFFFF3A2E333F";
    attribute INIT_17 of inst : label is "3F7F03330000C2C2000383A3FDFDC4C01333000233330C043331DCCCF33B333E";
    attribute INIT_18 of inst : label is "FFFD00000000FFFEFFFF00000000FFFF7FFF00000000FFFF0000BFFFFFFF0000";
    attribute INIT_19 of inst : label is "00000000000000003333000000003333CCCC00000000CCCC0000FFFF0000FFFF";
    attribute INIT_1A of inst : label is "0000FFFE0000FFFE0000FFFF0000FFFF0000FFFF0000FFFF0000BFFF00000000";
    attribute INIT_1B of inst : label is "0000000033310000000047D102801004000033324CCC000000008CCC0000BFFF";
    attribute INIT_1C of inst : label is "AAAA0000000000009C8C00000000340C323600000000301CB0240001180E4000";
    attribute INIT_1D of inst : label is "03030303333333333F3F3F3F3FFF3FFFFFFFFFFFFFFFFFFF00000000300C300C";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFF33333333CCCCCCCCFDFCFFFF3F7FFFFF000033330000CCCC";
    attribute INIT_1F of inst : label is "3F3C3F3C3330333003000300FFFCFFFC00000000000000000000333200008CCC";
    attribute INIT_20 of inst : label is "580F3B3F03230203F0E4DCD4ECE8C8C0333937770002C4C00FDEFDDDFEEE8CC4";
    attribute INIT_21 of inst : label is "033300010333BB99840C4CCCFCFCC31CBB99033200030000CC0C1C0CFCFC050F";
    attribute INIT_22 of inst : label is "12303337342CBB99CCC8CCC00000D1153C3C3B7F382E1C0C342CEDF8B4C03337";
    attribute INIT_23 of inst : label is "C6C6BFFF0000BB99C4C0FEEE0002C0003C3C3B7F382E1C0C0313FDDCB4C00000";
    attribute INIT_24 of inst : label is "2818200F0002213208400C80000010C4000000000000040C0000221000000000";
    attribute INIT_25 of inst : label is "1011030000000132904C08000000E40C0000102000000230104C000000000000";
    attribute INIT_26 of inst : label is "2818200F0002213208400C80000010C4000000C8000000000200000000000210";
    attribute INIT_27 of inst : label is "1011030000000132904C08000000E40C00000303380C00000400300800000000";
    attribute INIT_28 of inst : label is "FFFF7F5DBBFFC111CCCB444088885754000055550202BBBFFFFF7F5DBBFFC111";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "00000000000000003FFC302C000000001333020200000000FFFCB8AC0000C4C0";
    attribute INIT_2B of inst : label is "3FFF3A2E00000313C00088800000C4C02CCC3A2C000003133330002000000000";
    attribute INIT_2C of inst : label is "28F1888800001C30ECCC00000000000028F0888800001C300000000000000000";
    attribute INIT_2D of inst : label is "3E0C000000007FFC00002008000014443E0C000000007FFC0CC0022200000000";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "B7F0777CBBBF00000000000080000000B7F0777CBBBF00000000000080000000";
    attribute INIT_31 of inst : label is "FEF8FFDF21130000BFF8FF7C4840000072F4FFD7299300008DF4FF7468600000";
    attribute INIT_32 of inst : label is "00000000000200000FDE3DDDFEEE000000000000000200000FDE3DDDFEEE0000";
    attribute INIT_33 of inst : label is "FEF8FFDF21330000BFF8FF7CC840000072F4FFD72B9300008DF4FF7468E00000";
    attribute INIT_34 of inst : label is "000303073FEF0203C000F880C808C000280803073FEF300CE8E8F880C8082888";
    attribute INIT_35 of inst : label is "3F3F07073FEF340C3C3CF440C80828882B2B03073FEF20282828F440C8083C4C";
    attribute INIT_36 of inst : label is "280803073FEF2028E8E8F440C8083C4C2B2B03073FEF300C2828F880C8082888";
    attribute INIT_37 of inst : label is "141413133F2F00001404E4ECF8FC14043C0C07073FEF340CFCFCF440C8082888";
    attribute INIT_38 of inst : label is "10143B1B3F2F10141414C4C4F8FC0000101413133F2F20281404C4C4F8FC2808";
    attribute INIT_39 of inst : label is "3C1C13133F2F00001404C7C7F8FC00001014D3D33F2F0000343CC4C4F8FC0000";
    attribute INIT_3A of inst : label is "000303073FEF0203C000F880C808C000280803073FEF300CE8E8F880C8082888";
    attribute INIT_3B of inst : label is "3F3F03073FEF340C3C3CF440C80828882B2B03073FEF20282828F440C8083C4C";
    attribute INIT_3C of inst : label is "280803073FEF2028E8E8F440C8083C4C2B2B03073FEF300C2828F880C8082888";
    attribute INIT_3D of inst : label is "141413133F2F00001404E4ECF8FC14043C0C03073FEF340CFCFCF440C8082888";
    attribute INIT_3E of inst : label is "10143B1B3F2F10141414C4C4F8FC0000101413133F2F20281404C4C4F8FC2808";
    attribute INIT_3F of inst : label is "3C1C13133F2F00001404C7C7F8FC00001014D3D33F2F0000343CC4C4F8FC0000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "11112222010102025555AAAA5454A8A844448888404080800000000001C40288";
    attribute INIT_01 of inst : label is "04402EE804043F3D05411ED60440199405413FFC05410FC305413E3E15152A2A";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFEFE8888BFBF22225555AAAAFFF72AAADFFF2AAAFFFF2AAA";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF5555AAAA0000AAAAFFFFFFFF6009D557FFFFFFFF5555BEBE";
    attribute INIT_04 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5555AAAA0000AAAA";
    attribute INIT_05 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_06 of inst : label is "3ABA2008377C0A822BA9020227702AAA3B3E02023B3C28283030202025690A82";
    attribute INIT_07 of inst : label is "9484212912166848121668489484212910140000100200083F3D02023C3C22A2";
    attribute INIT_08 of inst : label is "277B0A823FFE08803F3E08082DE90A82266808803FFC0A8225692AAA00000000";
    attribute INIT_09 of inst : label is "2F690A821FD72AA21FD72A820C0C08081EC628A8030302023A3A20201FD70A82";
    attribute INIT_0A of inst : label is "1FD72AAA0FD72A280FC30A823A3A20203D3C02022FF928A82F692AA22FE92AA8";
    attribute INIT_0B of inst : label is "0000000050008222500088886C299C16322400083ABE28081B1E20201A962A28";
    attribute INIT_0C of inst : label is "4440DCDC2BAB00005555FFFF1111377F00000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000D4542BAB00004101D7F34000DD9411117677E8E800005551F7FB5551F7FF";
    attribute INIT_0E of inst : label is "E868000044448880700DA00A00000440341CBAAE00000110FEEC88883BBF2222";
    attribute INIT_0F of inst : label is "000000000000000015552AAA4404B8A8019004D5000040001111022200001517";
    attribute INIT_10 of inst : label is "0020000008800000C18082832CEDA89911140101000040401737222AE574A888";
    attribute INIT_11 of inst : label is "000000010028000041409A862DEDE89A019005C4000040004440DDDD02020000";
    attribute INIT_12 of inst : label is "022000000800000080800000064057107B38662A0243C2828880800001117777";
    attribute INIT_13 of inst : label is "ECCCBD9D9999747428000000064013507B78B62B0141D2A60111777700000001";
    attribute INIT_14 of inst : label is "C444A999666A80003F7F7FFFFDDD373FEAE8FBEF6AAA55552EEE08C817373F7F";
    attribute INIT_15 of inst : label is "EAE8FBEF6AAA5555FFF7EB3F11156F7B4150EAE86EEA8080FFEFCCCCDDD5FF7F";
    attribute INIT_16 of inst : label is "08080000F7762424EEECCCC877757777A8A800006809D5543F7F7FFFFDDD373F";
    attribute INIT_17 of inst : label is "111523334000C1C1000153535444C8880332012113372119333E6C68D7F73B3D";
    attribute INIT_18 of inst : label is "FEFE00000000FDFDFFFF00000000FFFFBFBF00000000FFFF00007F7FFFFF0000";
    attribute INIT_19 of inst : label is "00000000000000003333000000003333CCCC00000000CCCC0000FFFF0000FFFF";
    attribute INIT_1A of inst : label is "0000FDFD0000FDFD0000FFFF0000FFFF0000FFFF0000FFFF00007F7F00000000";
    attribute INIT_1B of inst : label is "0000000032320000000088224551A82A000031318C8C000000004C4C00007F7F";
    attribute INIT_1C of inst : label is "555500005555AAAA644800004440988C21190000011132264918820224618082";
    attribute INIT_1D of inst : label is "010102021111222215152A2A15552AAAFFFFFFFFFFFFFFFF00000000300C300C";
    attribute INIT_1E of inst : label is "AAAAFFFFAAAAFFFF222233338888CCCCAAAAFFFFAAAAFFFF000033330000CCCC";
    attribute INIT_1F of inst : label is "15142A2811102220010002005554AAA800000000000000000000313100004C4C";
    attribute INIT_20 of inst : label is "A6E3277311018193C8C8C8C06C6CC4C41636AAAB01002889ACECECCC76764CCC";
    attribute INIT_21 of inst : label is "0332031203234320189CACCCFCCC61284322013100120000DC1C6C8CFCCC0A2C";
    attribute INIT_22 of inst : label is "0112232B391D43209DD5C4C0400060083E3C3FBE37772C0C391D9E8E1004232B";
    attribute INIT_23 of inst : label is "B9B87FFF140443200000EAEA000140003E3C3FBE37772C0C2B2B9FDD10040000";
    attribute INIT_24 of inst : label is "2210101B00011204282C480C00044C4810000000000008080000220000000000";
    attribute INIT_25 of inst : label is "23020100000020280C8004000000408800002208000120012800000000000000";
    attribute INIT_26 of inst : label is "2210101B00011204282C480C00044C480080080C000000000010000000002020";
    attribute INIT_27 of inst : label is "23020100000020280C80040000004088000000010C0000000008040000000000";
    attribute INIT_28 of inst : label is "3FFFBEAC7F7F6E6AC4450808C888ABAB00002AAA111573393FFFBEAC7F7F6E6A";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "00000000000000003EBC1D1C000020082323011100000002FEFC5D5C0000E888";
    attribute INIT_2B of inst : label is "3FBF35750000222BC04040400000C8801C9C3464000022292230011000000000";
    attribute INIT_2C of inst : label is "1494044000002C2C0CC00000000000001094044000002C2C0000000000000000";
    attribute INIT_2D of inst : label is "732C00040000FEEC0808140400002888732C00040000FEEC0CC0054100000880";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "3B3D333A9D9D222A00008080004000003B3D333A9D9D22280000808000400000";
    attribute INIT_31 of inst : label is "F9F47CE7120322026FF4BD3484008800A9B8FECB564702026AE83FB895148000";
    attribute INIT_32 of inst : label is "00000202010000007CECACCC7676A88800000202010000007CECACCC76762888";
    attribute INIT_33 of inst : label is "79F47CC7120322026FF43D3484008800A9B8FCCB564702026AE83F3895148000";
    attribute INIT_34 of inst : label is "00012A2A1D5F01134000A888D4D4C88014042A2A1D5F20081414A888D4D41404";
    attribute INIT_35 of inst : label is "00002A2A1D5F10100000A888D4D4140414142A2A1D5F10141414A888D4D40000";
    attribute INIT_36 of inst : label is "14042A2A1D5F10141414A888D4D4000014142A2A1D5F20081414A888D4D41404";
    attribute INIT_37 of inst : label is "2808222A151F10142028B89CF454000000002A2A1D5F10100000A888D4D41404";
    attribute INIT_38 of inst : label is "2808362E151F00002028A888F45414042808362E151F00002028B89CF4540000";
    attribute INIT_39 of inst : label is "0000222A151F10142220AB8BF45428080888E2EA151F20280000A888F4541404";
    attribute INIT_3A of inst : label is "00012A2A1D5F01134000A888D4D4C88014042A2A1D5F20081414A888D4D41404";
    attribute INIT_3B of inst : label is "00002A2A1D5F10100000A888D4D4140414142A2A1D5F10141414A888D4D40000";
    attribute INIT_3C of inst : label is "14042A2A1D5F10141414A888D4D4000014142A2A1D5F20081414A888D4D41404";
    attribute INIT_3D of inst : label is "2808222A151F10142028B89CF454000000002A2A1D5F10100000A888D4D41404";
    attribute INIT_3E of inst : label is "2808362E151F00002028A888F45414042808362E151F00002028B89CF4540000";
    attribute INIT_3F of inst : label is "0000222A151F10142220AB8BF45428080888E2EA151F20280000A888F4541404";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
