-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "3C003C000F000F553C2D3D781E0A0B5E3C0F3D5E1E2D3C0F3C0F05783D0C255E";
    attribute INIT_02 of inst : label is "0000000000000000FFFF2FF8FFFF2FF807D0000007D000000140000001400000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "061800000924000000002800000000000BDF000AF500A800004305F7FD40A000";
    attribute INIT_05 of inst : label is "00000000F000E0000F000BFFF000BFFF0BFF0002FF8000001FF4FFFF7FD0FFFC";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "C000D555C000C000000355570003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "002A0000003F003FAAAA0000F400FFFF2AAA00003FC03FFF0002000000000001";
    attribute INIT_0D of inst : label is "00000000000000002AAA00000000000702AA000003FD03FFAAAA00000000FFFF";
    attribute INIT_0E of inst : label is "00000000F03CF000F0F0F000F03CFFF8F000BFFF3E0F3C0F3D503FFFF055BFFE";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "00000000FFFCAAA8FFFFAAAAA4C3A02800000000000000000000000000000000";
    attribute INIT_12 of inst : label is "02FF0000FA00000000030FFF0000FFC00BF30000FFC00000000007E500000000";
    attribute INIT_13 of inst : label is "023C0A800DA000A007F53C0337D0C03C0BFF0000FFE00000000107FF0000FFD0";
    attribute INIT_14 of inst : label is "000C000000000000000000008000000003FF0000FFC0000001500FFF1500FFF0";
    attribute INIT_15 of inst : label is "000C000240000000000000040000400000670000FE00000000000000025067E0";
    attribute INIT_16 of inst : label is "F000C000FFFFFFFFFFFFFFFF03FF0FFF00000000FFFFFFFCFFFFFFFF3FFFFFFF";
    attribute INIT_17 of inst : label is "00000000000003FF000003FF00000000000000003CFCC3F00FCF3F0F00000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "C240C00001830003C2400A55018355A0C300C30000C300C33015C300540C00C3";
    attribute INIT_1B of inst : label is "000000000000000000005555000055555555000055550000C015C300540300C3";
    attribute INIT_1C of inst : label is "000000C0000003005555000055550000000030000000000C0A55000055A00000";
    attribute INIT_1D of inst : label is "00D5000057000000000000C100004300002500005800000000C000C003000300";
    attribute INIT_1E of inst : label is "000000C0000003000180000002400000540000C000150300000055570000D555";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000540000C0001503000025000058000000";
    attribute INIT_20 of inst : label is "02FF0FFF00030000FA00FFC0000000000BF307E500000000FFC0000000000000";
    attribute INIT_21 of inst : label is "023C3C0307F50A800DA0C03C37D000A00BFF07FF00010000FFE0FFD000000000";
    attribute INIT_22 of inst : label is "000C000000000000000000008000000003FF0FFF01500000FFC0FFF015000000";
    attribute INIT_23 of inst : label is "000001000000000000000000000000000075000000000000FE0067E002500000";
    attribute INIT_24 of inst : label is "000A0D4E054000008CC0C00000000000000A030E010000008CC0C00000000000";
    attribute INIT_25 of inst : label is "000A00CE054000008CC0C00000000000000A05CE054000008CC0C00000000000";
    attribute INIT_26 of inst : label is "0000003317000000373B15000000002A000303313000000073B05000000002A0";
    attribute INIT_27 of inst : label is "000A00000000000AFF0000000000A0000000003335000000373B15000000002A";
    attribute INIT_28 of inst : label is "0000D55A0007000000000000D57000000017000000007D5AD55A001700000000";
    attribute INIT_29 of inst : label is "3000BA00E1E1555500030003E1E355570CEA0C1D0DE10D55CC0007A2E1E15555";
    attribute INIT_2A of inst : label is "7A805FF500000000000055F001400000015F00000000FD5AF555000100008000";
    attribute INIT_2B of inst : label is "000000000000B4B4000000000000B4B7000000000000FDB4000000000000B4B4";
    attribute INIT_2C of inst : label is "0FFF3FE007FF000040000000E00000000000FFFF005F00000000FF54FF800000";
    attribute INIT_2D of inst : label is "0FFF3FEA07FF0000FFC00000FF40000000003FE007FF000000002FF0FF400000";
    attribute INIT_2E of inst : label is "0696003C0000000096903C00000000000696003C0000000096903C0000000000";
    attribute INIT_2F of inst : label is "000000000000000000000000000000000BFFFFFF1FF40002FF80FFFC7FD00000";
    attribute INIT_30 of inst : label is "3FFF1FF001FF0A02FFFCFF04FF4080A03FFF1FF001FF2028FFFCFF04FF402808";
    attribute INIT_31 of inst : label is "3FFF1FFF01FF0A02FFFCFFF4FF4080A03FFF1FFF01FF2028FFFCFFF4FF402808";
    attribute INIT_32 of inst : label is "3FFF10FF01FF0A02FFFC0FF4FF4080A03FFF10FF01FF2028FFFC0FF4FF402808";
    attribute INIT_33 of inst : label is "3FFF1FFF010F0A02FFFCFFF4F04080A03FFF1FFF010F2028FFFCFFF4F0402808";
    attribute INIT_34 of inst : label is "0202630C0000000080A0330C00000000AA82818C0000000080A0330C00000000";
    attribute INIT_35 of inst : label is "8280CD5300000000A0280CC3000000002A02958C0000000080A0330C00000000";
    attribute INIT_36 of inst : label is "0BDF05D50043000AFFF87FFCFD40A8000BFFFFFF0000002FFC00FF5400008000";
    attribute INIT_37 of inst : label is "0BDF05DE0043000A40000000F800A8000FE03FFC07FF00002FC0FFF0FF400000";
    attribute INIT_38 of inst : label is "0FFF3FFF017F0028FFE0CF50C100A0000000AAAA000000000000FFFD00000000";
    attribute INIT_39 of inst : label is "20003FF8017F00000020B250C10000000FFF3FFF07FF0000FFC0FFF0FF400000";
    attribute INIT_3A of inst : label is "005F000A017F002AF7E0DF50C100A0002FC03FFC017F00000FE0DB50C1000000";
    attribute INIT_3B of inst : label is "0BDF05F70043000AF500A000FD40A80001BF0FEC01C00000F7F00FFC00D00000";
    attribute INIT_3C of inst : label is "005F000A017F002AF7E0DF50C100A0002FC03FFC017F00000FE0DB50C1000000";
    attribute INIT_3D of inst : label is "0BDF05F70043000AF500A000FD40A80001BF0FEC01C00000F7F00FFC00D00000";
    attribute INIT_3E of inst : label is "005F000A017F002AF7E0DF50C100A0002FC03FFC017F00000FE0DB50C1000000";
    attribute INIT_3F of inst : label is "01BF0FEC01C00000F7F00FFC00D0000001BF0FEC01C00000F7F00FFC00D00000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "15553EA805550FA815503C0F01543C0015543EAD01503D5F05540AAF05501AF5";
    attribute INIT_02 of inst : label is "00000000000000001FF4FFFF1FF4FFFF00000BE000000BE00000028000000280";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000001400000000000FF502FF0000FFE00000027E0000BFA0";
    attribute INIT_05 of inst : label is "00000000D000F00007FF0F007FFFF000BFFF002FFFF8E00001407FFF0500FFF4";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "C000C000EAAAC00000030003AAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "003F00000000003FFFFF00000000FF503FFF000000003FF40003000000000000";
    attribute INIT_0D of inst : label is "000000000000000001FF00000000000003FF0000000003FFFFFF00000000D400";
    attribute INIT_0E of inst : label is "00000000FFF4FFF8FFFFF0F07FF4F03C7FFCF000FDFD3C0FFFFF3EA07FFFF0AF";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000F0F00000F0F000F000F000F000F000F000F0F0F00000F0F00000F0F00000";
    attribute INIT_11 of inst : label is "000000005554FFFC5555FFFFA8690CC3F000F000F000F000F000F0000000F0F0";
    attribute INIT_12 of inst : label is "0BFF002BFF80A000000007D400005F400FF90002CF40FF800000000000000000";
    attribute INIT_13 of inst : label is "2F0F01E3347CF3D000001E08000078BC0FFF02BFFFF0FE800000005700005500";
    attribute INIT_14 of inst : label is "000000020000000000000000140000000FFF00BEFFF0FE0000000FFD0000FFD0";
    attribute INIT_15 of inst : label is "000C000CE000E000000000000000000000060BFF7F80A0000000000000400FF0";
    attribute INIT_16 of inst : label is "F000C000FFFFFFFFFFFFFFFF03FF0FFF00000000FFFFFFFCFFFFFFFF3FFFFFFF";
    attribute INIT_17 of inst : label is "0000C000000000FF000000FF00000000000000000F3CF0F003CF0F0F00000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "C300C02A00C3A803C300302A00C3A80CC300C30000C300C305AAC180AA500243";
    attribute INIT_1B of inst : label is "0000AAAA0000AAAA0000AAAA0000AAAAAAAA0000AAAA0000C000C18000030243";
    attribute INIT_1C of inst : label is "0000001A0000A4000000000000000000000005AA0000AA5030000000000C0000";
    attribute INIT_1D of inst : label is "00C2000083000000000000EA0000AB0000C000000300000000C000C003000300";
    attribute INIT_1E of inst : label is "0000001A0000A40000C0A8000300002A00000240000001800000AAAB0000EAAA";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000AAAA0240AAAA018000C0000003000000";
    attribute INIT_20 of inst : label is "0BFF07D40000002BFF805F400000A0000FF9000000000002CF4000000000FF80";
    attribute INIT_21 of inst : label is "2F0F1E08000001E3347C78BC0000F3D00FFF0057000002BFFFF055000000FE80";
    attribute INIT_22 of inst : label is "000000000000000200000000140000000FFF0FFD000000BEFFF0FFD00000FE00";
    attribute INIT_23 of inst : label is "020000000000000000000000000000000007000000000BFF7F800FF00040A000";
    attribute INIT_24 of inst : label is "000C05C000000000C540000000000DC0000C030000000000C540000000000DC0";
    attribute INIT_25 of inst : label is "000C00C000000000C540000000000DC0000C0D4000000000C540000000000DC0";
    attribute INIT_26 of inst : label is "002A353B15000000330000000000003302A333B0100000003000000000000330";
    attribute INIT_27 of inst : label is "001F00000000001FF40000000000FE00002A173B150000003300000000000033";
    attribute INIT_28 of inst : label is "5A0017D50000000000005A0017C0000000000000000017D517D5000000005A00";
    attribute INIT_29 of inst : label is "3000AAAABEBE30000003AAABBEBF00030C730EAABEBE0CC04C00AAAABEBECB50";
    attribute INIT_2A of inst : label is "5557001500000000A800FDC000000000000000000000FF5515FF0000000057A8";
    attribute INIT_2B of inst : label is "000000000000EBEB000000000000EBEB000000000000EBEB000000000000EBEB";
    attribute INIT_2C of inst : label is "3FF41FFE001502BF000000005000F000AFFF07FF00000000FEAAFC005FF80000";
    attribute INIT_2D of inst : label is "3FFF1FFF001502BF5400FE805000FA003E001FFE0015000002F0FFD050000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "00000000000000000000000000000000BFFF7FFF0140002FFFF8FFF40500E000";
    attribute INIT_30 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_31 of inst : label is "3F0F0FFF00053FEFF0FCFFF05000FBFC3F0F0FFF00053EFEF0FCFFF05000BFBC";
    attribute INIT_32 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_33 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_34 of inst : label is "AB8C070600000000330C91A400000000180C6A4600000000330C91A400000000";
    attribute INIT_35 of inst : label is "CC33C6A1000000000CC3A46900000000C0CC6A4600000000330C91A400000000";
    attribute INIT_36 of inst : label is "0FFF027F000002FFFFF4FFF00000FFE0AFFF0555000002FFFEAA50000000F800";
    attribute INIT_37 of inst : label is "0FF40278000002FF0000E0000000F0003FF01FFF001502803FF0FFD050000A00";
    attribute INIT_38 of inst : label is "3FFF0FEF00000BFFDFF0ED800000FF8000000000000000000AAA17B000000000";
    attribute INIT_39 of inst : label is "3F800FEF000000000BF0ED80000000003FFF1FFF001502BFFFF0FFD05000FA00";
    attribute INIT_3A of inst : label is "00000AFE00000BFF5FF0BD800000FF803FF00FEF00000B0037F0FD8000000380";
    attribute INIT_3B of inst : label is "0FF5027E000002FF0000BFA00000FFE00ADB07F0000000833FFC03F40000FE80";
    attribute INIT_3C of inst : label is "00000AFE00000BFF5FF0BD800000FF803FF00FEF00000B0037F0FD8000000380";
    attribute INIT_3D of inst : label is "0FF5027E000002FF0000BFA00000FFE00ADB07F0000000833FFC03F40000FE80";
    attribute INIT_3E of inst : label is "00000AFE00000BFF5FF0BD800000FF803FF00FEF00000B0037F0FD8000000380";
    attribute INIT_3F of inst : label is "0ADB07F0000000833FFC03F40000FE800ADB07F0000000833FFC03F40000FE80";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "3C003C000F000F553C2D3D781E0A0B5E3C0F3D5E1E2D3C0F3C0F05783D0C255E";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "061800000924000000002800000000000BDF000AF550A80001BF0FF5FD40A000";
    attribute INIT_05 of inst : label is "00000000F000E0000F000BFFF000BFFF0BFF0002FF8000001FF4FFFF7FD0FFFC";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "C000D555C000C000000355570003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "002A0000003F003FAAAA0000F400FFFF2AAA00003FC03FFF0000000000000000";
    attribute INIT_0D of inst : label is "00000000000000002AA800000000000702AA000003FD03FFAAAA00000000FFFF";
    attribute INIT_0E of inst : label is "00000000F03CF000F0F0F000F03CFFF8F000BFFF3E0F3C0F3D503FFFF055BFFE";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "00000000C1435557C3307D5FA4C3A02800000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0004000010000000005702115400200000800000400000000000001805F01800";
    attribute INIT_13 of inst : label is "023C0A000DA000A005F53C0317D0C03C0000000000000000000100027D400000";
    attribute INIT_14 of inst : label is "00F3000AFFC0A8000001000FD000FC0000000000080000000001000080000000";
    attribute INIT_15 of inst : label is "000C000240000000005A00AE9400E80000000000600000000000000000000000";
    attribute INIT_16 of inst : label is "F000C000003FC0FF003F0C3003FF0FFC0000000003FFFFFC3C0FFFFF3FF0FFFF";
    attribute INIT_17 of inst : label is "FFF0FFC0FFFFFC00FFFFFC000003000FFF00FC00C3033C0FF030C0F0003F00FF";
    attribute INIT_18 of inst : label is "000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_19 of inst : label is "0000AAAA0000AAAA000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FF40FFFF01FFFFFFFF400AFF01FFFFA0FF00FF0000FF00FF3FFFFF00FFFC00FF";
    attribute INIT_1B of inst : label is "0000FFFF0000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFFFF00FFFF00FF";
    attribute INIT_1C of inst : label is "000000FF0000FF00FFFF0000FFFF000000003FFF0000FFFC0AFF0000FFA00000";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF00002F0000F800000000FF00FFFF00FF00";
    attribute INIT_1E of inst : label is "000000FF0000FF0001FFFFFFFF40FFFFFFFF00FFFFFFFF000000FFFF0000FFFF";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFFF00FFFFFFFF00002F0000F8000000";
    attribute INIT_20 of inst : label is "0004021100570000100020005400000000800018000000004000180005F00000";
    attribute INIT_21 of inst : label is "023C3C0305F50A000DA0C03C17D000A00000000200010000000000007D400000";
    attribute INIT_22 of inst : label is "00F3000F0001000AFFC0FC00D000A80000000000000100000800000080000000";
    attribute INIT_23 of inst : label is "7FF4010000002AA0000000000000000000000000000000006000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000D55A0007000000000000D57000000017000000007D5AD55A001700000000";
    attribute INIT_29 of inst : label is "3000BA00E1E1555500030003E1E355570CEA0C1D0DE10D55CC0007A2E1E15555";
    attribute INIT_2A of inst : label is "7A805FF500000000000055F001400000015F00000000FD5AF555000100008000";
    attribute INIT_2B of inst : label is "000000000000B4B4000000000000B4B7000000000000FDB4000000000000B4B4";
    attribute INIT_2C of inst : label is "0FFF3FE007FF000040000000E00000000000FFFF005F00000000FF54FF800000";
    attribute INIT_2D of inst : label is "0FFF3FEA07FF0000FFC00000FF40000000003FE007FF000000002FF0FF400000";
    attribute INIT_2E of inst : label is "3FFF1FFF01FF0A02FFFCFFF4FF4080A03FFF1FFF01FF2028FFFCFFF4FF402808";
    attribute INIT_2F of inst : label is "000000000000000000000000000000000BFFFFFF1FF40002FF80FFFC7FD00000";
    attribute INIT_30 of inst : label is "3FFF1F0F01FF0A02FFFCF0F4FF4080A03FFF1F0F01FF2028FFFCF0F4FF402808";
    attribute INIT_31 of inst : label is "3FFF1C0301FF0A02FFFCC034FF4080A03FFF1C0301FF2028FFFCC034FF402808";
    attribute INIT_32 of inst : label is "3FFF1F0F01FF0A02FFFCF0F4FF4080A03FFF1F0F01FF2028FFFCF0F4FF402808";
    attribute INIT_33 of inst : label is "3FFF1F5F00FB0A02FFFCF5F4EF0080A03FFF1F5F00FB2028FFFCF5F4EF002808";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0BDF0FD501BF000AFFF87FFDFD40A8000BFFFFFF0000002FFC00FF5400008000";
    attribute INIT_37 of inst : label is "0BDF0FD601BF000A40000000FE00AA000FE03FFC07FF00002FC0FFF0FF400000";
    attribute INIT_38 of inst : label is "0FFF3FFF017F002FFFE0CFF0FE40E00000000000000000000000FFFD00000000";
    attribute INIT_39 of inst : label is "38003FF8017F000000B092F0FE4000000FFF3FFF07FF0000FFC0FFF0FF400000";
    attribute INIT_3A of inst : label is "055F000A017F002AF7E05FF0FE40A0002FC03FFC017F00000FE0CBF0FE400000";
    attribute INIT_3B of inst : label is "0BDF0FF501BF000AF550A000FD40A8003EFF0FEC01F000A0F7F00FFC03D00000";
    attribute INIT_3C of inst : label is "055F000A017F002AF7E05FF0FE40A0002FC03FFC017F00000FE0CBF0FE400000";
    attribute INIT_3D of inst : label is "0BDF0FF501BF000AF550A000FD40A8003EFF0FEC01F000A0F7F00FFC03D00000";
    attribute INIT_3E of inst : label is "055F000A017F002AF7E05FF0FE40A0002FC03FFC017F00000FE0CBF0FE400000";
    attribute INIT_3F of inst : label is "3EFF0FEC01F000A0F7F00FFC03D000003EFF0FEC01F000A0F7F00FFC03D00000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "15553EA805550FA815503C0F01543C0015543EAD01503D5F05540AAF05501AF5";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000001400000000000FF502FF0000FFE000503DFE0000BFF0";
    attribute INIT_05 of inst : label is "00000000D000F00007FF0F007FFFF000BFFF002FFFF8E00001407FFF0500FFF4";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "C000C000EAAAC00000030003AAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "003F00000000003FFFFF00000000FF503FFF000000003FF40000000000000000";
    attribute INIT_0D of inst : label is "000000000000000001FF00000000000003FF0000000003FFFFFF00000000D400";
    attribute INIT_0E of inst : label is "00000000FFF4FFF8FFFFF0F07FF4F03C7FFCF000FDFD3C0FFFFF3EA07FFFF0AF";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000F0000000F0F0000000F000F0000000F000F0F000000000F00000F0F00000";
    attribute INIT_11 of inst : label is "00000000AAABC283BEAFC330A8690CC3F00000000000F000F000F000000000F0";
    attribute INIT_12 of inst : label is "00410000080000000000002B0000A1000100000030002000000000010000A300";
    attribute INIT_13 of inst : label is "2D0701E33478F3C000001E080000783C00000000000000000000000700006A00";
    attribute INIT_14 of inst : label is "003F00BDFF00FF80000000071400F40000000000030000000000000200000000";
    attribute INIT_15 of inst : label is "000C000CE000E000000000FF0000FC0000000002000000000000000000000000";
    attribute INIT_16 of inst : label is "F000C000C00F30FFC03F0C3C03FF0FFF00000000C3FFFFFC3C03FFFF3FFCFFFF";
    attribute INIT_17 of inst : label is "FFF03FC0FFFFFF00FFFFFF000003000FFF00FC00F0C30F0FFC30F0F0003F00FF";
    attribute INIT_18 of inst : label is "000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_19 of inst : label is "0000555500005555000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FF00FFFF00FFFFFFFF003FFF00FFFFFCFF00FF0000FF00FF05FFFF80FF5002FF";
    attribute INIT_1B of inst : label is "0000FFFF0000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFFFF80FFFF02FF";
    attribute INIT_1C of inst : label is "0000001F0000F400FFFF0000FFFF0000000005FF0000FF503FFF0000FFFC0000";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF0000FF0000FF00000000FF00FFFF00FF00";
    attribute INIT_1E of inst : label is "0000001F0000F40000FFFFFFFF00FFFFFFFF02FFFFFFFF800000FFFF0000FFFF";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFFF02FFFFFFFF8000FF0000FF000000";
    attribute INIT_20 of inst : label is "0041002B000000000800A1000000000001000001000000003000A30000002000";
    attribute INIT_21 of inst : label is "2D071E08000001E33478783C0000F3C0000000070000000000006A0000000000";
    attribute INIT_22 of inst : label is "003F0007000000BDFF00F4001400FF8000000002000000000300000000000000";
    attribute INIT_23 of inst : label is "074000000000FFFC000000000000000000000000000000020000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "5A0017D50000000000005A0017C0000000000000000017D517D5000000005A00";
    attribute INIT_29 of inst : label is "3000AAAABEBE30000003AAABBEBF00030C730EAABEBE0CC04C00AAAABEBECB50";
    attribute INIT_2A of inst : label is "5557001500000000A800FDC000000000000000000000FF5515FF0000000057A8";
    attribute INIT_2B of inst : label is "000000000000EBEB000000000000EBEB000000000000EBEB000000000000EBEB";
    attribute INIT_2C of inst : label is "3FF41FFE001502BF000000005000F000AFFF07FF00000000FEAAFC005FF80000";
    attribute INIT_2D of inst : label is "3FFF1FFF001502BF5400FE805000FA003E001FFE0015000002F0FFD050000000";
    attribute INIT_2E of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_2F of inst : label is "00000000000000000000000000000000BFFF7FFF0140002FFFF8FFF40500E000";
    attribute INIT_30 of inst : label is "3FD70F8200053FEFFD7CF8205000FBFC3FD70F8200053EFEFD7CF8205000BFBC";
    attribute INIT_31 of inst : label is "3DF70FAF00053FEFDF7CFAF05000FBFC3DF70FAF00053EFEDF7CFAF05000BFBC";
    attribute INIT_32 of inst : label is "3D7F082F00053FEFD7FC82F05000FBFC3D7F082F00053EFED7FC82F05000BFBC";
    attribute INIT_33 of inst : label is "3FFF0C0300053FEFFFFCC0305000FBFC3FFF0C0300053EFEFFFCC0305000BFBC";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0FFF3DFF005002FFFFFFFFF00000FFE0AFFF0555000002FFFEAA50000000F800";
    attribute INIT_37 of inst : label is "0FF43DF8005002FF0000E0000000F4003FF01FFF001502803FF0FFD050000A00";
    attribute INIT_38 of inst : label is "3FFF0FEF00000BFFDFF0EF7C0500FF8000000000000000000AAA17F000000000";
    attribute INIT_39 of inst : label is "3F800FEF000000000BF0EF7C050000003FFF1FFF001502BFFFF0FFD05000FA00";
    attribute INIT_3A of inst : label is "00000FFE00000BFF5FF0BF7C0500FF803FF00FEF00000BC037F0FF7C05000F80";
    attribute INIT_3B of inst : label is "0FF53DFE005002FF0000BFF00000FFE00FD307F00000027F3FFC03F40000FE80";
    attribute INIT_3C of inst : label is "00000FFE00000BFF5FF0BF7C0500FF803FF00FEF00000BC037F0FF7C05000F80";
    attribute INIT_3D of inst : label is "0FF53DFE005002FF0000BFF00000FFE00FD307F00000027F3FFC03F40000FE80";
    attribute INIT_3E of inst : label is "00000FFE00000BFF5FF0BF7C0500FF803FF00FEF00000BC037F0FF7C05000F80";
    attribute INIT_3F of inst : label is "0FD307F00000027F3FFC03F40000FE800FD307F00000027F3FFC03F40000FE80";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
