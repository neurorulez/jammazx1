-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "60A7C66AE1C8E920AAB4B8F8B8C0101494E352438C45C488080240710901C4A0";
    attribute INIT_01 of inst : label is "37D7D4675D9F3E7F59859C7F55A93010187581C75818693038DF3A11DAFFB61A";
    attribute INIT_02 of inst : label is "845028401F4FC11ED9E7273DDA3E836E8084043900392CF9B64DD30EB3871A4C";
    attribute INIT_03 of inst : label is "B64CC86BA984F242179CECC9449933212AA613C9085E63B2F71594F9C33823E1";
    attribute INIT_04 of inst : label is "22B31337A3B51B64CC86BA984F242029CECC9449933212AA613C9080A63B3B51";
    attribute INIT_05 of inst : label is "A75908420000601E800EACEEC0628F39FD24444244404046404641FDA3CFA38B";
    attribute INIT_06 of inst : label is "064B0FA199DD5C3B55DDEAABD1D99C18CD7417B15E2BE9D2C57A248A28A2800A";
    attribute INIT_07 of inst : label is "9FF58606FE44FE6343E38F75F71EE21F471F738FEE1C0EBC7A70E9C183B8F70E";
    attribute INIT_08 of inst : label is "171B8986E26C26E26C29804CB1FAC7CB9FAC7CBA17BF2583CE287E6BD64F9F97";
    attribute INIT_09 of inst : label is "387670C259C3816700A59771418F11393DF69DBFFFF878007879E661E660C336";
    attribute INIT_0A of inst : label is "E608EB7132CADC4CBAB7132CA55B8997429BA98052CBAC65CC05D53B4C099C32";
    attribute INIT_0B of inst : label is "A2DC290B18530545BBA49EE6310E0241C98B7212621C0486AC927D440A8C998B";
    attribute INIT_0C of inst : label is "C92AB87169B4E9A4C80626401004C164A27E78B04868B67BB4D121920C838C82";
    attribute INIT_0D of inst : label is "B9249EEC98581AA345A850AAA32675464CB3AA3265DD51932EBE763A493A6162";
    attribute INIT_0E of inst : label is "3260A8C9875F19D2CF3DDED24F765C2C1D5122C452AAA32635464CB2D8E39E7B";
    attribute INIT_0F of inst : label is "765C2C1D5122C452AAA3260A8C9865B1D42CF3DDC924F764C2C0D51A2C452AAA";
    attribute INIT_10 of inst : label is "9107DC305ACFCDBB28CF1ACB3384BAECF1ACB3384BAEF1050144F3CF3DDED24F";
    attribute INIT_11 of inst : label is "D6E2596F5D0FAA338F448748D06175A25CDCFD3FEBFB64F98555489E77FC90E3";
    attribute INIT_12 of inst : label is "1B426C25A0550BCF3D8044A114802383887C30E8415032820880461F12A3D6B0";
    attribute INIT_13 of inst : label is "F72DCF52D4B52EFDE5FB7DFCABCED1401A610F5A2AD55D0B7147F3273249925D";
    attribute INIT_14 of inst : label is "000076C924014992482974D692EC3401E6F2BD79474FC1E9192824C4A0723FAA";
    attribute INIT_15 of inst : label is "9216511C6A2C5E992BE1CB1C6EA29570E492439092C8E1566600055555566600";
    attribute INIT_16 of inst : label is "4AF4A1BD92C9AFE5DE4B64A0BDD2E9F2FA57A501EC965CC96C940C1ED8B97537";
    attribute INIT_17 of inst : label is "18FB773E25CB17F2902CD7D9ECF133B592E6C964B9AF3A5D2575774BAE064DDF";
    attribute INIT_18 of inst : label is "7FCAFF1E77E2B21BDFE733EDBA4F954B64509F4F672DD07F9AC73E6EFDC05327";
    attribute INIT_19 of inst : label is "0D0D0B29D805118853729514736D36190002A200325E5DCADABEF6D55B59FB84";
    attribute INIT_1A of inst : label is "3AA5DC9A2B8382DF0586348090FF0002A02A9CE7BAAD1007C031287B6BEFFDFC";
    attribute INIT_1B of inst : label is "66E99D864C5573E299B54CDD11EE6C08F33684799B367126DEEDAE3BA12D9F9F";
    attribute INIT_1C of inst : label is "0004000C0C0C0C200000000000000C1FF83FFFFD7A20361757FFFFD41AF15D4E";
    attribute INIT_1D of inst : label is "BF5971A7FCF5D33B0EA2A2A2A29A483050BBA8EEEE05B6AC2C0C2C0C2C0C2C00";
    attribute INIT_1E of inst : label is "A7D6A4850FA58575555554437F8FFBBF0A5D362F9ADD2E3BF686E359E648D6C7";
    attribute INIT_1F of inst : label is "0608AC043490DF9E42BC1D08411794E2060010064006D667EBA9FAEA6EBA9FAE";
    attribute INIT_20 of inst : label is "545400200004BAEE4000000000FFFCFEBFBF521621431298E77CB23C4EE3A0CB";
    attribute INIT_21 of inst : label is "70C80F22F3C8490112481820060879611D4408E0000441011044383CEE3C5119";
    attribute INIT_22 of inst : label is "71C80808F24841251008092112485B7B76C83FFFFFC841191008093012484301";
    attribute INIT_23 of inst : label is "62C43018C1844C21006408800A5C432170340F00F24849231048186012C879E1";
    attribute INIT_24 of inst : label is "71DCC6339E595DF00BDCBBEC87FFE600F87F0017B9370000000000318304582D";
    attribute INIT_25 of inst : label is "A013ED4B7028A9388A90A6365155EBE3170AAF735F0A0E6C924E7FC1FF6318CE";
    attribute INIT_26 of inst : label is "8ECE030C9E029F2F945515455054552549525415255154551705415147815497";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF5A450E07333929DA9E8D4FF9CAAB93D507672A";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "EDB1372C7E9E14029BB9B39BF32F635F26802020202023110243CCD92C90A208";
    attribute INIT_31 of inst : label is "8256493EC12D8DA1150B8570810A0ECA5266DB6B0EAB3709AEE648893FC9E4C7";
    attribute INIT_32 of inst : label is "82228280A80405B0D89140892DC04063492131AC00005000F32448880B6E6A50";
    attribute INIT_33 of inst : label is "312281125965B3EC490031414297635914111AA142862FF496CD111111111947";
    attribute INIT_34 of inst : label is "6EECD9A6975C47F936D71145022496CFB10066DC82CEB6CD8B389A028BA4B6DD";
    attribute INIT_35 of inst : label is "2772806CC999BBA7773A76E59CE0F4E32626CC2753806CC999BBA77C9B913626";
    attribute INIT_36 of inst : label is "BBA7773A74E59CE0F4E32626CC2753806CC999BBA777B876C59CC0E4E32626CC";
    attribute INIT_37 of inst : label is "2AB9ED2550B8E0929C0A371479012D97B876C59CC0E4E32626CC2772806CC999";
    attribute INIT_38 of inst : label is "DC00880FB4D34660237D007407666F68AC161AC5464CACB35519309D5010E0CC";
    attribute INIT_39 of inst : label is "2C9361A65F85B1A851606F924D93A16B096AC2AE30CB32D9481302867CAF7B04";
    attribute INIT_3A of inst : label is "99BBA7749EC933CF77DA49EEFB0F121433DD37896AB393214A4B5617797096AC";
    attribute INIT_3B of inst : label is "BEB9DFB42ADC90237FEE4F00C07D9A7624B278419CC0F4E32626CC2753806CC9";
    attribute INIT_3C of inst : label is "D5E080B9A114A22D409C9F5CAEEFB5B264A36F67515FAFE4A4CD3671D99D35A6";
    attribute INIT_3D of inst : label is "FFFFFDCCD6DE829D50703345263B814ED2D26826004D52B34B9A4C4B14C02E08";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "8B884DBC2E8E7F805554A1A32C3CDDC92AB0A4BAC29963E66EE49758F25D635F";
    attribute INIT_01 of inst : label is "5CBCBCD3804B4A01E270A30BFEC7C5BAA30A2A70A2A70AC54609BEA020EE7DA7";
    attribute INIT_02 of inst : label is "60AF561DC88C6A03A441425603915C139561A9064B083E46F59274E14528C2B1";
    attribute INIT_03 of inst : label is "C9BB369007730DB0151219137B22644A400CC412407E4864BF5A4D5530ED008C";
    attribute INIT_04 of inst : label is "93C1AD7FB4DCA59BB36B107730DB0001619377962644AC40CC412402A58644CA";
    attribute INIT_05 of inst : label is "649264D56DB6D5F6DB96E96E9AA7F06491B641864387844386438400F41F50D9";
    attribute INIT_06 of inst : label is "8214C05B283262D75D7D5D57254AB9D22BEAA065E160136597854D263C63C597";
    attribute INIT_07 of inst : label is "2D810602BEBABEBC779054C8E8A990CEAC40885519690512265C916058054CB4";
    attribute INIT_08 of inst : label is "E4A0D5E81581C83583C9325FBD24DC93D2CFCB376156C92E0067E0B20547E018";
    attribute INIT_09 of inst : label is "564AA4B9E2B2EFAAC47DA4AB733A8B94548D3657FFF87878007E0786078094C1";
    attribute INIT_0A of inst : label is "149F548C46952713A548C46B1EA4E2759F44C2733CD00B485B6837A497642924";
    attribute INIT_0B of inst : label is "6504721CD7382CCA004939DE1319B5B497E725FEE6336B6B7CE18AFBE073225C";
    attribute INIT_0C of inst : label is "327DC5D6B2CD164E65F1C2A4326306882490A214E021D5A00E1ACC2611046B16";
    attribute INIT_0D of inst : label is "02C928001B8313C08E48E4C01CC8B03991AD81CC8D6C0E646900A48A9283432C";
    attribute INIT_0E of inst : label is "CC8807323584568F34D2216DB4888DC389E0C774EED01CC8F03991AC269028A0";
    attribute INIT_0F of inst : label is "889DC399E04774EED01CC8807323480D69F1450032494001DC199E0C734E6C01";
    attribute INIT_10 of inst : label is "1E8845926223FA045F3CEF1A473BCEB3DE73AC779C6959C266232734D2232DB4";
    attribute INIT_11 of inst : label is "2C1CB69218E13C8631A1D5B47B5E5B538027FD7F3494A90025555AA113282A0E";
    attribute INIT_12 of inst : label is "40F81E147AEAA24E6A3677772DD906261A3F1461C9E02B940ACA068365BB092F";
    attribute INIT_13 of inst : label is "1000A5200A120344D6C9B492BF446DB5B05B708570C7DDC2782E8102101080DC";
    attribute INIT_14 of inst : label is "00110BB6DB2F972492C7A00404AD4202AA6F7417AF05B4628816C1F7EF1DC5FF";
    attribute INIT_15 of inst : label is "B85EAFBF8E497F53D468D8EF05754A361964B02F2413886C3B0A2D4454443B00";
    attribute INIT_16 of inst : label is "B98BBBF22613AA09109889BBF26E37048DC8DDDF9331913313376BB9877B8B9F";
    attribute INIT_17 of inst : label is "25469871C933A28529552863C60ED77CF7AD1309EB396DC6EE55D0B849DA0200";
    attribute INIT_18 of inst : label is "B8050FBFFC7E51A02718FA02009C2204888126918E63252A2CAA60100025AB5A";
    attribute INIT_19 of inst : label is "3218DB84E3748A2737E8CB76CD04D2CE4002280016ECD41B111F964B69140B1F";
    attribute INIT_1A of inst : label is "0FEBB237BB9D980F3B994E5DCDFF0008A08A408AFFF0BF6F8FCFCF9A6A183971";
    attribute INIT_1B of inst : label is "05AE18ACD2FAC81D640AA2039BD9038DEC8146F4408412B8122BF30A390CBC00";
    attribute INIT_1C of inst : label is "A880A0090909A9A000000000000009BFFA3FFFFA9A0053F25FFFFFDDFC8B27B3";
    attribute INIT_1D of inst : label is "FEB25E0381F35C315ACC44CC4CEAAD4CA768CCA3E8CE42E02020000020200008";
    attribute INIT_1E of inst : label is "D9BDDAC99636499AAAAAAEFFB7A2F01F1CF2D27565965455215CBCD2E0540A4E";
    attribute INIT_1F of inst : label is "39A17CFFD16F6C0FBBFCEB99AB325C54052814A044A214B9A4F6293D8A4F6693";
    attribute INIT_20 of inst : label is "986500000000BFBEBFBBBBBBBBAAAA015A01104B509B260367CCF44606A76757";
    attribute INIT_21 of inst : label is "0108220060881C10070820708828100007052C4088250804220D2894AA2D6181";
    attribute INIT_22 of inst : label is "808820906008041881281B6376E80000000812426488041C0128239878E80410";
    attribute INIT_23 of inst : label is "A145000000050800014D2310702D04000100221060081C7200E8208078081040";
    attribute INIT_24 of inst : label is "B79F6D634E79DA7E95573EFCC9879E7FAEF5DD2AAE3D20000000082522452814";
    attribute INIT_25 of inst : label is "C0394BEF8166E3406B8924F6956C2280C5018AF250F4EDBCEDADA196007DB5AF";
    attribute INIT_26 of inst : label is "164A0003948197189445014451140521405214850150501507014052A80D6A17";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF7029EA3529A84D57D5CBEAA9418DB2C34B2506";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "2490961B43477EADAADAADAAB50AFC496C822222222203E4F67E21192590D90D";
    attribute INIT_31 of inst : label is "6FF66B64AE737B6FA7DBAB717E65F8EBA58EDA4EC53C7A76696A933A5544F360";
    attribute INIT_32 of inst : label is "F7CA2A8AAAC7923E191AFA8B24AB2D8814DF8FF110040004E22CFD25FE10C6FF";
    attribute INIT_33 of inst : label is "CEB5F51AD925964AAEDBEAA8FD68A271B7DA137EEDD9D40A40300000000008FF";
    attribute INIT_34 of inst : label is "4D509AC24824FC8053484F6BEA3592592F3ECD06774E96595C15EFFB892C966E";
    attribute INIT_35 of inst : label is "00463218020004C0856D58578155F80A24080000473208020000C01F13FE27F8";
    attribute INIT_36 of inst : label is "04C085EF5A778175E80A24080000663208020000C0056F58738175E81A240900";
    attribute INIT_37 of inst : label is "FFE43EF9F517D5FF00FFE32FE0CBE3E5ED5A538155F81A240900006732180200";
    attribute INIT_38 of inst : label is "FA65EBCF6BEFB9054CA4ACDD5699F5B9B63B0C865AF73589996BDEAAADC27DD4";
    attribute INIT_39 of inst : label is "65D6F3F5192EFF5ED8B2B1BAFA56CBBB760CD60DFD5FCC9CB106E77911EEE2AD";
    attribute INIT_3A of inst : label is "0004C0971326CD34882DB6910FF36CBBC8EE776E9C5A86CBB3B066B21FCB60CD";
    attribute INIT_3B of inst : label is "4F2AAC4A15712854360AFC2A1564BFD95B8DC6088175F81A2409000047321802";
    attribute INIT_3C of inst : label is "16B2524F763E276091110A9527F259258396E06A0B004008D896C4A0220924DA";
    attribute INIT_3D of inst : label is "FFFFFA31FDE1E5E2B6A41CA80A698D125480A56BB4E6FBD7F875BFB033654891";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "2AAB6EBF3C027055145585C631B9C8C8AAC6E2AB1AB18DCEC644556371558D51";
    attribute INIT_01 of inst : label is "666B6EE3E055781A59E01E04AB9F95DD9E04F9A04A9A179734318EC112471645";
    attribute INIT_02 of inst : label is "93299989F05B6C1493323B18CBE0E44CED9A7C4934089B88A64C9340B7C684A5";
    attribute INIT_03 of inst : label is "A3446D563CC6B360AA386C698E8D11B558F31ACD82A8E1B07F5C25D341ADC23E";
    attribute INIT_04 of inst : label is "BBE9AD7FC5A63226649563884BA40B5B86C69DC89992558E212E902D6E1B1A77";
    attribute INIT_05 of inst : label is "EF197B59B6DB5BD0E1B0AD0AFCB5F13958D85A185A181A581A5A1A015D1F68D2";
    attribute INIT_06 of inst : label is "C6BB013D188968F57557D5578142314308E32E547E4969D151FB3DD369A4CD35";
    attribute INIT_07 of inst : label is "4B32060042D842EC3A400E208C1C40E8F4EBDC0C44898F060E0C1870FC64E244";
    attribute INIT_08 of inst : label is "36533D84C74CF4EE4E6BA76CB1B2CECBBBAE6EBA78432183E4C6592AC94FE016";
    attribute INIT_09 of inst : label is "3C6670C999C326478661DBA03092438500073F07FFFFFFFFFF8067F867FDDE26";
    attribute INIT_0A of inst : label is "061820E070C8381C320F078C190783C60C87038332E9CC61FE7E9633446D1E32";
    attribute INIT_0B of inst : label is "45CCF83E186C2C8BDD74D6B44008383249129228401070644061EA64DC8CCC9E";
    attribute INIT_0C of inst : label is "3DB171C642CD47A64ED25324262F467726E73925FA4BF6399B5D359A2C0B0C16";
    attribute INIT_0D of inst : label is "99A6CF7491BD3B02DF35F2E723334C6744B2723335939199AE7B1650EC895304";
    attribute INIT_0E of inst : label is "3335C8CCD73D19CC671CCCD367BA48DE9D816F91F0E633A24C6744B9ECCACE39";
    attribute INIT_0F of inst : label is "32C8DC9D81EFD1F8F633A258CE8963919CC479EEC9A4732C8DC9D816FD1F8F72";
    attribute INIT_10 of inst : label is "0BCC4D0360CFC2064C4E304B138C1AE6F306B9BCC1AE50C3777747479EEC9A47";
    attribute INIT_11 of inst : label is "D8EF2DEC7105798E7224F644DF667119B217AB6AB2D6ED80322A9BBD05A46F2E";
    attribute INIT_12 of inst : label is "EA4159738ABAE8E1CC44FE380DE480A08A3F946085737A8CDA862E8D3B62DE19";
    attribute INIT_13 of inst : label is "00148509020210B12126C92EB1B3F1DBD61371028CB6498249636B8AB41584AC";
    attribute INIT_14 of inst : label is "FD9424CD2686499A4D865448A98F82F94515E19AEF271563DA9251E72D55C255";
    attribute INIT_15 of inst : label is "B4EEC63FA60D7F1BC56CD9992531583E369240D1D06C26708A80054454408AFF";
    attribute INIT_16 of inst : label is "4E241D2C93C8BB26EA4EA41D2CDBEC1B5B75B0ED66DF6E6DC6C38C96D47A69CF";
    attribute INIT_17 of inst : label is "3193233466C2F151B159928BE2631337DA646DF699253379A3B5724F36461CEA";
    attribute INIT_18 of inst : label is "017C07AF38B85180E66B7C3C20DC1346E4D1B4DA2F0997C592470AF77F059333";
    attribute INIT_19 of inst : label is "B9E4C82D0E75AF73A40CC9660C8A8AC94002800016E6D4DB023E052904442893";
    attribute INIT_1A of inst : label is "9F60603F30F3F291E4F21C2F0CFFAAA2082052295D513E4F8E286F16DA8E295D";
    attribute INIT_1B of inst : label is "F663042F5A67DDDBCEE9F7721D3BBB2E99DD174EEE18A3385A4E345339042CCD";
    attribute INIT_1C of inst : label is "2088000829290920000000000000093FFFFFFFFFDF40840ED2AAAADF5F33FBFE";
    attribute INIT_1D of inst : label is "FEFFFF2035F4C6085A6666EEE6BAF4E8F7FECDFBEA8B74E82828282808080801";
    attribute INIT_1E of inst : label is "FDEFFEF4E7B771DFFFFFFBBADFDBFB9F16FFF45DB7FFFB6EFFDBFF9B8659DECB";
    attribute INIT_1F of inst : label is "05535C08591CBD1C597C1E80991346D56F1DB462947266ECFF7F3FDFDFF7F3FD";
    attribute INIT_20 of inst : label is "BA6D00300005FBEBFFEBEBEBEAFFFFEFAFFC60187180364283801C02AE83A0F7";
    attribute INIT_21 of inst : label is "800809B03A6841819068000000084D8192600C30000561919865102844156995";
    attribute INIT_22 of inst : label is "00680C003B6861B11808001820086C3C38680939326861959808082822086181";
    attribute INIT_23 of inst : label is "42852814A14560318005080023556031802D09803B6841039808000023084D31";
    attribute INIT_24 of inst : label is "BAB15CE62E10B17166E262E836619FE7917222CDC48500000000200000005029";
    attribute INIT_25 of inst : label is "E01AE72E4820E7240BF2425D21DDAB9357162F4230A91AB8649AA61E80D57398";
    attribute INIT_26 of inst : label is "140E008D1E045D0F5C4711C0701C0721C8701C0701D0741C0501C0718F01D805";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF551D8E07A2B995CE1FC70F75D60503AC0A0758";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "36D81A4F431537669B51B51BA32E93C92CAAA8A8A8A88B8C9B7323196595C01C";
    attribute INIT_31 of inst : label is "B6927924B32DEB4D964AA3407145CCDB916DBE7B1431A3992C467609D544A0E2";
    attribute INIT_32 of inst : label is "8020A2282A86571F100263992CB3645C54927973755DE67D14551E6692F98263";
    attribute INIT_33 of inst : label is "E884C73E496C924A224D2CB4E46707DDC6583E3060E317F6FB7FB33B333B3BF7";
    attribute INIT_34 of inst : label is "CCAD98AFDBC8C2EFE4BEE9098E7C96492879987F7A04B259693644609BE4B246";
    attribute INIT_35 of inst : label is "F2C74D767E2BDD732B3973E93C65E5E51A1266F2C64D767E2BDD7335B32B6656";
    attribute INIT_36 of inst : label is "D973AB3973ED3C65F5F51A1366F2C74D667E2BD973AB3973ED3C65F5E51A1266";
    attribute INIT_37 of inst : label is "EFA549259F97D9DCDDEFA026588B29CB3B73C93C45F5F51A1366F2C74D667E2B";
    attribute INIT_38 of inst : label is "9C45CC87A4DA2D19C70CE8E15C2F4643BD7C9B4C464466D3B11912DDF0AAE2E5";
    attribute INIT_39 of inst : label is "667B533ED05F239CDDE2F0CF6C1397CB9A24E66E1367165DE91BAF8D18EB41CE";
    attribute INIT_3A of inst : label is "2BDD7328B4CD19C732D26CF75330797C689825898EF11B97C4D1273273E1A24E";
    attribute INIT_3B of inst : label is "FD3BB66E1D99B877361749DB55C3D266749B09B03C4DF5E51A1266F2E74D767E";
    attribute INIT_3C of inst : label is "DAA2626DBC5B35E1CBCE1FFFA7737D37C23088A62BFCFDDE6CEB77787739E76F";
    attribute INIT_3D of inst : label is "FFFFF9EFDE84C589E9A63669537DCF0F70553664DAB39B1A4D936CD1319B4499";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "22A22D0654BD9450004410CA14A22665A25296894A50A7113312D129CB44A731";
    attribute INIT_01 of inst : label is "774A4AD0C9146A1648910926234A11DC8924D8924D8902111252C4EB9211C7E4";
    attribute INIT_02 of inst : label is "CB399DBBDACBAEBEB9B3B38AE8B5E65EE9DB4E9DB61A8EDD2BEB91349AA26086";
    attribute INIT_03 of inst : label is "266CECDB1DFE3360000E7DED8C99B3B36C77F8CD802A39F7402C968BE1B5D766";
    attribute INIT_04 of inst : label is "55E2D967F3B77A76CC8DB19BC3240008E7DED8E9DB3236C66F0C9002839F7B63";
    attribute INIT_05 of inst : label is "23ABBB69B6DB739475740D40FCD1257CE89E56085602025C025C01441288735B";
    attribute INIT_06 of inst : label is "AE13851D928AB8AA0A222800B4D27DC13CBF36941EC9E996507936FACF2CA002";
    attribute INIT_07 of inst : label is "423279FC40644072B4452A2A165454617646892845DD5D438F1A3C2A4D20A2EE";
    attribute INIT_08 of inst : label is "D2DFEEF7FA7F27D27D3688F7969C5271C947251E5AB9D8B96556990CC8581FE6";
    attribute INIT_09 of inst : label is "AF3B567DA559F6B56F78F65D2F1C8B63E72B95E7FFFFFFFFFFFF980798035FBF";
    attribute INIT_0A of inst : label is "4ABF166D34759B4D1D66D347DAB369A3ED73E9E6BE7D152E86FE9AD34EC6579C";
    attribute INIT_0B of inst : label is "54CF4FD3FF1C02E99D35BF6A421535B64D71932E642A6B6E60B8CBEEE89D9B3F";
    attribute INIT_0C of inst : label is "59B1BCCE51E8EBA2EFD2633466E7666B02F63C4A9ED53F9D970FAA9FAFEBFF83";
    attribute INIT_0D of inst : label is "D975C764B79FB576C97697722766C46FCD56337F7AB19BFBD573B3BC68855B14";
    attribute INIT_0E of inst : label is "7F7A89D9AAB94E6DE70CECBAE3B2DBCFDABB64AE977237E6C64EEF55CE77CE19";
    attribute INIT_0F of inst : label is "3ADBCDDABB64AE97732777A8DF9ABBD4E6DC70CECFBC33A5BCDDABB64AE97733";
    attribute INIT_10 of inst : label is "23A6C0AAD2EFE20375EB354D7ACD5B7CA356DF28D5B7A171C6C7E2C70CECFBC3";
    attribute INIT_11 of inst : label is "B0EEA9DC715516D4A63712C6A32EBD939C1AFF3FD262E5C89555419254280A14";
    attribute INIT_12 of inst : label is "45AFB509414140550044CC5B0CE48080883E98604451588052002B0CB67C9D51";
    attribute INIT_13 of inst : label is "8CE718EE399C75997B72CB6DD5833EF9DF07A40AAD9AA2C25BEBBB03B01D8083";
    attribute INIT_14 of inst : label is "654074ED24C6E9DA49269544A8BE93FFDFD4D11A47C43041D81268EF5DB99311";
    attribute INIT_15 of inst : label is "F467D33D8064DF4951E4C89127319C3B64936199D04832B9CC0005445441CC76";
    attribute INIT_16 of inst : label is "623D1A1FD8FB19EDFF633D1A9F90DFFEF21578D4FC86DFC865E3654F8C260847";
    attribute INIT_17 of inst : label is "7C93AB3676EC797CBC0BFBA93173B3A1B6E5CC6DB96F3B1F63620F63EE943CCF";
    attribute INIT_18 of inst : label is "85BDF8A987FCCDB1D41655EBB39B5182D460BE5EA5DEB545D6756BF755309971";
    attribute INIT_19 of inst : label is "D096D7B9EF3AA22193594EB2A82A834D00000000245AAB569BBF490F8146F339";
    attribute INIT_1A of inst : label is "13631E137C3B1BD0761B0A676DFFAAAA8AA89A0245141707E7A40FC592550501";
    attribute INIT_1B of inst : label is "BC43D8B69E779D93CEC9F7676EF3B25779D92BBEEC5161DECCC7D4B1DE143DC7";
    attribute INIT_1C of inst : label is "0908000809090900000000000000091FFA9FFFF89A810D5497FFFFDFE92A4A5C";
    attribute INIT_1D of inst : label is "BDEBB3281888C7B16E2222AAA330E72A73D6BB581AB7F5818181818181818189";
    attribute INIT_1E of inst : label is "2E632D2E5DE72FFEAAAAABE9CFC9F9AFC669F4BADF496EBB95B76789EABD5695";
    attribute INIT_1F of inst : label is "36510CA9705AC809693CD018991146902B00A4005012426F494BD252E494B925";
    attribute INIT_20 of inst : label is "000000000002501115104510440000045057381871811A50F18E0C082A0306A0";
    attribute INIT_21 of inst : label is "00000582B9602C000B0000B000002C000B0200B0000000000000000000000000";
    attribute INIT_22 of inst : label is "01600000B80000000000292132600C3C386029213260000000000580B9600180";
    attribute INIT_23 of inst : label is "000000000000000000000580B800000000020580B8002CB201600000B8002CB0";
    attribute INIT_24 of inst : label is "231042120E1010700B9C20E807FE6000700E0017384000000000000000020000";
    attribute INIT_25 of inst : label is "E010630028200F140580084A00848950120824459F02083852483FE1FE410848";
    attribute INIT_26 of inst : label is "1C2402804A000B2D000000000000000000000000000000000000000048040402";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF004984125090848649C32434880709100E1220";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "5B68097740B1A66483C03C03806EB2C924802222222200B493BD810B24905415";
    attribute INIT_31 of inst : label is "2796D924F32EE49EABCB62397D89F6FFB16DF65D0517A91F35006A11AA801680";
    attribute INIT_32 of inst : label is "A08082A20222AB9A49C3A80324E66A6956DAB9B900045004101445A493D284E1";
    attribute INIT_33 of inst : label is "E8875006C924924E234939E0AE7B00E8A2AB0654A853196C92488888888080AF";
    attribute INIT_34 of inst : label is "17502F76DB69FB496C97490EA00D92493CBE885F1A009249E90C4460836C9242";
    attribute INIT_35 of inst : label is "FB626F7F6E3F9DFB3BB12DE96BE0EB6FF71267F3624B7E6C3F9DF32085D40B82";
    attribute INIT_36 of inst : label is "99FB3BB12DE96BE0EB6FF71267F3624B6E6C3F99F33BB12CE96BE0EB6FFF1A77";
    attribute INIT_37 of inst : label is "495BEDB4B4D4999CB5494B3AF8ADCABBB12CCD6BC0EB6FFF1A77FB626F6F6E3F";
    attribute INIT_38 of inst : label is "D904D8ADE7D63C1A76D8623876FF53715B2776F44ECDB6F199BFBCFF7F7F3E7B";
    attribute INIT_39 of inst : label is "24363F2C8EC9E31DEAD3B686EF95727378175205D9E2FFCADB5564FC0D4ECFCE";
    attribute INIT_3A of inst : label is "3F99F3B70E9D31E3B39E78677B9C7727E09B575CF56F157279C0BA9051CF8175";
    attribute INIT_3B of inst : label is "9A13B22709889C27B6376BD3CF6FDA7474920DB06BC0EB7FF71367F3624B6E6C";
    attribute INIT_3C of inst : label is "4963737DAF471134589D84C9D9192E92FA0C04CC317226456469636B11926B2C";
    attribute INIT_3D of inst : label is "FFFFFEB5DEF5D6F8ED757E2519681D0637D1A6E6D9F79D7B6FD64FC090FA7F91";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "4F40880430A48C1A4416580404022220281000A0402020111130140800502005";
    attribute INIT_01 of inst : label is "48A8A88887456E58900D00C0A002AD6280C9380C9380C2A701A1488621545085";
    attribute INIT_02 of inst : label is "10A2502DE08648612002542088C11411080050800005C101C0802019242031E9";
    attribute INIT_03 of inst : label is "DC20A085300841014246B3162B70828214C0210405231ACC00487C5200C90C08";
    attribute INIT_04 of inst : label is "512684001058ADC208485344A40214846B3162B70821214D1290085091ACC58A";
    attribute INIT_05 of inst : label is "9186A480CB2C852C155C39C3B29D12CC0890560A5C08025E085C005750001344";
    attribute INIT_06 of inst : label is "98FC00D22345A688082822A86131214CA698AA204354366C910D126492591242";
    attribute INIT_07 of inst : label is "A425000372637250252411114022228408895410A23133CF9F7A75F9D0551118";
    attribute INIT_08 of inst : label is "B1B0DC6C36C36C36C3658C330D8C363058C163046050C86905C4A28095300020";
    attribute INIT_09 of inst : label is "441A80356A00D588155C242A2A1B89C25217B857FFFFFFFFFFFFFFFFFFFAC661";
    attribute INIT_0A of inst : label is "01D68ECB6633B2D98CECB663D6765B31EB765B3BAE11031A0ABA618DB346220D";
    attribute INIT_0B of inst : label is "670A4390A70124CE110050040A56E625060A41A114ADCC4943AC80993542449C";
    attribute INIT_0C of inst : label is "16CD01428ACC12DA8008E4BC7E6C570006C46048959929C11006D80111C45310";
    attribute INIT_0D of inst : label is "56D0104703E080F8C8508454400008A1008455091422200021C141C406854B34";
    attribute INIT_0E of inst : label is "0917100010E0072B2C20AB68082301F0407C6428845540112AA12287043C5841";
    attribute INIT_0F of inst : label is "A381F2407C6428845440007500450E007AB0C20AB6828A301F2407C642884555";
    attribute INIT_10 of inst : label is "60E9DE280FB8218813098C1042630C3098C30C2630C34758E7E7000C20AB6828";
    attribute INIT_11 of inst : label is "2204E09114EE850840B970972E080813E4C2AA2A9902C5A008800335D17C8214";
    attribute INIT_12 of inst : label is "8EBEBBBEDEBBEEEAE2006751A8C016165102020DEEAD2D534B683441243609C1";
    attribute INIT_13 of inst : label is "4852358D210AC3669E8936990F4E8865659210018D41E892DE4C0800801400F2";
    attribute INIT_14 of inst : label is "E5801B041015B6082035C81D03100307FE20502000CC0000C004D82AED814050";
    attribute INIT_15 of inst : label is "4C612096014E00DC350001A6084520000000006D0004820DE40005445445E416";
    attribute INIT_16 of inst : label is "8C5A930263345581018D5A93826330808C62C49C13199031BB126181E30527C0";
    attribute INIT_17 of inst : label is "254422B1090E61449135238B41080CD6699B319A6658CC669A5FE98CC9786289";
    attribute INIT_18 of inst : label is "3CFB062CA620C92C9C015534944869B2DA6CB44E2C4225A52D988B045604C0C4";
    attribute INIT_19 of inst : label is "48B89C9636A2255201200281823220062A8800554104CB8079810102A1818D38";
    attribute INIT_1A of inst : label is "1B6A030554381922731D03F6C9FF000AA2AA5B4C4451C17011C60CB7DB986DD9";
    attribute INIT_1B of inst : label is "6CC370A3199C558E28C70561C2CA39C36558E0B08EE3631BDBCFD5B31A152FD7";
    attribute INIT_1C of inst : label is "6000000928006060000000000000007FFA9FFFF838220998D555557DC12EDA4E";
    attribute INIT_1D of inst : label is "00DB7343D009C6E1406666666630E42930BE0AF016032C882808280808280800";
    attribute INIT_1E of inst : label is "24E7250A13830ACEAAAAABA8D85B0BC026196C1996D96208B1D2E719471CCD83";
    attribute INIT_1F of inst : label is "B8338298F1E31BD98102E05D32A46A59A5A696834680E64CDB4936D24DB4936D";
    attribute INIT_20 of inst : label is "ABAA7FC7FFF84110514104145100001440456178E38980F8FBAF5D68E535D700";
    attribute INIT_21 of inst : label is "0007000400070006200700062007000623080006238A2E16ABAA3E1EEFBA2E16";
    attribute INIT_22 of inst : label is "00070010000700182007049C89070C3C3867049C890700182007001000070182";
    attribute INIT_23 of inst : label is "FDFA2FD6BD7A03C63C2A0186183A000600280006000700062007000600070002";
    attribute INIT_24 of inst : label is "642AC0055E492AF0100055E4880000000480802000AA0FFFFFFF2FD6BD783FDE";
    attribute INIT_25 of inst : label is "EE218C21A54A0852A073672BB4A8084890112090300495648015600000AB0015";
    attribute INIT_26 of inst : label is "808002420080003003C0F03C0F03C0E0380E0380E0300C0302000002A1842A90";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF047021C08E001018000C00C011282062404044";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "3FF91BFB604849DB0EE0EE0E41D988900077757575757628240C3202400B1BE1";
    attribute INIT_31 of inst : label is "D96492000A52148270B05A454E013093658B2414EE8420C6418224089FC8BE04";
    attribute INIT_32 of inst : label is "AA0A002A0A60B2240568999A410E4F1093014202AAAAFABAABAAA14125290288";
    attribute INIT_33 of inst : label is "82D1333482012000B4B24289890A86A0708635061C38D4080D90CC4C4C4C4C0F";
    attribute INIT_34 of inst : label is "01AA02510412B012000482A26669208000715120050704801411634D1A4904A4";
    attribute INIT_35 of inst : label is "C2850198707415C2284D1B1271101F04A50047C2850198707415C23F407F80D7";
    attribute INIT_36 of inst : label is "11CA284D1A1271101F04AD0857CA852589727411CA284D1B1271101F04A50047";
    attribute INIT_37 of inst : label is "B2F532C864440529B8B2E00982AAD6284D1A3271301F04AD0857CA8525897274";
    attribute INIT_38 of inst : label is "631C7280C040B00291846019DAD841BFD321A43880005162A200003F57771E14";
    attribute INIT_39 of inst : label is "2124CA69D4884A56BA9ED424B7246214600412618D31ED12956464301C48842B";
    attribute INIT_3A of inst : label is "7411C23D43700308226C051444D8E62180330476DD4C646219002092658E0041";
    attribute INIT_3B of inst : label is "BB3BB66E9D99BA763610B0119DA66D9B4081400071381F04A50047C285018870";
    attribute INIT_3C of inst : label is "488FEFE6E2181D00D9986CD995532CB2C9244AB0A0146CCD2671338E33304125";
    attribute INIT_3D of inst : label is "FFFFF8006A4B1166C104CDAA04406E00A5204149270060CDB6002500106210F5";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "44E14CC5B3A5A50A5512FAB5AD00000000B40002D02D68000000005A0001680D";
    attribute INIT_01 of inst : label is "1D5554C4B46B42A1C009008354C020768089100891008022012DFC9225DCF190";
    attribute INIT_02 of inst : label is "34A6535AEC0A69238044AA4191D814839534B9E24928AD622D96701104602008";
    attribute INIT_03 of inst : label is "DD993205B7634593485693372B7664C816DD8D164D295A4C885B4865126D240B";
    attribute INIT_04 of inst : label is "5716820810DCADD991205B76344934A5693372B76644816DD8D124D0B5A4CDCA";
    attribute INIT_05 of inst : label is "14D72482D964C5349994394392B70AC41AD24E164E161E461E4E1EA4A0C01749";
    attribute INIT_06 of inst : label is "A8B44AD75A322682882A880163497B4056D9E9285150176CB145002618619048";
    attribute INIT_07 of inst : label is "10C080028E028E212416ACC8015995901D9532AD193553970E58B060D2DACC9A";
    attribute INIT_08 of inst : label is "85A0C32830830830830D00996D0DB436D0DB436CC456E5630855804102900040";
    attribute INIT_09 of inst : label is "B6D965B52D96D496554B621A2259B88C5CC5024FFFFFFFFFFFFFFFFFFFFC9441";
    attribute INIT_0A of inst : label is "AD92020B05B082C16C20B05B5210582DA930582AA5B20B580AB975ACB1565B6C";
    attribute INIT_0B of inst : label is "FC345314A6868BB8361B0000029C242537284DA50538484942AA949B323932BD";
    attribute INIT_0C of inst : label is "926D452942CC325A436DC0A43AA89E8CA488832AB255698361B6DA6C110453C7";
    attribute INIT_0D of inst : label is "26CB20D815A216D4EA52A5CD9EDDAB1CBB6548E4CB2ACF6EDB4985E436916344";
    attribute INIT_0E of inst : label is "EDD923932DA4570930419365906C8AD10B6A7522A5CD9EDD8B3DBB6D26BC6083";
    attribute INIT_0F of inst : label is "6C0AD10B6A7522A5CC8E4C923932DA4570910419365906C0AD10B6A7522A5CD9";
    attribute INIT_10 of inst : label is "80C86660A80001109331AC9A4C6B2EB31ACBACC6B2EB55542E6B101041936590";
    attribute INIT_11 of inst : label is "200C81901005652948A1349426C95915A024ABAAB410E1A0222A8DD51B4D02C4";
    attribute INIT_12 of inst : label is "95511584055411450D95EEF328C92405104220C9CCDBE992FA486E11E4223903";
    attribute INIT_13 of inst : label is "63084630C633980000049249240ACF2D715709F3B224CDA3CC484C22C0561086";
    attribute INIT_14 of inst : label is "B8AA9BB24924B76492548C0780C42B000020CE001880C008E02DCC2A558121AA";
    attribute INIT_15 of inst : label is "5D697586D45A20D4B2214218446506518924926D6C93CD4FFF8005445447FFC9";
    attribute INIT_16 of inst : label is "B19952026C33995889B19952826C336C4D8CCA9413618936332A59018365B628";
    attribute INIT_17 of inst : label is "652E64794892E685244326104A8A46482449361913846D864A2839B0C4A61191";
    attribute INIT_18 of inst : label is "425BFB36F54D39289180EEC2C61400A2A028A49040537D9A2456768CBAF1A648";
    attribute INIT_19 of inst : label is "04009B14C6AE14CAC0C2920DB013001A08A00044122CF80540006D8230C04A50";
    attribute INIT_1A of inst : label is "279D11815BB1914D6090210649FF0000000072C3E6A9CB703B421D9EF822B875";
    attribute INIT_1B of inst : label is "409A538050C836241B120C88D606CCD903266C819136127A122AFB0A7E1E6C48";
    attribute INIT_1C of inst : label is "0001000040600020000000000000003FFF5FFFFDDFC40E1F02AAAAA0B6469692";
    attribute INIT_1D of inst : label is "40925AE0240974A70266664444AE800AA5235685142A09402000002000200000";
    attribute INIT_1E of inst : label is "48B54A4C9292488800000402985B0BA074D04951049041802530B412D4D2892A";
    attribute INIT_1F of inst : label is "2A37909DC42943D4A540A49933254FD37D25F486F48484A892D224B4892D224B";
    attribute INIT_20 of inst : label is "661D00000007FEBEEBFEAFEAFEAAAAEFAAF9FA586185608E77EEFC517E660524";
    attribute INIT_21 of inst : label is "78E802024088100004081C4007081070040700400005180C661D180C661D180C";
    attribute INIT_22 of inst : label is "7888001040080018000816DECD8813C3C78816DECD8800180008021040880200";
    attribute INIT_23 of inst : label is "60C5180C60C50000001D0200401D0380781F02004008104000881C7040E81040";
    attribute INIT_24 of inst : label is "77AAC0055E492AF7910855E6EFFFFFFBE4BE8F2210AB00000000180C60C7180C";
    attribute INIT_25 of inst : label is "0E00002A010AA000AA0000540140028015002A0014D69576A495600000ABFFD5";
    attribute INIT_26 of inst : label is "808A00001400140017C5F17C5F17C5E1785E1785E1705C170501405000054015";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF50000BC50028014014000A0140202280404500";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "B6DA7F41046C4CD98E70E70EE19B0C4924D757575757572926DA2649249A9EE9";
    attribute INIT_31 of inst : label is "4B3249248AF139176DBA1AC95A11684B6D84924AAAE4C4D669C204881553F000";
    attribute INIT_32 of inst : label is "8028800A0265DA14B10C9889248ACD92C2258627AAAEEABEBBAAA94926A52258";
    attribute INIT_33 of inst : label is "9699311249249248A4B2628AD94882572CB613265C9854090D80CCC4CCCCC44F";
    attribute INIT_34 of inst : label is "6BFED65100929092082097326224924923333700870492491C11615989249266";
    attribute INIT_35 of inst : label is "84B59394A1F236C648ED5A33B3311B8E6304C884B59394A1F236C65FDAEAB5D7";
    attribute INIT_36 of inst : label is "32C648ED5A33B3311B8E6304C884B59384A1F232C648ED5B33B3311B8E6304C8";
    attribute INIT_37 of inst : label is "34D736DB24646D6B9034ECC982A85668ED5B33B3311B8E6304C884B59384A1F2";
    attribute INIT_38 of inst : label is "371436A45925B0254584E25D59D189BFF2A964491C9949CE6472673F57F7CCB6";
    attribute INIT_39 of inst : label is "2B6DCADBF48A5AD2BB96CC6D930C629CE055B2FB8515E90B95C455303ED9B469";
    attribute INIT_3A of inst : label is "F232CE57D376C4106C6DB20D8E58E6298177ACC2CDCC44629902AD96EEBA055B";
    attribute INIT_3B of inst : label is "B3B3366299598A647611982B159425DB5BA4F349B3311B8E6B0CD88CB5B785A3";
    attribute INIT_3C of inst : label is "58AE6E627219B7189939489135D329B2996E5AAEA2746CCE6DE36F3A335BEF6D";
    attribute INIT_3D of inst : label is "FFFFF9086B6B1026C2D545AB02662E4025301B4B661A76C49C2C930295655091";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "24234407648CD0150545D86A58800005816216058852C4000002C0B10B02C430";
    attribute INIT_01 of inst : label is "33EBEC48ECC57A3F1D89D8AEAB88108C58A4958A49588812B15B4B4993579740";
    attribute INIT_02 of inst : label is "82198828DAC9D49E3B727918CDB5E25E408204D9241686D8834DCB14B7D62204";
    attribute INIT_03 of inst : label is "264CC8CA5CC67240AAB96CC884993323297319C902AAE5B2E82ECE99C19A9324";
    attribute INIT_04 of inst : label is "11C0094843221264CE8CA5CC67340A0396CC8849933A3297319CD02A0E5B3221";
    attribute INIT_05 of inst : label is "0F68124924DB308368826C26CD51253A7088580058080850085001FD50084208";
    attribute INIT_06 of inst : label is "0607070832CC18220A800AAB93C10001082616B8DE0BE892E37865D041042AA0";
    attribute INIT_07 of inst : label is "46B2000642464243B0E59B322736606263468999669A0E04004489120DA5B34D";
    attribute INIT_08 of inst : label is "3A33188CC6CC6CC6CC75A244119046411904641238572A8CE7463918C948000E";
    attribute INIT_09 of inst : label is "6820D8418361062D84609E6FA71E8D9504371B07FFF80000000000000004F766";
    attribute INIT_0A of inst : label is "625844603041180C10460304182301820C030182304914A5D82E8A534C063410";
    attribute INIT_0B of inst : label is "CDC95856081D7DDBD92439CE1865B1B0C8073201F0CB63660820EA748DDECD0A";
    attribute INIT_0C of inst : label is "4D903884E5A7C9A04C9342142326667542F73800B00162399F0920909C27043C";
    attribute INIT_0D of inst : label is "99248E6591B811020B18B06377B316EF6618B77B30C5BBD984721A3248004100";
    attribute INIT_0E of inst : label is "7B3099C88239A86CC71CCC924732C8DC08810590B06377B336EF6611C9478E39";
    attribute INIT_0F of inst : label is "3248DC08810590B0626722099C88239A86CE71CCC92473248DC08810590B0637";
    attribute INIT_10 of inst : label is "00536D0038CC02634ECE3065B38C114CE3045338C114A040020342E71CCC9247";
    attribute INIT_11 of inst : label is "C59732E2DB057294A716AB62D434A481B81D5755D2F2E5F615554BBF31EC0182";
    attribute INIT_12 of inst : label is "41115150044440440C48545986A4D898EDBC9236E23924624D31244238B98E65";
    attribute INIT_13 of inst : label is "42108000000215BB7376DB6C51B9A0988300276EE13A4A9463A3798191ACC107";
    attribute INIT_14 of inst : label is "C0006449A4964893490635448888830000B0B448388602F448D2488301F09755";
    attribute INIT_15 of inst : label is "7049C72D872DA19AEDD688712310B82264924190906820A0000005445440001C";
    attribute INIT_16 of inst : label is "4624187D91C99927DE4624187D91C913F23120C7EC8E7CC8C483067E8E470D08";
    attribute INIT_17 of inst : label is "98D9A3B677EAB979B3D8DA897273B12392E4C8E4B8AF123921EA9E473E3C9CEE";
    attribute INIT_18 of inst : label is "01260E0CA4F04D9A54276C3D804E9386E4E1BADA258CC065DBCDBEF77D8F9133";
    attribute INIT_19 of inst : label is "B04EC8340C224A21BED94803680E82430A0000512CB548C1C660C30860443821";
    attribute INIT_1A of inst : label is "9A68911418A28341448285352CFF00000000C663555E2E881E630F7248E7E85E";
    attribute INIT_1B of inst : label is "24C3C8849E219910CCA866466D73AA46B9D5235CEA92291E5E4E5D1318163CCD";
    attribute INIT_1C of inst : label is "2020200000000000000000000000003FFABFFFFA1A28101FCAAAAA80B61EDADB";
    attribute INIT_1D of inst : label is "42DB7BA0748987910C2222222330C920B1B846E9160B6C604060404060406060";
    attribute INIT_1E of inst : label is "6EE76E64CB5B60ED55555556D85B0B9036596C5D96D9665DBD96F659421C458B";
    attribute INIT_1F of inst : label is "8C81526A48B19826C1423ACC88DB224924C49B124313164EDB5BB6D6EDB5BB6D";
    attribute INIT_20 of inst : label is "FFFF7FFFFFFF55405400055500000050005721830C273359123253B8A53051D4";
    attribute INIT_21 of inst : label is "FFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFF";
    attribute INIT_22 of inst : label is "FFFF7FFFFFFF7FFFFFFF7FFFFFFF73C3C79F7FFFFFFF7FFFFFFF7FFFFFFF7E7F";
    attribute INIT_23 of inst : label is "FFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFFFFFF7FFF";
    attribute INIT_24 of inst : label is "67AAFFF55F6DAAF7910855E6EFFFFFFBE4BE8F2210AA7FFFFFFF7FFFFFFF7FFF";
    attribute INIT_25 of inst : label is "F1FFFFA1FEF01FFF01FFFF43F03FE07FC0FF81FFB4D69566A495600000AB0015";
    attribute INIT_26 of inst : label is "7F01FFFF03FF03FF001004010040101405014050140D0340D0F43D0FFFF43FC0";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFF0FFFA000FE07F03F03FF81F03FDFC07FBF80FF";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "6490D304109322341B09B09B136C464924A8888888888B94903191092494C10C";
    attribute INIT_31 of inst : label is "26824924F184E24CC36730667301C64FD8249249147323199626CA1B3546B08A";
    attribute INIT_32 of inst : label is "A8208800088643921CA2719924E024E9449319104551554145550CA490D28663";
    attribute INIT_33 of inst : label is "4844E3324924924E1269186024632648830D3258B143096DB24A2222222222E7";
    attribute INIT_34 of inst : label is "F411E925B258C65B25934889C664924938B8884E184C9249E13C0C241924924C";
    attribute INIT_35 of inst : label is "3B426C6F4E1BD93B3710A5C898C720E31F1A763B426C6F4E1BD93B28BD117A20";
    attribute INIT_36 of inst : label is "DD3B3710A4C898C720E31F1A763B426C7F4E1BDD3B3710A5C898C720E31F1A76";
    attribute INIT_37 of inst : label is "E59CC920909092840EE587274C03299710A4C898C720E31F1A763B426C7F4E1B";
    attribute INIT_38 of inst : label is "8904981B249A0C10264CA020842646411C2C9BE4CE44A4311339108282806348";
    attribute INIT_39 of inst : label is "245263141B6B210808E0238A48D39AC11804422430C612C8E11B858C134E4B84";
    attribute INIT_3A of inst : label is "1BDD3B20BC9939C7339248E6790639AC6088C70834731B9AC2C0221210418044";
    attribute INIT_3B of inst : label is "BC33362609989827362E4180C8499224249A082098C720E31F1A763B426C7F4E";
    attribute INIT_3C of inst : label is "6947677919165124688ECCD9DD5B2EB2C100476E21FE2EC66C5B62F91118616D";
    attribute INIT_3D of inst : label is "FFFFFD8C849401981868320512200DAD5AD1043698738132439348C011902ED7";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "A4E12239480822BAFAAE81A86B80000781AE1E06B8435C000003C0D70F035C20";
    attribute INIT_01 of inst : label is "154142232CC4343D6E83E83E00A850546836968369682852D04A850FDA208900";
    attribute INIT_02 of inst : label is "101081288ACFB0FABFA23A288D15A35A801000D0001F9C5065055D06D65A0A14";
    attribute INIT_03 of inst : label is "000881C96442A0015FD5A2A50000220725910A800555568AC832834D80B61FA2";
    attribute INIT_04 of inst : label is "1202004822940000881C96442A0015FD5A2A50000220725910A800555568A940";
    attribute INIT_05 of inst : label is "557500409249601FA88E3CE3C474068BE0C4580850000858005001FD01008108";
    attribute INIT_06 of inst : label is "1C8A068518441477F5555FFF51C03100804512D06A2FA54B41A821420820D555";
    attribute INIT_07 of inst : label is "0FA0000640C640C3A2A18D10A71A242A570A018C22063A81024489120594D103";
    attribute INIT_08 of inst : label is "1D1E0907827827827838A20820E083820E0838210BAA3357C544703C8138001C";
    attribute INIT_09 of inst : label is "305060A10182840604410255A51514A425320A27FFF800000007FFF80004733C";
    attribute INIT_0A of inst : label is "655156C160A5B058296C160A10B60B0508560B0220811AD790225C6928041828";
    attribute INIT_0B of inst : label is "CE8950540034799D1100AD6A100BA3A28115A002A01747423904040201080119";
    attribute INIT_0C of inst : label is "44A0280041A3A890580100142224454762545000A00140511D1400008822003C";
    attribute INIT_0D of inst : label is "100014469150120A0A38A08042007084002B8420015C21000AA87D7E00004100";
    attribute INIT_0E of inst : label is "200054A4455435688A2888000A2348A809050500A08042005084002AA1AF1451";
    attribute INIT_0F of inst : label is "23C8A809050500A0815291054A4455435688A2888000A23C8A809050500A0804";
    attribute INIT_10 of inst : label is "0043692039DC002B8088202EA2080BA88202EA2080BAB2080202018A2888000A";
    attribute INIT_11 of inst : label is "17D47A8BFFAFE210851A6D234C50D581585954556B664CF00555422F30D40000";
    attribute INIT_12 of inst : label is "0EBFEBBECFAFAEBAAF2845E504924A8AA83E1052405900A24010220B22FB88F5";
    attribute INIT_13 of inst : label is "42108421084007FFF7FFFFFC63FFC1085303050A215C42B0F7857903980C8055";
    attribute INIT_14 of inst : label is "400040800014010000045C0D818C02028AB08468380602D04C00100201701F00";
    attribute INIT_15 of inst : label is "0048142404A5A00A81E0E1D80620B03040000100000002C0000005445440005E";
    attribute INIT_16 of inst : label is "0E001155038166008C0E0011D50381006070008AA81C0881C0020AAA88402188";
    attribute INIT_17 of inst : label is "204A22304088816093E9028883C22207004081C0118620700035540E0476288C";
    attribute INIT_18 of inst : label is "85F008810BE0951A542508058002F9127E449A4A2201542508463F447C8F5205";
    attribute INIT_19 of inst : label is "801688B428240000BA15A114242A422F2000000025B05141CAA0450020C2F830";
    attribute INIT_1A of inst : label is "14339204186B4B40D44A027428FF555DD5DDC623080C280818E70C6000F7C00C";
    attribute INIT_1B of inst : label is "2449C943CD57558BAAE5D57534EAB10A7558853AACB221164E456D1111061CCD";
    attribute INIT_1C of inst : label is "0000000000010100000000000000011FFFFFFFFD5FD01FE017FFFFD5F72E484D";
    attribute INIT_1D of inst : label is "404929E0740093928622222223927F60909C4471020924410101010101010101";
    attribute INIT_1E of inst : label is "26422654A9595067FFFFFFFE48090180120B2448B24B3659948653CB02484489";
    attribute INIT_1F of inst : label is "5C01510018F3900FC14172A80149060120448102410172C64909924264909924";
    attribute INIT_20 of inst : label is "DDF77FF7FFFFAAAAFFFFFAAAAAFFFEFFFFAB4081000B515D101202B92223CB94";
    attribute INIT_21 of inst : label is "830F6DB7BB6F6DB7BB6F61B7B86F6D87BB6F6DB7BBEF77BBDDF767B399E777BB";
    attribute INIT_22 of inst : label is "836F6DB9BB6F6DBDBB6F6DBDBB6F6000000F6DBDBB6F6DBDBB6F6DB9BB6F6C33";
    attribute INIT_23 of inst : label is "9F3F77FBDFBF6FF7BF776DB7BB676C3783776DB7BB6F6DB7BB6F6187BB0F6DB3";
    attribute INIT_24 of inst : label is "742AC0055E492AF85EF755F48800000416C0F0BDEEAA6FFFFFFF77FBDFBF67F3";
    attribute INIT_25 of inst : label is "0000001400034000340000680A8015002A0054007B24D574DB557FFFFEAB0015";
    attribute INIT_26 of inst : label is "0014000028002800281A0681A0681A0681A0681A0681A0681A0681A00006802A";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFA000140A005002802800140280000500000A00";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "4000011600DA04008FA8FA8FD1FF4A4924F777777777751002458009249A8AA8";
    attribute INIT_31 of inst : label is "00124924D0B686C1040D00204701164F08A4D26DAFA22010BAA2480920001280";
    attribute INIT_32 of inst : label is "FFD757D5F57405900884008924C00561C0005122AAAAAAAAFAAEF88003C20242";
    attribute INIT_33 of inst : label is "000801124924924C000030404043E269041113E3C78E0F6C9FDFDDDDDDDDDDC7";
    attribute INIT_34 of inst : label is "78EAF1F6FB788BFDBEDF01100224924930A001EC0BC49249AF1838008924927A";
    attribute INIT_35 of inst : label is "E30001C4783D11E23E28D681A98701C5220046E30001C4783D11E235DE3EBC57";
    attribute INIT_36 of inst : label is "11E23E28D781A98701C5220046E30001C4783D11E23E28D781A98701C5220046";
    attribute INIT_37 of inst : label is "840CA081105008001E8402401E02141E28D681A98701C5220046E30001C4783D";
    attribute INIT_38 of inst : label is "1084000C00001C00246A8140C0FC40011028A060840080F00210001D5557478C";
    attribute INIT_39 of inst : label is "204062100DAA00000882050801602A8038048208E0847F488120051C05840D50";
    attribute INIT_3A of inst : label is "3D11E23DD800228A230001446A0A22A8E00162005445202A8FC02410020B8048";
    attribute INIT_3B of inst : label is "9B11122C0C88B032363C0D05CC0D004000800100A98701C5220046E30001C478";
    attribute INIT_3C of inst : label is "31674750151D74047090C64CEA29671648040764404E264624A9254111210424";
    attribute INIT_3D of inst : label is "FFFFFD8C001A01145018E10701158835037012024AD112200F0001C0110036D5";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
