-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9797979349294A02942528493FE22AAA6AAAAA712E050080A16135DFDEA3B3FD";
    attribute INIT_01 of inst : label is "210130DF1E20023F9E010DB2F915D4929A4CC000CE6575AA0AA098CE19679797";
    attribute INIT_02 of inst : label is "B4E1150552009416A045530284C0AA502861184C1B6A12EC39272882019A4C9B";
    attribute INIT_03 of inst : label is "7336492C92A3A8EDD893242211518A8C7473A39127F6F4ADF0521F62B642CFA8";
    attribute INIT_04 of inst : label is "8454F73EE5B7DE7BFDF79EBF79E7BFDE79EBE12ED77000888888888888C44091";
    attribute INIT_05 of inst : label is "D7680F5FBFC804C965E135DA64D4449A9B06CB0F616C3FDF7B25BB4959FE610A";
    attribute INIT_06 of inst : label is "44444444473CC8022202FB9B9412B26B27D8093A3684542D88C106142D94A466";
    attribute INIT_07 of inst : label is "0A5439DBB363C55BBCB8BF14E6675399DD4E6675399D725995F97F9CBEC08144";
    attribute INIT_08 of inst : label is "D868A044966B8888A4909EB010A0A00220002BB4ACACACA68C993060C281C685";
    attribute INIT_09 of inst : label is "4D140902E9024B2DB3EC49003129388DA450451A4CA8A28162965965D6E10161";
    attribute INIT_0A of inst : label is "6D9B27B24999FC4018B980C0840101010208808000C4CFAD9A00011644C4088C";
    attribute INIT_0B of inst : label is "7BF6B75FB5A7ACDBB5AADDAD3D76FDADD7ED69EB36ED6AB76B4F5CA4B267AC1C";
    attribute INIT_0C of inst : label is "6A1BFB0DDED08404B4A424B0A249437EB13191017208034007D7559575586205";
    attribute INIT_0D of inst : label is "0DFAB61BBDA10985A5212586124A1BFB086930DBCA586EE4C6262535B1258613";
    attribute INIT_0E of inst : label is "1446A0018EF3C0F03C0F00063776F99D3D99959994017AD892C226D437FC0DB1";
    attribute INIT_0F of inst : label is "FFFFD2048A95555111139234D34D34B0FFFFFFDB6DB6D2766E44B88C522C0561";
    attribute INIT_10 of inst : label is "A4E8C49286FEA661BCEE8CA380CEEC63CC718BACBA83AE967B6B0924B9CA2E19";
    attribute INIT_11 of inst : label is "7B89B50DFDCCC7F4992D18D210DFD449286FEA665F36E8C4DA86FEE667A54D37";
    attribute INIT_12 of inst : label is "F70E051233D19DDD5555AAA753A74517541295100454BA70A3DE6DDAD18DB61B";
    attribute INIT_13 of inst : label is "5A934244926CDDB64DDB64D6E94D3EC89B93BB847813E343E342E242E242E4DC";
    attribute INIT_14 of inst : label is "3EFC7DF8DBF1B7E1951477EF8FDF1FBE3F7C6EF8DDF2038A2B95C47B13FDDC50";
    attribute INIT_15 of inst : label is "02040810265BBAC39D9718EEB0E765C60DB614535E189EB0548E7EC9CFBF1F7E";
    attribute INIT_16 of inst : label is "02D1CC6633148C623118B558E73239114A5191A20A52ADB6924444000000B211";
    attribute INIT_17 of inst : label is "265D9B899666E265D60C652E8BAA6BA31EB31EBB1EB31EBBC220BE08C500002F";
    attribute INIT_18 of inst : label is "273DEC106002164A9D90CB041800869C925D440A8C98D519316697B9B899666E";
    attribute INIT_19 of inst : label is "0F692B4938E19965889FC63E6277EC5D86EE49928A516D903BA2945B64C0FEE9";
    attribute INIT_1A of inst : label is "CD0AA1BBBA2222720E9A69A696C373772490DDBAC8B345156B5A0BBA21F0E262";
    attribute INIT_1B of inst : label is "A3260E2A8C9938AA3264E3F363271DD3D8EBC8A496A496A495490D526A20BAF3";
    attribute INIT_1C of inst : label is "675464C59D5193161B9CB7186EE4921BBA60632BAB02C514555464C2A8C9830A";
    attribute INIT_1D of inst : label is "B14535551932AA3264EAA8C9938FCC538C377B490DDF7032B995316F0A4AAA32";
    attribute INIT_1E of inst : label is "DC0C2C654C5B8282AA8C98D51931635464C586E72DC61BB92486EE9818CAEAC0";
    attribute INIT_1F of inst : label is "FF9009E339662013847AEE40278CE598804E11EBBE2454C5B4F3E30DDED24377";
    attribute INIT_20 of inst : label is "90E91A0617742BC23287640ED650CE054AC21D68872FCC2AAA44F9FA7FCCF6C9";
    attribute INIT_21 of inst : label is "0AD3D1091E8DD34900103CB6A261427CA794EF24E05C27849B498DD152E3A8E8";
    attribute INIT_22 of inst : label is "48971A4A82DD6215A3744A0A0C42B468A8E89C38D68E8869A4DA3A258D146243";
    attribute INIT_23 of inst : label is "9921D149F5251500AF5217F8045A114802381887C327420A8819410440230C4C";
    attribute INIT_24 of inst : label is "1748C9084461236B5293739E8903CCDAD4A49CE19207997EBE6DF72133327324";
    attribute INIT_25 of inst : label is "E4B2591C8E4725D0E8F47A3D0C30C30C225DDDDD9111113AC5BEEEB7D9D1B761";
    attribute INIT_26 of inst : label is "485944715458BD32574E375164CB24921E96198B24924925DB6924324870C849";
    attribute INIT_27 of inst : label is "1EC9E4D7F3EF2732509EE9F4F9FD3FD286F64F3E64EE4A066F254585FB9597DE";
    attribute INIT_28 of inst : label is "3CB9BBA7D3A7D08EC9E4C9E4233A7D3A7D08EC9E4C9E4233A7DF133EFFA7BA50";
    attribute INIT_29 of inst : label is "1013E9DCF60FFB5E73FEEFE038731EDE7C6B971FFA901C6BDCFE38993C9AFBD9";
    attribute INIT_2A of inst : label is "BA6C3679705ACFDEDAAB6B37708F315FE3CEDEA0E1C0000E9E67DA3527DA92DB";
    attribute INIT_2B of inst : label is "0484F3CF5568803E039943EDAFFEFE064A85F4F40288C529B002A800252A28E6";
    attribute INIT_2C of inst : label is "D023CCEA11E674D9C49B7BB2B8EE84B67E7CD5FA7F0CA6F4D15C7C76F8EC51B5";
    attribute INIT_2D of inst : label is "34B460A17B51EDDC0B6D600000AAB7C575319BA6761D315DCE8E675733B447B9";
    attribute INIT_2E of inst : label is "1FF77E14BA6C5F35BA5C77ED0DC7B3CC91AD8F7EB2E34FF9EBA6761D45454545";
    attribute INIT_2F of inst : label is "3FFFFFFFFFFFFFFF667EBA9FAEA6EBA9FAEA7D6A7FF90A1F4B0AEF7777777EFF";
    attribute INIT_30 of inst : label is "0D71030008032003A6AE45191E25EF5596E1F897BD56E1D59F4251082B089A09";
    attribute INIT_31 of inst : label is "9615E1E8022044088150A3008C4208A8A71DD0404040007FCEE8200650214167";
    attribute INIT_32 of inst : label is "1DA91D00182051EA0190C1604CC00026535CEF964789DC601CA1C1158085963B";
    attribute INIT_33 of inst : label is "41F9FDFFD114662E62C444019F8BF1500C22E7A8001F188B89414787A2FAB333";
    attribute INIT_34 of inst : label is "00000101F4516E00000000020000000C0000009001000000001C550467F2AF15";
    attribute INIT_35 of inst : label is "33FFFFFF4927D3A76F400000000090080C30030E00007000024803C3EFF00000";
    attribute INIT_36 of inst : label is "DCF5D4000235E817EDF55DFDBD74FA4927FFFFFE633EE74E9FDF07F7DD3A7DC6";
    attribute INIT_37 of inst : label is "AE6540B4023E6A177028E9388E90A61F61D4F1F1C000F4E0F8C5C2ABDCD1393D";
    attribute INIT_38 of inst : label is "751D4741D0761D07C7FEC1FEB87FAA5FFF2EA97A41E9077D3B49DF6EDDBF705A";
    attribute INIT_39 of inst : label is "A7569DF6EFDB81CCCE4A77D3B53D1A9C06193D507672AAE4E551D9E029F2F9D4";
    attribute INIT_3A of inst : label is "A1958850FFF50078F001FEF17C3DDFBF800F00001E3FBFD50FFA87F6A5FBF2EF";
    attribute INIT_3B of inst : label is "4DCDE4264B944EB0BA0124C521442424000000000C000C004C4100000AA0A803";
    attribute INIT_3C of inst : label is "00000000122AA2D351A6A54D4772AA884128A21031C44411114A522294A44529";
    attribute INIT_3D of inst : label is "FFF1C01BFFEB8AA70F470D6E26AE349C5B1CD1B8D6BFD76337FAEC64B4023E6A";
    attribute INIT_3E of inst : label is "DEEDBD97CEB3C279B8EEDCD239CDDA4639CDDA44076D38027FFC7006FFFAE009";
    attribute INIT_3F of inst : label is "D2ED45C1871FC3334E5CAC382553A070F845AD0152D7F602B8222771009F8000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "ADE5ADE0024FDF5FBE9F7D00802643334CCCCC29F2162C04B3289E7E7E66E3F7";
    attribute INIT_01 of inst : label is "63AD7C2502529340216CB264A5B200240C999B6D99DA40145145111C8095ADE5";
    attribute INIT_02 of inst : label is "4E5FEB53A9CF9FBCDAFDA437D53BFF73FF6577A8043A4EDA8DC36DB0AABF5E23";
    attribute INIT_03 of inst : label is "8846C92592DCED326C2CD949E6223113888C449B3774EBD697F7B104473EBFEE";
    attribute INIT_04 of inst : label is "6EA49203392920AE165829C5960AF12482980B2480A000808080808080F93D9F";
    attribute INIT_05 of inst : label is "D2745BEADA82C92C9F4E4D24A9A99D3562F192D45E8B4349801926868464085D";
    attribute INIT_06 of inst : label is "8C8C8C88CC104003497FE431BB7FB36B6C95A76DEDBE9F6ED4C2F4CBF1D75ACE";
    attribute INIT_07 of inst : label is "DDF9E746CDB2343D726446E900F8A423A2900E9A423E04DE29333FA1BE3CB3CC";
    attribute INIT_08 of inst : label is "396D7D45926956520A6FC7C0000AA88938458201141414012FDFBFFEFFFB1B6C";
    attribute INIT_09 of inst : label is "EDAFA8A24DDAC92D964AAEDBEAD6C209D69F68129F6F36D45D4C0698448C9E7C";
    attribute INIT_0A of inst : label is "8002552494665BCFB20CEDAD93FFFFFFFDF3B3EDED90E92CB20002480D3ADA0A";
    attribute INIT_0B of inst : label is "156A5DAA526ACB6AD66F56B3564D7A97EB949AB25BB59FDDACD596DCCF2AEBAA";
    attribute INIT_0C of inst : label is "9D8486C20139CB2B4949D90E34939010E4652B6B969B50757205C760CC7209FA";
    attribute INIT_0D of inst : label is "C265D98406E316D2DADEC871A5BC8086F696E4061DB2011B8C4B5ACA4E5831AC";
    attribute INIT_0E of inst : label is "4688D77D2979E97A5E97A7B1649905AA4237765629540D6F2C185B7B090796DE";
    attribute INIT_0F of inst : label is "BFFFFFE7D7C26262626027496CB25B5FFFFFFFB6DB6DB6EDD8027419CE6D9F18";
    attribute INIT_10 of inst : label is "C997892520200A0810B50B42509333302604C2C808EC4B04E886404127296983";
    attribute INIT_11 of inst : label is "C116DAC24094384B76D2D12DE4060896D20204A0A249B38B2561200A1A71B240";
    attribute INIT_12 of inst : label is "4CB48BF0C02A83355555D544B84D96A076B28BFC86D924E46725B76D6516DD84";
    attribute INIT_13 of inst : label is "A7C4B6692CBBF66D9F2ECA83BFB248B24445065F46CA9A1A3ABA9A1A3ABA9E01";
    attribute INIT_14 of inst : label is "A35BC3B2AD6F4EC87B2F94B5793A52D5E4E95B57B3A75097C2C0B1258527660F";
    attribute INIT_15 of inst : label is "24599166A9226CBAF364D699269CC974AB2D61A66DB32D16D75C939728D6F0EC";
    attribute INIT_16 of inst : label is "CF2671985C79718DC263CAB0BF4BEA4D85DAE2DCEC2EF2597C8989919191C9E2";
    attribute INIT_17 of inst : label is "89D2E46235B9389D60AB4B92A06CD249E925EB25E92DEB2C9B936F131E64E45B";
    attribute INIT_18 of inst : label is "6F7BDCB35DBDAC9F7B27EF24D76F6B4CE1AAFBE0732240E644D8F8EE46234B93";
    attribute INIT_19 of inst : label is "609F8302655A824D69242099B73336E72000962D9CB39722A0672CE4C94A8116";
    attribute INIT_1A of inst : label is "9E9B3A4C4C4C4C04D92D964B6B2CB000496C223A35CDAE7E1EF3E687D269F186";
    attribute INIT_1B of inst : label is "1CC8BB2073236C81CC8F940A4A4C4B24B6B15F6B2D6B3D6B3ED67EF89E47F4B4";
    attribute INIT_1C of inst : label is "8B0399172C0E644DA4D2488200092D844C6E992EE8B72DB938039912073226C8";
    attribute INIT_1D of inst : label is "CDAE5E00E64581CC8B96073226D22B2CC30884B2400437449734CBB2DD9D01CC";
    attribute INIT_1E of inst : label is "9DD1EEDD1EEFD77F40732340E646DD03991F283596208006CB61123BA7DD9A75";
    attribute INIT_1F of inst : label is "7CCDF3BDE3498BEF7BCEB137CE739D622FBCE71A56BD37BD7B0730C2236C9001";
    attribute INIT_20 of inst : label is "3AB68F4DE59ED47E59F59ED04B3EB1DE1B6FD2D4E800012AAAD50FFAFE602952";
    attribute INIT_21 of inst : label is "5326645719126DB6332B8069C83CB0195B7B6A4916E3DB3B6D8032652D411F34";
    attribute INIT_22 of inst : label is "E365A59161E290E6489915F47E89E4499111023935511196C01544566AAE90B0";
    attribute INIT_23 of inst : label is "0809C4ADFB678811AFCC06A3677772DD906241A3F1030E4EF01DCA0565034106";
    attribute INIT_24 of inst : label is "CF1C406F0E2BFC2100402154B274300840020A4D24E8607D52F43E6580102101";
    attribute INIT_25 of inst : label is "894C82D328B0C82E328B4CE2E10C10C11E26A6A6A62626052C2DA185B03C2418";
    attribute INIT_26 of inst : label is "E17ABEFEBC92FEA7A8B782BA8A14CB2581788370C965B2C86592CBCCB20C13B7";
    attribute INIT_27 of inst : label is "79361BD50498D80DDDF9120982424026EDC8B0498B10BBB5FC843B9FD7ABAF7E";
    attribute INIT_28 of inst : label is "C1266CC864C8663B361B361B86C4824482639160B160B864C8645D0000C88CDD";
    attribute INIT_29 of inst : label is "2524D231DBA54D91A6010025860CA930E3B267AA8D29539431EBC762C17AA222";
    attribute INIT_2A of inst : label is "49A594B3526333F2C96D229963F7D0A1F7FFEF1BF7FBFED601F4054A4E213924";
    attribute INIT_2B of inst : label is "AE680205FF8DF97C7A5E7C69A81CB8999C6DE271BA55139BF80222081196ED9A";
    attribute INIT_2C of inst : label is "4E3632251B1112104AE048A9CC28E432F0003E2BFF2DEF91FDDCCCE0799CC8F1";
    attribute INIT_2D of inst : label is "D55A994ED99967D19C85F00000BBF84C9EC416B862B34BEB2275912A888E6C64";
    attribute INIT_2E of inst : label is "45E03E39E5A4EACB2CA8AA42B979A5C0A8149DFD64BC0703E6B862B598899899";
    attribute INIT_2F of inst : label is "7FFFFFFFFFFFFFF94B9A4F6293D8A4F6693D9BDD8005932C6C93357D7D757F6F";
    attribute INIT_30 of inst : label is "595803940A5022508D652CA15EC35639CBC47B0D58E7C460BF68DE2D3287EC40";
    attribute INIT_31 of inst : label is "D59FE55CD44A89532A2547371CCD598AE2AA904040432497D70466A9C59A1448";
    attribute INIT_32 of inst : label is "40883FA4C82A2BCB26130AF4D1E99268C0ECF99E88F0D4CA5565342F9FFA25AD";
    attribute INIT_33 of inst : label is "0A061201E14209D19D5051EA60741441021D185000008274664450781D052121";
    attribute INIT_34 of inst : label is "3019CB971FFFFB973C30B394E1859CFFE187DC28609EF830FF1E502A184D5794";
    attribute INIT_35 of inst : label is "7200000069A453A000A0CF3C73C427039EFB87BB97DFF5F394D1C86E3119C86E";
    attribute INIT_36 of inst : label is "0B82A888828AB26AD15FF7E002748A69A4000000E722074E821000841D3A440E";
    attribute INIT_37 of inst : label is "EE0986F8074C5F138166A3406F8924D61D6C1D7208FCAD04E035C06BBC944442";
    attribute INIT_38 of inst : label is "7ADE77ADC372DCB737FE69F5225FCC97D54F327C09F037B23D916C8B2A38EA94";
    attribute INIT_39 of inst : label is "578B56CAB5AB8DCA6E137993AFBB97DC00073C34B270636CE0C2C9C819F189E7";
    attribute INIT_3A of inst : label is "B722D424910AAF85156A2115C00004043F10F8BE21E23FAB6FDEB5F42D7516F7";
    attribute INIT_3B of inst : label is "49F689B493E50E9F920200DC04650D0900444441454D49416D61AAAAA0A0089E";
    attribute INIT_3C of inst : label is "00000000034C835BF9B7F76FE69B0B25156AA9453CC51505414A528294A50529";
    attribute INIT_3D of inst : label is "FFF97FE2C03390D7037516AA15EE591C03956628C73B6100276C2006F8074C5F";
    attribute INIT_3E of inst : label is "2996C208B3E57D92442F5A353C0040243C00402607893C057FFF5FFAB00EF011";
    attribute INIT_3F of inst : label is "4122CA4597EE6BA3AC35C4B8C4E50C2562204A2241C34C803A00257E0B300000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "BFFFF7B9548B1B86372C6E40DFC233C390F0F04252F48950210C2A2E2E77C91E";
    attribute INIT_01 of inst : label is "522A5F02E0108302DFB58DBFD984B508A926649265712DE79E79EE5F48CFF7B7";
    attribute INIT_02 of inst : label is "CB55ED7A230C552694E58C73C307BE1FBE215738E0001CE3F9E36DC802FFFF48";
    attribute INIT_03 of inst : label is "48C6D96595CF5C4CD1D13563C3331998ECC766385C0986C329898A28863AEFEF";
    attribute INIT_04 of inst : label is "A72EB37DCB8AEFFD2EABFF0BAEFF52EBBFD4FB64FDDB333BB33BB33BB3E326DC";
    attribute INIT_05 of inst : label is "F24CF58FBFA76976B57335CE67B304F67DB4CD39A33462FFFDBDBCC8C4B638F1";
    attribute INIT_06 of inst : label is "155115511145105799A49E619DB493D92496DDC3AD36592A44A0EE8B89B7338D";
    attribute INIT_07 of inst : label is "9366CD9B364CD9A2448911CDAAFF36ABFCDAAFE368BB64DB8D933FB5BF729455";
    attribute INIT_08 of inst : label is "104131CC96D966C72A492DC400000E4CB40DC8852D2D2D2B099326CC9B326CC9";
    attribute INIT_09 of inst : label is "28263D86FCCE4B64924A224D2CC6171F2759623E7B0C32EEF15F6BBFB6DEBC3E";
    attribute INIT_0A of inst : label is "C4CB9292DCCE821E675EF6B6F80101010100E73676B84B64B25042EE04AB6F1B";
    attribute INIT_0B of inst : label is "76AE7A3473672CF1F7C387BB396387BA1C3DD9CB0D1CD468E6CE5D1A6D870EB4";
    attribute INIT_0C of inst : label is "66195D0CCCDDECCE647476134E68C32B31B9C94B134A5D395E175DD7719D2E62";
    attribute INIT_0D of inst : label is "8E8E631DD9BBDD1323A320DB7B471D5D1CED38EAE66C7666EF767323A330DB72";
    attribute INIT_0E of inst : label is "E71CE379CE69AB6ADAB6AF39B724131B6EB8971C8C5791D1D04CF68E3AA89DA3";
    attribute INIT_0F of inst : label is "BFFFCE6CC563773BFFB9933692493666FFFFFFFFFFFFFD896DB4B62EB5AF3922";
    attribute INIT_10 of inst : label is "B4C98CD18645C6A541E55E0781E4E6C2D85B0B0D9675B5975E63996DB99B1A0D";
    attribute INIT_11 of inst : label is "571DA38E8B8D6E269D1D91DA38E8B8ED1C745C6B7134CD8CD18645C6A758DB7B";
    attribute INIT_12 of inst : label is "F344C995F0D98CC2AAAA8AAF2D3668AC18A04999A65CB0FA2B8269D1D31DA71D";
    attribute INIT_13 of inst : label is "6562B3649B4C1D0745D9731C44DB7AE77EE319A686E434B49494941434343B38";
    attribute INIT_14 of inst : label is "366EEDDDD3B1A364FB266ECE8D8D1B9B7776ECE8D8D359930703C1F303DCCC37";
    attribute INIT_15 of inst : label is "D1336688ABFB38CBB9C65DCE32E671D72FF6F2103801989897D664E9DD3B1A36";
    attribute INIT_16 of inst : label is "CF835CAED77C5AE5763BE3DFCF613308EE5837664772E536F767771B391BE3CC";
    attribute INIT_17 of inst : label is "0E1D8783C761E0F1D3EE72C779ACF3B31C3B1C3B1E3B1E3A7B391331DF064EC4";
    attribute INIT_18 of inst : label is "8421080149C9834A10D102005272665061CA66D8CE88B91998723E987038761C";
    attribute INIT_19 of inst : label is "6E6ECF59ECD9A87589BD86552FAA85F5867661D83E07C592BD0F81F1608AE75D";
    attribute INIT_1A of inst : label is "9A9C186EE77FF7324ED24926CCCF233B36D0CEB2E3E05F0794ABB33A1929B7AC";
    attribute INIT_1B of inst : label is "33A26E9C8CCC3A633A20C323731CC18C58C72C4EC84ECA4ED49D90AC56532535";
    attribute INIT_1C of inst : label is "36C674499B9199B6191C62186766DA19DE4664738AEF9B7CDEC67449C8CCDBA6";
    attribute INIT_1D of inst : label is "F6DFA7319D13723334CD8CE89B0CCE310C33B3698ECF233A398577CDBE6F7233";
    attribute INIT_1E of inst : label is "48CCCE6179FA6FD39C8CCDB19D1266E46669C76718C71D99A4C767919D9CC2BB";
    attribute INIT_1F of inst : label is "BD10CDE62D722193CC52C4632798A588C66F314B171E3BDEE747638ECCD3433B";
    attribute INIT_20 of inst : label is "DEEC93D76622C8D270C622C80E18C45D13CB1846648C019154DDEF56D56CADDB";
    attribute INIT_21 of inst : label is "1B8ED239099F9245545551239C79C240E05C0F36FB5AE01C76C977D331040E64";
    attribute INIT_22 of inst : label is "6B82324B90F8CC7719F48E2AAE3DA0C099DDF23181999DC7649777630334CA64";
    attribute INIT_23 of inst : label is "584C4EB3010F6914ABFBADD44FEB80DE481A38A3F903042A39BD466D4317438E";
    attribute INIT_24 of inst : label is "4B1ED44D0A3FFC4290E55ACCB3777410A42B14A936EEE8C532F8E07960B8AB41";
    attribute INIT_25 of inst : label is "341B0D148A61B09269B65369345965145A73BF73FB377396C8BFE717FCECBF38";
    attribute INIT_26 of inst : label is "D3BB18FECC1AFE378ACC9298A2EDB49204922D59B69349B0DA49B49B489068E8";
    attribute INIT_27 of inst : label is "1468F65D9A65A31B0E9468F60D2D1AD876A367A6366B41C76A25238997B3A73E";
    attribute INIT_28 of inst : label is "9ED8B9B3D1B3D30E68F668F6C39A3D9A3DB2E6CF46CF4CB9B3D3130665B31A0E";
    attribute INIT_29 of inst : label is "30369B55E2FCB36A78A667E5B8573B576CC9CAF151B15AED55F139CD9E8BBD8D";
    attribute INIT_2A of inst : label is "35159E9A5360CFC0A520888512606F80F5E715188506108C04F870246E0981B9";
    attribute INIT_2B of inst : label is "386288C2AA81F27C7773785B6B14AEDC266436853AC7BAD2000282201990EC19";
    attribute INIT_2C of inst : label is "8CBBE7545DFBA0628CE1693ED14CE410B3366F23FE2DFB01E8879FB48F2792E3";
    attribute INIT_2D of inst : label is "75E9D1EFF19BC7D516E9F55555EBFF4FEFF3D98C10BD699F746F3A27DD0877EE";
    attribute INIT_2E of inst : label is "B7F73E2DFFE8BB6FFFF6DDFFB7FF370CB3BD97FDFFFE406BE98C10B4CCCDDDCD";
    attribute INIT_2F of inst : label is "7FFFFFFFFFFFFFFE6ECFF7F3FDFDFF7F3FDFDEFFC005E9CF6EE3BFD57FDFF5BF";
    attribute INIT_30 of inst : label is "92E8B78EDA314A388D4949654035D65F518000D7597D80693F4E03A1AAA1BC00";
    attribute INIT_31 of inst : label is "AE8BE3F4664CD9B9332667199C04C88636A29AE8CAE3202FD7042154031626FE";
    attribute INIT_32 of inst : label is "083001203B6E022301C0C6840D089006C81070038045D0423F63AA6B81082FF7";
    attribute INIT_33 of inst : label is "B5FBEFFFFD69362EEA8F5A159F8BFC623162E7A800004D8B98C44007E2FAA121";
    attribute INIT_34 of inst : label is "2011366C1041226C13CF6E6F9E7B73249E7913F79E6083CF005F96D16FBAAFE5";
    attribute INIT_35 of inst : label is "DC000000B6D82C5890010413C103FCEF659679626CB28B2E6FBF365820973648";
    attribute INIT_36 of inst : label is "8B8080A0A81770DDF57D5542408B05B6D8000001BDC118B16020800822C5823B";
    attribute INIT_37 of inst : label is "0A0E08FC035239164820E7240FF24254A15CD1F92400FC92E4D1C583D08DDDD8";
    attribute INIT_38 of inst : label is "5C1745E1585415058500C14A08504254212BC17E51F815862C9161AB42BE8860";
    attribute INIT_39 of inst : label is "D7B75E38FAA381E8AE657A4B9C3F8E1C011A3AC0A0758140EB0281E045D0F578";
    attribute INIT_3A of inst : label is "2D061C61000054020AB4010E45862040E1E00F43C00038002E2B970941CB40F1";
    attribute INIT_3B of inst : label is "4B070000060FE120760408FC414F4A4C020005414745454D4848FFFFF0FAAE23";
    attribute INIT_3C of inst : label is "0000000033093455FAABF157EC180BA51128894460055455544A52A894A55129";
    attribute INIT_3D of inst : label is "4001602A800B9D570517128E700A491438152AA8E0AEF1A055DE3408FC035039";
    attribute INIT_3E of inst : label is "244D090FBC50DB731100C3E02840698A2840698807A0BC0577F97FF8EFF0BFF1";
    attribute INIT_3F of inst : label is "10001090118BEAE0E9B298609120A219003142C8847F468ABAAA947F01550000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "72323239548B9DD73B8E7740CA0203FC00FF005A44EB8955010448C8C9D6584E";
    attribute INIT_01 of inst : label is "3A0674104A121D42FBB1AD96DAACB508A937679EECA924C71C71DDCACCDA7A7A";
    attribute INIT_02 of inst : label is "DF306E1BF586C57610FAF65A7595255D25450FDEE2220989C15434F8A941A360";
    attribute INIT_03 of inst : label is "E042CB24955445C8919125BCB111888C4462232A0A03577961A5A2A22E1ED7EA";
    attribute INIT_04 of inst : label is "262492A50B0CB3B54F2CED53CB3B44F2CED13B24A82A2A2AAA22AAA2A2AD24EF";
    attribute INIT_05 of inst : label is "B27A88B525412512653366B606AD08D5B4D55148290526FBCDFC940E499230C1";
    attribute INIT_06 of inst : label is "D9999DDD9B6DDF696924D4A0393CB6D9249ED94F927AAF2D4672FB13FDFF628F";
    attribute INIT_07 of inst : label is "200000000000000000000D85FA4E17E93C5FA4F17E93BC438FD1083C817C7799";
    attribute INIT_08 of inst : label is "C9C1D4019259CCDA2B6D5EE00444472E780CA8D52929292A5020400100040010";
    attribute INIT_09 of inst : label is "383A83A0DAD6C924924E234939E7DA03F28AAD0669D5D65431FBEFBFB2741F34";
    attribute INIT_0A of inst : label is "C6C97292CEEDA72FA23E36F693FCFCFCFDF72B7676D0292492EBBB42008F6A06";
    attribute INIT_0B of inst : label is "2B95EE5CAF45F71C2B70E15A2FB8C15B060AD17DC70ADC38568BEBBCFF85F59C";
    attribute INIT_0C of inst : label is "6619190CCEFDFDCD6C76741B66ECC3239514B44A2822503476DB9EE6B9EF266D";
    attribute INIT_0D of inst : label is "0C8C6E199DFBFB9B63B330DB3766191D1CDDB0CAC6E86677ADEC7B63B320DA37";
    attribute INIT_0E of inst : label is "63EC77BCA596D5956D59579BAAE413917C98AB4B8D1D31D9984C6ECC32389BB3";
    attribute INIT_0F of inst : label is "3FFF88317FE5111D99999BA4926DA475FFFFFFC92492493692491094B5815BA0";
    attribute INIT_10 of inst : label is "34CD8DD98646C42F55755755C17EEEEBDD7BADEDB26FBEF2B72D4B6495DF7E09";
    attribute INIT_11 of inst : label is "5B1BB30C8D885E369D9991BB30C8D8DD98646C42D1B4CD8DD98646C42FB8493B";
    attribute INIT_12 of inst : label is "A2ECAEB0918928A08888200ADD275D942CC6AFB1DB8516562AA369D9931BB619";
    attribute INIT_13 of inst : label is "EFE23ABCD36E0F93E4F03D8EF249735A344251761660B0B0B0B0B03010101750";
    attribute INIT_14 of inst : label is "D5AD2A5A54B4A96C8E3AAADAB5F5EB6A96952D2A5A54F95D6566589602B8B81F";
    attribute INIT_15 of inst : label is "F9E2C58AD2CD1E71C8F38E479C723CA3B492D36B2379A10EE80A9054B56B6BD7";
    attribute INIT_16 of inst : label is "F4F5EAF57AA7EF57AB553F4F5FAD976D4BAF1F23EA5D5DA49B544445C767BCBC";
    attribute INIT_17 of inst : label is "A68E3369A38CDA68FA352FD709366524559C559C559C559FCF75D7DAA9F65D77";
    attribute INIT_18 of inst : label is "FFDEFCE2B9BDB34B8CD13B38AE6F6E70B8EBEEEC9DDF19BFBEAD7E03369A38CD";
    attribute INIT_19 of inst : label is "67EDC149A4E90FAEA0BDCF22D4CCDA9BA7767AD653CA7BB03D94F29FEE40F649";
    attribute INIT_1A of inst : label is "090F1AA223B333336C924DB48EE7C3BB3EB0CC96B13CE9EBBBD7F7F959F0E3A5";
    attribute INIT_1B of inst : label is "37E6D5CCDFDFD7237E6F77A93D6D4AB4AA5B5584C984C984D70993FC443B4723";
    attribute INIT_1C of inst : label is "6E64EEFEF99BFBFBBD4E6E3866779F1DDEDE7E7D7AC4B2A5EC64EEFC89D9B572";
    attribute INIT_1D of inst : label is "2CA97B91BF3622766D78C9DDF5DEA7371C333BCB8ECD6F3E3AFD725DD2D62276";
    attribute INIT_1E of inst : label is "5BCDCEBF5C9774B5CCDFDF91BF37BE44ECDEEF539B8E19DDF5C767B79F1F7EB1";
    attribute INIT_1F of inst : label is "BFB8D967A9AF71B2CF535EC3659EA6BD86EB3D4D6B2F1ADEA7E2C70CEEFAC333";
    attribute INIT_20 of inst : label is "E258DC42EAE3DDD27B52E3DC8F2A5C7F81ED4B64E70644AAAA0C95FE7FA4C5CB";
    attribute INIT_21 of inst : label is "35B4922FA08900054551410368117FD0AA15413E3B68AA17FB7FA1931C4515C6";
    attribute INIT_22 of inst : label is "5EA25656BB78CC6F6C6483A2A3C9210308CC9160ACCCCD5FBFE2222551115660";
    attribute INIT_23 of inst : label is "D808345EAAD0D5AE405051144CCDB0CE48181883E9C3022278AC402900158503";
    attribute INIT_24 of inst : label is "CE0EC05DEBE3B95214C01A9D3BE06454852244A0B7C0C84926280B2E81B03B01";
    attribute INIT_25 of inst : label is "36130994CA41A0D349A65369B6114514015D5111DD51119A599B44336899DA20";
    attribute INIT_26 of inst : label is "D19F4CF600C9BE92A3489398E347249A0E934D9D34936D209249B692483068EC";
    attribute INIT_27 of inst : label is "CDE9FF8CFFFFA71F8D0DE9FFFFFD3EFC686F6FFFF6EBF1B2A6AC61190261611F";
    attribute INIT_28 of inst : label is "3FFB57A5F7A7F777E97FE9FFD5FA5FFA7FF57ED7FEDFFDDFA7FF6A1677A79E8D";
    attribute INIT_29 of inst : label is "1C17CBD4BEA8BACF56B66550987F93566CE9D0797CBC1FFDD498F9DD3FB19FFD";
    attribute INIT_2A of inst : label is "55069A6AAAD377E921F028D66730BFBF1530DF5B873BDEE80EABDF39CDB8E0B7";
    attribute INIT_2B of inst : label is "7B6CC80488A0B83F3D207E16488280E8CB6BDCFD9D5111C9A0000080329D4550";
    attribute INIT_2C of inst : label is "C95DE774AEFBB94587FB331F52C7F850F71C4C485F9890F88AE1F8DE83F0F85A";
    attribute INIT_2D of inst : label is "61EA54E7AD76A0356FEB255555ABD2292972F10F62DE79D6764B3B25DD9DBBCE";
    attribute INIT_2E of inst : label is "93F35F8CD3E975BE92DD772B6ECE13D57AAD2B7BD7665031118F62DC44455546";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFE26F494BD252E494B9252E632FFFA5CBBCE5FFFFFD55D7B9F";
    attribute INIT_30 of inst : label is "08A515805200280985280C203E00C11705A27A13055C22411F040B8181899A00";
    attribute INIT_31 of inst : label is "2B49E680E59CA394768E533944C4C880348010404260840FCA804444A59EB6A0";
    attribute INIT_32 of inst : label is "019C098451481B432182C0A0CE4142274A5E31C1812540586A06CA21952D0B59";
    attribute INIT_33 of inst : label is "A00DFDFFF680C1D33505A000607402DCC095185000003054650D280015052121";
    attribute INIT_34 of inst : label is "CFE673E5E4104CE5D7DF26E4BEF937493EFA672FBFC103DE005F6A80B7F557DA";
    attribute INIT_35 of inst : label is "1000000010402040100175D7DD7F25E2E8A2FA2CE5148946E4D3718BCE637193";
    attribute INIT_36 of inst : label is "D5DFFD77D81557D53422A0004008041040000000210100810020780802040202";
    attribute INIT_37 of inst : label is "0ACFEAFC025818122820AF140B80085F01444160A4FCAC52F405C20B91655557";
    attribute INIT_38 of inst : label is "5F1785C14050140505FEC570C95FF017D70BFD7E05F8056CABC5590A883ADA01";
    attribute INIT_39 of inst : label is "95085592A48B85D42E217B0B8CBB865C0500B900E17201C2E40385E001F2D17C";
    attribute INIT_3A of inst : label is "53061C600008040010200000024200000000000000002FC42BDA95F3857072AD";
    attribute INIT_3B of inst : label is "0107E492420FBA6AA40848F4404E40464044480E0A080A08446855555F00585A";
    attribute INIT_3C of inst : label is "000000003067B78000000600041BB00C5062831420C00154550000AA00015400";
    attribute INIT_3D of inst : label is "60154002C02283150B550F2A48AA3C544154F8284A2A146655428CCAFC025818";
    attribute INIT_3E of inst : label is "62B0C68A3AF53D42AC2A56602B191B8A2B191B8A07A0ABF958055002B00AA005";
    attribute INIT_3F of inst : label is "500C040C018BF2A44998A16AA40808801A25283814600C88900A007D94978000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "363636319115846919D611970AB57C001F00000EC3E200A15A53C02C2D440D07";
    attribute INIT_01 of inst : label is "42D5461A8751505284C9280D1420285506181201810FEDBEF965B0D88CB63636";
    attribute INIT_02 of inst : label is "017603608C59E83550C82824921249124917BC9102854088896C061400C16286";
    attribute INIT_03 of inst : label is "0C808240011451332526CE052333199AEED7764690001112052122B760A53063";
    attribute INIT_04 of inst : label is "D9A30502161140241050090414024105009002002088088088808800888A0902";
    attribute INIT_05 of inst : label is "20002A2A8ACED96D8718D860221A0443201330C0180303498043609607FE31F4";
    attribute INIT_06 of inst : label is "444440004114050050492A41A6CB2490400336805209C2C0348A90024126DB09";
    attribute INIT_07 of inst : label is "000000000000000000000244E2CD13AB344E2CD13AB310C36D63003DC0604004";
    attribute INIT_08 of inst : label is "05544CCD20121494418080054505039F944CD068404040488000000000000000";
    attribute INIT_09 of inst : label is "AA899926909490012000B4B24290A41A11C21A3420618E380D2480006D883248";
    attribute INIT_0A of inst : label is "C8884AB6DA88901C540019196155555555516ED95920500901FBA88004019418";
    attribute INIT_0B of inst : label is "668C6AB563D8213063458B1EC109A31AAD58F6084D18D56AC7B042586C382134";
    attribute INIT_0C of inst : label is "9401900089319908494952002492803286CC274E8CBA71255830B02C0B42204C";
    attribute INIT_0D of inst : label is "00CA48011273B2124A4A1001249401945492400E84A00449CECA524A4A100024";
    attribute INIT_0E of inst : label is "80B0122461451765D97454804092072378B0024221560525082049280322924A";
    attribute INIT_0F of inst : label is "7FFFC2343403333BBBB164DB6D924942FFFFFFA4924924804924820B8C637612";
    attribute INIT_10 of inst : label is "4920092500650846F81AC1B07811919232464840084E9340CCD874DA07127106";
    attribute INIT_11 of inst : label is "D4124A00CA108D0922542324A00CA0925006508448492009250065084440DB62";
    attribute INIT_12 of inst : label is "001A8267802A30175F5F7540A0C892AA12ED0270C1838EC46670922548324801";
    attribute INIT_13 of inst : label is "A4000C1B2491C2609C270A1808DB62142AA4600F1EA8F878F878F8F878F87121";
    attribute INIT_14 of inst : label is "F1E1E3C3C7878F08A209EE3E7C3C7878F0F1E1E3C3C51104C851144504644424";
    attribute INIT_15 of inst : label is "264C99321D230410582082C1041608208DB6E0A431A173120FF1B6183CF8F8F0";
    attribute INIT_16 of inst : label is "542B1A8D46A118D46AB50ADEC80DB26CCDC2BB77666E136DF6EEEF7575F50D23";
    attribute INIT_17 of inst : label is "6CC2B65B30AD96CC22010A411446C04D220522052205220585D53955A85D754E";
    attribute INIT_18 of inst : label is "B50D42CA3F393936D64D98B28FCE4B63ACA09B3100012200030BBA8B65B30AD9";
    attribute INIT_19 of inst : label is "E13E4620882A301861B54822C4C4789E6055BC4310E21E62058430869E081440";
    attribute INIT_1A of inst : label is "198193777777762CB36DB2492845C02ADA0828A7310CC8728004548D1894862C";
    attribute INIT_1B of inst : label is "401143D542450745080434920850AC2A821563806C806C806D00D88000AAE626";
    attribute INIT_1C of inst : label is "0488000C32200031A4824920054948015C0E86107CE43B218AAA122D542450F5";
    attribute INIT_1D of inst : label is "0C8872AA008A55091619542458D241249002A4A0008C0743083E621910C54400";
    attribute INIT_1E of inst : label is "81D2C30F9C876439554245A284020E88000869209248015250004603A1061F31";
    attribute INIT_1F of inst : label is "BC689110E618D12221CC31A24443986344A88730D3EF9B9EE7002400A92820A3";
    attribute INIT_20 of inst : label is "6E36EDD1808BB46C58308BB41B0611728168C204E92100440019A5545520058B";
    attribute INIT_21 of inst : label is "B328669689986DB40011100A5025B902D84B02DA0CB2D85B0DA440662C501137";
    attribute INIT_22 of inst : label is "9B69A59978E69D665019A5AA20B048D09999E11939999990D266667673359500";
    attribute INIT_23 of inst : label is "4008A850500140105544140006651A8C0141451020106F74F696A9A5B41A2204";
    attribute INIT_24 of inst : label is "CC0600CD8B86B410043010CCFB2754061185063AB64EA844CC29616460800801";
    attribute INIT_25 of inst : label is "00010090482090492410880400030C1009333333B33333113FF6C4FED89FF621";
    attribute INIT_26 of inst : label is "31848258029C01B86A1304228A3C00010258261010012490492400C000883680";
    attribute INIT_27 of inst : label is "4110082AC98040244941100844C207224A08A0580A0C8931A0A5985540585C01";
    attribute INIT_28 of inst : label is "03240440284028A110081008284402040208114081408284402C8C295440A549";
    attribute INIT_29 of inst : label is "999689F598B0AC9180A845448005A174663242694C9102B5F5A80C4603455046";
    attribute INIT_2A of inst : label is "04400012280EA82020543029A7074F60C594A512B556B5D010AA60122414DCB2";
    attribute INIT_2B of inst : label is "B64ACD08828E0B80880064DF6E36ECA4144E0B095112A8409A88020140072304";
    attribute INIT_2C of inst : label is "E70C15638202338D8C6F6F3956CC6854BF5C6E0D005000103BA180891318A815";
    attribute INIT_2D of inst : label is "618452617C15F02C065910000010413B6921B30DC28466695634A31A15C70828";
    attribute INIT_2E of inst : label is "B617804C32D8332DB2C41163A5CD328E399B0601B6E687A0138DC280CCCCCCCC";
    attribute INIT_2F of inst : label is "7FFFFFFFFFFFFFFA64CDB4936D24DB4936D24E724002142706159AAAAAA081B0";
    attribute INIT_30 of inst : label is "6E03D2D34B41A3412438963AFFACA1C4B5357CA28612B55F10B52B11D9551360";
    attribute INIT_31 of inst : label is "60081402B43786D0DA1B40AD02E9952B52C284040403568028A354CF3963C600";
    attribute INIT_32 of inst : label is "7EB0A356ED282F1AB64B288AF005AB781FDF75EBAD2CA6A540140670531F3003";
    attribute INIT_33 of inst : label is "8A161201E8A40E2DDAF2280B9F8BFDAA844AE7A80001032B93F208004AFAA121";
    attribute INIT_34 of inst : label is "281473E4038E00E437DF26E4BEF937003EF8072FBEFFFFDFFFDE222C584AAF88";
    attribute INIT_35 of inst : label is "000000000000000000010C37830725F2E082F820E4107106E493724829937250";
    attribute INIT_36 of inst : label is "FD5D75D7581FF75575F777600000000000000000000000000000500000000000";
    attribute INIT_37 of inst : label is "01E00A1DC4036101A54A0852A07367231428041A93FF014812240448240FFD55";
    attribute INIT_38 of inst : label is "806018060180601810FF2036000F8603C000012ED4BB504002201000000002A4";
    attribute INIT_39 of inst : label is "003C01200300702380040060300018000484062404044A080890100800030201";
    attribute INIT_3A of inst : label is "9E8E38E000000000000001044240000000000000000007C601C100FCE0360008";
    attribute INIT_3B of inst : label is "B2AC1249255FFF4CC61001B400050006010E0001030301010541AAAAF0AAF7DC";
    attribute INIT_3C of inst : label is "000000003C000820044008800AB44452AA9554AA55F2AAA9AAB5AD556B5AAAD6";
    attribute INIT_3D of inst : label is "201000004020020008C0080024802200470080008600050F5000A1EA1DC40961";
    attribute INIT_3E of inst : label is "0224A4BCF2604B9AA8D5C00107BD420A07BD420A000200000804000010080000";
    attribute INIT_3F of inst : label is "C9562AAD54000A302020300295012A28420C080C04990AAA2A8200FC8AB28000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "24242426C225AECB4C9299C03D266000000000D94A0C2BE5130035D151660B8F";
    attribute INIT_01 of inst : label is "6760EE079650964DC8DB292483210C2784D55B6D555A4934D34D2B01B6942424";
    attribute INIT_02 of inst : label is "20D5372D9CC38C3050996B0D32C0D300D3042588EFE802E5EFFC7C1354C1E399";
    attribute INIT_03 of inst : label is "899249249095491225244C0823331112CCD4441614828192412126466A8D9057";
    attribute INIT_04 of inst : label is "5CA4934001104024841009200002480000920124AA00800088880000884A49B7";
    attribute INIT_05 of inst : label is "9272232FBF87F87F9B9ADD60201A4403241114E69CD39820104000A7342442D6";
    attribute INIT_06 of inst : label is "44444444011045065249E948925992492491339CE45DB6E83592BC22F096CB24";
    attribute INIT_07 of inst : label is "00000000000000000000066DA608B69826DA609B6B8246026928002001A5C040";
    attribute INIT_08 of inst : label is "11464C4492491594E912E095455003E54048184C6C6C6C600000000000000000";
    attribute INIT_09 of inst : label is "A8C98B224A9249249248A4B262948489CCB2DA1200596D998500824120097229";
    attribute INIT_0A of inst : label is "C192D726439490CCCCC10989E40202020208AA495BA44924931550984401BC88";
    attribute INIT_0B of inst : label is "64894A244A765B204A410253B2D9025208129D96C812904094ECB6594CD65B34";
    attribute INIT_0C of inst : label is "B4C3A461B361194A5B5B4927ACB69874AC45675AC4BAD6A55925A5695A1640C8";
    attribute INIT_0D of inst : label is "61D058C366C23292DADAC93D65B4C3A4D496E61F05A30D9B4AC852DADAC93D65";
    attribute INIT_0E of inst : label is "949296A52B4D374DD356DCCCED9B27180103225629564D6D649ECB69874692DA";
    attribute INIT_0F of inst : label is "3FFFA132B5322222222226DB6DB6DB4BFFFFFF800000000000000009CE4152C9";
    attribute INIT_10 of inst : label is "DBB3C96D30E9668A40B10B42C0B3B3B676CEDADA60480825A44AD2012C2A4893";
    attribute INIT_11 of inst : label is "E592DA61D2CD141B76D6792DA61D2C96D30E9668A0DBB3C96D30E966884C924C";
    attribute INIT_12 of inst : label is "CC9AB265C269A3280AA00005A65DB2E912BD3263CD91E40CA321B76D67B2DCC3";
    attribute INIT_13 of inst : label is "95300ED92C9B16C5B56D5A5994924CB4E993464E87B4B4B43434B4B4B43439AC";
    attribute INIT_14 of inst : label is "A149429285250A490049849429285250A4A1494292840224D2DDB66C93132244";
    attribute INIT_15 of inst : label is "264C993234020DB6D06DB6836DB41B6DC92444ECAB656B62788DD8B5685250A4";
    attribute INIT_16 of inst : label is "952A52A954A952954AA548968049A04C9992A25464CC92491488880505054823";
    attribute INIT_17 of inst : label is "60B610582D84160B640B587812EC1ADC1B6C1B6C1B6C1B6D4AA52A552A6B694A";
    attribute INIT_18 of inst : label is "400420A2E92928BF422DA828BA4A4B42AAB499323932A472645AB9010582D841";
    attribute INIT_19 of inst : label is "699C6200000583CF292670D525AA84B070C9B42D14A29078C24528A51A231D86";
    attribute INIT_1A of inst : label is "C351D24444444444BB6DB6DB6964A864D9661B1521480A464004584498849445";
    attribute INIT_1B of inst : label is "8E4C8B523932AD58E5D8981C5AD2916916B4A9036D036D037E06DAA6016A6044";
    attribute INIT_1C of inst : label is "D8B3DBB562CF6EC4C0D659C30C9B24C320570A2AD48520291991C99523932AD4";
    attribute INIT_1D of inst : label is "480A566CF6ED59EDD8B567B76A606B2CE1864D9661B02B84116A529494ACD9ED";
    attribute INIT_1E of inst : label is "0AE1455A90A40523367B76A4F6655A91C99130359670C326CB30D915C288B521";
    attribute INIT_1F of inst : label is "3CE59635F759CB2C6BEEB39658D7DD672C91AFBAD4284118C31038619365986C";
    attribute INIT_20 of inst : label is "66B68CF5959A9626CC959A9789D2B352E13A564570090111546EA957556A21C3";
    attribute INIT_21 of inst : label is "B7296FA60DD86C96232ABCA6522534B69ED3C2D94DC61EC30012486ECEF2A934";
    attribute INIT_22 of inst : label is "EC78849660869F6E521BE9FC7CB27870BBDDE41427FDDF10095FF76C4BBD189B";
    attribute INIT_23 of inst : label is "610DE9FFFFFAECAEFFAAABE95EF7328C9270610422064E666DF4C97D24370A44";
    attribute INIT_24 of inst : label is "4C470155AB0232CE77A7AD85B103C8B18D69EB6A1407918DB29AF21D62C22C05";
    attribute INIT_25 of inst : label is "5B2C965B2D924967B3D9ECF67927965973222222AAAAAA216C249884910C24C2";
    attribute INIT_26 of inst : label is "75A5D61BC8B441A96CCC22329A144924932C9616CB6C92496DB249649244B6B6";
    attribute INIT_27 of inst : label is "813799CCA544DE8CA9813799B2A6F4654C099CD499D1952DC0AE1B16E65B5BA1";
    attribute INIT_28 of inst : label is "F3132CDE64DE674B37993799DACDE64DE674B33993399D2CDE6A6318D8DE8CA9";
    attribute INIT_29 of inst : label is "0C1492381CB34C8C6778CBB1A325A5F8F6B172EE8D2464B7382DCD66F3399166";
    attribute INIT_2A of inst : label is "46003C32E0A9100DB04618114A08DB7F66DECA938723188C81DD858D0A2060AC";
    attribute INIT_2B of inst : label is "324BAB57D54E5B81DE30ED7BE15C3A82084DCA73570A642068A0000005263B60";
    attribute INIT_2C of inst : label is "53650CA9B28654D849E848AFEC29F879B12093AA40F450940ADDCCCA6B84C113";
    attribute INIT_2D of inst : label is "5D6C154A4EAD3A285412B00000EBAFFA5A5902694E0D4338DA9C6D4E32E35A1B";
    attribute INIT_2E of inst : label is "B61740E9A092A2092083004A616B25A9A512548124B5C04812E94E04CCCC8889";
    attribute INIT_2F of inst : label is "3FFFFFFFFFFFFFFE4A892D224B4892D224B48B5480049925249115555555FD30";
    attribute INIT_30 of inst : label is "6ED0BE92FA437A4221789E2C3F9DA1CEB764FC66863AE4D7003F23B197B19241";
    attribute INIT_31 of inst : label is "4D2A0724BD76AED5DAB95D2574C999207E9004040403A488399645CFBD7AF7D4";
    attribute INIT_32 of inst : label is "7EFD3224EBE8732F27738844D899D26C118EFDDF8A3FCCE2724746F213BB8D68";
    attribute INIT_33 of inst : label is "35F9EFFFE28B31D66520A3F4607408220B2518500000CC946828807FA5052121";
    attribute INIT_34 of inst : label is "EFF72449F4516E49E38E4C491C72626D9C7372471C40038E005EA0D367BD57A8";
    attribute INIT_35 of inst : label is "0000000000000000002079E39E7E48F44D34734E49A68A6C492627D3EFF627DB";
    attribute INIT_36 of inst : label is "F557D5FD581F5557FDD7D7C00000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0BEFE2A1C0000012010AA000AA000054014001400000A000A005400A8007D57D";
    attribute INIT_38 of inst : label is "505415054150541505FE0170005F8017C00BFC50C54315822C11608B02A80200";
    attribute INIT_39 of inst : label is "45815608B02AF1400A005002802800140000280404500808A010114001400141";
    attribute INIT_3A of inst : label is "263618600000000000000100000200000000000000002F800BC005F0017000B0";
    attribute INIT_3B of inst : label is "AAAC36DB655AAE70F820019608040004010601010303030307035555055500BA";
    attribute INIT_3C of inst : label is "000000002D7FBFE3FDC7FB8FEAB8007003801C0055F7C00300AD6A015AD402B5";
    attribute INIT_3D of inst : label is "6011602AC0229055004510AA008A4154011502A8022C800F159001E2A1C00800";
    attribute INIT_3E of inst : label is "A192632C21E33B82447F40202FFC00022FFC000205002C055804580AB008B015";
    attribute INIT_3F of inst : label is "4A040488242000240820800005282081048D0000100102888A8220EA9ECD0000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "36363639449A19B4336866469FF1A000000000384E0190B0C8642BEDEDE23939";
    attribute INIT_01 of inst : label is "20682C004F02E13FB3208CB2488CB4688D2EE492EDA36DC71C71DC4A48E63636";
    attribute INIT_02 of inst : label is "DE466D9B75AEA1B706F6D6B9658B965B9672874E1888006AB8C0C4C8518142C8";
    attribute INIT_03 of inst : label is "6442492491C15CE89191A4259999CCCC6663332C5ECBDE4B6D8D9BB3243A6846";
    attribute INIT_04 of inst : label is "3204922421249212492484924921249248492124AAA088880000000088E5240C";
    attribute INIT_05 of inst : label is "9248239AEA800000656322926CB50D969256E308610C2592C92C92084CB7A089";
    attribute INIT_06 of inst : label is "0000000001004113292434A199341249249ECC4389330D9DE0CCE6038C9FB084";
    attribute INIT_07 of inst : label is "000000000000000000000BCDA24E368938DA24E36A93644B8C81093484705104";
    attribute INIT_08 of inst : label is "3C3138CC9249C04A22499C414555595000012894383838230000000000000000";
    attribute INIT_09 of inst : label is "0627188648C24924924E126918463A19220C3532CB06184430B24B6DB2643924";
    attribute INIT_0A of inst : label is "46CD32B6DCC8CE2E223C367610000000000083362450C924935551420D86421E";
    attribute INIT_0B of inst : label is "22C42316210D84162118B1086C209108448843610588462C421B0904270D8416";
    attribute INIT_0C of inst : label is "4219130CCC853C69642424101E48432253129D0132680C3086BA328CA3292161";
    attribute INIT_0D of inst : label is "0C896619991AF8DB21212080F242191302C910CA9618666429E34B21212080F2";
    attribute INIT_0E of inst : label is "4A094A72D4F7D3F47D3F4E53026418F36C9CCBA9CE21B0909041E48432385921";
    attribute INIT_0F of inst : label is "FFFF90B16BC111111119D9A492492436FFFFFF80000000000000008EA5241830";
    attribute INIT_10 of inst : label is "24482C9086469CA154C14C0314CC4C4188310524B363249A13250925D0CD0F0C";
    attribute INIT_11 of inst : label is "5A59210C8D3942648909059210C8D2C9086469CA3324482C9086469CA1B24933";
    attribute INIT_12 of inst : label is "B34D09D011872CCAA0002AA679A24816380F89C0C346185201C6489090792219";
    attribute INIT_13 of inst : label is "4AC61836D364691A4290A12E6249734A344E19A0D04606060606868686868E53";
    attribute INIT_14 of inst : label is "346468C8D191A32481A71666CC8D191A32346468C8D009D3AD334CD20EB8980A";
    attribute INIT_15 of inst : label is "9122448956CB1041188208C4104620820DB63A262D318D1908A643468D999A32";
    attribute INIT_16 of inst : label is "059188C4622C8C4623116458C065B1AC46691A2362334B6D82CCCC0101016598";
    attribute INIT_17 of inst : label is "060823018208C0609214A78DAD1465247410741074107412C881BC188B22606F";
    attribute INIT_18 of inst : label is "1EF39E3C25858E427B9007870961641820CA748DDECCDBBD99A454223018208C";
    attribute INIT_19 of inst : label is "6E4B864B21C30830D0B98608959112B286664691D63AC68799758EB0A15E6649";
    attribute INIT_1A of inst : label is "0B3C18222222233B64924924869613332490CC9085616B1B3B71217053665334";
    attribute INIT_1B of inst : label is "77B3142DDECCD0B77B334723A5294294294A34248024802484490178C0632121";
    attribute INIT_1C of inst : label is "316EF66685BBD99A39296618666492199646E32D021585AC6C6EF662DDECC50B";
    attribute INIT_1D of inst : label is "632B1B1BBD99B77B3346DDECC51C94B30C3332490CC9237196811AC65616377B";
    attribute INIT_1E of inst : label is "C8DC65A042B0B58D8DDECC53BD10A14CE4428E4A5986199924866491B849408D";
    attribute INIT_1F of inst : label is "7F32C9C628A665938C514CCB2718A299964E3145298B0C6B1B42C30CCC924332";
    attribute INIT_20 of inst : label is "9548529A4A614991634A61486C294C290D8D29206E0FB0AAAA5DFAAEABACE5CB";
    attribute INIT_21 of inst : label is "739490581CC9DB600114147B2872C249612C27243209612CB249A19030514CC2";
    attribute INIT_22 of inst : label is "2187334991B840E72864162A06490CD9CCCC903984CCCDCB249333272993CB60";
    attribute INIT_23 of inst : label is "CC10F41155511045440145C48545986A4D998EDBC911B710DC9231269892250E";
    attribute INIT_24 of inst : label is "2FA2460183E129631CCD189833006658C73A46203600CC2DEA1AE0260998191A";
    attribute INIT_25 of inst : label is "241209148A4120904824120904534514451111111111119CC4B6E496DE84B720";
    attribute INIT_26 of inst : label is "C1271CB66E5B4335D3389188614B24930C820909249249209249241248384848";
    attribute INIT_27 of inst : label is "3EC8E4CC92EF23520C7EC8E48979189061F6472E646241823F2C726D14727421";
    attribute INIT_28 of inst : label is "1CB8532193239034C864C8E40532193239014C864C8E40D323970E4E6723520C";
    attribute INIT_29 of inst : label is "39375B54A10CB37BDBEF77CFBC5A1A5768CF8EB171B3CB4954B131991C999B99";
    attribute INIT_2A of inst : label is "3D0486542038CC18610C0887042024C1C1949C58489AD6BB6ED87A422749C9B9";
    attribute INIT_2B of inst : label is "A96639C6AAF17440F3187BC923F42F5827641A041125139F62000001329006D0";
    attribute INIT_2C of inst : label is "A91AE7548D73AA48A4797939744C6058F3366C48A0796480A0C5141A0A241420";
    attribute INIT_2D of inst : label is "61B64163708DC22C16D8C00000016D1B6B6C930F2216788E644732A39919B5CE";
    attribute INIT_2E of inst : label is "B617206CB2D8BB2DB2CCBB7B2DEDB284388B1685B6F740E9130F221844444446";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFB64EDB5BB6D6EDB5BB6D6EE76FFFCC996B6C1DAAAAAAA05B0";
    attribute INIT_30 of inst : label is "1B6192624D892189C5647DF960C6D16D49BB831B45B5BBC8909CCB07C185BB80";
    attribute INIT_31 of inst : label is "160A11D640580B01602C0ED03A6446CB124FF62626233B5C3DC5B3650B162F67";
    attribute INIT_32 of inst : label is "0190CDBB39310B6B99C8F0374C7E9DA66B62464A7714A60B9D59902A4D491633";
    attribute INIT_33 of inst : label is "8007FDFFE8A0C7799F8228019FDFE088B09AE7A80000306B862888001AFAA121";
    attribute INIT_34 of inst : label is "EFF776EDF7DF6EEDF7DF6EEDBEFB776DBEFB776FBEFFFFDFFFFE82009FF7FFA0";
    attribute INIT_35 of inst : label is "000000000000000000217DF7DF7F6DF6EDB6FB6EEDB6FB6EEDB777DBEFF777DB";
    attribute INIT_36 of inst : label is "00A880AAA00AA282A802A8000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "A010181E3FFFFC01FEF01FFF01FFFF43F43FF03FF0001FF81FF03FE07FE80282";
    attribute INIT_38 of inst : label is "00000010240902400001F40FFD007F403FA0010F243C907C83E41F20FC87FDFF";
    attribute INIT_39 of inst : label is "907E41F20FC8003F81FC0FE07E07FF03FFFE07FBF80FF7F01FEFE03FF03FF000";
    attribute INIT_3A of inst : label is "4140C308000000000000010000020000000000000000007FA03FD00FF40FFA0F";
    attribute INIT_3B of inst : label is "5AAC36DB65551580FE400195000501050107000200000000050100000000008E";
    attribute INIT_3C of inst : label is "000000000CCD655D54BAA9754ABFFFFFFFFFFFFF557D5555555AD6AAB5AD556B";
    attribute INIT_3D of inst : label is "1FE41FC83FC86F90FF90EF21FF21BE43FE42FC87FC837FF0C06FFE181E3FF7FC";
    attribute INIT_3E of inst : label is "5A24B5029A914C508855DFD00003FFFA0003FFFA00FE03F907F907F20FF20FE4";
    attribute INIT_3F of inst : label is "817A7AF5C787E3D3E7ACF8FE74C7ACF9FAF5CBE9C7FD220280AA80E00A080000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "12121211C0010A8215042AC05FE2A000000000380E055008812221C7C6913829";
    attribute INIT_01 of inst : label is "226868002E02823FB2900D92D90CBC018404400044D124820820884508A21212";
    attribute INIT_02 of inst : label is "5D2680C0402805A6068310A1041A105A10420C6E1A802AE03084C825053E1C28";
    attribute INIT_03 of inst : label is "E0024924918558A1020280051111888C44622370CA594A8925050AA002212004";
    attribute INIT_04 of inst : label is "0404926C6165963059658C165963059658C16124800088888888888800440090";
    attribute INIT_05 of inst : label is "925A0310300490494502175624440488B2DA2204408815B6592496102C922080";
    attribute INIT_06 of inst : label is "00000000011401162000908090009249249A45061B041034804082021C9E1004";
    attribute INIT_07 of inst : label is "000000000000000000000B04AA2512A8944AA251288920314480F69479409140";
    attribute INIT_08 of inst : label is "286200449269800860001C85411114000000385C6C6C6C600000000000000000";
    attribute INIT_09 of inst : label is "0C40080248824924924C000030043809641045124208208060B64B24B2603120";
    attribute INIT_0A of inst : label is "C28EB2924888DC28003812D2815555555551821212C04924935551060485280C";
    attribute INIT_0B of inst : label is "22C4631623068A162318B1183450B118C588C1A28488C224460D140C66868A16";
    attribute INIT_0C of inst : label is "00111208880F68695200000034000222EA8B500829004020C29D1344D1342141";
    attribute INIT_0D of inst : label is "08895411101ED0DA90000001A00011168780208AB53044407B415A90000000A0";
    attribute INIT_0E of inst : label is "0C018E235ABAE1B8EE3B8C4AA55208D92A845AB54A30A8000001400022347000";
    attribute INIT_0F of inst : label is "3FFFB1A38FA1111111114A1249249210FFFFFF80000000000000009A00381016";
    attribute INIT_10 of inst : label is "928038000446570154A40A0294AA2A21442886AD97416D9D33269B6CE9EC2D05";
    attribute INIT_11 of inst : label is "597000088CAE0652500007000088CB8000446570329280380004465701EADB6A";
    attribute INIT_12 of inst : label is "D10310043145844000002AA57495201210079000842228280145250000500411";
    attribute INIT_13 of inst : label is "2FA20242492A749D2749D03226DB2BA8100B4880C02606060606868686868D4A";
    attribute INIT_14 of inst : label is "1830306060C0C18080C0132346060C0C18183030606001602EB7ADE90B54540C";
    attribute INIT_15 of inst : label is "020408116249E0A28F05147828A3C145049308422611062110AC43A3468C8C18";
    attribute INIT_16 of inst : label is "051188C462288C4623114448604518A844311A23422189248244440101014511";
    attribute INIT_17 of inst : label is "2C14760B051D82C1421AD74584B81690D828D828D828D82848819C188A226067";
    attribute INIT_18 of inst : label is "0A5294304505040A29000D0C11414219040402010800421000D4726760B051D8";
    attribute INIT_19 of inst : label is "442B42C91081E05158950419B53336A604440200D41A8207913506A0811E4440";
    attribute INIT_1A of inst : label is "82121022222222290A49249242553222000088908D432A0C3FF0132A51405234";
    attribute INIT_1B of inst : label is "42001A210800E8842003A283D6A1075075A9182000200020144001F440421010";
    attribute INIT_1C of inst : label is "010840074421001D14355410444000111244412682350CA83008400210800688";
    attribute INIT_1D of inst : label is "412A1C021001842003A610800E8A1AAA08222000088B222093410A8254180420";
    attribute INIT_1E of inst : label is "C88865D042A0B50E010800CA1089D32A5227450D55041110000445911049A085";
    attribute INIT_1F of inst : label is "7E02810425D40502084BA80A041097501408212EACC184290A01820888000222";
    attribute INIT_20 of inst : label is "4DA4699D0D518543538D5184EA71AA309D4635604607802AAA1172A8AAC4CC99";
    attribute INIT_21 of inst : label is "51104850088949211000146A20228249412822006959412896C98148210008A3";
    attribute INIT_22 of inst : label is "69052109109400E62052142A2C402C588888821B10888C8964C2222221128804";
    attribute INIT_23 of inst : label is "C800D04441551450504405D2844E504924988A83E1029202CC80512008110404";
    attribute INIT_24 of inst : label is "2A826001026121D6B181189821014475AC60462012028829B856C00701903980";
    attribute INIT_25 of inst : label is "00000010080000000000000000C00820861111111111111844924492488492A0";
    attribute INIT_26 of inst : label is "01205090694B4015036C03105122000108002100000000000000000000A80000";
    attribute INIT_27 of inst : label is "2A8040B300460100086A80408030080043540204402001051504420104020420";
    attribute INIT_28 of inst : label is "08106A010201003A804080400EA010201003A8040804006A01020B0C46010008";
    attribute INIT_29 of inst : label is "919349544384A10B63EC47CF105C0854608104816093C9815441211008166110";
    attribute INIT_2A of inst : label is "348452404038CC08A00418470610660110211C50408A52AD0A100A42014C8C99";
    attribute INIT_2B of inst : label is "A14638C600614040C108638003E0064007443A0C1200035D000000002B422848";
    attribute INIT_2C of inst : label is "A4285552142AAAC884593913B444441873344558C061448020C33A3A06623000";
    attribute INIT_2D of inst : label is "24B6C1213488D2041248900000542C19212C91272507354D5526AA135514D0AA";
    attribute INIT_2E of inst : label is "1203002416489164966CB3290CA59604908912809253C0E80127250C44444447";
    attribute INIT_2F of inst : label is "BFFFFFFFFFFFFFFB2C64909924264909924264227FFCA952B2A0C80000000490";
    attribute INIT_30 of inst : label is "9121902240812081414C38BC40431E285E49810C78A149C180184A0502852480";
    attribute INIT_31 of inst : label is "120A089520640C819032040830400A4A30000404040121283146000001020526";
    attribute INIT_32 of inst : label is "01A045A139001A6B09D0D0144C2890A62B2202405714445A0940802A20011212";
    attribute INIT_33 of inst : label is "8A1A1201EA8C0CAEEAAAA20A212A002804600800000103803800000060002121";
    attribute INIT_34 of inst : label is "EFF776EDF7DF6EEDF7DF6EEDBEFB776DBEFB776FBEFFFFDFFFDEA22C684AAFA8";
    attribute INIT_35 of inst : label is "000000000000000000017DF7DF7F6DF6EDB6FB6EEDB6FB6EEDB777DBEFF777DB";
    attribute INIT_36 of inst : label is "AA0000AAA808880A20A800000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "340003400000014400034000340000680280068004004003400A80150018888A";
    attribute INIT_38 of inst : label is "AF2BCAE298A6298ACA00068001A00068003400A002800A005002801400500000";
    attribute INIT_39 of inst : label is "0A002801400502801400A005005000280000500000A0000140000280028002BC";
    attribute INIT_3A of inst : label is "60204000000000000000000000000000000000000000500034001A0006800340";
    attribute INIT_3B of inst : label is "02AFC924955545FF0080009C000C000400040008080808080C0055555555558D";
    attribute INIT_3C of inst : label is "000000001A000000020004000AB0000000000000556000000000000000000000";
    attribute INIT_3D of inst : label is "80068005000D000A001A0014003400280068005000D000000A00000140000001";
    attribute INIT_3E of inst : label is "5A2495068A914ED08800400450000000500000000A005000A001A00140034002";
    attribute INIT_3F of inst : label is "D30E0E1D54A02A54E8AE8D0A9560AE0D0E14585850052228A80080680A0A8000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
