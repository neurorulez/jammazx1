library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity berzerk_program2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of berzerk_program2 is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"F3",X"AF",X"D3",X"4D",X"ED",X"47",X"DB",X"61",X"CB",X"47",X"C2",X"00",X"02",X"CB",X"57",
		X"C2",X"A7",X"06",X"CB",X"5F",X"C2",X"5B",X"06",X"DD",X"21",X"73",X"00",X"18",X"0F",X"04",X"00",
		X"F8",X"C8",X"00",X"01",X"00",X"00",X"0D",X"20",X"FD",X"10",X"FB",X"DB",X"66",X"3E",X"01",X"01",
		X"41",X"01",X"11",X"47",X"82",X"ED",X"41",X"0D",X"ED",X"51",X"0C",X"0C",X"ED",X"41",X"0C",X"ED",
		X"41",X"0C",X"0C",X"0C",X"ED",X"59",X"0E",X"51",X"3D",X"28",X"EA",X"01",X"00",X"00",X"0D",X"20",
		X"FD",X"10",X"FB",X"DB",X"67",X"AF",X"D3",X"40",X"D3",X"50",X"DD",X"E9",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D3",X"4D",X"F5",X"3A",X"04",X"40",X"B7",X"C2",X"BC",X"04",
		X"C3",X"04",X"1A",X"1E",X"04",X"DD",X"21",X"00",X"10",X"01",X"00",X"10",X"26",X"00",X"2E",X"FF",
		X"DD",X"7E",X"00",X"57",X"A5",X"6F",X"7A",X"84",X"67",X"DD",X"23",X"0D",X"20",X"F2",X"10",X"F0",
		X"3A",X"1E",X"00",X"FE",X"FF",X"28",X"2D",X"7B",X"FE",X"02",X"C2",X"A1",X"00",X"DD",X"21",X"00",
		X"C0",X"B7",X"F2",X"A9",X"00",X"7D",X"3C",X"28",X"04",X"7B",X"BC",X"20",X"17",X"7B",X"CB",X"07",
		X"DA",X"CC",X"00",X"1D",X"20",X"C3",X"ED",X"57",X"A7",X"C2",X"3D",X"01",X"DD",X"21",X"00",X"00",
		X"1E",X"80",X"18",X"B5",X"ED",X"57",X"A7",X"C2",X"02",X"01",X"18",X"FE",X"DD",X"21",X"D3",X"00",
		X"C3",X"23",X"00",X"C3",X"3D",X"01",X"EA",X"3E",X"01",X"ED",X"47",X"C3",X"73",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"D5",X"01",X"C0",X"08",X"21",X"00",X"00",X"16",X"08",X"7E",X"09",X"AF",X"ED",X"4F",X"32",
		X"00",X"10",X"15",X"20",X"F5",X"0E",X"7F",X"16",X"20",X"7B",X"E6",X"20",X"47",X"ED",X"78",X"CB",
		X"0B",X"0D",X"15",X"20",X"F4",X"3E",X"80",X"01",X"57",X"80",X"ED",X"79",X"05",X"0D",X"CB",X"0F",
		X"30",X"F8",X"0E",X"47",X"ED",X"79",X"0D",X"CB",X"0F",X"30",X"F9",X"18",X"C5",X"2A",X"1F",X"00",
		X"ED",X"4B",X"21",X"00",X"36",X"55",X"2B",X"ED",X"A1",X"E2",X"4F",X"01",X"23",X"18",X"F5",X"16",
		X"AA",X"31",X"FF",X"FF",X"ED",X"4B",X"21",X"00",X"7A",X"2F",X"AE",X"20",X"16",X"72",X"2B",X"ED",
		X"A1",X"EA",X"70",X"01",X"7A",X"FE",X"55",X"28",X"25",X"31",X"01",X"00",X"16",X"55",X"18",X"E4",
		X"39",X"18",X"E5",X"57",X"ED",X"57",X"CB",X"0F",X"38",X"01",X"76",X"1E",X"12",X"7A",X"E6",X"0F",
		X"CA",X"02",X"01",X"1D",X"7A",X"E6",X"F0",X"CA",X"02",X"01",X"1D",X"C3",X"02",X"01",X"ED",X"57",
		X"CB",X"0F",X"1E",X"20",X"D2",X"B1",X"02",X"C3",X"02",X"01",X"21",X"C1",X"03",X"11",X"01",X"00",
		X"78",X"A2",X"C2",X"C1",X"01",X"79",X"A3",X"C3",X"C1",X"01",X"EB",X"29",X"EB",X"D2",X"A0",X"01",
		X"11",X"00",X"40",X"1D",X"FD",X"7E",X"00",X"C2",X"B3",X"01",X"15",X"C2",X"B3",X"01",X"C3",X"B8",
		X"02",X"08",X"7E",X"23",X"D9",X"6F",X"D9",X"7E",X"23",X"D9",X"67",X"11",X"1F",X"00",X"06",X"03",
		X"08",X"B7",X"28",X"07",X"36",X"FC",X"23",X"36",X"3F",X"18",X"05",X"36",X"84",X"23",X"36",X"21",
		X"19",X"10",X"EE",X"06",X"24",X"B7",X"28",X"07",X"36",X"FF",X"23",X"36",X"FF",X"18",X"05",X"36",
		X"80",X"23",X"36",X"01",X"19",X"10",X"EE",X"D9",X"C3",X"AA",X"01",X"FF",X"A8",X"04",X"B6",X"04",
		X"01",X"48",X"10",X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"0C",X"ED",X"78",X"0C",
		X"ED",X"78",X"0C",X"ED",X"78",X"0C",X"3E",X"01",X"ED",X"79",X"01",X"48",X"00",X"ED",X"78",X"0C",
		X"ED",X"78",X"0C",X"ED",X"78",X"21",X"00",X"50",X"11",X"00",X"70",X"06",X"10",X"78",X"3D",X"D3",
		X"4B",X"3E",X"80",X"77",X"12",X"4E",X"CB",X"0F",X"30",X"F9",X"AF",X"DB",X"4E",X"3E",X"08",X"32",
		X"00",X"50",X"32",X"00",X"70",X"AF",X"DB",X"4E",X"23",X"13",X"10",X"E1",X"06",X"0D",X"11",X"00",
		X"A0",X"21",X"FE",X"5F",X"3E",X"80",X"25",X"77",X"4E",X"24",X"37",X"CB",X"15",X"CB",X"14",X"19",
		X"CB",X"0F",X"10",X"F2",X"21",X"11",X"11",X"11",X"11",X"11",X"31",X"00",X"88",X"0E",X"10",X"06",
		X"10",X"E5",X"E5",X"E5",X"E5",X"10",X"FA",X"19",X"F1",X"3B",X"3B",X"0D",X"20",X"F1",X"DB",X"4C",
		X"AF",X"DB",X"4E",X"AF",X"DB",X"61",X"CB",X"4F",X"28",X"FE",X"21",X"00",X"50",X"11",X"00",X"70",
		X"3E",X"F0",X"ED",X"47",X"01",X"4B",X"00",X"ED",X"57",X"ED",X"79",X"0E",X"00",X"79",X"70",X"12",
		X"48",X"2F",X"46",X"47",X"B1",X"20",X"F6",X"ED",X"57",X"D6",X"10",X"ED",X"47",X"20",X"E5",X"18",
		X"FE",X"DD",X"21",X"B8",X"02",X"C3",X"23",X"00",X"21",X"FF",X"5F",X"11",X"00",X"00",X"DD",X"21",
		X"C5",X"02",X"C3",X"95",X"03",X"01",X"00",X"00",X"21",X"00",X"40",X"DD",X"21",X"D2",X"02",X"C3",
		X"76",X"03",X"21",X"00",X"40",X"11",X"55",X"00",X"DD",X"21",X"DF",X"02",X"C3",X"95",X"03",X"21",
		X"FF",X"5F",X"11",X"AA",X"55",X"DD",X"21",X"EC",X"02",X"C3",X"95",X"03",X"21",X"00",X"40",X"11",
		X"FF",X"AA",X"DD",X"21",X"F9",X"02",X"C3",X"95",X"03",X"21",X"FF",X"5F",X"11",X"00",X"FF",X"DD",
		X"21",X"06",X"03",X"C3",X"95",X"03",X"79",X"B0",X"C2",X"9A",X"01",X"DD",X"21",X"12",X"03",X"C3",
		X"23",X"00",X"21",X"FF",X"87",X"11",X"00",X"00",X"DD",X"21",X"1F",X"03",X"C3",X"95",X"03",X"01",
		X"00",X"00",X"21",X"00",X"80",X"DD",X"21",X"2C",X"03",X"C3",X"76",X"03",X"21",X"00",X"84",X"DD",
		X"21",X"36",X"03",X"C3",X"76",X"03",X"21",X"00",X"80",X"11",X"55",X"00",X"DD",X"21",X"43",X"03",
		X"C3",X"8F",X"03",X"21",X"FF",X"87",X"11",X"AA",X"55",X"DD",X"21",X"50",X"03",X"C3",X"8F",X"03",
		X"21",X"00",X"80",X"11",X"FF",X"AA",X"DD",X"21",X"5D",X"03",X"C3",X"8F",X"03",X"21",X"FF",X"87",
		X"11",X"00",X"FF",X"DD",X"21",X"6A",X"03",X"C3",X"8F",X"03",X"79",X"B0",X"C2",X"6C",X"03",X"DD",
		X"21",X"E1",X"03",X"C3",X"23",X"00",X"16",X"00",X"72",X"7E",X"AA",X"B0",X"47",X"23",X"72",X"7E",
		X"AA",X"B1",X"4F",X"2B",X"15",X"C2",X"78",X"03",X"36",X"00",X"23",X"36",X"00",X"DD",X"E9",X"D9",
		X"01",X"00",X"08",X"18",X"04",X"D9",X"01",X"00",X"20",X"D9",X"7E",X"AA",X"B0",X"47",X"73",X"7E",
		X"AB",X"B0",X"47",X"CB",X"43",X"C2",X"AA",X"03",X"2B",X"3E",X"23",X"78",X"41",X"4F",X"D9",X"0D",
		X"C2",X"B7",X"03",X"05",X"CA",X"BB",X"03",X"D9",X"C3",X"9A",X"03",X"D9",X"78",X"41",X"4F",X"DD",
		X"E9",X"8D",X"50",X"4D",X"4A",X"0D",X"44",X"CD",X"56",X"15",X"44",X"55",X"4A",X"95",X"50",X"D5",
		X"56",X"89",X"50",X"49",X"4A",X"09",X"44",X"C9",X"56",X"11",X"44",X"51",X"4A",X"91",X"50",X"D1",
		X"56",X"21",X"00",X"60",X"16",X"01",X"42",X"AF",X"4F",X"5F",X"ED",X"47",X"ED",X"57",X"D3",X"4B",
		X"36",X"FF",X"72",X"36",X"00",X"7E",X"BB",X"20",X"FE",X"ED",X"57",X"3C",X"ED",X"47",X"FE",X"10",
		X"20",X"0B",X"CB",X"12",X"30",X"E0",X"DD",X"21",X"26",X"04",X"C3",X"23",X"00",X"79",X"CB",X"1F",
		X"CB",X"18",X"CB",X"19",X"59",X"ED",X"57",X"FE",X"08",X"38",X"D1",X"3E",X"08",X"CB",X"08",X"CB",
		X"13",X"3D",X"20",X"F9",X"18",X"C6",X"1E",X"00",X"DD",X"21",X"69",X"04",X"21",X"00",X"60",X"01",
		X"01",X"01",X"7B",X"D3",X"4B",X"78",X"32",X"00",X"40",X"71",X"79",X"DD",X"E9",X"AE",X"20",X"FE",
		X"77",X"78",X"A1",X"28",X"02",X"3E",X"80",X"57",X"DB",X"4E",X"AA",X"17",X"38",X"FE",X"CB",X"00",
		X"30",X"E0",X"CB",X"01",X"30",X"DC",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"3E",X"10",X"83",X"5F",
		X"30",X"D0",X"DD",X"21",X"99",X"04",X"C3",X"23",X"00",X"00",X"18",X"D1",X"B0",X"18",X"CE",X"2F",
		X"18",X"18",X"AF",X"18",X"21",X"A0",X"18",X"C5",X"78",X"18",X"C2",X"A8",X"18",X"18",X"2F",X"18",
		X"EB",X"2F",X"18",X"0F",X"A8",X"18",X"B6",X"78",X"18",X"0C",X"A0",X"18",X"09",X"AF",X"18",X"AD",
		X"2F",X"18",X"E2",X"B0",X"18",X"00",X"2F",X"18",X"A4",X"ED",X"5E",X"3E",X"01",X"ED",X"47",X"DD",
		X"21",X"D0",X"04",X"3E",X"FF",X"D3",X"4F",X"47",X"31",X"FF",X"43",X"DB",X"4E",X"1F",X"CB",X"10",
		X"78",X"EE",X"55",X"28",X"03",X"FB",X"18",X"FE",X"D3",X"4F",X"06",X"FF",X"31",X"FF",X"43",X"DB",
		X"4D",X"DB",X"4E",X"1F",X"CB",X"10",X"78",X"EE",X"20",X"CA",X"23",X"00",X"DB",X"4C",X"18",X"FE",
		X"F3",X"31",X"80",X"F8",X"21",X"80",X"F8",X"01",X"48",X"00",X"CD",X"40",X"06",X"21",X"00",X"40",
		X"01",X"00",X"04",X"CD",X"40",X"06",X"CD",X"66",X"00",X"CD",X"A6",X"08",X"21",X"6E",X"40",X"11",
		X"1B",X"F9",X"06",X"3C",X"CD",X"44",X"08",X"DB",X"49",X"2F",X"21",X"59",X"40",X"77",X"23",X"77",
		X"31",X"80",X"F8",X"AF",X"32",X"56",X"40",X"CD",X"2F",X"05",X"CD",X"A9",X"30",X"CD",X"A6",X"08",
		X"CD",X"86",X"0C",X"AF",X"32",X"56",X"40",X"CD",X"99",X"10",X"CD",X"84",X"11",X"CD",X"86",X"0C",
		X"CD",X"C2",X"11",X"CD",X"86",X"0C",X"C3",X"EE",X"0F",X"CA",X"00",X"05",X"C3",X"47",X"05",X"F3",
		X"AF",X"32",X"07",X"40",X"3D",X"32",X"5E",X"40",X"CD",X"C2",X"16",X"CD",X"77",X"20",X"3E",X"55",
		X"32",X"C7",X"F8",X"CD",X"97",X"13",X"C9",X"31",X"80",X"F8",X"21",X"56",X"40",X"CB",X"FE",X"CD",
		X"2F",X"05",X"3A",X"56",X"40",X"6F",X"CD",X"D1",X"0C",X"CB",X"4D",X"3E",X"01",X"28",X"05",X"CD",
		X"D1",X"0C",X"3E",X"02",X"32",X"21",X"40",X"FE",X"02",X"28",X"07",X"0E",X"03",X"CD",X"0F",X"08",
		X"18",X"0A",X"0E",X"04",X"CD",X"0F",X"08",X"0E",X"05",X"CD",X"0F",X"08",X"0E",X"05",X"CD",X"0F",
		X"08",X"CD",X"11",X"06",X"01",X"0C",X"00",X"11",X"07",X"40",X"21",X"50",X"06",X"ED",X"B0",X"2A",
		X"64",X"40",X"EB",X"2A",X"18",X"F9",X"19",X"22",X"64",X"40",X"22",X"08",X"40",X"DB",X"60",X"E6",
		X"0F",X"32",X"11",X"40",X"AF",X"32",X"5E",X"40",X"32",X"9D",X"F8",X"32",X"12",X"40",X"3C",X"32",
		X"9C",X"F8",X"21",X"07",X"40",X"11",X"13",X"40",X"01",X"0C",X"00",X"ED",X"B0",X"3E",X"02",X"77",
		X"3A",X"21",X"40",X"FE",X"02",X"28",X"04",X"AF",X"32",X"18",X"40",X"FB",X"2A",X"53",X"06",X"22",
		X"0A",X"40",X"3A",X"07",X"40",X"CD",X"A5",X"1E",X"CD",X"39",X"10",X"3E",X"5A",X"CD",X"0E",X"18",
		X"CD",X"77",X"20",X"2A",X"64",X"40",X"22",X"08",X"40",X"21",X"0C",X"40",X"35",X"CD",X"29",X"06",
		X"20",X"D9",X"CD",X"29",X"06",X"20",X"D4",X"3E",X"FF",X"32",X"5E",X"40",X"CD",X"B6",X"1A",X"CD",
		X"D5",X"27",X"CD",X"29",X"06",X"CD",X"D5",X"27",X"31",X"80",X"F8",X"CD",X"2F",X"05",X"C3",X"13",
		X"05",X"21",X"00",X"00",X"22",X"68",X"40",X"22",X"6A",X"40",X"22",X"6C",X"40",X"22",X"5B",X"40",
		X"21",X"A7",X"30",X"22",X"9A",X"F8",X"C3",X"B6",X"1A",X"E5",X"21",X"07",X"40",X"11",X"13",X"40",
		X"06",X"0C",X"1A",X"4E",X"EB",X"12",X"71",X"EB",X"23",X"13",X"10",X"F6",X"E1",X"7E",X"B7",X"C9",
		X"79",X"B7",X"48",X"47",X"28",X"01",X"0C",X"AF",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"01",X"00",X"00",X"1E",X"74",X"03",X"06",X"00",X"5A",X"00",X"00",X"21",X"00",X"44",X"54",X"5D",
		X"36",X"01",X"23",X"73",X"23",X"01",X"FD",X"1B",X"EB",X"ED",X"B0",X"21",X"00",X"45",X"54",X"5D",
		X"06",X"20",X"36",X"FF",X"23",X"10",X"FB",X"01",X"80",X"02",X"09",X"EB",X"01",X"7F",X"18",X"ED",
		X"B0",X"CD",X"B2",X"0D",X"CD",X"70",X"09",X"21",X"00",X"44",X"11",X"01",X"44",X"01",X"FF",X"1B",
		X"36",X"FF",X"ED",X"B0",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"07",X"36",X"11",X"ED",
		X"B0",X"CD",X"70",X"09",X"C3",X"5B",X"06",X"F3",X"DB",X"4E",X"AF",X"D3",X"4F",X"D3",X"4D",X"31",
		X"80",X"F8",X"CD",X"1A",X"11",X"CD",X"B2",X"0D",X"21",X"38",X"07",X"11",X"20",X"00",X"CD",X"10",
		X"07",X"11",X"20",X"80",X"CD",X"10",X"07",X"11",X"08",X"10",X"CD",X"10",X"07",X"11",X"10",X"D0",
		X"CD",X"10",X"07",X"21",X"A0",X"47",X"CD",X"11",X"11",X"21",X"A0",X"55",X"CD",X"11",X"11",X"11",
		X"08",X"20",X"DB",X"61",X"CD",X"16",X"07",X"DB",X"60",X"CD",X"16",X"07",X"DB",X"62",X"CD",X"16",
		X"07",X"DB",X"63",X"CD",X"16",X"07",X"DB",X"64",X"CD",X"16",X"07",X"11",X"08",X"90",X"DB",X"48",
		X"CD",X"15",X"07",X"DB",X"49",X"CD",X"15",X"07",X"DB",X"4A",X"CD",X"15",X"07",X"C3",X"DF",X"06",
		X"06",X"00",X"C3",X"85",X"08",X"2F",X"0E",X"08",X"1F",X"21",X"80",X"07",X"38",X"03",X"21",X"82",
		X"07",X"F5",X"D5",X"C5",X"CD",X"10",X"07",X"C1",X"D1",X"F1",X"21",X"20",X"00",X"19",X"EB",X"0D",
		X"20",X"E6",X"21",X"00",X"0F",X"19",X"EB",X"C9",X"5A",X"50",X"55",X"20",X"44",X"49",X"50",X"20",
		X"53",X"57",X"49",X"54",X"43",X"48",X"45",X"53",X"00",X"56",X"46",X"42",X"20",X"53",X"57",X"49",
		X"54",X"43",X"48",X"45",X"53",X"00",X"31",X"20",X"20",X"20",X"32",X"20",X"20",X"20",X"33",X"20",
		X"20",X"20",X"34",X"20",X"20",X"20",X"35",X"20",X"20",X"20",X"36",X"20",X"20",X"20",X"37",X"20",
		X"20",X"20",X"38",X"00",X"30",X"3D",X"4F",X"46",X"46",X"20",X"20",X"31",X"3D",X"4F",X"4E",X"00",
		X"31",X"00",X"30",X"00",X"AF",X"D3",X"4F",X"DB",X"4E",X"31",X"80",X"F8",X"CD",X"81",X"09",X"20",
		X"FB",X"CD",X"1A",X"11",X"CD",X"F0",X"0D",X"F3",X"21",X"EA",X"08",X"0E",X"FF",X"0C",X"79",X"FE",
		X"0A",X"CA",X"D4",X"07",X"CD",X"6C",X"08",X"C5",X"06",X"00",X"11",X"00",X"CF",X"CD",X"85",X"08",
		X"C1",X"CD",X"6C",X"08",X"CD",X"DF",X"07",X"CD",X"81",X"09",X"28",X"0E",X"CD",X"99",X"08",X"CD",
		X"81",X"09",X"20",X"FB",X"CD",X"99",X"08",X"C3",X"9D",X"07",X"CD",X"7B",X"09",X"28",X"E8",X"CD",
		X"FB",X"07",X"18",X"E0",X"CD",X"81",X"09",X"20",X"FB",X"CD",X"99",X"08",X"C3",X"D0",X"04",X"C5",
		X"E5",X"CD",X"34",X"08",X"EB",X"21",X"00",X"00",X"E5",X"E5",X"E5",X"39",X"CD",X"44",X"08",X"11",
		X"CF",X"00",X"CD",X"5F",X"08",X"E1",X"E1",X"E1",X"E1",X"C1",X"C9",X"C5",X"E5",X"79",X"FE",X"09",
		X"20",X"01",X"0C",X"CD",X"34",X"08",X"2B",X"04",X"36",X"00",X"23",X"10",X"FB",X"18",X"E9",X"F5",
		X"C5",X"D5",X"E5",X"CD",X"34",X"08",X"16",X"00",X"58",X"1D",X"19",X"0E",X"10",X"1E",X"00",X"7E",
		X"E6",X"F0",X"81",X"27",X"77",X"38",X"02",X"0E",X"00",X"2B",X"83",X"5F",X"10",X"F1",X"73",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"21",X"C9",X"08",X"59",X"16",X"00",X"19",X"19",X"19",X"5E",X"23",X"56",
		X"23",X"46",X"EB",X"C9",X"E5",X"D5",X"C5",X"CB",X"28",X"1A",X"13",X"E6",X"F0",X"4F",X"1A",X"13",
		X"07",X"07",X"07",X"07",X"E6",X"0F",X"B1",X"77",X"23",X"10",X"EE",X"C1",X"D1",X"E1",X"C9",X"C5",
		X"D5",X"E5",X"53",X"1E",X"00",X"CD",X"53",X"2E",X"E1",X"D1",X"C1",X"C9",X"C5",X"D5",X"E5",X"01",
		X"C0",X"19",X"11",X"00",X"44",X"21",X"00",X"46",X"ED",X"B0",X"EB",X"01",X"00",X"02",X"CD",X"40",
		X"06",X"E1",X"D1",X"C1",X"C9",X"EB",X"CD",X"B6",X"2D",X"EB",X"4E",X"CD",X"EE",X"2D",X"13",X"23",
		X"47",X"7E",X"B7",X"78",X"C2",X"8A",X"08",X"23",X"C9",X"06",X"00",X"DD",X"E3",X"DD",X"E3",X"DD",
		X"E3",X"DD",X"E3",X"10",X"F6",X"C9",X"0E",X"00",X"CD",X"34",X"08",X"2B",X"7E",X"E6",X"F0",X"08",
		X"16",X"00",X"23",X"7E",X"E6",X"F0",X"82",X"57",X"10",X"F8",X"08",X"BA",X"C4",X"FB",X"07",X"0C",
		X"79",X"FE",X"09",X"38",X"E3",X"C0",X"0C",X"18",X"DF",X"CA",X"F8",X"02",X"CD",X"F8",X"08",X"D6",
		X"F8",X"08",X"DF",X"F8",X"06",X"E6",X"F8",X"06",X"ED",X"F8",X"06",X"F4",X"F8",X"0C",X"01",X"F9",
		X"0C",X"0E",X"F9",X"0C",X"1B",X"F9",X"06",X"1B",X"F9",X"3C",X"43",X"72",X"65",X"64",X"69",X"74",
		X"73",X"00",X"43",X"68",X"75",X"74",X"65",X"20",X"31",X"00",X"43",X"68",X"75",X"74",X"65",X"20",
		X"32",X"00",X"31",X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"47",X"61",X"6D",X"65",X"73",
		X"00",X"32",X"20",X"50",X"6C",X"61",X"79",X"65",X"72",X"20",X"47",X"61",X"6D",X"65",X"73",X"00",
		X"54",X"6F",X"74",X"61",X"6C",X"20",X"50",X"6C",X"61",X"79",X"73",X"00",X"54",X"6F",X"74",X"61",
		X"6C",X"20",X"53",X"63",X"6F",X"72",X"65",X"00",X"54",X"6F",X"74",X"61",X"6C",X"20",X"53",X"65",
		X"63",X"6F",X"6E",X"64",X"73",X"20",X"6F",X"66",X"20",X"50",X"6C",X"61",X"79",X"00",X"54",X"6F",
		X"74",X"61",X"6C",X"20",X"53",X"65",X"63",X"6F",X"6E",X"64",X"73",X"20",X"47",X"61",X"6D",X"65",
		X"20",X"4F",X"6E",X"00",X"48",X"69",X"67",X"68",X"20",X"53",X"63",X"6F",X"72",X"65",X"73",X"00",
		X"CD",X"7B",X"09",X"20",X"FB",X"CD",X"7B",X"09",X"28",X"FB",X"C9",X"CD",X"8B",X"09",X"CB",X"67",
		X"C9",X"DB",X"65",X"CB",X"7F",X"C9",X"DB",X"65",X"CB",X"47",X"C9",X"3A",X"22",X"40",X"B7",X"DB",
		X"48",X"28",X"02",X"DB",X"4A",X"2F",X"E6",X"1F",X"C9",X"D9",X"C5",X"3A",X"BA",X"F8",X"47",X"E6",
		X"F0",X"4F",X"78",X"E6",X"0F",X"47",X"D9",X"06",X"02",X"CD",X"BA",X"09",X"06",X"02",X"CD",X"BA",
		X"09",X"06",X"07",X"CD",X"BA",X"09",X"D9",X"C1",X"D9",X"C9",X"21",X"1B",X"80",X"C5",X"E5",X"CD",
		X"CB",X"09",X"E1",X"C1",X"11",X"0F",X"00",X"19",X"10",X"F3",X"C9",X"7E",X"F5",X"E6",X"0F",X"20",
		X"02",X"F1",X"C9",X"01",X"01",X"00",X"09",X"87",X"4F",X"09",X"5E",X"23",X"56",X"EB",X"7D",X"B4",
		X"28",X"05",X"CD",X"19",X"0C",X"36",X"80",X"F1",X"E6",X"F0",X"20",X"08",X"21",X"FF",X"FF",X"19",
		X"ED",X"42",X"35",X"C9",X"62",X"6B",X"2B",X"2B",X"ED",X"B8",X"23",X"0F",X"0F",X"0F",X"4F",X"EB",
		X"21",X"0E",X"0A",X"09",X"7E",X"23",X"66",X"6F",X"EB",X"4E",X"23",X"46",X"EB",X"E9",X"2E",X"0A",
		X"57",X"0A",X"4D",X"0A",X"2E",X"0A",X"39",X"0A",X"61",X"0A",X"71",X"0A",X"2E",X"0A",X"43",X"0A",
		X"81",X"0A",X"91",X"0A",X"2E",X"0A",X"2E",X"0A",X"2E",X"0A",X"2E",X"0A",X"2E",X"0A",X"EB",X"AF",
		X"77",X"2B",X"77",X"2B",X"7E",X"E6",X"0F",X"77",X"C9",X"EB",X"05",X"78",X"FE",X"04",X"38",X"EF",
		X"C3",X"A1",X"0A",X"EB",X"04",X"78",X"FE",X"C8",X"30",X"E5",X"C3",X"A1",X"0A",X"EB",X"0C",X"79",
		X"FE",X"FC",X"30",X"DB",X"C3",X"A1",X"0A",X"EB",X"0D",X"79",X"FE",X"08",X"38",X"D1",X"C3",X"A1",
		X"0A",X"EB",X"0D",X"05",X"78",X"FE",X"04",X"38",X"C6",X"79",X"FE",X"08",X"38",X"C1",X"C3",X"A1",
		X"0A",X"EB",X"0C",X"05",X"78",X"FE",X"04",X"38",X"B6",X"79",X"FE",X"FC",X"30",X"B1",X"C3",X"A1",
		X"0A",X"EB",X"0D",X"04",X"78",X"FE",X"C8",X"30",X"A6",X"79",X"FE",X"08",X"38",X"A1",X"C3",X"A1",
		X"0A",X"EB",X"0C",X"04",X"78",X"FE",X"C8",X"30",X"96",X"79",X"FE",X"FC",X"30",X"91",X"C3",X"A1",
		X"0A",X"70",X"2B",X"71",X"EB",X"60",X"69",X"CD",X"19",X"0C",X"36",X"80",X"DB",X"4E",X"07",X"D0",
		X"36",X"80",X"22",X"00",X"40",X"1B",X"C5",X"CB",X"38",X"CB",X"38",X"CB",X"38",X"CB",X"19",X"CB",
		X"38",X"CB",X"19",X"CB",X"38",X"CB",X"19",X"08",X"3A",X"22",X"40",X"B7",X"CA",X"DA",X"0A",X"21",
		X"FF",X"87",X"ED",X"42",X"C1",X"08",X"3F",X"C3",X"E0",X"0A",X"21",X"00",X"81",X"09",X"C1",X"08",
		X"DA",X"F4",X"0A",X"7E",X"E6",X"F0",X"FE",X"70",X"CA",X"05",X"0B",X"D9",X"B9",X"D9",X"CA",X"D7",
		X"0B",X"C3",X"21",X"0C",X"7E",X"E6",X"0F",X"FE",X"07",X"CA",X"05",X"0B",X"D9",X"B8",X"D9",X"CA",
		X"D7",X"0B",X"C3",X"21",X"0C",X"1A",X"E6",X"C0",X"28",X"1F",X"2A",X"00",X"40",X"CB",X"AC",X"7E",
		X"26",X"90",X"CB",X"51",X"28",X"02",X"26",X"09",X"08",X"3A",X"22",X"40",X"B7",X"CA",X"24",X"0B",
		X"3E",X"99",X"AC",X"67",X"08",X"A4",X"C2",X"2F",X"0B",X"01",X"57",X"0B",X"C3",X"32",X"0B",X"01",
		X"97",X"0B",X"1A",X"E6",X"F0",X"0F",X"0F",X"6F",X"26",X"00",X"09",X"1A",X"E6",X"0F",X"B6",X"12",
		X"13",X"23",X"1A",X"86",X"4F",X"12",X"13",X"23",X"1A",X"86",X"47",X"12",X"60",X"69",X"CD",X"19",
		X"0C",X"36",X"80",X"32",X"91",X"F8",X"C9",X"00",X"00",X"00",X"00",X"20",X"01",X"FC",X"00",X"10",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"80",X"03",X"01",X"00",X"60",X"01",X"FF",X"00",X"50",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"40",X"03",X"FF",X"00",X"A0",X"01",X"01",X"00",X"90",
		X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"01",X"FC",X"00",X"10",
		X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"80",X"04",X"01",X"00",X"90",X"FF",X"01",X"00",X"A0",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"FF",X"00",X"50",X"FF",X"FF",X"00",X"60",
		X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"E6",X"0F",X"12",X"AF",X"13",X"12",X"13",X"12",
		X"CB",X"51",X"11",X"F0",X"0F",X"28",X"03",X"11",X"0F",X"F0",X"3A",X"22",X"40",X"B7",X"28",X"03",
		X"7A",X"53",X"5F",X"7E",X"A2",X"57",X"3A",X"BB",X"F8",X"A3",X"B2",X"77",X"78",X"E6",X"FC",X"67",
		X"79",X"E6",X"FC",X"6F",X"CD",X"19",X"0C",X"EB",X"21",X"66",X"40",X"7E",X"C6",X"01",X"27",X"77",
		X"32",X"90",X"F8",X"21",X"80",X"0C",X"C3",X"6F",X"15",X"C5",X"06",X"90",X"CD",X"B6",X"2D",X"C1",
		X"C9",X"1A",X"E6",X"0F",X"12",X"3E",X"18",X"DD",X"21",X"AD",X"40",X"08",X"DD",X"CB",X"00",X"56",
		X"CA",X"76",X"0C",X"79",X"DD",X"96",X"09",X"3C",X"FA",X"76",X"0C",X"FE",X"0A",X"30",X"37",X"78",
		X"DD",X"96",X"0B",X"3C",X"FA",X"76",X"0C",X"FE",X"1E",X"D2",X"76",X"0C",X"DD",X"66",X"0D",X"DD",
		X"6E",X"0C",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"CB",X"7A",X"CA",X"68",X"0C",X"EB",X"29",
		X"29",X"29",X"94",X"EB",X"23",X"5E",X"23",X"56",X"14",X"14",X"BA",X"D2",X"76",X"0C",X"DD",X"CB",
		X"00",X"F6",X"DD",X"CB",X"00",X"EE",X"11",X"0E",X"00",X"DD",X"19",X"08",X"3D",X"20",X"AC",X"C9",
		X"01",X"04",X"60",X"F0",X"F0",X"60",X"06",X"05",X"CD",X"B1",X"17",X"36",X"1E",X"E5",X"CD",X"43",
		X"0D",X"CD",X"27",X"0D",X"C2",X"47",X"05",X"E1",X"7E",X"B7",X"20",X"F1",X"10",X"ED",X"CD",X"E3",
		X"17",X"C9",X"E5",X"21",X"00",X"00",X"39",X"CD",X"B5",X"0C",X"77",X"06",X"02",X"11",X"78",X"D5",
		X"CD",X"53",X"2E",X"E1",X"C9",X"3A",X"CB",X"F8",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"4F",X"3A",
		X"CA",X"F8",X"E6",X"F0",X"B1",X"C9",X"CD",X"B5",X"0C",X"FE",X"99",X"C8",X"C6",X"01",X"27",X"18",
		X"08",X"CD",X"B5",X"0C",X"C6",X"99",X"27",X"18",X"00",X"C5",X"32",X"CA",X"F8",X"4F",X"07",X"07",
		X"07",X"07",X"32",X"CB",X"F8",X"E6",X"F0",X"81",X"E6",X"F0",X"32",X"C9",X"F8",X"C1",X"C9",X"DB",
		X"64",X"B7",X"20",X"06",X"C5",X"E5",X"06",X"01",X"18",X"25",X"7E",X"B7",X"C8",X"C5",X"E5",X"35",
		X"C5",X"78",X"C6",X"00",X"4F",X"CD",X"0F",X"08",X"C1",X"E1",X"E5",X"06",X"FF",X"DB",X"64",X"5F",
		X"21",X"5B",X"40",X"ED",X"78",X"86",X"04",X"77",X"93",X"30",X"FB",X"78",X"B7",X"28",X"05",X"CD",
		X"C6",X"0C",X"10",X"FB",X"E1",X"C1",X"C9",X"C5",X"21",X"57",X"40",X"CD",X"B5",X"0C",X"F5",X"01",
		X"62",X"02",X"CD",X"EF",X"0C",X"23",X"0C",X"10",X"F9",X"CD",X"B5",X"0C",X"C1",X"B8",X"C4",X"A2",
		X"0C",X"C1",X"C9",X"CD",X"86",X"09",X"C8",X"CD",X"C6",X"0C",X"CD",X"86",X"09",X"20",X"FB",X"C9",
		X"CD",X"0A",X"0E",X"00",X"00",X"0A",X"20",X"99",X"CD",X"0A",X"0E",X"40",X"01",X"04",X"20",X"33",
		X"CD",X"0A",X"0E",X"C0",X"01",X"01",X"20",X"77",X"CD",X"0A",X"0E",X"E0",X"01",X"1F",X"0A",X"22",
		X"CD",X"0A",X"0E",X"EA",X"01",X"1F",X"08",X"11",X"CD",X"0A",X"0E",X"F1",X"01",X"1F",X"0F",X"33",
		X"CD",X"0A",X"0E",X"C0",X"05",X"0A",X"20",X"77",X"CD",X"0A",X"0E",X"80",X"06",X"04",X"0A",X"AA",
		X"CD",X"0A",X"0E",X"96",X"06",X"04",X"0A",X"EE",X"C9",X"CD",X"0A",X"0E",X"00",X"00",X"13",X"20",
		X"99",X"CD",X"0A",X"0E",X"60",X"02",X"25",X"20",X"BB",X"CD",X"0A",X"0E",X"E0",X"05",X"04",X"20",
		X"44",X"C9",X"CD",X"0A",X"0E",X"00",X"00",X"38",X"20",X"FF",X"C9",X"CD",X"0A",X"0E",X"E0",X"05",
		X"04",X"20",X"33",X"C9",X"CD",X"0A",X"0E",X"E0",X"05",X"04",X"20",X"66",X"C9",X"CD",X"0A",X"0E",
		X"00",X"00",X"08",X"20",X"BB",X"CD",X"0A",X"0E",X"00",X"01",X"10",X"20",X"66",X"CD",X"0A",X"0E",
		X"00",X"03",X"04",X"20",X"FF",X"CD",X"0A",X"0E",X"80",X"03",X"1C",X"20",X"AA",X"C3",X"88",X"0D",
		X"CD",X"0A",X"0E",X"00",X"00",X"2F",X"20",X"CC",X"CD",X"0A",X"0E",X"E0",X"05",X"09",X"20",X"AA",
		X"C9",X"CD",X"0A",X"0E",X"00",X"00",X"34",X"20",X"55",X"C9",X"E1",X"5E",X"23",X"56",X"23",X"E5",
		X"3A",X"22",X"40",X"B7",X"20",X"06",X"21",X"00",X"81",X"19",X"18",X"05",X"21",X"FF",X"87",X"ED",
		X"52",X"EB",X"E1",X"4E",X"23",X"08",X"7E",X"23",X"08",X"B7",X"7E",X"23",X"E5",X"EB",X"20",X"11",
		X"11",X"20",X"00",X"08",X"47",X"08",X"E5",X"77",X"23",X"10",X"FC",X"E1",X"19",X"0D",X"20",X"F3",
		X"C9",X"11",X"E0",X"FF",X"08",X"47",X"08",X"E5",X"77",X"2B",X"10",X"FC",X"E1",X"19",X"0D",X"20",
		X"F3",X"C9",X"CD",X"0A",X"0E",X"80",X"06",X"04",X"20",X"77",X"CD",X"88",X"0D",X"21",X"85",X"0F",
		X"01",X"07",X"00",X"3A",X"12",X"40",X"08",X"08",X"BE",X"38",X"06",X"08",X"09",X"7E",X"B7",X"20",
		X"F6",X"23",X"7E",X"23",X"32",X"0E",X"40",X"7E",X"23",X"32",X"0F",X"40",X"7E",X"23",X"4F",X"32",
		X"BB",X"F8",X"7E",X"23",X"32",X"A2",X"F8",X"7E",X"23",X"32",X"BA",X"F8",X"7E",X"32",X"B9",X"F8",
		X"3A",X"22",X"40",X"B7",X"21",X"00",X"81",X"DD",X"21",X"00",X"44",X"28",X"07",X"21",X"80",X"81",
		X"DD",X"21",X"00",X"46",X"3E",X"34",X"08",X"06",X"20",X"DD",X"7E",X"00",X"DD",X"AE",X"20",X"DD",
		X"B6",X"20",X"57",X"E6",X"0F",X"20",X"03",X"79",X"18",X"1B",X"FE",X"0F",X"20",X"15",X"DD",X"AE",
		X"00",X"E6",X"0F",X"20",X"05",X"3A",X"A2",X"F8",X"18",X"0B",X"FE",X"0F",X"28",X"05",X"3A",X"BA",
		X"F8",X"18",X"02",X"3E",X"77",X"E6",X"0F",X"5F",X"7A",X"E6",X"F0",X"20",X"03",X"79",X"18",X"1B",
		X"FE",X"F0",X"20",X"15",X"DD",X"AE",X"00",X"E6",X"F0",X"20",X"05",X"3A",X"A2",X"F8",X"18",X"0B",
		X"FE",X"F0",X"28",X"05",X"3A",X"BA",X"F8",X"18",X"02",X"3E",X"77",X"E6",X"F0",X"B3",X"77",X"23",
		X"DD",X"23",X"10",X"A5",X"11",X"60",X"00",X"DD",X"19",X"08",X"3D",X"20",X"99",X"C9",X"21",X"AD",
		X"40",X"CB",X"5E",X"C8",X"CB",X"9E",X"2A",X"AB",X"F8",X"11",X"AD",X"F8",X"01",X"1F",X"00",X"3E",
		X"05",X"08",X"1A",X"13",X"77",X"23",X"1A",X"13",X"77",X"09",X"08",X"3D",X"C2",X"21",X"0F",X"C9",
		X"CB",X"DE",X"11",X"09",X"00",X"19",X"5E",X"23",X"23",X"3A",X"22",X"40",X"B7",X"7E",X"28",X"0A",
		X"ED",X"44",X"C6",X"D0",X"08",X"3E",X"F7",X"93",X"5F",X"08",X"CB",X"3F",X"CB",X"3F",X"67",X"6B",
		X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"01",X"00",X"81",X"09",
		X"22",X"AB",X"F8",X"3A",X"BC",X"F8",X"4F",X"11",X"AD",X"F8",X"3E",X"05",X"08",X"7E",X"12",X"13",
		X"71",X"23",X"7E",X"12",X"13",X"71",X"79",X"01",X"1F",X"00",X"09",X"4F",X"08",X"3D",X"C2",X"6C",
		X"0F",X"2A",X"BD",X"F8",X"C9",X"01",X"00",X"50",X"33",X"44",X"55",X"01",X"03",X"01",X"46",X"99",
		X"44",X"55",X"01",X"05",X"02",X"3C",X"66",X"44",X"55",X"01",X"07",X"03",X"32",X"AA",X"33",X"99",
		X"02",X"09",X"04",X"2D",X"CC",X"33",X"99",X"02",X"0F",X"05",X"28",X"55",X"33",X"99",X"02",X"10",
		X"03",X"19",X"AA",X"55",X"44",X"03",X"11",X"04",X"14",X"44",X"33",X"22",X"04",X"15",X"05",X"0F",
		X"55",X"33",X"22",X"04",X"17",X"05",X"2D",X"DD",X"44",X"77",X"04",X"18",X"02",X"0F",X"66",X"44",
		X"22",X"04",X"19",X"03",X"0A",X"AA",X"33",X"44",X"03",X"1B",X"04",X"05",X"44",X"55",X"99",X"02",
		X"1E",X"05",X"05",X"55",X"66",X"99",X"02",X"00",X"05",X"05",X"33",X"44",X"66",X"05",X"CD",X"C2",
		X"20",X"11",X"5F",X"40",X"CD",X"2E",X"10",X"2A",X"64",X"40",X"E5",X"21",X"59",X"10",X"22",X"62");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
