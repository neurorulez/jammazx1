-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity INVADERS_ROM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of INVADERS_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D85108AC4F29B72B38BB46CE3B38AC62B74ED8A638ACA3B7D504A255035500C0";
    attribute INIT_01 of inst : label is "0000000000000000EE7A91838A8242EB4E1BB924B56D04AC61B38AC62B007551";
    attribute INIT_02 of inst : label is "1524260A5893964A49B538A2B38C2309D050B748E733412FFABBDA7B3B294B89";
    attribute INIT_03 of inst : label is "2512A5366B071278F9EC32499559DB9118DF621552B2256577C9CC7CF23E4BAE";
    attribute INIT_04 of inst : label is "C5986F4157B5DBB8BBB93B9A8E819C19D614565AB19489A4667AE9E36BD95969";
    attribute INIT_05 of inst : label is "FBC1A7AD3B2CACB8D9B65DC1338C644A92C41048AF9D828860BC7FBAD9FDBD07";
    attribute INIT_06 of inst : label is "2885B6D07AF6FC7FEBDB1BECECE6CCFB60408E53EDDED6421C1BA4EA2E89B510";
    attribute INIT_07 of inst : label is "8EC0C12D5D7CD2414E8A4AECAAE98EC6927BE9FAFC2D07FC663F39F88FCE3E61";
    attribute INIT_08 of inst : label is "08AE94F4984A95A308E0E188EE41A9ED45241BCD2C64A31851B425495410C128";
    attribute INIT_09 of inst : label is "4AA481C5E1708AC8E229D18A08A4585182329AC81C5E1709D18A08A458542CA1";
    attribute INIT_0A of inst : label is "C22CDE188658A36BE36BE34E422A92071785C22B2498A746282291E15ACA2992";
    attribute INIT_0B of inst : label is "31AA63A1382B38626A378694E26B29053CA34EE9F964B4A38ABBB03B6B180ED6";
    attribute INIT_0C of inst : label is "22ED147B459CE31A975046065BBA416E7E4F99CE57E58977239398E1BA8EAA8E";
    attribute INIT_0D of inst : label is "4DE4072C81E3C8BEE9D1A66698A2712AF89AB85292716788ABBB7B29EE34A094";
    attribute INIT_0E of inst : label is "8D2F4D655C139ABF73391C7204AFB4D1F91F9295423AD9FC89144A18664EBDA3";
    attribute INIT_0F of inst : label is "1916D462481451A9ACDB9E15575918E3855D75508205D3B0E2B6F89CDB4E2053";
    attribute INIT_10 of inst : label is "C6C20E9FDBFCB1BDC8DA403C1BD4921A5C415797B291759849254576D2B39D1B";
    attribute INIT_11 of inst : label is "539D35B8F244CA4AE18A7BAC73513B3B121D56422308223352CE36B1D52CE00B";
    attribute INIT_12 of inst : label is "912C86E2F46D11412490558642D9248AD8EF45BA546CE68561182187B2755C98";
    attribute INIT_13 of inst : label is "453991B855884948B9C894101CE3E955E55EFF5D997EEFFAFFE7291B319970B2";
    attribute INIT_14 of inst : label is "496FC8D9112488B39E19AA5BA530822AA50D174345509AEC2F26B9D9CEA9CE39";
    attribute INIT_15 of inst : label is "88DC29765FFAC896AC20AFEC5BB0BBB18B6F2BCAF05B9EA420B93651B9B3AC6A";
    attribute INIT_16 of inst : label is "F696F585D19A975146D785DB799A4DAF65869D65869C61A65EB0A9165B5DB49C";
    attribute INIT_17 of inst : label is "EAB0DB67FB5D3D9D881261A75E882A49C7EEC127136B5E8823711491946FE946";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "A5BEF9465417BF3FFBF394100000119507E539505FFD410465417BCFFEF39404";
    attribute INIT_29 of inst : label is "4886E96A0CA4B218A18642541DD09505E4661A7CFFE4661A7CE51B050950529F";
    attribute INIT_2A of inst : label is "7199C9129C951466C2040213E2B18812084D6C6E4E276DB492E546609DCA6448";
    attribute INIT_2B of inst : label is "C7BB1955E5417F3FFF395045E7BBB97C5154538A0819A85617B1948873B503F1";
    attribute INIT_2C of inst : label is "E85D9246DDD1A18AEA71985460B1461982C62C6AB38C60B81386738963462959";
    attribute INIT_2D of inst : label is "5DAA524811BC1DD573B669B6A94679B8D94D0AECEE5B4A9366CA46BEA2AF8AEB";
    attribute INIT_2E of inst : label is "65EB197209389BFBDB29E0449DB0B44D02E936D8864EB27FE2CA506D97FADD9D";
    attribute INIT_2F of inst : label is "E2B96D2241DD29B259204CA0ADB5FACE17C81E4F8451BC6C8BEB2813ADFFA8A9";
    attribute INIT_30 of inst : label is "222820AD5B097FBEFBCFA5B70951492C1097650C1389642A358D04B63BFB819C";
    attribute INIT_31 of inst : label is "202412A9CCD3AB38996481ACD2B509860986188AE0AA92C414E601FED14E4108";
    attribute INIT_32 of inst : label is "DD76B19A745F4517556615C16C538FD55E5FBBB9705704F84927338D7C17E17C";
    attribute INIT_33 of inst : label is "0D24945C816B57C2021FD198631B6AB0C3DBDB42A7282A9D2CA003F9935B7464";
    attribute INIT_34 of inst : label is "599505B9FE95B88C815CB8A9F7CE5DBBBB9A9FEDDC6342E1B1B25839C0A895A6";
    attribute INIT_35 of inst : label is "901AA1AB39C1AA9BC6903F8DA6F1A40F26B6103E91A02CC00808C017E5567536";
    attribute INIT_36 of inst : label is "07103E0F02014003C0064280C0844080C08000A0F04003C004001E8000020001";
    attribute INIT_37 of inst : label is "40C0C0003104000019A67030F030018000C3301024018C0C020104201211003D";
    attribute INIT_38 of inst : label is "4C7FFFD03FFFFFF0009006000894588002D28780006699000180090005A28A50";
    attribute INIT_39 of inst : label is "04F208A080000006E608880801862490F3020D3891C86A2D2EBD218710FFFED0";
    attribute INIT_3A of inst : label is "48000B8282E000450041146C11FFFFFFCCCCCCCCCCCFFFFFEA3866CE275E715D";
    attribute INIT_3B of inst : label is "0B4BA3B4BA713823C6129A12B000200429314A2383C00000A6FAEE0081A06240";
    attribute INIT_3C of inst : label is "000C09580C0C0C0C055C060C095801D00C0C0D58000C055C095C0958095C0C0C";
    attribute INIT_3D of inst : label is "095803000958055C01D00958055C00C00C0C0E2C0260095800C00958060C0658";
    attribute INIT_3E of inst : label is "18610592AE903ECA640F89AC0C0C08C800000000009001800254095800300958";
    attribute INIT_3F of inst : label is "0000B8E4A8A40F800008430CCCC0004019A640C0B31BDBEAC94AAD2424018030";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "32C30024CC20D401080BCC4A313824A239C844EB2824A1B27D0003550C550900";
    attribute INIT_01 of inst : label is "00000000000000090820E3300FC8C83E08234D9C00CB000C2113824A0300A002";
    attribute INIT_02 of inst : label is "231803128AF202C41170DF119184292AA02034C4A25AB01D5D4C061D1B1961C0";
    attribute INIT_03 of inst : label is "D7070080200201961611C404E2110540244D1F10B1C110E44EC6E60191BB1AF1";
    attribute INIT_04 of inst : label is "8731488C243194C21C12340BEFC011F20806C2B01095E440003300C4320E3323";
    attribute INIT_05 of inst : label is "A02B3C2D18E4E39E779BE7909384EBC6318005C4A211620C823442BF00292201";
    attribute INIT_06 of inst : label is "00DB9EB20E4254CC3B0B3804E4A1801C120020B92F62F9C8D2039C431004F070";
    attribute INIT_07 of inst : label is "4A741391514104D34FD65831A328E70272042108308DC15441CC2338E308CEBA";
    attribute INIT_08 of inst : label is "280888008C1C207118CCE31D23F3A359044D3A04527809093234E01355341322";
    attribute INIT_09 of inst : label is "C28C4081811284A9631930060064FC40C21388040818112930060064EC488987";
    attribute INIT_0A of inst : label is "42125629C24070209020900C881A310206044A12A59C64C0180193B1070630D8";
    attribute INIT_0B of inst : label is "9092729F2039288D4B304A5D141C2732447008E7562C7C40C669C23959088E5A";
    attribute INIT_0C of inst : label is "842B210AC8505C31D65308F1750F489479C5D646D4B5BE7D92A0042114074BCA";
    attribute INIT_0D of inst : label is "1B4C0414C8D17ADAFD2FD9836AF21F210C851C42721F17AC261C7119E7003088";
    attribute INIT_0E of inst : label is "A37C009EB9000E081C13C4D32064AC461381302AA1137306ABCC1D3803B35F90";
    attribute INIT_0F of inst : label is "27BEF1CC3289C330CC730C8C73E710433027AE7308027210A339794A3B247832";
    attribute INIT_10 of inst : label is "8A4A90B60DC6BBBCA63A00B2745EB5AAB7EB9DFB90AB4EB6EB18C33C38B18F03";
    attribute INIT_11 of inst : label is "2830BD8D81B04E8CB2C2844A86ECAB19C1A23AEC590803B50FC68FE082F46024";
    attribute INIT_12 of inst : label is "F0A048F1A8EBC6F01A3541DBEB2B1AA4967A8EFD380803428708B298492AAC5C";
    attribute INIT_13 of inst : label is "1D1A723BEA8F84ABF70508C88C6B2627D27DFF5A3ACD315B3532090390AB89C8";
    attribute INIT_14 of inst : label is "8019840EF8AE6B93AF1A82B9AB9080382B9033E49C720E2F91F3833075FD4610";
    attribute INIT_15 of inst : label is "1C44E8E8D038340A842020F92ABABAB08024390C802832CC201CBE6039929003";
    attribute INIT_16 of inst : label is "E2AD236CF00CB3C31EF323B13A79DB91238E3E238E38238E4A13A79E3BFC8F8A";
    attribute INIT_17 of inst : label is "F1C828AE88F8B2747CCBE38F4A0CE9EBC224AF9FCBCC0B0CE8F0C3EB8C0E0AC4";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "359017944801724C172495700000261200665120011D5709448014930524945C";
    attribute INIT_29 of inst : label is "50CA558FA4241B2839C69C4805E6120050037949305003694925035E71200730";
    attribute INIT_2A of inst : label is "410E4D72ACD174A63134732C50311D71184060438034EBBC5274C4711F4A4E42";
    attribute INIT_2B of inst : label is "379D04E14480124C124955C94461D58E3175210E2230F45F4513A48791BC0159";
    attribute INIT_2C of inst : label is "B842B18EBE63331D2FC38448C0538C10E14D84E49384604C03C6918E12030261";
    attribute INIT_2D of inst : label is "2772BAD5B1390A234339E78EE4E0C69E78EFB56C6958DE481A4E8CC0D8DC61AA";
    attribute INIT_2E of inst : label is "20691A412A21C66E7909320447929F480A06CD60C68CDCC14A5E0E32BA26BEB4";
    attribute INIT_2F of inst : label is "0238E3713CA720DC675404A94A2898C6244C8DB3448134350DDD1C812501CC28";
    attribute INIT_30 of inst : label is "E50AA8A4BC40918E18E7E88F3986C5A2FA7F23A279A7F0CB8DF082811C59C460";
    attribute INIT_31 of inst : label is "406930860C41A832E71C5092F1C08046A84601CCF00E31800883010AB10480A0";
    attribute INIT_32 of inst : label is "279D430D0BE4BE3AE7AEF8048302A0E107B34C4E032022091CF8B18451B00080";
    attribute INIT_33 of inst : label is "DB1B39BC70A908040620E20EF80F31C8282E4E075233054AC4E0080EC824A80B";
    attribute INIT_34 of inst : label is "EA1200A30596B0F0508477A1FDF16C4CC4E8106D6BF06C74055AC76248640A87";
    attribute INIT_35 of inst : label is "5D4C14C39594C17C11462E6BDF04418BD365462D45D716830CCEC024D409DD9B";
    attribute INIT_36 of inst : label is "36462D8B000000C3031D0100031C014003D00140F10B0080000CDCC022A80000";
    attribute INIT_37 of inst : label is "B070F000340000002BAEA6402B1001C0008322802EFBA190C300001234A3403C";
    attribute INIT_38 of inst : label is "01B3C4043FFFFFF000BBEE000EFFFEC00AFEBFA000AEBA000BFFFF800ABEBEA0";
    attribute INIT_39 of inst : label is "08B38C34C30C31D7F69181890A1001282800980531053083BDA6FFFB84A5E218";
    attribute INIT_3A of inst : label is "40007DF7DF7D0045004114E511FFFFFFFECCCCCCCEFFFFFF269546588A012404";
    attribute INIT_3B of inst : label is "00EF6D0EF6D842D9FBB7BBF3FCECECFEF041E54322C0A800AEEAAD082B48DDE8";
    attribute INIT_3C of inst : label is "02AC0C0C0D8C0C8C000C006C0C0000C00EAC050C02AC02AC0C0C000C06AC0D5C";
    attribute INIT_3D of inst : label is "0C00075C0680029000C00C9C009000C001900CCC0C0C0C0C00C006A002EC0C4C";
    attribute INIT_3E of inst : label is "0000007B19462DA5418B74D9019001D005540000090000180EA006A4009006AC";
    attribute INIT_3F of inst : label is "0AA851CEC7418B7B04C00304CEC000C02BAEA0C04843C9CACBEC504E2EFBA030";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "40008EF40CACC8029C0304AB22AC0ABAE42B80C7AC0AB241438AF39300930500";
    attribute INIT_01 of inst : label is "00000000000000022FBCC8F10FE3C03EA28AAE000000A812322AC0ABBE003C60";
    attribute INIT_02 of inst : label is "8B12338F76F8A32310223F18EACA32AC9388E512232E52140E2E8CAEAE8E72E2";
    attribute INIT_03 of inst : label is "859088C89C891033B38908A0C8008F220AAB2F88432388044F134A01C4D11CC8";
    attribute INIT_04 of inst : label is "B3300041A62AA6602E33C203CFE631C21494F18028CCE24238612184310C305C";
    attribute INIT_05 of inst : label is "AECC00D3AC8A322D862214E32ACAB501C45666126138FAFEBAE0E33FA02B0117";
    attribute INIT_06 of inst : label is "9CDC41C98101040804049C8AB273832E3A8030011C31C127C79E32BB8142CC83";
    attribute INIT_07 of inst : label is "27F40C3BFBEBA50C83CCC8380330CB990A4003802268780272C89F23F227C87C";
    attribute INIT_08 of inst : label is "BAF7E3AE2E0820B28E2A28985BE89C066A50C72A303232AD4AE2B61424C40CAC";
    attribute INIT_09 of inst : label is "E371224448ABEF4C97BC8BE7BEF12E10E32AE712E744BABC8BE7BE313ED2E80F";
    attribute INIT_0A of inst : label is "AF388CACE300BB9C0B5C0BAF26B9C4995126AFBD735EF22FBEF8C479632EACC0";
    attribute INIT_0B of inst : label is "2AC57BC8BCBCBEF127B82F33802E50B4ECFBAE87833122E22E12E78C12BDE300";
    attribute INIT_0C of inst : label is "251CB9472E3088BCFEFBAE58C20FEE0C60CEC6AB08024F6209CBCEF9D14B15EF";
    attribute INIT_0D of inst : label is "900001AEE68201C07F94C0DB36F88C8CAE212E25084C304E322E029C0B8838E2";
    attribute INIT_0E of inst : label is "CC077611CE39CDC44C89E73F9910722700300BAAA28F10623515808AF3530408";
    attribute INIT_0F of inst : label is "0401C22EBBE400BEF84BEF10C214AAAAF094618BAE090AE2B8E43084C44449BA";
    attribute INIT_10 of inst : label is "A22310410CC1424050C740110171C0004604310228C071051C850C00434AC08E";
    attribute INIT_11 of inst : label is "4305314108D8A32FF4E30084843604AE6821C00C228E3F37672B301D98EAB000";
    attribute INIT_12 of inst : label is "DA7127F3A510F719413A8BF21F80400850BA50F9426A33088F99F8DC10A6A8A4";
    attribute INIT_13 of inst : label is "23AC4AE3014F4125DB8E22E6E2B310402C0200DCCC8AB9E39E3ABABE2BC024E4";
    attribute INIT_14 of inst : label is "2A3B8EECCC70032ACF9C10400428E3F10400020040C9ECD3FBEB139AF2FAABAF";
    attribute INIT_15 of inst : label is "036AB334046702204A38C40982464348CC84310C0981044E38CD3148E028C633";
    attribute INIT_16 of inst : label is "8C104C5008CC420021CBC412BC43100F8C00844C00874021502ACC50C01911D2";
    attribute INIT_17 of inst : label is "021054400119504CBEA50021510EB31C60105051430F620EB31598103238012B";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "78404B14008BA119BA1161C00000070021D060022BBA1C010008BC466F116070";
    attribute INIT_29 of inst : label is "45E301D3CA3747AC30EB10008C850022FEB372C466FEB362C458AE7070022709";
    attribute INIT_2A of inst : label is "08CC9548C9414A3504757014C8EACD84A8E242B323751C10DCB42B3A98AB6277";
    attribute INIT_2B of inst : label is "872F05094008B119B11627010262D189C50A88E38F8CF143A728C5D02AEC000D";
    attribute INIT_2C of inst : label is "76D8035108C9FAB99FEA8EA2B1902BACC6410AB52ACAB32E63E72AC83A838F70";
    attribute INIT_2D of inst : label is "9460470149EE30141AE10C101998842D830CD1D2B4A1119890A351E5D5D05506";
    attribute INIT_2E of inst : label is "56629C1E9C9CCEEE628C798E662AD8E607014C70EB23D4199D01A778063109C8";
    attribute INIT_2F of inst : label is "79E3040D9DD49CD40408CA708410512B01EE68520E69EF361C2CEE69D4191E36";
    attribute INIT_30 of inst : label is "228D4E3042E22104208FC010AC07107105440C61075472B3311999C02E02E242";
    attribute INIT_31 of inst : label is "7E7038C092AAC88CD4202330C2F640A770A78CEFF8CDC44662330149C8A24D42";
    attribute INIT_32 of inst : label is "10518ACDC51071461851472E332ACC672022AE65CB9CB8C666424AEA51402206";
    attribute INIT_33 of inst : label is "D0463DC119722067A7148ACE011042106300D98FE19F37858A700311D8844237";
    attribute INIT_34 of inst : label is "060022609F6050F8E20AFB409E700A22E64706DC000556AC000015ACC892E1CF";
    attribute INIT_35 of inst : label is "A61061070A6106815291019020549440649A91029120001D856FC00028B63F22";
    attribute INIT_36 of inst : label is "399102400130904301440000018400C0018000C0F03950C001E60C0033FC0040";
    attribute INIT_37 of inst : label is "D09090001C0000001EFB470011400004006359C01EFB45C0614000001465A03C";
    attribute INIT_38 of inst : label is "00223040055FD540007BED0001EFED000FEBEBF0007BED000DEFEDC00FEBEBF0";
    attribute INIT_39 of inst : label is "08070C78C32E74C9F41899180090018041E48018010841940259FFF4100A1080";
    attribute INIT_3A of inst : label is "880007FFFFD0001457154155D437FFFFFFFFFFFFFFFFFF730000000000000000";
    attribute INIT_3B of inst : label is "050096500965152ED61E1A1A3484868685010A00500001B95555560105E17FD0";
    attribute INIT_3C of inst : label is "0C0C0C0C0C1C0E6C000C024C0C0000C00C0C000C000C000C0C0C080C0C0C0624";
    attribute INIT_3D of inst : label is "015C039009000C0800E00D0C0900091809180C0C0C0C0C0C00C0080C0C0C0C0C";
    attribute INIT_3E of inst : label is "000000802691026A9440992600C009D805540000018000900C0C0C0C09000024";
    attribute INIT_3F of inst : label is "0000851009944099856901054FC009081EFB7918901368685800A5101EFB5E46";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "31C32001C330072E20B2C78C1E30B8C321CC0C3B3078C1C33C3048FF0BFF03C0";
    attribute INIT_01 of inst : label is "0000000000000003CC303003C3C00F34C001472CB1C700B0C2E30B8C1200FFF0";
    attribute INIT_02 of inst : label is "010C00011CD011C01C52CC0011380E13C03023C000E700040F4403E511030E40";
    attribute INIT_03 of inst : label is "0C0010F103000CD91910F0303F3C000034493100F04000F0B14D792C53532CD1";
    attribute INIT_04 of inst : label is "101C0700FF13F442E41D942FFF400C70F0CF3C71E23C00008120C48300C33CC3";
    attribute INIT_05 of inst : label is "04470C331038C0E4F1E0CFC0E33843C0300000C002C01100412700FD32C01C01";
    attribute INIT_06 of inst : label is "00031C300B0B03C72C2C0078C40002E401003C30C73C73C80D022C4000C00CF1";
    attribute INIT_07 of inst : label is "C040C300000031C3F3430330333CF93C30071C071C0610000307001CD1C007F7";
    attribute INIT_08 of inst : label is "00003D048F0700DE2080821077420300001C30C00F3C0E10B0180FC7FC30C300";
    attribute INIT_09 of inst : label is "080C041071210410F31071041001F04CC8E130C00007021071041041F00C00B9";
    attribute INIT_0A of inst : label is "84038B10CC3ED10301030104C410301041C4841040CC41C4004107C131C41003";
    attribute INIT_0B of inst : label is "E1033107121110433E10C41C0734C31306D1044D4D1F0C40440E4E312E138C4B";
    attribute INIT_0C of inst : label is "41C310B0C41F87100001043071CD04C3137241440B02CD1D30310C4020C30CC4";
    attribute INIT_0D of inst : label is "0F1C033648CE0CC7340FCCFF3CD203220483E48C320300CC82E40E103923323C";
    attribute INIT_0E of inst : label is "0F03003C7C020032032041D920070C80C73C730010210C00E0410120C03F0702";
    attribute INIT_0F of inst : label is "0F2C73CC3040CF30C8F30C3CF3C730C3100F0C330C007308C3281CCCF3070003";
    attribute INIT_10 of inst : label is "C0400C32C072C1C0E0F2000C331CF01C70CF0C33E20B3C30CF03CB3C31C10F32";
    attribute INIT_11 of inst : label is "33C33F00F0038CC4CCC8CCCCB3C03C10002C33CB3E30C83C00043C0403C4400B";
    attribute INIT_12 of inst : label is "C83C08C000CB30C401C00340F90F01CCC3900F703C8080003923700330F00430";
    attribute INIT_13 of inst : label is "3F10F320F3DD003CCD000CCCC043CFCF3CF300F4B4B51149149F3332E30FCCCC";
    attribute INIT_14 of inst : label is "C40100C4753C11E33F031C71C7E30C01C70CF3C30CF2003101CD0C0843734413";
    attribute INIT_15 of inst : label is "C008C2F2CCE0C0CCF8C30B0032C1C2C307CF83D07132C0B0C3033CF322E30CC0";
    attribute INIT_16 of inst : label is "871CCF0CF30033CF3C730F1E30F2CF020B2CF30B2CF20B3C81E30B0CB3C82CC3";
    attribute INIT_17 of inst : label is "00000B0C32C83CF4C4C2CB3CC3CCC2C320F0C71C83C002CCC3C8000B2CC8B1C0";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "1F1CCDC7300D833818333C70000030CC004F0CC0311BC70C3300D8CE06333C1C";
    attribute INIT_29 of inst : label is "0EC04C7F7800DF033CC0CF3007B2CC036C402ECCE06C402ECCCF121F1CC031C0";
    attribute INIT_2A of inst : label is "72034C7034C47401C3E2E00FC020003013001C00C003C31C0392C00107401D0E";
    attribute INIT_2B of inst : label is "03E400FCF300D3381333F1CCF01E40B8FCF030000100333C82E032CCD112A804";
    attribute INIT_2C of inst : label is "20C0F00CBB3013107743000C0CCFC000333C7801E3380E440FC0D1030133213C";
    attribute INIT_2D of inst : label is "0F3C73C0F02C02CF3323CB2C0800F3E4F2CF40B04002C0800F8C1C404B8B2CB0";
    attribute INIT_2E of inst : label is "002E2333232000441E20D23081E1070803C0FC0CC0CC430038408210F1F0B8F0";
    attribute INIT_2F of inst : label is "8222CB0008CF200F0F00388CCF3CCF0433648C3F30822602CC35348202C0B880";
    attribute INIT_30 of inst : label is "C330B8C4F40CE1041073CF2D13F0C30C7C730B0C70C720403C0800F0E40E483C";
    attribute INIT_31 of inst : label is "888CC20330C10F30073C002CF0003CC42CC43004C20030304CC000FC330C002C";
    attribute INIT_32 of inst : label is "C73CF10073C70C70C30C70CC2C030F20002D4444330330F3000CC10C2CF3C0CC";
    attribute INIT_33 of inst : label is "4F03C434043C0CC8880FB3000000000003C0C0337300DDCCB80003C0800F2CC0";
    attribute INIT_34 of inst : label is "F1CC031C063F1DD000F4CD1C4510F5444470C04C00000000000000033AC44CF3";
    attribute INIT_35 of inst : label is "000000000000000000000000000000000000000000000000080EC00F3033D3E0";
    attribute INIT_36 of inst : label is "300000000000003300C0008000C0008000C00040F000808000010C8830440000";
    attribute INIT_37 of inst : label is "000000020400000001F401002CC0000000230A8001F4004002001000040C403C";
    attribute INIT_38 of inst : label is "00402000000740000007D00000901800015FF5400007D00004901840015FF540";
    attribute INIT_39 of inst : label is "000B4C30CB8C30C1219181890109181000000000000000000002484849401081";
    attribute INIT_3A of inst : label is "8000001554000000000000AA003337FFFFFFFFFFFFFF73330000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000C80C0C0C3001000100000000001555400000000248940221";
    attribute INIT_3C of inst : label is "0154015004040404000404040400015004040550055405540154015001540040";
    attribute INIT_3D of inst : label is "0554010005540150004001500554040404040404040404040554015001540150";
    attribute INIT_3E of inst : label is "0000000000000000000000000040004000000000001001000150015005540540";
    attribute INIT_3F of inst : label is "0000000000000000080300882EC0015001F40404000330101000000001F40101";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
