-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu1 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "833A3A2830855FFFFFFFFFFF3C6E1E930855D38FF5C5FF7B92FD510FF7EEF8C1";
    attribute INIT_01 of inst : label is "05AA56AF42C24249F029E25E260411E25E26D5727508AE9B619832954EE8BA29";
    attribute INIT_02 of inst : label is "DFA99476559BE0B4242493B89D3C2C4B92B73C26A95ABD0BE8EA97E8EAF7E8EA";
    attribute INIT_03 of inst : label is "85E50557F2CECA14B9C896999B8D54B9ACC2142C2D555552DFA9947655555552";
    attribute INIT_04 of inst : label is "F041488266D86D5412FEC85E5070FFFFCEB5F535542962D421584E262E8AD541";
    attribute INIT_05 of inst : label is "ED6C50B1CF2B063C72BC819C499181205144956B594513561644D8597C107443";
    attribute INIT_06 of inst : label is "BCABAAA9A8A84ED8DAF83446855705C6E78FDF425157D7EEEF0F53B4B8F0B57E";
    attribute INIT_07 of inst : label is "18D1902E529190939559C4B1082CA6347FD69C8DD5A94D5F5E5DEFED8F8D5C5F";
    attribute INIT_08 of inst : label is "8CF369495D79382C208EF7B93789561D84B612A79DD67B51FFFE4A9350890D96";
    attribute INIT_09 of inst : label is "6055366A0A08202B81C7519A5DDBF6552FE182B45264263422C6956909D55351";
    attribute INIT_0A of inst : label is "4D3B6A3480AC40400012675A653756575E46427A7554D63767D09365D2F8A778";
    attribute INIT_0B of inst : label is "15BC1EEA07810954636234282460B786608E984BEF29755555D8422C682C2755";
    attribute INIT_0C of inst : label is "B0BCAC18E6F0B3F6B4F08DD55771C67962F264279AB4DD4906666F9F82420167";
    attribute INIT_0D of inst : label is "0FC9985CF0810153CA0F20B5E5619DDC3499141256E2E2E2C2C1E7DC75CAAAB8";
    attribute INIT_0E of inst : label is "DCF091551D7B5579716CAC12127105092773099082FBE6831BECED7B9F6C1C75";
    attribute INIT_0F of inst : label is "93492234BC95DE786F283C25D5C70977741524150226C4BFCC9504569C579255";
    attribute INIT_10 of inst : label is "2B3C27D9A3635DDF7A8D8D77E4F2B3C28F59634922234BC95DE5B55193333F79";
    attribute INIT_11 of inst : label is "563F4CA49415CA73492E0293CACF0ADA7AB7FFB767D9A3635D2DF7A8D8D77E4F";
    attribute INIT_12 of inst : label is "73C206A57A5D5155F952FC02D5029C4B691075FFCB52505CA45072C1CB729250";
    attribute INIT_13 of inst : label is "09755F19635055F7D53393C2872A1098D669E65E71B6DC7A1CF0A1865F527172";
    attribute INIT_14 of inst : label is "55C8DE55723755615F7DE5D572A1098DE71B6DE65C79E48204A875A94CEE5979";
    attribute INIT_15 of inst : label is "15EAD1EF9792A9E697909755F5CEE0B994A859A49DE6B18D81579C8DD557237D";
    attribute INIT_16 of inst : label is "712FF2ED219CBFCAEBA155E4D0717524558EE0B5C64929ECA727414A554242CA";
    attribute INIT_17 of inst : label is "FCF7B8A1210FCFE0D308CFBA221C985F84DB87928373C21502C8DC888CF2F1EF";
    attribute INIT_18 of inst : label is "EED779A7CE0D571703333D075E2795F7583993971E5C4BFFF1857FFEDFF7FDF3";
    attribute INIT_19 of inst : label is "33D075E2795B0F2D2CE45357C592CBD60950954451059274B38179B63755C5FA";
    attribute INIT_1A of inst : label is "1441649D2CE462355C5F7694D79B63755C5FAEED779A50C4355C5F74B4793E33";
    attribute INIT_1B of inst : label is "00CCCC888844454BB8465406543CACF0B8152DE79590E026538ED088E8258951";
    attribute INIT_1C of inst : label is "4492F4F36DDB760944A3BBA3FBF6A591555D58551049D04BD245548888444400";
    attribute INIT_1D of inst : label is "762791558155541D7B6DE4BD9CBD075EDA7075ED92C1D7B61349E2F7792F6615";
    attribute INIT_1E of inst : label is "57DD55FD2D97DB894BFBFBFE21B2D8947D4A41F47141E56154455549D24BC1D7";
    attribute INIT_1F of inst : label is "8D2A35000012AE29F4B2860DCDCA6D24B55557167679D25B0B22D248F0A0B551";
    attribute INIT_20 of inst : label is "927971CA053D283A4B855CD90F90F9A77D76552CDB4D461375504B7FF7B96919";
    attribute INIT_21 of inst : label is "11111000000000154549D45795C70BB02E4B0B9445871971E5115D6A0808CD95";
    attribute INIT_22 of inst : label is "1152F9FF9B7415635A8DD088E663A39C9479F41CF089B92F4647E5373C215505";
    attribute INIT_23 of inst : label is "79654AD58BD06D846715C6579A79A5115649649C72BD8AE5D7A05566379A2919";
    attribute INIT_24 of inst : label is "4BD685506372F5109BA354514514514514514514514508000200000080000014";
    attribute INIT_25 of inst : label is "15649F72341D71C957236967BE7921949F4B9D425DA846B234A929F6492F8AB4";
    attribute INIT_26 of inst : label is "B5925079E59D4987B25929769F4B9D59D70B98C70B90E6E8D020828288D08D11";
    attribute INIT_27 of inst : label is "E49341F934B9D7984327D2E6155155F59C70BD82E49415172B49445841867054";
    attribute INIT_28 of inst : label is "9D958554DA59C708609B908639989415172B49445841867054B59255A5941E49";
    attribute INIT_29 of inst : label is "DF57351CB49A415C6332E15FD4248288D482C0288D88D820820000000792D78E";
    attribute INIT_2A of inst : label is "455927F7146FC9F79B695CDED89584BFE76424A7D2D5D209097A353752505652";
    attribute INIT_2B of inst : label is "A5E798D2E02756579A7F7195BCE4A636FC65421E69F194274A359279A5D5A084";
    attribute INIT_2C of inst : label is "7D2D4BDBB6712FEE426E8D00000000040C7584DD08272405C70BD82E7197DE6D";
    attribute INIT_2D of inst : label is "6D6B084455927D445C79A67E5479C8DE796796F6D9E4BF8D0F2E46424246424A";
    attribute INIT_2E of inst : label is "70B392D593902E4D24B8D27DA635C6579A7DC8D4435CC539BBDA43548D7962F7";
    attribute INIT_2F of inst : label is "19293929190909C8DD34D34D34D34C5B1080449D1141CA0859259271CAF62B9F";
    attribute INIT_30 of inst : label is "954B370224D04154D9C70BD82E5D68E23A34F8DC2111672D6490F9000C9A4349";
    attribute INIT_31 of inst : label is "49249249249249105D673482C8D651E594D2FFF24235115E696491F19755F1DD";
    attribute INIT_32 of inst : label is "6792FCB9B736712E329CEEE5737362E579A4C2298D5A34003000412492492492";
    attribute INIT_33 of inst : label is "0808DC6579A6340848D4455927F4A8AD1690971AEE17A556A363E726A5B09397";
    attribute INIT_34 of inst : label is "46705279575E5495C2E72375E6099C8D6B6E180B98099E68267979A2F6E76D5B";
    attribute INIT_35 of inst : label is "279C6579A71445592416ED24A53C325BE9095B44559271C6579A41D505BB59A9";
    attribute INIT_36 of inst : label is "957D4BC551DDCF095814F5A3298DC659F9A5115649CBF2E2797D00CC0CC6C1D5";
    attribute INIT_37 of inst : label is "124C37EF381DC4BD04FBC41C8D0507C104BF1714DD5575E56065FDF65555DCF0";
    attribute INIT_38 of inst : label is "0C40E6804D8537D83031023213103023203003614DF60C0C4C888D8537D83012";
    attribute INIT_39 of inst : label is "4DA0594DA855555640C04040408C84C40C08C80C00D8537D83300023614DF60C";
    attribute INIT_3A of inst : label is "790495E94366666CB9ECD1CEC064263EBBB9594DA3555D8F0B1556D5554F0A59";
    attribute INIT_3B of inst : label is "179C5B127823B902CF78EA51D3A947EC2A1618EEE2F8EA523068EA51270A316C";
    attribute INIT_3C of inst : label is "B8DCC930DCAEA2909D3C235A095975A1551BD0987414A31A41D90491C74B30C7";
    attribute INIT_3D of inst : label is "954D35C8D3416BD17234907A8D055543F420621E383DE0FF2032495945A555CC";
    attribute INIT_3E of inst : label is "7142711105851CDFB63750E3015FDF15DDDC8308408091BF88CDC190FBAED555";
    attribute INIT_3F of inst : label is "6964909E6914DF6985A5383774229A42764964944D43C2058555CA59703EC473";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C1091EA590805555555555550087225908056618530055A4E12CA3C15A135030";
    attribute INIT_01 of inst : label is "100F003A0601C1C441B843C43F1C7443C43FA331A00803D2811C109C003E2411";
    attribute INIT_02 of inst : label is "0000110002C281381C1C623C48382ACF73CC18203C00E8193236C13236A13236";
    attribute INIT_03 of inst : label is "F3B321DFF1C2CF84E48C470109C0929E924203BB380000040000110000000004";
    attribute INIT_04 of inst : label is "7000C842B4A04CCC316DFF3B3223EEEE42F39311DE3D33A1311C67038904CCC3";
    attribute INIT_05 of inst : label is "39131B4C462B008AF238407BC4C10010100C85583C403016450C09111C4038F0";
    attribute INIT_06 of inst : label is "10B3B0B1B2B320D3D12052A063425103632338D2302486139A2059CE6E04E361";
    attribute INIT_07 of inst : label is "74B87E33E17179707EF48CEF000C1F2D8F30FACBB9B220909392727352525251";
    attribute INIT_08 of inst : label is "5D360F844BD6003441001C4F5C5F5D760058017D34C5FD80AAA3C5F5EA5F25F8";
    attribute INIT_09 of inst : label is "6A5D97C4A58699B1802310CA407C1F901D5192E2210003FC038CDB07079EC111";
    attribute INIT_0A of inst : label is "0423732D2952BD04146132F58FFE33DEB8E1C1C1E7B0492C1C71F5F981C465F4";
    attribute INIT_0B of inst : label is "80428923EAC01BBE12E12C8C688231083204E507150946FBEF0CC038CC0C1E7B";
    attribute INIT_0C of inst : label is "64E498061E60A951C2E0849EC32F14B77101001F7DCFF9C033032A0A84060000";
    attribute INIT_0D of inst : label is "24040C82E088004B82AE10AB8CF03D301C7C0C001F819BA3A380FFF4D749D7E2";
    attribute INIT_0E of inst : label is "C2E0B4EF88CEBDE3AB37B80331303207120918C000D4DE69F984ACDFFFF804D7";
    attribute INIT_0F of inst : label is "F1C711F84AF2B5FE8E0AB826702301CEA80018048B3CCC7564F5014C723B7DEF";
    attribute INIT_10 of inst : label is "09B82872D2F2EBA1D64BCBACF4E09B8261D7B1C7113F84AF2B7E1C76F66661D5";
    attribute INIT_11 of inst : label is "D6804462F2356681C71F61D3826E0871F71D54C1F873D2F2EB5A1C64BCBACB4E";
    attribute INIT_12 of inst : label is "0B8232EA73EC80CDF681D5E310A3E2074720047FC76BC8D46BE9F1A7E6998BC8";
    attribute INIT_13 of inst : label is "07337EFCD2C1738E37129382BF000174BBC7DFFEF7BEF8CF32E0BBFF75001433";
    attribute INIT_14 of inst : label is "E72CB339CB2C8DEF38E36CCDF000174BEF7BEFDFF8CEDDC000000F0747ADC4DB";
    attribute INIT_15 of inst : label is "23A388A3BB7707DE4DB07337CF2FD08BCC002F1C4CDE6F4BC5CDF2CB339CB2C0";
    attribute INIT_16 of inst : label is "A01FF17230A07FC7AB722F0F79C8EF92370FD087A7EF10A0410F60863F448682";
    attribute INIT_17 of inst : label is "70C0331DFEDBB980F000A06031A47C87680EA1E1D00B821183C4BA8C628BABFF";
    attribute INIT_18 of inst : label is "889FC73D6D4DCB05EAAAA49D739DF65FFE8CF37B01E007EEE188FF032C8F22C8";
    attribute INIT_19 of inst : label is "AA45C735CF7CC15E1CE02379C0770DB39DD85C5D731177E87380430D0372C150";
    attribute INIT_1A of inst : label is "1CC41CFA1CE000B72C15FFC6633CD0372C150889FF7FDA60372C15FDD5F73DAA";
    attribute INIT_1B of inst : label is "44000000000002804DC6E286E23826E084B49E38F8FA3A33E30CC8D4EC6741C7";
    attribute INIT_1C of inst : label is "CC81DA41F27CDF274C43F74BB45F5DF2378735D73108E004B3C8DC4444444444";
    attribute INIT_1D of inst : label is "1F1FF13762378F79C9FE204AF6DB1F737F4DE727E1C7DCDF30001B6F8812FD75";
    attribute INIT_1E of inst : label is "1E3D7900180BB4C087E396789199E6E037A780DC9000F8D75CC41EC0E40747DC";
    attribute INIT_1F of inst : label is "CB232D00002E1DEAE07B2BD999829AD070000BB193B4D1840F27AD06E098F8D0";
    attribute INIT_20 of inst : label is "77E2F00303B30A13C800724F33B337B5F79F801D7DE7CA302871071D1C4F07C7";
    attribute INIT_21 of inst : label is "40C840000000002302C44C44770CA19C11DC0C71C76679F91D75EBD5ADAFC4F9";
    attribute INIT_22 of inst : label is "3221C754F02841F2C4CB767110A371EC4C37CC42E0844E1DCA31F000B8211558";
    attribute INIT_23 of inst : label is "DF5E27BA24B304DDDD375D7A7BD77D75E9EF5DF0C3C38F1EBF537B1D2F733777";
    attribute INIT_24 of inst : label is "24B31C7412D92C007232C20C00420C004308100308103C488F32230488C3222B";
    attribute INIT_25 of inst : label is "5E5DFCC12D71F322C592C73CCEF7FE7275E67CC5D732C3D12CC7279F9C1D461F";
    attribute INIT_26 of inst : label is "2F7FD5EF7D74D45CC5DF175CF5E67CDF9C8EFA9F0DFE7C6CB636A3C384B8CBD7";
    attribute INIT_27 of inst : label is "5EF423D79E67CDF5D85D717D75E2075DF0C3C38F1EF234701ED8DF7DC060F818";
    attribute INIT_28 of inst : label is "F0175D7805DF0C3DC27183DC171AF2347092D81C71C060F8182C73CD5DF57BEF";
    attribute INIT_29 of inst : label is "C7D69B0C62F1235259B18B90063A634CB623A834CB04B4514D2003939BFFBD45";
    attribute INIT_2A of inst : label is "D7977ECF301C07DEFDEF34327D5E70753D9C9C5D79CD7B1707632E720BC8D881";
    attribute INIT_2B of inst : label is "BCDED4B36B9337D977ECF7DE70DCDD2DC5D783E5DFB7DF8F412F7FF7FEBC52F5";
    attribute INIT_2C of inst : label is "D79CEE7C9F941D13C1DCCB00100010040493527CAFBC1C070C3C38F1D75F7BF7";
    attribute INIT_2D of inst : label is "ABC42F5D7977F3DF7CE7BD8EEBD026B51F5F73DF7E607F4B4ED3C1C1C9E5C5C5";
    attribute INIT_2E of inst : label is "C2D9F9CDF976B7C71D74B3F7FD375D7977F324B019725D1F1B7FF37E4BBF3120";
    attribute INIT_2F of inst : label is "370797171717070CB8E28608E28605394A70006071E765AFB7FC73C3030E0C75";
    attribute INIT_30 of inst : label is "EA079F67BE09FA766F0C1C3871EBF68BA92E84B63D75CF0B5DFB3B999EC3E427";
    attribute INIT_31 of inst : label is "0C72CF0C72CF0C69E0FDDC6B24B7EF7D7A01C75BE92D75E9EF5DFA279FAC2A27";
    attribute INIT_32 of inst : label is "FA81FF4F1D1FA81E0474313CD0C5FDA1F7347A07CBB32C0031541032CF0C72CF";
    attribute INIT_33 of inst : label is "0FECB9E7A7BF2D0F8CB5D7977ECC283880741EEE26273E8B12E0EEE73EC17071";
    attribute INIT_34 of inst : label is "E0F015CF8D392C47E3BD32D3910DF6CB90380A86F085F46E35EFBF310130ABD5";
    attribute INIT_35 of inst : label is "5CF9E7A7BF05D7977C0B073C1FB997EC0741EC5D7977F09E7A7BD71E02C1CF07";
    attribute INIT_36 of inst : label is "B0901F6ED0B42E0B0D20E1A0474B9E73E7BD75E5DFA3AA65CF4D3804804B171E";
    attribute INIT_37 of inst : label is "DD2B02319D0EB076828E0105C002C9C01077D08BF8CDEB8D9A0D1E731EEF42E0";
    attribute INIT_38 of inst : label is "0220340042121021000881099099098088088084840840022000021210210FCF";
    attribute INIT_39 of inst : label is "C4533DC85937EFBD001313131342642642602202202121021000001084840840";
    attribute INIT_3A of inst : label is "EBD3E0499EF61CFB43403C03AFC22A00C44E3DC4533EF42609BBE33EFC0E0BFD";
    attribute INIT_3B of inst : label is "F826FE4FA3B1A8DF6B21B26886C9A2BE76225BBC768BB2646932B264459C9BF9";
    attribute INIT_3C of inst : label is "566835980C75C9C8D0B82104863DC812372371A4E80040C1909110C8223DA663";
    attribute INIT_3D of inst : label is "DDC4336CB10CD7700B2CC132CB03779072763A0BBD93D6FF1823CE3DC0135C81";
    attribute INIT_3E of inst : label is "9AD8F88003290A6AA0AA82A98063F7E08888AC882959E10C0799B1A8A1E1E333";
    attribute INIT_3F of inst : label is "CF3C7AF7D70E74D3833C40CCCFB873E0F3C73C740CDB823393775E0A0AAAA2AA";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "DA8DAD4CD4E2B00000000000108B20CD4E2B04D3021200A6518538DB02990323";
    attribute INIT_01 of inst : label is "888E6239A343C34C44B443C4373CDC43C43782803E0E33AE38DDA8CBA33BE78D";
    attribute INIT_02 of inst : label is "00000000009E78E03C34C8FCE6323D0C037082323988E68FB3B19BB3B19BB3B1";
    attribute INIT_03 of inst : label is "ABB986E40E936EEAE6AE271312E2302C33538BB3B00000000000000000000000";
    attribute INIT_04 of inst : label is "E12242932B8E3A6CC882BABB984A0000938BA986E7BABB88B89CCB8AF9E3A6CC";
    attribute INIT_05 of inst : label is "9842440D208E008D28ECC26C0E299638B4B8080A5AD2E02250B80962980CAE36";
    attribute INIT_06 of inst : label is "5AABAAA8AAA9583A39E88A2A0939393809214F3884608699B255CAE2C552C9A9";
    attribute INIT_07 of inst : label is "DC1CD33348D4D0D0D71A60F08E3836048938D281D8AB59696B6A59585B5A5958";
    attribute INIT_08 of inst : label is "88138D0E64006D31B4D3340D340D34DD6935283769E06F52CCC144D37C4D28D0";
    attribute INIT_09 of inst : label is "7534A34040404CB8EE1A88EB20DE374A1429C48A83AA33523360C80D0D52D984";
    attribute INIT_0A of inst : label is "668E02040000011000038900245183310733634354B6630434DCD374614A734A";
    attribute INIT_0B of inst : label is "4000B01328128DC5A04A05CE32BAE9E739E7D085204C821C71E523360E3A354B";
    attribute INIT_0C of inst : label is "4280322100C8CAE1E288E652D9B0000073A3A834C47145258A7679D9E363E200";
    attribute INIT_0D of inst : label is "1E8EAEA288EAE209132808D0726A6A9B341E6659A62906280A22E1020000CB01";
    attribute INIT_0E of inst : label is "2288D271E60D031C34F1222FE021880D398A8E28E384300A9C8A311784322200";
    attribute INIT_0F of inst : label is "D3C33EC46058817C444CA23840AA636E200934A5333DB80028F6C6E0DAB0CC71";
    attribute INIT_10 of inst : label is "4CA230F7F0F0C8C3C7C3C321F644CA2313C5F3C33EEC460588343CF0D88883C4";
    attribute INIT_11 of inst : label is "246A353488094723C3EB1EC913288CF0CB3C02E3F0F7F0F0C81C3C7C3C321F64";
    attribute INIT_12 of inst : label is "8A23A888D34A13EE0B614310BA37DA8587506E0038422025700215C84311D220";
    attribute INIT_13 of inst : label is "0D9999C50068D953C928CB23329820D01934210F3CE3460CC2CAC8304409902A";
    attribute INIT_14 of inst : label is "582C1B960B06A64C953C026669820D01F3CE3421060C01EE0A60A40DEA730240";
    attribute INIT_15 of inst : label is "9B022A0080070D312400D999A4232AFC5260A4D0E6311C01A36542C18960B066";
    attribute INIT_16 of inst : label is "4A140E39BAD8503B00BAA4B043C6504A99632AE47FCF990268DA81664C6666A6";
    attribute INIT_17 of inst : label is "3AE63A9100033330F0003000FECD3EACB41C2AD1788A23BA6BA0132FBD8B3BF0";
    attribute INIT_18 of inst : label is "2211279CA2DFC3832CCCC2BEFBAEB8D1349EF7F38A1485CCC9E6FF9BAE63BAE6";
    attribute INIT_19 of inst : label is "CC2FFFBEFB80DB091639BBF3E079AC3887E2BEBEFE02BAE458E6AFBE57F0E0D2";
    attribute INIT_1A of inst : label is "FF80EFB91639B4BF0E0D1346B2FBE57F0E0D22211279CAB37F0E0D1240B702CC";
    attribute INIT_1B of inst : label is "91919191919190D664A7286728913288D24A4830F0F2727BC8E38CC2332F2FFF";
    attribute INIT_1C of inst : label is "FA9002A7FAFE7F0FFE08C90A323F2CB9BB10B3CFE025148611E6ED9191919191";
    attribute INIT_1D of inst : label is "BFADBABB19BB2EFBEBF1686276C3BDF9FC8BEFAFD16F7E7FE029AA0C5A185CF3";
    attribute INIT_1E of inst : label is "33C892AA22A1066605C30B70E9DE44D9800366001812F2CF3F806DC917852F7E";
    attribute INIT_1F of inst : label is "814204E4E4C9C29D24A333D2122611885EE040033B4E650CDCC7D884C8C8D274";
    attribute INIT_20 of inst : label is "926B3223085098A35C08D28D408400374D375215D34DE7E6A6904000348D0DCD";
    attribute INIT_21 of inst : label is "CC88882003000009D14111E019E0F8CD504DDF075D20D34804D34410FCCF28D4";
    attribute INIT_22 of inst : label is "E0000100D4A41A60548100000027EAD88F4B521288ED2114E7498088A23B8000";
    attribute INIT_23 of inst : label is "0515201520105A34348D34D4514924D35145249E0CF433C04008D23704030D0D";
    attribute INIT_24 of inst : label is "201375D0A0490428D4206186186082080104104000003C000F30330000C33300";
    attribute INIT_25 of inst : label is "3514540A05D7481B20A05145020030D0D34013034D31D3CA05010D375214A737";
    attribute INIT_26 of inst : label is "5892550D14511675C60D1D74D340130D34ECD134ECD3363413313F33281641CD";
    attribute INIT_27 of inst : label is "54868055740131D75861D576DB516974DE0CF433C0880958805634D34239A066";
    attribute INIT_28 of inst : label is "D51DB6D41A69E0CC8D58DCC8D58C88095880D63CF3C239A06658B2EEA6954355";
    attribute INIT_29 of inst : label is "00C5AE45748C80461AD5F02AA33133241573573241681041041113FEA0C34209";
    attribute INIT_2A of inst : label is "4D49264082101D34D34D9D98DC25785034343434D030DF0D8D62045742202360";
    attribute INIT_2B of inst : label is "3600E8129F08C36492640D3540343605034D33D2498D35DA5204514924410CF3";
    attribute INIT_2C of inst : label is "4D433CDE375E14236350813A223A2220200448D8CF34759DE0CF433C0D34D34D";
    attribute INIT_2D of inst : label is "B411CF34D4515034D20105C20016201485140734DD7850812423474743734343";
    attribute INIT_2E of inst : label is "4DCCD430D4D3734D04A4134D358D34D451502410B4D134CD8CD348D6810C73BA";
    attribute INIT_2F of inst : label is "4D0D4D0D8D0D8DA8104104100000003FF4000071D74D84CF4515967837D0DF03";
    attribute INIT_30 of inst : label is "D585363335A364D28DE0DF437C040113400500133CD35A96249508555523540D";
    attribute INIT_31 of inst : label is "08238E38E28A28821615365B2013401455A141035804D3514524960D3456860D";
    attribute INIT_32 of inst : label is "7561408D7477561500D232367663704A4072A70D81420400300010638E38E082";
    attribute INIT_33 of inst : label is "DF64134D492504CF24134D4926426422A0D2755D1DDD35A72050214335C1D1D7";
    attribute INIT_34 of inst : label is "39A46659244594193B34904458ECD24138A223D4D7D0D237B14D0C739BBAB411";
    attribute INIT_35 of inst : label is "65934D4927134D4924171D7434B0A75C0D275C34D4927134D4925D7505C75D0D";
    attribute INIT_36 of inst : label is "D6102C170916288D6398C9D00D8134D68924D352494310B55500208008C71D75";
    attribute INIT_37 of inst : label is "64DB6E882D117850EF240126C048D7B2042602A1463310733C9AB860A4716288";
    attribute INIT_38 of inst : label is "2102010000000000108400C00C00C00C00C00000000004210220000000001545";
    attribute INIT_39 of inst : label is "1608951A099971C4800303030330030030030030000000000108000800000004";
    attribute INIT_3A of inst : label is "516555A1674445041041D41451944365E264951E0897166C8C5C69C7166C8D05";
    attribute INIT_3B of inst : label is "54755495448511255042485109214445844691455B11485896044858A5611552";
    attribute INIT_3C of inst : label is "C2BDBCADA130CCEDE8A2398040951208998D88CA24A535D3419542D914554946";
    attribute INIT_3D of inst : label is "525E892835A241094A0E1990C38BB916E1B23C8070A92100E20340951A09A6DA";
    attribute INIT_3E of inst : label is "35CCA3C10BD7D0B4C76A4D0AC24ABAC22220D0D0364EC9A6AB12398D661089B9";
    attribute INIT_3F of inst : label is "4F2CB0D14534D34D8936492EECC853C9A2CB1450224A23899BB96C0889530F4C";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "024024000810FFFFFFFFFFFF2CB92C00810FFB7DF2E0FFF44037F0C1FF11F1D0";
    attribute INIT_01 of inst : label is "407981E51000C0C07C2072C72D0C3072C72DC110FF8100410410241FD0041041";
    attribute INIT_02 of inst : label is "000000000361442C0C0C34321CDD02D0B00C1D01E60794414078614078514078";
    attribute INIT_03 of inst : label is "534343FC0F2009009009040C0E50C3E70020431F1C0000000000000000000000";
    attribute INIT_04 of inst : label is "60106DE0D0410BFCB33315343402333360534343FC240241241339410410BFCB";
    attribute INIT_05 of inst : label is "1F010000074300F2E42C2072E1C4140833EC0F0608CFB03D80EC063338043C30";
    attribute INIT_06 of inst : label is "14151515141614373714171717171727273C31C433FC0F11EC00024070007FF1";
    attribute INIT_07 of inst : label is "3CF430F1F430303030C42C0B81080F3C4F20704F271614070606363615150505";
    attribute INIT_08 of inst : label is "08B107E1C2C3D2070C341CC71CC70C34C0D3031D7BC2D13C3331C071C0C7487C";
    attribute INIT_09 of inst : label is "000C21C000000024100700DC0C741D0406340F773871003D082C0B03832DC404";
    attribute INIT_0A of inst : label is "10423D3C00000000003870B0C73CF02CF2D0F0C0CB710F3C0C7871D0404D01CD";
    attribute INIT_0B of inst : label is "201C1C730760403233C13C0D0D042614041041013080F2C30C40D082C10A0CB7";
    attribute INIT_0C of inst : label is "F070DD02CF7402434074102DC70B00CB0008700C700CF2D041898525109050C0";
    attribute INIT_0D of inst : label is "4421C50074106001E007040F2FF37B311C758D853EC1C3C1C1D03CB1C70CCDF0";
    attribute INIT_0E of inst : label is "C0740C0C83C0F2CBCB01DD00B0104303870241C420831C02403902C0F2ED01C7";
    attribute INIT_0F of inst : label is "71CBF3700C7C32F037801D0FC072C0CF304F000F031CAC1A087F6140373C700C";
    attribute INIT_10 of inst : label is "801D0C7B33F3C371CDCFCF0EC07801D0C1CBC1CBF33700C7C31F1C78733331CC";
    attribute INIT_11 of inst : label is "FC0004DCBC7F4DC1CB310341E0074072CD1C0041DC7B23F3C3371CD8FCF0EC07";
    attribute INIT_12 of inst : label is "01D040C071C4F1FF4D30680073034701CF011C403DF2F1F4D0F3D34F4DD372F1";
    attribute INIT_13 of inst : label is "8373FC71E3F03F1C7FE401D03F50083CF1CF0C72C73CB2C0F0750F0C3C053024";
    attribute INIT_14 of inst : label is "C304F630C13D8FCFF1C72DCFF50083CF2C73CB0C72C32C10A1400B03C901C3CB";
    attribute INIT_15 of inst : label is "533DDC3C7CB0031D3CB8373FCB0335031D40073E1C1D078F80FCF04F630C13DC";
    attribute INIT_16 of inst : label is "0C040F512500103D3CD50F2C30C3CB073F03350302C7533D4C1EC014CBD414D4";
    attribute INIT_17 of inst : label is "74D1377000033330F0202C0F7F74C544D00F0E404501D0430304F2DFDCC1C2CF";
    attribute INIT_18 of inst : label is "CCF2C71D03CCF3CF0333371C711C7CD2F00C7333C0CC01333514FF766D9B55D5";
    attribute INIT_19 of inst : label is "3371C711C7CBC10805843333F07004FCF0F00F1C7B0071F01618C71F0F3CF3D8";
    attribute INIT_1A of inst : label is "1EC01C7C05843033CF3D2F109C71F0F3CF3D8CCF2C71F09F33CF3D2C1DFB9333";
    attribute INIT_1B of inst : label is "33773377337733C045D43014301E0074000C0B0C7C703031F61882CD83C300C7";
    attribute INIT_1C of inst : label is "ED406081D0741D031E00CC01C01D1C753FC3F1C7B014C500C1D4FF7733773377";
    attribute INIT_1D of inst : label is "1D1C753F053FFC71C1DC500C704F1C7074F1C70740471C1DB014013F14031C71";
    attribute INIT_1E of inst : label is "2C7FFF03DDCC7454C1B8CD4EF51F7B0407DD181CF03CCFC71EC0FCC0C501871C";
    attribute INIT_1F of inst : label is "CF1D3EFFAA7423403010034CCCD4FC4012AEBCF0DD0873C00CB344037400DFF3";
    attribute INIT_20 of inst : label is "71F3F80310075021C70030873C73CB01C71D000471C714B333F001A61CC70303";
    attribute INIT_21 of inst : label is "CCCCCC200200303FCCC03CCC7F1C241C31F00C71C70071C01C71F2C03C0D0870";
    attribute INIT_22 of inst : label is "B0004BA870300FF3CB4F000000F332442C8D0D4074104406141380501D040000";
    attribute INIT_23 of inst : label is "C71C04F004F0000C0C031C7071C71C71C1C71C71C0C7031F2C003C0F3CB00303";
    attribute INIT_24 of inst : label is "04F01C7033C13C8833D3C30C30C30C30C30C30C30C30CC0C0333300080031330";
    attribute INIT_25 of inst : label is "1C1C71C13C71C703FC13C71C71CB003031CCB0C0C700CB013C07031D0804D01C";
    attribute INIT_26 of inst : label is "5C71F3C71C73C80CB2C7031C71CCB0C70C0C700C2C702D0CF0B0070B04F04F47";
    attribute INIT_27 of inst : label is "1CB207471CCB0C70C72C731C71C03F1C71C0C7031CBC7F2013C81C70C00DE031";
    attribute INIT_28 of inst : label is "73C31C7001C71C0DC0B400DC0B40BC7F2013C81C70C00DE0315C71FF1C7CF1C7";
    attribute INIT_29 of inst : label is "693C2734DCB207F002534FF030700F04F00F00704F04F0C30C3334000CB02C38";
    attribute INIT_2A of inst : label is "C7071F1C7003031C71C7FC30743C001A1C0C0C0C730C7C03831D3F19F2F1F040";
    attribute INIT_2B of inst : label is "1F2C38F0423C31F071F1C71C0C0C0F3C31C70F41C7C71C1E3D3C71C71F2C00D1";
    attribute INIT_2C of inst : label is "C730F0741D080631E0CF4F333333331010CF10780C1C0C031C0C7031C71C71C7";
    attribute INIT_2D of inst : label is "42C00D1C7071C71C71C71CB1F0CC04F3071CB01C742010CF0731C0C0C0F0C0C0";
    attribute INIT_2E of inst : label is "C2C0B30C7830B1C72CC8F1C71C031C7071C704F000300C0B4071D0304FCB0E51";
    attribute INIT_2F of inst : label is "4303430303038304F000000000000A955003012C71C34C0D071C71C7031C0C71";
    attribute INIT_30 of inst : label is "40011E031CC0C030871C0C7031F2C0731D3C7CF0B471DE571C71C7000C01C303";
    attribute INIT_31 of inst : label is "1040000000000033C01D1CF304F1C31C70C06101C13C71C1C71C72C71F0032C7";
    attribute INIT_32 of inst : label is "D00040C71E1D00047030331FF0C1D003CB009003CF2D3C043C00104000000104";
    attribute INIT_33 of inst : label is "0D04F1C7071F3C2D04F1C7071F1D41DDC0300C08C84B1C82D3C71C331CB03031";
    attribute INIT_34 of inst : label is "0DE031C7FCF00C0F031C13CF003C704F043D008C708C750032C7CB0E726182C0";
    attribute INIT_35 of inst : label is "1C71C7071F81C7071C82C71C0C1C21CB0300CB1C7071F81C7071C71C20B1C703";
    attribute INIT_36 of inst : label is "04F00300C1C407404443770703CF1C77871C71C1C71DC791C700304004C2C71C";
    attribute INIT_37 of inst : label is "00CF0711E78C301BC90B038C00E3C190003E01CCF3F2CF2FF3DF1BE0FF0C4074";
    attribute INIT_38 of inst : label is "100100223000000000400C000000000000000400000000100222200000000221";
    attribute INIT_39 of inst : label is "F80432F8063F0C31010000000000000000000000010000000004CCC000000000";
    attribute INIT_3A of inst : label is "000003C00000D000300380380000EF004447F2F80430C40740032030C4074072";
    attribute INIT_3B of inst : label is "00D000000C00000000F00003C0000F00000D000000340000000D000000034000";
    attribute INIT_3C of inst : label is "109C0027860400C2701D040003F2F0043F40343C300C303000F301300C00000F";
    attribute INIT_3D of inst : label is "2FF84304FE10C034013D04034F43FFF06000341C30233000F071C3F2F80FFFC0";
    attribute INIT_3E of inst : label is "30C1EE4003C30F933F3300C240F11478CCCEC02031C1F400DECCD43C0080BFFF";
    attribute INIT_3F of inst : label is "C71C7071C71C71C7631CBC0CCC00B1C1E1C71C7010C1D04363FFC0063CCCF933";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
