-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D352A0B57FEA2A4977BB18080082410493A17FCFB718695F95FEA7A3D3F3EAB5";
    attribute INIT_01 of inst : label is "208B53050688596AA38094500A24F28449614EA8FBC4F2612971B05C07AC02D0";
    attribute INIT_02 of inst : label is "FC616582249E4F061E45A982F781CB31445F03C419E84F03FF2289804DBFC109";
    attribute INIT_03 of inst : label is "89B63410344D9CAFED990C5043700EA7DC55555ED5E67E73C262E38A88145499";
    attribute INIT_04 of inst : label is "51A089270943A937BBA93780076A8522A21166842AD64C1728AB834419386F50";
    attribute INIT_05 of inst : label is "F34F2110D2108910805499B883E2D415122286315E25C47E8BC50451075D544E";
    attribute INIT_06 of inst : label is "4250545C512B4B32A602B64F14BA4DFDB349E492C9BD50493C0A4D0060B24174";
    attribute INIT_07 of inst : label is "829D5134F22CF4224501505499A48FD17E8F9C7A14936A1964B02AA294A2545C";
    attribute INIT_08 of inst : label is "830615731605408A9A97523A1128A7118145084A0E87140824926D50CB94E216";
    attribute INIT_09 of inst : label is "54CA121CA721674943381D902702F8AD58C58A4236918946074DE28A00013802";
    attribute INIT_0A of inst : label is "0124C9D65DF6D4EBED1FB80AFE698E58E738922B18201AA08422A43896244542";
    attribute INIT_0B of inst : label is "E5EB397467B396ACE5D199110A51D6846A3DD99A0867819214870E9F122A1D00";
    attribute INIT_0C of inst : label is "6B64AA0978053234FBB84E2BE5E79653807D913E85137D246FA142D79E5651EC";
    attribute INIT_0D of inst : label is "0065F7E9E00041882DCCBD13E898CBF13E89886EA5A11A3AD6B1955950B5A7F2";
    attribute INIT_0E of inst : label is "85B548468F01009124598E6A22882AD59ADD56D23D4A4ED952BA0284EDB65400";
    attribute INIT_0F of inst : label is "F4A295C73B654AE89C589DB05B731885559263340305B27CBA5FD229C587F434";
    attribute INIT_10 of inst : label is "27D74148A8F2C9B6D28C5AD2B138C30E8DB55592F44F98D5564BF13E621BA97F";
    attribute INIT_11 of inst : label is "EF7F119E3768C5EE6CFBDFF11A5D76E27AF816A69B46E37D78F97539621A8572";
    attribute INIT_12 of inst : label is "0B1A0B4C50962510C48201547BBC4D10C674809C069A3A2A10AB50F7389A30C4";
    attribute INIT_13 of inst : label is "084546A0EB0C98394CB61EBBB0BBBBBBBEBBEEB734C2F3E330000EAA465AAA44";
    attribute INIT_14 of inst : label is "8D0918952320E8076376325A8341C4A881AE9CC930E60660D74F76216C736985";
    attribute INIT_15 of inst : label is "8BC8E48A2FFE4E880F51E6212262E221589B4358CA17429C88993C46D35C0290";
    attribute INIT_16 of inst : label is "ABCF40838708A302315814F5635D52D15505BA343749AA2A41A13C9263A14808";
    attribute INIT_17 of inst : label is "088D11C7AA801570B003B7378DF741A66D0AF7DBC646754A7661364651397DDF";
    attribute INIT_18 of inst : label is "06845ADA168B448DC8AA48A4CCE8D70C5F2D812B88F7399239CD38191C264767";
    attribute INIT_19 of inst : label is "2E7BFF822726DCCCE49B8C34294A3010D7DC0BC7E82692858267E886AC18A310";
    attribute INIT_1A of inst : label is "51100284406842221250C068413619260C34CC01030D25967F30100000C02B02";
    attribute INIT_1B of inst : label is "232032823232520204400104A798668B10FC11028CBAFEA0114670029ED2FE3D";
    attribute INIT_1C of inst : label is "0A78EF5A24BC6E930D0D10402032C320EC4A2C458A8D5406EC19E94100801669";
    attribute INIT_1D of inst : label is "0000000054000000E2000000000200000014204404AD120482E8110842108421";
    attribute INIT_1E of inst : label is "3605E90BAC185C70E5656D284000000488A0A003FED2B5BF001F644F4603930D";
    attribute INIT_1F of inst : label is "FFFC32C8F9764B4AF9AB8889161222B8AC5A1681AA680632A8755570AA7424E5";
    attribute INIT_20 of inst : label is "7BF7A77B4826D648F836A54A89FFC719E08ED558FD7FC8763CABA0288D3AA281";
    attribute INIT_21 of inst : label is "994F3A2F708DAA1734B67BED3EE806D34DB687E687CB6FC2D77BEBD03C25B01E";
    attribute INIT_22 of inst : label is "75537FC410400154D0D151EA3B56A3D92E0B48F8B7CFC9E23418CA7F49226965";
    attribute INIT_23 of inst : label is "C9DC67004569C57DC8E3861C248D9BA9E0888AF75D71749C679F44EAA312E843";
    attribute INIT_24 of inst : label is "C40C0048EF0681103A36F19F8CFAE300304038400C000E1003000364BAD5A573";
    attribute INIT_25 of inst : label is "716E254B123DB4AA403695E4CDA07F3FDCF4FE196E9E0F6E87C0E8012A3517C6";
    attribute INIT_26 of inst : label is "7BAB3B0CD8273514654040B8B6736B4A0D20DD01216F54B0D0870C1742121A69";
    attribute INIT_27 of inst : label is "64433292727D3EFCE6BCAEC1BFF72B63001D74F6020AF470A5AA916ACAF5F1DE";
    attribute INIT_28 of inst : label is "2B1CA28A551C6D442D924980EB25D92062821141095000205A89071852840D93";
    attribute INIT_29 of inst : label is "9433C2259EE8763B7A99499840F1129331F81E11D5637ED3D00C17CDFF008049";
    attribute INIT_2A of inst : label is "6C3DD3ECF742DBDB390CAA1E51F95B7BDE0D6DDD8AA6FA4C6FCE2A99EA4C57E6";
    attribute INIT_2B of inst : label is "0000FFBBB3BDEBDDDCF1F7FD488BF2D13277D6260DBBAEF5C357AFBC99DFFBF1";
    attribute INIT_2C of inst : label is "7128C632EEFDB8992AB2376948CC666CAC92666955799999098C4D8C9999C64D";
    attribute INIT_2D of inst : label is "0E574E3675B6E694668474AF6BD92ADB6EF0DD4CB446D282EF8C9E71933D2BCC";
    attribute INIT_2E of inst : label is "EA74A8FB752A2D915E7CDE8C1FBD504BBB660C139B984E26A2A262A24CA37ED1";
    attribute INIT_2F of inst : label is "2B26736CB3FE8621E770B081A7B81971813D5CA93F9E7FD19500009104F5BA7A";
    attribute INIT_30 of inst : label is "9FE89F986AD69F5124932A3A6AFFED67D457F409724DDC27100255CD0F527F22";
    attribute INIT_31 of inst : label is "2AEB23645AA133269A5000000002BB8BB88FAFF8C5BDB9C92D38DA63D2BF9FCC";
    attribute INIT_32 of inst : label is "095B0F79B2DC0B2707DE3634EFF3F4D4EEE135A55D22BFA84B926E6138B9FFAB";
    attribute INIT_33 of inst : label is "7BFC4678DD398B028B4FF84FC72A3F068D28EFE1370CF319AF9A180D045E687D";
    attribute INIT_34 of inst : label is "A0083522E19CE0F7309A17786664131F5BA49620255777D1D19C7BB8451C43BB";
    attribute INIT_35 of inst : label is "BCA9ECC46657CD2B4750AA755CDC6B0EB1E19CA8AF725DEC273D30005403632C";
    attribute INIT_36 of inst : label is "EFD2B1D2AC71844E35A3D956A09D722C404F81BBB09F8B335514BA49659BCA20";
    attribute INIT_37 of inst : label is "B274C99A00140C99895A5990301F259E503B567D5FCF64F3BE3CFB767E000CEC";
    attribute INIT_38 of inst : label is "73AAF24D3751684351162623A6D5F3DA164CC4D05E44203345E57F4ADA2D29F1";
    attribute INIT_39 of inst : label is "DBDF4A66944FEE7F73E111D1D12F2599953004C8908182935429FCFECF9ACE7C";
    attribute INIT_3A of inst : label is "A3A3A27474744A515BCDE97CDE9FCC695BE6F4A752114428EEB6A6B6A797A540";
    attribute INIT_3B of inst : label is "F0046400FF8E38E38E38FF5C3C0A5A952C03FFE2AAFB52D2FFFFFFF82BFBE7A3";
    attribute INIT_3C of inst : label is "030CAA209154C300030C551022A8C3000304AAA01554C3000300551022A8C300";
    attribute INIT_3D of inst : label is "9BFFD7FF4F7D51C4A5001FF4400C540AA00CB414803580AF625FFFFD0177E500";
    attribute INIT_3E of inst : label is "000AFEAA5D545C5A55A1B0A42A962DFCFF7577FABF7577FFFF7577FABF7577FF";
    attribute INIT_3F of inst : label is "7F8000E03003C0383FC7FFC1F9FFE307882DDD5510A4F55745FE195D488527D2";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A480EAC280DD640080263924B2C96C90016CC03D91B5A32013FBCD6603636BD3";
    attribute INIT_01 of inst : label is "6400615610D5FA3944364C9B2D5143EAAE9FE14B6405A52B5A83597D393D67CB";
    attribute INIT_02 of inst : label is "4D17E8104A28E0228F0030ABD7019C420C06030CCA5306031F8502F9012225BC";
    attribute INIT_03 of inst : label is "B2405B74058EE5E07ABFAA00496000CDF89FC6B8C908800548000735662AF04E";
    attribute INIT_04 of inst : label is "862D9050B4EE2C0160AC013DB6644885AC7A8B16F01A855B41300868EB9A0050";
    attribute INIT_05 of inst : label is "27164A2D02D76622DDF04E00E8001D59845DB2BCF468AA84B405010400A28A46";
    attribute INIT_06 of inst : label is "D59785D26A604788D4B56DA2004D14D84DB68A0BD51B2A9C599832ED0607840D";
    attribute INIT_07 of inst : label is "BCF36A71645925D189B25DF04E05549680E63AE14A0907F80E06E52FFD2C85D2";
    attribute INIT_08 of inst : label is "B7297D25E74BA7FBC1983362683C97B8AB2146E1C8F734BB0E112038C02796AC";
    attribute INIT_09 of inst : label is "AA92C6EB2C7E0B90F0D2B6E47AD45F5AA8A07BF426FD0DB5EC1FEBF9E9EB8164";
    attribute INIT_0A of inst : label is "677385ECA40002F651392CA91EB695AAB0855FA723523B26B6B542C70F12AA86";
    attribute INIT_0B of inst : label is "0110004E100004400178452A93EFDF7274A04C435AEFA3FDFBE8D83F23F9F527";
    attribute INIT_0C of inst : label is "9C9AC883DF781CA74802204C592B3B8D08965A0B3DA11653A2CF3BA4ACED9D00";
    attribute INIT_0D of inst : label is "B2D16D424CB2C2F9743200208BD1200208BD11CCDE3C50AB0847462A63AF4F86";
    attribute INIT_0E of inst : label is "44C9AF142AFDB95E9092E6ADB6D171464910BD23F63D222DBBD3471E9252B6CC";
    attribute INIT_0F of inst : label is "A25E7A18C8B6EF4D84E3D240E50C617622A90540542E880054BFC5E32E4800E2";
    attribute INIT_10 of inst : label is "4079E3A31100F7D1665B66464A87EA2BB42622A8008211188AA00208457337A8";
    attribute INIT_11 of inst : label is "22142FAF7A81F03E9A108252FC968284E221388B65689FFFB23B8204CDA10E08";
    attribute INIT_12 of inst : label is "74E3D4A285CB57AF6A75CCB9484621A294FB3FC49B38C45D291DAA90CC435B72";
    attribute INIT_13 of inst : label is "AD6AB1595634D765D7FD8D4175501501111105B6A814ED5A80000058BD234D5B";
    attribute INIT_14 of inst : label is "D64F4A47B56D794CF3C8C4DD03D1E47EE3F23FD378F62D51F91EFBB868FEFF6D";
    attribute INIT_15 of inst : label is "7749CD6F4154DCDF512281DEFD2905DFFF7F1F8C4D485BD6D5509EAC2CE9BBDA";
    attribute INIT_16 of inst : label is "4A1B9533BB15566118A0ED258369665E6DAF5DEDCA729EACFC7FC9979CBDADBC";
    attribute INIT_17 of inst : label is "51225E6B54B02F2111622CF3A39DC6F9927B114471B108ADBD9A78897672504C";
    attribute INIT_18 of inst : label is "20C8C9495CEF7295C3CF3CCC919B9CC5A0524A48C359E642CE36A5ED6C5C8BA8";
    attribute INIT_19 of inst : label is "0D3BFF3FD0CB26221B2CC186ADBC20CB1F2CD86E143A20CE234E14E840D83BB2";
    attribute INIT_1A of inst : label is "DE315720857211C628E40572123098668D1EC45551F17EA8FE54AE4292845E7D";
    attribute INIT_1B of inst : label is "86B2FBB044C04B6521E525B26FAA2E1AB444555118CFF3C233887A498B61A3E0";
    attribute INIT_1C of inst : label is "BD1B208FC9B8A1874345821EE4A5CA72BC944788F3929C992E583FF7F04B6E20";
    attribute INIT_1D of inst : label is "00000005401C0000FC3E0000003DFFFC0022E56092E19EA7AB1C8F7F5BD6DEF7";
    attribute INIT_1E of inst : label is "4EAD985B2A9A038F09B986649FFFBFF7330F0F03AF467B57EF53A89FD38F3874";
    attribute INIT_1F of inst : label is "FFED10FFE2EADD190F4F1CFC3F290018045705C1775C000E1AB031B418B0622E";
    attribute INIT_20 of inst : label is "2E7FABFE6B29492BAA31158CB50011231AD81F92081FCFAA8970964EDE2396BA";
    attribute INIT_21 of inst : label is "25D1BF1163D31C8D3FE8C4DA502AA03CA2482FD080031E85CF2273F8807FC440";
    attribute INIT_22 of inst : label is "3FE7B2A0120000200C5AEA35702094126A4C777DF00C462525C84E101B680214";
    attribute INIT_23 of inst : label is "AD14AF00E15D40FBCAE41520AC4893D83AA0A05F5F6291882FFE2DFB995C6DD9";
    attribute INIT_24 of inst : label is "76F3F52B1F49CED9BD12C07E03E5E2BFB01FD80FFC07FE13FB09FDC87400876A";
    attribute INIT_25 of inst : label is "CEF9DFF7FD7FD1991B6A325C11AC8CC01157FE5BC4008BA12FC5132A536FBFCD";
    attribute INIT_26 of inst : label is "B5D01F62A7DFD62B45E52BF1191D3D991DC97C1600AA7361442360D93084A2B7";
    attribute INIT_27 of inst : label is "2CF755A9B13DDACB4ED1965A033EB5F5002F91AE0ADB7FEEEFCFE7D16E3DD8AB";
    attribute INIT_28 of inst : label is "CF6D43CF69AED26B7CB6F52D299226D4E4D933CD189AD295FB9888A7ADCB265D";
    attribute INIT_29 of inst : label is "E137B6AC6DD4F339F1AB183A03F7567077FBD783BDFC29C9C4043818FEB5FED9";
    attribute INIT_2A of inst : label is "C66F36017FEF4B2E9DBF532F7FE0E91FCDDFA5BA57C7FC18A4015F1FFC189201";
    attribute INIT_2B of inst : label is "0000FF6BC73188BAF5A8633C17A465283600E913A689533AE9FCDE403BCC9F7D";
    attribute INIT_2C of inst : label is "46DC56FD4EAA13968B5E1FC5F4EAE86BEF58EADCFFCE78B19D1B00F1AE142F71";
    attribute INIT_2D of inst : label is "E5B81D09708B5B330261C9E77630E36F311B46D368884643C592069D084665DD";
    attribute INIT_2E of inst : label is "B18B97E3B8C45006270751EBD79F55560770128848422020C4C4AC4421E68C28";
    attribute INIT_2F of inst : label is "7745A52023FC0A5C009DDDEAC28EA002AA1B95747E04FF826A0000063A6D48D1";
    attribute INIT_30 of inst : label is "BFFCD7A3D4BB6CE34C0A0CCC04BFC48123ABC1AAC8A401107255395475E8FC04";
    attribute INIT_31 of inst : label is "C5B04388E880E4CAECC8000000010671A99673CD6E4847824847909D3D1FA696";
    attribute INIT_32 of inst : label is "FBE552B3F4015500A9AFCF51BFD7F325218886CCB46C5E15564521088116FF0C";
    attribute INIT_33 of inst : label is "10AABF3DEA17E027371FFFDFEF508359294D218886A2015E4438A2DAEBE0E292";
    attribute INIT_34 of inst : label is "D2915AB4D539CE904443480CFFF28856D48D06455D3B84662539480214AA1B75";
    attribute INIT_35 of inst : label is "5190F5088988F665E9EFAC8081FAE7516D80F81316B4540110563010E8E5747B";
    attribute INIT_36 of inst : label is "76664F66419D211C4CC0EA62C4A64E50BA863FB0D445E437091A0DA0553D1900";
    attribute INIT_37 of inst : label is "19A8D838001565BB41023C4025AF6928C8FD28938FD3AA95C4F17E6DE0000175";
    attribute INIT_38 of inst : label is "B6355C34CD8F6210626ADEE4CB0C214AAADDA000E8D26E360E8CA1990AC66538";
    attribute INIT_39 of inst : label is "2A4199EA3347C3C3548CBF4767E0E3C47AE5AFF488980000AAB33190962FA6C2";
    attribute INIT_3A of inst : label is "33333226666644C1753BDF13BDF13ADFE89DEF857E7DDD3EEE9E9E8E8F676D60";
    attribute INIT_3B of inst : label is "F7FD5000FF8000000000FF60350C0CE60C0200E7FFF99CE0FFFFFFF6AA346933";
    attribute INIT_3C of inst : label is "5659FFFFEEAAAAAAABAEFFFFFFFDD7555555555FFFFE69AAA8AAAAEFDD551455";
    attribute INIT_3D of inst : label is "DEAAA3FE8A021096000001FFF002AA800AB41FF7C01FF000A2000002C1555FFF";
    attribute INIT_3E of inst : label is "00000155F7FFF7FAAAF0FC80556A02A8FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03803C0383F87FFC1F9FFE307D300A0005F138AAA1000DB7DE76FB0AE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B6D02A0085B16A1BA59A10000002090400207FF083A1835F81F94D7719690A81";
    attribute INIT_01 of inst : label is "62680570D0025A10412486004930C06B44554158A6C4438230F5085D1E2F01C0";
    attribute INIT_02 of inst : label is "91016801061827128E3402B83180448007430087540D43008700E9BD409AA128";
    attribute INIT_03 of inst : label is "8C641017A40B156251A2A8120030040DB89D540B544E02263A1A0004A7855407";
    attribute INIT_04 of inst : label is "81204C382523E90251E9020484400021A0518604AA0395C3444868007B1A2EAA";
    attribute INIT_05 of inst : label is "C10C3994C294A7809054070328DA05400709A2F85628EBFA86C4185001659386";
    attribute INIT_06 of inst : label is "1314F514504867A0A700FFED1FF6E925B6C9759910820AC0312A04081A813D10";
    attribute INIT_07 of inst : label is "A7945010C330C521E120505407057F50D8202AD2D281C01D0250A9AB7BA8F514";
    attribute INIT_08 of inst : label is "550C054514382FF902D65AFA030801BD3A8BC6F1C4F5140AC8003848E83CA098";
    attribute INIT_09 of inst : label is "A05AA4A1AA4A87E4F14551FAE8E8522923A3A1534850D142881FE1DF51720047";
    attribute INIT_0A of inst : label is "66414DB7B0D466DBD90DB8B6D9DB36BA71105A03441218A2A42092824F00382F";
    attribute INIT_0B of inst : label is "23F148EA22148FC523E88D0498B009823690BD0A023FB2401006903F297F442F";
    attribute INIT_0C of inst : label is "5EC2E80BF7557691297204666DBDAEE48C9FE66FBF66DF5D9BEB8EF6F6B7F485";
    attribute INIT_0D of inst : label is "A2CFB77F68A2C7817B599FB37BFB99FB373FBDB67B824C9BBDF6B3B3733BCFE4";
    attribute INIT_0E of inst : label is "616EF0932648D1906CFAFFE8A8897BF339B8F591DBA8DAAAC21A05DFDB2C1448";
    attribute INIT_0F of inst : label is "CE6051AD6AAB08689CB3FB71F2CE7B837B36D67E5E2B666FB7C3FE18AF4DDED2";
    attribute INIT_10 of inst : label is "665963DDDDA8DCC106967D06B619A9A61B83FB367ECDFB8FECD9FB37EF6D9EF3";
    attribute INIT_11 of inst : label is "BBD770F36C85613E8ABEF77716A96C86D3E1B4FDB7ADCBFFDFBBC3336A318F37";
    attribute INIT_12 of inst : label is "7A120A50052497F092DE1DAD2936050A52245004838066617F96C2526C0A1B7E";
    attribute INIT_13 of inst : label is "08413C998A690A159ED80AC0A105405411110501505784891000018A69520156";
    attribute INIT_14 of inst : label is "868ED68420BB0EC2A57A668A08A15991165030A6C0A8D88B2818415796492005";
    attribute INIT_15 of inst : label is "D0950B68C4A61984DA73FC91A74AAC915A3762EAA8D552148051E486C0F8C210";
    attribute INIT_16 of inst : label is "2C41052BAC524B25A8D5A9052369449541484CA8AA51830F0821F10401214834";
    attribute INIT_17 of inst : label is "9950940330A048FAB22324BBA5DC263504135550110841297512B500543935FA";
    attribute INIT_18 of inst : label is "E040524A40E0708156AA2AC4808F58046011462C809064A8C324A9695078CFFC";
    attribute INIT_19 of inst : label is "4DF2AA2A127DB6864DF6C11429A820C84722D02207198A47BB02066002551AFF";
    attribute INIT_1A of inst : label is "A50637605AF618A0D6EC5AF61190C873E715C02370C168A0DF54B0F69A64CB21";
    attribute INIT_1B of inst : label is "E07A97A03BB00009002101242FBA040D741023704E03F0C6112212008260004C";
    attribute INIT_1C of inst : label is "190A209551B86387D3C40002A455C5D15C2645D8B980CC0F43B8046120004E28";
    attribute INIT_1D of inst : label is "000000100401B6DAE701FFFC0011FFFC0004210084C80DA1286C018843188C63";
    attribute INIT_1E of inst : label is "E02A0054284A1C70E1C1D06ADD552A8AAAAAAA003F06821CCE7BFCC4A0D6E130";
    attribute INIT_1F of inst : label is "FFE91F2AE3CE4C1A30248E781A0C2050144E1384EF38013560A2C0A160A1006F";
    attribute INIT_20 of inst : label is "3EFFAAFE0A0B6D4AAB11A442A142D23AFA8C5D68433FB82AA452047FDE3B8438";
    attribute INIT_21 of inst : label is "0C8209051241A3A20660C1E05A83E84145142FE4E902222D592053D0A875C650";
    attribute INIT_22 of inst : label is "0AA7EB2480000074DC91AD255A44A05B4A6C0CFF5068C1C12511461E124E2A55";
    attribute INIT_23 of inst : label is "11E1A2806038CB1D0CF24F126F9709B9AFFF57028200810C2B410DF0285A2D29";
    attribute INIT_24 of inst : label is "A20E150A2F52D1DA5A24C9AE4D78D23F681F944FDA27E503F281FBDF18C2AB01";
    attribute INIT_25 of inst : label is "6B0D6058162EC1A15140344C737DFDCFD747FC5BCA9F8BAEAFC57A341A2597CF";
    attribute INIT_26 of inst : label is "58924B4338E5477D286118F1BC343C1A1C097615C5A35161042B44E830A4FC80";
    attribute INIT_27 of inst : label is "1462890270443E2186C1A450B88142020002818704AAF4818C6633192CE71092";
    attribute INIT_28 of inst : label is "02205A0045004A02392485C0081649254400118E08929084788CC9294AD2285E";
    attribute INIT_29 of inst : label is "152004411000AB90C910103003062060630083A7A888A80984002819FE00008A";
    attribute INIT_2A of inst : label is "27712401C00D984183A8A3B82000A0603610CC0034C30D1F9000D30A0D1F8800";
    attribute INIT_2B of inst : label is "0000F40267421000108074414D2A1294960918456166B09618B930C030112280";
    attribute INIT_2C of inst : label is "49D5CF6150A8716A04BAAA211F9CB708C889A32055598B0A8128822028DA0839";
    attribute INIT_2D of inst : label is "A3A9981B511809356461ACC2A8CCD30683F70D1E40CC0685A2380BE481406A22";
    attribute INIT_2E of inst : label is "F0FF7CBAF866DB3330D9C1264F97D5DD2C521A8159520512EE66C666058C5764";
    attribute INIT_2F of inst : label is "7CE697F9B2A988E1CFD9F9CFBF78F377CFFDFBD4753ED507770000332DFBC8C9";
    attribute INIT_30 of inst : label is "B57D6F748269B6B5EFFC667E2FEA8371A1FFC0BBAB4C9902629F5FBF12A8EA6E";
    attribute INIT_31 of inst : label is "EFD061CCFEE0CFEC60D000000003BB58791358E10F6F6A4F6F6A5ED4AD1575D6";
    attribute INIT_32 of inst : label is "85F297836FFC78FF3F14AF51BAB6AFF5A4C8160D4A1EFE0DDD5A644811BFAA0F";
    attribute INIT_33 of inst : label is "DEB1C3CDF202C2279C1AA45A967B6D6DA565A4C81403F0A7E83CF105BC60F3CA";
    attribute INIT_34 of inst : label is "12FB7C1684A5B252E40A2450888E8467BC8FFCF9F23D4777F4A5297210B43489";
    attribute INIT_35 of inst : label is "41A17F8EDFDE306B2F31C6FFDC3014DC464137FFFF5E44B902632030FDFF1790";
    attribute INIT_36 of inst : label is "A906A4068564A15AF396FF7C797F78F9E3FF2221740E8696140DB659798C1A00";
    attribute INIT_37 of inst : label is "0A02580A0001421480433D00380829A0D081DDFA8ABBFE46B36ECB04D20001FF";
    attribute INIT_38 of inst : label is "842FAC34CF810214773C1C2809150050B50A430960D4AA96160D049A02926A10";
    attribute INIT_39 of inst : label is "17401A88358FC3A277C00151718033D0143803A2BB2220800002391E1C690084";
    attribute INIT_3A of inst : label is "484848890909048129D1001D1001D080B0E8800660215033A4ACACACAC1C0540";
    attribute INIT_3B of inst : label is "F000833FFF8000000000FF7E3D0C83CA4C0200E555F87964FFFFFFF881162C48";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "21555C015F55FA29555554000A95555555514002954005554855555514000000";
    attribute INIT_3E of inst : label is "0000000000000005555A01FAFFFF5557FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03003C0383FC7FFC1F9FFE3074CFF555553731999100068EC647279BA";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "924488E0854024AF76D20822820820D4410C5410826BC16801FE64D6D87889E1";
    attribute INIT_01 of inst : label is "28225067448048026804948001A280505444505B0FC60A0210940140252C200A";
    attribute INIT_02 of inst : label is "404920A0545101400211283330806004151100D5086C1100F10BA5A41450A800";
    attribute INIT_03 of inst : label is "B0FE105308C95962C19284000330044484F5B8CD5CD7836A30A8A82601255529";
    attribute INIT_04 of inst : label is "014668A0042A6D0130ED01029F260441451D14203895419D0102A24070081C01";
    attribute INIT_05 of inst : label is "8828AD5686D201240055291B2088911D024101404E205000BFC40B048430C282";
    attribute INIT_06 of inst : label is "1A1249E21A82EA009C2EB6DB0DB65B6697EDBEF40811A960A00A12080C281042";
    attribute INIT_07 of inst : label is "92231A828BA2848848059855291A0017FC045A3852A4420C50742125482649E3";
    attribute INIT_08 of inst : label is "5F2295922A752A1CAAD75ABEDF8E1C9E11EA0263A96E3DC9F4448808629118D0";
    attribute INIT_09 of inst : label is "28407241272CB76540C55D9AB06973AD3B49A87EF81D9866E60DF182713D5047";
    attribute INIT_0A of inst : label is "CEAB57B239F06BD9DB649C926ACBC234C11A53853498296C9DA63508D400546A";
    attribute INIT_0B of inst : label is "62C318B823318B0C62A08F708A139894A73DD00A63279B0310B62C1F132A68D0";
    attribute INIT_0C of inst : label is "46C22A217757F73473FC07332CACCC69F74DBB2696724D08C9A1FE32B332F9CC";
    attribute INIT_0D of inst : label is "AA66DBA9AAA27315198C89113709C89113F09872738A9D3EC721919153D8E7C3";
    attribute INIT_0E of inst : label is "D16C62A74F4AD88726489ED1049D189996CF6B9D098E4CC6CECA59B86F2764AC";
    attribute INIT_0F of inst : label is "95A51CC6331B3B294A3F0DF6B2631491191262B747233234AE55924C83066430";
    attribute INIT_10 of inst : label is "234D22CC88A25A63A2D55882F3B787DE49D119122444C9C664489113271C9CE5";
    attribute INIT_11 of inst : label is "CB6692304C6A804085CA592922EDB6C6D0D1A07EFA9E4E04CCB8F11923188B12";
    attribute INIT_12 of inst : label is "B254E808028016120262520E73B80538C724D6806DC0222961B0DCE7300AF84D";
    attribute INIT_13 of inst : label is "69CC0E13626F9B90394100D2235405404444500848D0018310000E8962027148";
    attribute INIT_14 of inst : label is "9916042DA6238AD204922229801020D1219C119808142890CE88CC490C240015";
    attribute INIT_15 of inst : label is "9890A443136C0B6258152695AC1036944053AE2439814ED69A6C42D52448DEF2";
    attribute INIT_16 of inst : label is "259B39A8314862B4645D4C0CC3AB32120C3526A2A09D0B16682528CA23652947";
    attribute INIT_17 of inst : label is "01107300B090820B2566360810503644821D451118084E2549D685E1984FA796";
    attribute INIT_18 of inst : label is "E14C48C101E7129D00B30FC718812A836A1168B6054C60A46304EF2D30214666";
    attribute INIT_19 of inst : label is "48FBFF0E77AD9806F7B30414A54E309987922890255D8F4D591024622528435D";
    attribute INIT_1A of inst : label is "CDA3A6828CA811B464D00CA8198144B0601D615240C1693C5E308228CCDF6A34";
    attribute INIT_1B of inst : label is "766AE6383FE400010129A800011034DB58595A400DC2F8A8A3023068D590206A";
    attribute INIT_1C of inst : label is "0A61E1413886404A0205041220D8CD0342A514B294D4A0D6F32C8C6900020922";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000010A9401145401003D6AB5ED6BD8421";
    attribute INIT_1E of inst : label is "389430282D4500000E0E2A2C5FFFBFFFBBAFAF015182D2EEAC4E646410C3A1B8";
    attribute INIT_1F of inst : label is "FFF0150BF5CFF60BF0038E4A19190340D00601806718050080E100E080E10073";
    attribute INIT_20 of inst : label is "2B67E4794124AD7352B1B9A91942D3B183B871A6413FCA82991A847B8C919210";
    attribute INIT_21 of inst : label is "00A3844E6711B0AD83144BD24CE02924D34D042F504414942A8F03D8C966A16A";
    attribute INIT_22 of inst : label is "233300000000019EB722A104327131C9555A4CFD3050B37589DC258B88029A19";
    attribute INIT_23 of inst : label is "C388E6004618441908C1450A2C02218880AAAAAA2AB0940A333E0428863D9CBD";
    attribute INIT_24 of inst : label is "AA5AD4398F189B7B53FD680F4072C13F601FB00FC807E403F201FBE8129A1140";
    attribute INIT_25 of inst : label is "2B45699A67A560BBE11C17203E5F1CE25390BF3133D3E90DEBD11AB6147557A1";
    attribute INIT_26 of inst : label is "029F490520C1C118F863083AE636068B1A01829402D4B101D00900CB60233052";
    attribute INIT_27 of inst : label is "567EE95BC340E4268460B84572D9D5D70024F8D808C9779C42050281814A0029";
    attribute INIT_28 of inst : label is "184068734B316B922059810BC6034926460019884EE2118C18CA8D294A63381C";
    attribute INIT_29 of inst : label is "5C264C4DB81C008069134092034626C12740C085D5555490800C0F8DFF0E208C";
    attribute INIT_2A of inst : label is "BB3271E0CCDFD575E792D999041839E67B33E80302350F08C7C408D20F08C3E3";
    attribute INIT_2B of inst : label is "0000F9B5F294210318C09F652C00DA00822DAEAAFFFF1FE3DF2FF03C133DE38E";
    attribute INIT_2C of inst : label is "97D690F3AAFDB111BBB6621B19999B13EC6C24C4AAA1C9C99AEC7766FB09992A";
    attribute INIT_2D of inst : label is "FD0F8BB34F152C17D6C026502143B5AA528B819D5D4582C4EB2C18FB81B82E01";
    attribute INIT_2E of inst : label is "4AC60D1AC56259911C48CA1F3FB7FFDF98A62B01D3DC0696AAAA42220605B2F4";
    attribute INIT_2F of inst : label is "5C24364C93FC8425657377BB671CB9558FA4C99C299A2AF5110000912C98FC6E";
    attribute INIT_30 of inst : label is "8A8C7FF6B24EFAF4E6D5222AAB557DB29C67C0FBFA59DE0342964C9D0738532B";
    attribute INIT_31 of inst : label is "224EA056B221C22C745800000002A95915915829696564C1656CCADBC8BFF461";
    attribute INIT_32 of inst : label is "153A99C1364B5A252C1248F0AFF3F8BBCEF01B4582433E0FDFD2CEF0188955F2";
    attribute INIT_33 of inst : label is "5B3648C131AD0035AC0550C55B19B6379CF5CEF0198490D17B9D3414C4DE74F8";
    attribute INIT_34 of inst : label is "921B8DD7339EE5E7380AC140888701098F87D4ADE93DE351139EF3BC12941E8E";
    attribute INIT_35 of inst : label is "20BA4CD444473A2C2C2D4AA5561702595E00DECAAEBF49DE03256833CCC61696";
    attribute INIT_36 of inst : label is "A4A2C0A2CCDBC06EA023995420755D5D43E9871BB80E8382140CDF6FA2C60B20";
    attribute INIT_37 of inst : label is "C61608E600100250861750006170A690580A47C85FFE65E2A13A0A1A7C000ACC";
    attribute INIT_38 of inst : label is "E165AA2CBA52A8051114103B4455B1B81D284186B0574F823B05D20B80E82C90";
    attribute INIT_39 of inst : label is "91CE0B0417B83C8A26604591D1437500936170C6020202A185488C4429316D2C";
    attribute INIT_3A of inst : label is "3F3B3E2767E762402E54B5A55B5A54352D2A5AC0292E6314462E2A2E2AE2D720";
    attribute INIT_3B of inst : label is "F000033FFF8000000000FF7AB10C803E4C0200E555F807E4FFFFFFF0AA850B3B";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "015554015F555000000000000015555555500002800005554055555500000000";
    attribute INIT_3E of inst : label is "5555555555555555555000AAFFFF5555FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03803C0383F87FFC1F9FFE3073D11111114A7A5A5055147E94F8285AE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "2490381AA55504A6D36A132CBA936DD8518E9560A2A5802A8AF96C444D6D71EA";
    attribute INIT_01 of inst : label is "804813E09021701340125A2DA5451011414050412035146B5AA2452061B06419";
    attribute INIT_02 of inst : label is "690DC00908A28A02082409F0100013811A40001AD423400034014AAB40582ED8";
    attribute INIT_03 of inst : label is "1218D92480B10F2C44B61E0925800A4C049190A208DC53EE9A12001406876830";
    attribute INIT_04 of inst : label is "0385514594A4CE05604E0516910C4885061A28BB62074F82042A5811C9101644";
    attribute INIT_05 of inst : label is "14514AA5146206876968302F61D20700450583307840510110001C8301A68A84";
    attribute INIT_06 of inst : label is "9462B0C61808BC111B074DA61B49B4984892012897C2259145B48C2812846D01";
    attribute INIT_07 of inst : label is "1507184515451881A2D609683028222203F101614B04093108E245442145A086";
    attribute INIT_08 of inst : label is "A4204A452048B5B0035E6B94C24D30082035103595E479B120608128886A34A3";
    attribute INIT_09 of inst : label is "019FC089F40891FF8707E41F403C8010AC80807E401B942C02981D0127600156";
    attribute INIT_0A of inst : label is "F6001636B3F2CB1B9A6DB2D6FCC9C6304111534C625463CD18C45E017820A8B4";
    attribute INIT_0B of inst : label is "E40F390022F3903CE4008A629E32A99BC617A08C52A84F40226AC430554126B4";
    attribute INIT_0C of inst : label is "970AFD7C802A86182FA845767DCDACC0B3999E6CB1A6D9669B2C3B3736B7D0BC";
    attribute INIT_0D of inst : label is "EFCFFE63FBEF5B119B19BB77ED199BB77ED1982675060C15AC60B77731FBEC6A";
    attribute INIT_0E of inst : label is "EB705183046AD9C26DD8B2E1051399F33C9A5BED598CDA52D47451A8EBCD78FF";
    attribute INIT_0F of inst : label is "0D66198C694B51D13A351D68FCC635973776CEE156AB66EDC26BC65AA90CCC11";
    attribute INIT_10 of inst : label is "EE79A6DFBBD79A4100707100527901141B47B776EDDF999CDDDBB77E66099D43";
    attribute INIT_11 of inst : label is "261CB2B3ECB80080D61983CB37BFFF44C411313FDA9CC400DC04C373E1F19B7E";
    attribute INIT_12 of inst : label is "BA70D10004085A330BC66ECC2FE8462842A392279DA26665A5D2C05F908C5C5A";
    attribute INIT_13 of inst : label is "318998D5CDF93055A2480EC0D145110450504199D84130E110000312A944458A";
    attribute INIT_14 of inst : label is "12A6D6A8C4D9344AB5B666E30C307117705203B41838CBB82901D9DC920DB6CA";
    attribute INIT_15 of inst : label is "D370016300E100E65C376C529D5A14522180282A91D18C63114F3608D002D463";
    attribute INIT_16 of inst : label is "6075B038399144B9A08E0888A02A24A2082044C8EA12294640360D0002463175";
    attribute INIT_17 of inst : label is "4132620331110113C64B28D0169126A59651186451BB5884E08A74A92266D368";
    attribute INIT_18 of inst : label is "2849924AD2E9153640E38D58311948066053706404016664CB32C72E2879CEEC";
    attribute INIT_19 of inst : label is "498000846FC49845FA930C18C50C00A948388028969E8A4AA908976002040A02";
    attribute INIT_1A of inst : label is "E8BB1492EE49039770906C480BD8681A7408A751C8C16838E122B3EED8774CBC";
    attribute INIT_1B of inst : label is "D70AE0B833A42DB501A5AEDB669833D3004751C9EFFC0F3022F6306D7B91BF62";
    attribute INIT_1C of inst : label is "7DDFE5753982F0810300419A40E02E0B8094B686F01280D9A3947FED904B2D08";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000002C510144C6DDB70E6873DEE7BFDFF";
    attribute INIT_1E of inst : label is "28AA145411E81C70E0001004C0000000445050037100727ABDDAECD41CF2E1B0";
    attribute INIT_1F of inst : label is "FFE80833E707E40102728F000B0B250943D8F63D8060048B1206250512058441";
    attribute INIT_20 of inst : label is "40C04400210DE021FF1410A4124480A0853001A6101FC022A052956EC1851330";
    attribute INIT_21 of inst : label is "8AB3DC01A7041B8FD900081642720F2CB2CB10265521109428A48019F30611F7";
    attribute INIT_22 of inst : label is "0AB74B200004118B04026515002212D8C50195041244E8D29098B756D24E0900";
    attribute INIT_23 of inst : label is "3D3D1BD88961C8BA56B53CA9E3909ED01A2222202226DF131434402A2D5F67B7";
    attribute INIT_24 of inst : label is "2A423471708F08590324645F22E5F800FDC07EC03F601FB00FD8051355180D02";
    attribute INIT_25 of inst : label is "638C7A1CC668401091C802E4D76B2F549D1A00A035648C71302B56F6D04E7811";
    attribute INIT_26 of inst : label is "18DCCE033CF1A33420E72903D02C34011E09441529B61621749A05E9F264BC86";
    attribute INIT_27 of inst : label is "1AF4CD69A120D0238840142659080A020022F99808D1079E084422112D128040";
    attribute INIT_28 of inst : label is "006150418A20930A510402C1C022B6DCAC492BD8538A539C8152FAB5BD4B689E";
    attribute INIT_29 of inst : label is "080524CA400620D01133D103022667A20722EA058280A88108002804FE251292";
    attribute INIT_2A of inst : label is "4A1324000A4C2012A50029010620A4A5241210005315E40380014C57D4038001";
    attribute INIT_2B of inst : label is "3EEEF480004210002100241255682442D0126D98F04498031C2841000290448A";
    attribute INIT_2C of inst : label is "7E817FF40057E141414A5F504A5A50FAE942A055AABEA1F4B452F5E1450F0F85";
    attribute INIT_2D of inst : label is "102881F55C101802B3E4084556AA9100802B0A9849CF0048B9387AC091000400";
    attribute INIT_2E of inst : label is "CACD1A3CC5665B3338D8C5140FC2281A061E2A110F88459EEEEE466644C4ED0E";
    attribute INIT_2F of inst : label is "DE225ED9F0038924CCCF6B4B8D36B3330B6CD9D4063600733B23C8336DB9C026";
    attribute INIT_30 of inst : label is "000348389FE8963861B86EE6D6C03B719CCFFF034137F4224FF78D9C8BA80C67";
    attribute INIT_31 of inst : label is "67CE61DFB660CE6D6008000000019F3A377F3E77A9FCF949FCF979E0E0A03CC9";
    attribute INIT_32 of inst : label is "18791BB006DB5E6CAD21C8B1E0200AD1BFA1120088C67FF01A09BFA111BD00E6";
    attribute INIT_33 of inst : label is "30EECA0FB2F801B5BC4000A018BBFC369475BF211083F125BBB53C9F8CFED4E0";
    attribute INIT_34 of inst : label is "5E5DAC561094B95F908C704CDDD210439C81B875783C5673B094AFC852E02001";
    attribute INIT_35 of inst : label is "40135D9CDCCC30062E39CEEDDD328C5E4E2197DBBFEE67E422674010CED79712";
    attribute INIT_36 of inst : label is "B90072007CB0840AFB56BB7C33333058E2DB050FE0886ED80013049241440100";
    attribute INIT_37 of inst : label is "480B4048001901200445E080582C4B200808ECDC501AEC463A2C8D8C54FFF3DD";
    attribute INIT_38 of inst : label is "E56DEE7DE6533E4C333C5C50080A564C80900206200307D83200840108500600";
    attribute INIT_39 of inst : label is "435E191802B8380EEEC4A22262C1DE08E3D82986002201230892BB5F3D392CA8";
    attribute INIT_3A of inst : label is "A1A1A434B43402C0AC17358163581734AC0B1A8229688B04800C0C0808E0DA20";
    attribute INIT_3B of inst : label is "F000073FFF8E38E38E38FF0738C38001CC0200E000F8001CFFFFFFFAAF56ADA5";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "015554015F555000000000000015555555500002800005554055555500000000";
    attribute INIT_3E of inst : label is "5555555555555555555000AAFFFF5555FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03003C0383FC7FFC1F9FFE30757EBEBEBEAA2FF0055454017AFFD55AB";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B6D24C5A9B546640412911A69A4924DC0626FA40C42188318BFE82666BEB618B";
    attribute INIT_01 of inst : label is "A4E92042F24B285144924E6DA5410144540144499025040EF2872D2320112509";
    attribute INIT_02 of inst : label is "012CA1172820802432F49021490090924F4A010F5CF54A0131676A254E0F26D1";
    attribute INIT_03 of inst : label is "9910C93794AD0533245A00000120042025B894A80E0B6504BA5A44944B933C08";
    attribute INIT_04 of inst : label is "3365104094A60740E207489090856A9525CA081B524801090CA969258068C144";
    attribute INIT_05 of inst : label is "041042210C424B936B3C0808B27A49889F2D4C412D6144109000082800A68A8B";
    attribute INIT_06 of inst : label is "8402FCF7C9C9260633242000090000490012490814CAC110409E01293A943529";
    attribute INIT_07 of inst : label is "1752C94104410096E6D2CB3C08428012023348614B82837D282265C42144ECB6";
    attribute INIT_08 of inst : label is "ED6C4C852868A09611CE39B44A0C141D34AF0877A5683881F0C05228E9389420";
    attribute INIT_09 of inst : label is "0C68690E8690D244C0181092E3015118AB8D992ECA4FB32250C215423DBC2B57";
    attribute INIT_0A of inst : label is "0F0436A62480CB53D6292B948012442C03614905225329471084F23BCC45FDEE";
    attribute INIT_0B of inst : label is "08090200EC9020240803B62292020810A4042030508063197668408071123480";
    attribute INIT_0C of inst : label is "808A4A280A0234000820997669A988D044181E6C25A6D8429B097BA6A6269024";
    attribute INIT_0D of inst : label is "AA0925485BEE3217D21112225511112225D116144A4E85492848222221AD401E";
    attribute INIT_0E of inst : label is "524803A1522AC9364A94409B6F1FD1222C121D0510A4938288C071688208388A";
    attribute INIT_0F of inst : label is "490749084E0A2301D62D104AA08424122224944164B244493480105222488902";
    attribute INIT_10 of inst : label is "4428A691112A56C530442910729411451202A224488951088891222545851292";
    attribute INIT_11 of inst : label is "2A5483ACEAA20C109D129248219248D494B5252024A884029486822253A11A24";
    attribute INIT_12 of inst : label is "B9365024941052020A40424808008828088696EC152044452110881041105C21";
    attribute INIT_13 of inst : label is "6118A05546AB094004F0BAC8E114514555005501D82080002000031A8548550A";
    attribute INIT_14 of inst : label is "12A75E9184E1384835A444A10031681768A0833018B40BB450C199DA490DB6DC";
    attribute INIT_15 of inst : label is "00CA50191FE2088454B36CD3B57A64D2611424AEF3D388C6135C2C1D822AC8C6";
    attribute INIT_16 of inst : label is "6C41301811534EB565450830A06426C6DB61846C6B4207D7249301C0CF0C63A2";
    attribute INIT_17 of inst : label is "47324636B2120C54078CA4647368DE54925B28A22C994AA4C48A54A9AA520800";
    attribute INIT_18 of inst : label is "E749DB6B9DEEB634E869044D9199DC5C6453526C4A0892684592852438508AA8";
    attribute INIT_19 of inst : label is "5012AA045001201A00241020848420A96822A16816B8964BBF2816E44A4496FF";
    attribute INIT_1A of inst : label is "A0B6AE86D8E86216D5D0DAE86BBA5D366CB5CD6B42C16822217C828C08264EA4";
    attribute INIT_1B of inst : label is "156E56922AB32DB564A7A6DB411056D558A56B42120D096BAA08036DC204D350";
    attribute INIT_1C of inst : label is "810C324A0C02D4522A2C934A6681281A129572AE5552AAD082B934ACB1692869";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000026724D5E8DF97E10E900421000010";
    attribute INIT_1E of inst : label is "51A2F145C1D9600010001304E4CB0CC000000003211072D64AD2A890B0C0C631";
    attribute INIT_1F of inst : label is "FFEA7F21E2C88C4106E00EC90F0D200803C0F03C0000000002040404020709E2";
    attribute INIT_20 of inst : label is "26886E84695B7129AADA158D955D0C44C039E8CDB4DFFFFD5EA7B57DC365B6A3";
    attribute INIT_21 of inst : label is "3EC4A8714A1A14B0A42A0C33E32A00E38E389C3FD51A774E73D69009F31250F4";
    attribute INIT_22 of inst : label is "B541D6200000134A4D321495132494105C1577043D994EE424B556765B68DA6D";
    attribute INIT_23 of inst : label is "030006180000C0180180048020000080057D7D7D7D66F12A5C756E1BB85A2657";
    attribute INIT_24 of inst : label is "6E73952130D95E5BC17FC00E0060C00021C010C0086004300218010030000100";
    attribute INIT_25 of inst : label is "4A895A54D4C944191558824533FD48C9035481E8A949A0E3601DE6F256C6C83A";
    attribute INIT_26 of inst : label is "D0DC2D1B38E5E22C11EF7B4150C444C11E692452D622D9CF45451AED15142C9E";
    attribute INIT_27 of inst : label is "1EF0CD699114CB368DCC11C60E1A9ADA0025141E8841039C8C562B1520A70981";
    attribute INIT_28 of inst : label is "7AD35AD10A30E38A698D9AC98C0A2CB6D4DB7BBE5BAA57B5A3DEE8EF2BEAF83F";
    attribute INIT_29 of inst : label is "480E65DED3B56CB6617712064142EE640C46DE31DDD75E06B00C1146FE2512BE";
    attribute INIT_2A of inst : label is "CA17760C1C8E6936AD1A69032FE34F2E6D173476347115439C18D1C225438E0F";
    attribute INIT_2B of inst : label is "3AFAFD20805AD6767399412650A94409BAD2CC8B76891B239DACCE8187148F1E";
    attribute INIT_2C of inst : label is "FFD4005FFFAAA1540155AA055AA5500542BFF005FFEA0155EAFFA01FEAF50AFF";
    attribute INIT_2D of inst : label is "AF51C38D5E21B9833A2ACEDA88CAB73C9A331D94588A10440211C6B02601073B";
    attribute INIT_2E of inst : label is "90AB56AA884452222895050307DF5DD434101226684099804444C44498C5E92A";
    attribute INIT_2F of inst : label is "D206049122A90804889B59DACA28A2228A489125042400222216D422292D4E24";
    attribute INIT_30 of inst : label is "20174028B49124A94128444484801255288BEFBA8D24204C23B58911C14A0844";
    attribute INIT_31 of inst : label is "54944089A44006646608000000011252275A565BD8495008495812B0610028AB";
    attribute INIT_32 of inst : label is "9CAD9AA84496D44B6A71C994502C092521826660CBC55F75D469218261100054";
    attribute INIT_33 of inst : label is "52AC0F33AA90186D100004B008D34B690145218265F9230A5007A09C80A01EB0";
    attribute INIT_34 of inst : label is "52110894B000101081306000AAA62662D4A12C59502996222000086080A660ED";
    attribute INIT_35 of inst : label is "4C10550888AB33072B3984488906865458018111175404204C626031E8C59596";
    attribute INIT_36 of inst : label is "39306430611009005394AA2873222CD0A2920708513484B2CC002090496CC100";
    attribute INIT_37 of inst : label is "44DAEB4C00151B76CE493030192CEA2608C088908012A804D306CF9E06000155";
    attribute INIT_38 of inst : label is "CDE564164483A2A222295978698F616A91BB671B6613A6B266609CC1165306D9";
    attribute INIT_39 of inst : label is "6A604188839811B44496A34B2B051303871928048A8AA98548D2D16B15B168B9";
    attribute INIT_3A of inst : label is "25252164242428710D973759737597B74ACB9BE66F6EAB36A4C8C8C8C8F4DC20";
    attribute INIT_3B of inst : label is "F00000C0FFB1C71C71C7FF01B24F7FFFBDFFFFE000FBFFFBFFFFFFF6BE76ED25";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "015554015F555000000000000015555555500002800005554055555500000000";
    attribute INIT_3E of inst : label is "5555555555555555555000AAFFFF5555FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03803C0383F87FFC1F9FFE307AAABFEABFFF7FFAAAAAABFFFAFFFFF00";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "002921387F45729964B63C924924924448D23FCBD30DB19F98FF46E2C97994B8";
    attribute INIT_01 of inst : label is "111481090924D10C30492124906180145111050CA27D86210C194C818C419124";
    attribute INIT_02 of inst : label is "069344C48C30C18B6D0A40846D80D868B0A301F0AB5AA301CE9093A2A120924C";
    attribute INIT_03 of inst : label is "C82736804A6F6434F2B2000003100804A6CF6B35E345FF22452530439048C44B";
    attribute INIT_04 of inst : label is "481198634210511010511046CF732650D0730C491D220426223484923DD58850";
    attribute INIT_05 of inst : label is "861863318129804924C44B982445242640909A24D3041401C240008206186044";
    attribute INIT_06 of inst : label is "C62802082474A00D4890B24B0592DB2D92D92592CC900058636232840146028D";
    attribute INIT_07 of inst : label is "4028246186618A64124824C44B8280384E24301C2088E4928C19109084130208";
    attribute INIT_08 of inst : label is "A7972273871615B1CC638CD12171C629836530A3986782140E111C8094C14631";
    attribute INIT_09 of inst : label is "1AEAC718AC618BCC012002B204031CC61893C5C26D7098972D8A115E83639C8E";
    attribute INIT_0A of inst : label is "BEF1A736B890C39B188DB0B6D2DB16B2C9DC2E729D0A94104A531044401A0220";
    attribute INIT_0B of inst : label is "20890821B39082242086C8980C9868CA17BCB06D18E86724892E7A10755E8C34";
    attribute INIT_0C of inst : label is "C67020282220B7B7799827336D8DAC4D88D95F2CA9B259D6CB3A793636B6DDE4";
    attribute INIT_0D of inst : label is "C6A5B679718283CBD98CC9196159CC9196159966633078B0E625911111B9C42E";
    attribute INIT_0E of inst : label is "4364CC1E2D80A089245A5CC41043D89198D859B1593A4E2CE50D0D8ACB66C344";
    attribute INIT_0F of inst : label is "243074C638B3943409B15974B66310C11112722CF67B332DE6D6B30B838664BB";
    attribute INIT_10 of inst : label is "33C706C88882DB5B430B16630B924B2D89719113246599C4444C9196665998C9";
    attribute INIT_11 of inst : label is "FBF618B2AC61985035DE7B21935B6EC441F1106DB72ED282DF96F1996C189B92";
    attribute INIT_12 of inst : label is "3481188203C70A98E15328AF79983697F6E8D92499B02230A9D4E6F3306D352D";
    attribute INIT_13 of inst : label is "94A62F017029DC704B4F09730DFFFEBAFFFFAA6624425DBBD0000CC4E0A530A0";
    attribute INIT_14 of inst : label is "4916214A530DC34E4236221C86C08C5887D014CB60426C43E88A662324F24922";
    attribute INIT_15 of inst : label is "0DC18C04301EC28B5B116F0C4895A30C8624B2B9042C252D4C2CC4602C20E529";
    attribute INIT_16 of inst : label is "83CA00C0C70C30300424044A40BA9128209E330306AB12069068601F31D29482";
    attribute INIT_17 of inst : label is "93CDA9C2DD440F87F80FB3A87D0F0F8B6D8DCF3DCB66B6331B718B66898B6CB7";
    attribute INIT_18 of inst : label is "30662C6C6072394C6114B8306E6B2B84BB8C1B9783F72D93786C58BA842C4667";
    attribute INIT_19 of inst : label is "02E95533332DB83665B704DA52BA100CA08C1CCC607B4160418C61F3057A5300";
    attribute INIT_1A of inst : label is "3690C192435908520A32415908984C122486A50D08C169A4407EE9425EE23025";
    attribute INIT_1B of inst : label is "719119C8445464909A10924936CD0AC9803D0D0800590E6299004F2452910618";
    attribute INIT_1C of inst : label is "334AF7D5088E30C1212248211E352358D2605C0B81CC0E42C854E21341248714";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000191093C856401004B64635AD6B5AC6";
    attribute INIT_1E of inst : label is "661D1C3A46492000100024306B34B33000000000B1630B1B29DE645CC28D99B6";
    attribute INIT_1F of inst : label is "FFEC8096F12DB58C991D96002A381FF7FC3F0FC3FFFFFFFFFDFBFBFBFDFA2243";
    attribute INIT_20 of inst : label is "24A87EC794E04D94A879CA104D724633E14A0F16C97FE222BC50C8EA8B31CA04";
    attribute INIT_21 of inst : label is "48DA88870425C142800449DE8E240338E3CF68002AF59E81A7A3D031F01D70FD";
    attribute INIT_22 of inst : label is "ABA2C8800004811A18084A60F499495A04071D843A44D9884A0206DC48070482";
    attribute INIT_23 of inst : label is "FCFFF9E7FFFFBFE7FF7FF37F9FFFFE7FF02A802A8038708B386B955CC8AA3513";
    attribute INIT_24 of inst : label is "C718CF94E0E6633C3C023FF9FFDF3FC09E204F30279813CC09E604FFEFFFFEFF";
    attribute INIT_25 of inst : label is "6B6D659B263B58CE412319CC49259D32449140F2E34302E1C40F58298138F01D";
    attribute INIT_26 of inst : label is "6707922586DA11136F5AC648CF35A10C1B87D81000621A21C81220D32042B621";
    attribute INIT_27 of inst : label is "624D3092424924C8F050CE0921E36F67000E80E306340C61630582C1C2DAF03E";
    attribute INIT_28 of inst : label is "850C251CA08608610676E0247303DA4207B6C90940E00D6326409F188420641C";
    attribute INIT_29 of inst : label is "9831B6217C4CB0981D89281901BB125031B84A41A08A8A51400C2889FF91C841";
    attribute INIT_2A of inst : label is "30290018636D92C9D104900CB226A4D19258C98994530C0CA436514A0C0C9219";
    attribute INIT_2B of inst : label is "2AFFF24F72A529898C609ED99C14B62091B67EA9FB76FDDF7EC331C318FB30E3";
    attribute INIT_2C of inst : label is "002BFFAAAAAAA155540000AAA555500015555FFA000001FF55000AAABFFFA000";
    attribute INIT_2D of inst : label is "4E288C972B9A4A18464063675F30A14B25DB665B64446303658E4ACD890630C4";
    attribute INIT_2E of inst : label is "DAC58B38ED63599116D9BE6CDF8822598BF20809B99826322222222224661651";
    attribute INIT_2F of inst : label is "D923B64CB15486726467653B6492B9913B2CD9D02B97AAF111E87F91ACB9C05E";
    attribute INIT_30 of inst : label is "EAD5D8B2C6E9B6B66493222272D57B61BC47D14B365CDC131A76CD9F37A05723";
    attribute INIT_31 of inst : label is "22DE2046B2212227686000000004CB58B13B5B6D696F6EC96F66DECD95AAB2D3";
    attribute INIT_32 of inst : label is "C2B25B91564B5B25ED8A45C0957D5DB9E6E09A8634623E8A59B2E660989955F2";
    attribute INIT_33 of inst : label is "DFB6624AB18F30BD8B155675655D6D6DEE75E6E09A05B0F36C1DB242A64076CA";
    attribute INIT_34 of inst : label is "0A9D4E574DEF6EF3704D0A10888E691B9C05962F67AE71111DEF799806981F13";
    attribute INIT_35 of inst : label is "10C8CCC44445B431ADA523246598C3596100EC888E371CDC13113812AEE65659";
    attribute INIT_36 of inst : label is "C2430943244D80762CE3991764B1935C4ECBB1F9204B63912105B6592C950C20";
    attribute INIT_37 of inst : label is "332646B60010248903A5006044970088602E46DAD55E64E324D97061BC0008CC";
    attribute INIT_38 of inst : label is "923598A696D8E009111303068261E1B8064480C1A858D0910A86610CC1243120";
    attribute INIT_39 of inst : label is "B3E18C23186C3D4966F238989822500628448CFA6446668CB64D1C848E058242";
    attribute INIT_3A of inst : label is "4E4E4F09C9C9E400F2C8C8AC8C82C9C9A1646443B1322419DE666666671F2280";
    attribute INIT_3B of inst : label is "F7FFFFFFFFBFFFFFFFFFFF1FFACFFFFFFDFFFFEFFFFBFFFFFFFFFFF050D3A64E";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "015554015F555000000000000015555555500002800005554055555500000000";
    attribute INIT_3E of inst : label is "5555555555555555555000AAFFFF5555FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03003C0383FC7FFC1F9FFE30755515554000800555540000050000055";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "802020307F04629B6CB028000000000D00E07FD9CA85101F91FE0391C8789091";
    attribute INIT_01 of inst : label is "2010010100001C08200004000061801051540558A64586000035080104010100";
    attribute INIT_02 of inst : label is "0C0070800C30C3020A8800802C805800048100C4A84A8100CD40934081698008";
    attribute INIT_03 of inst : label is "8A6E92100C626032962000000330044322882C1D8345FF224424200204001C09";
    attribute INIT_04 of inst : label is "2021986100024308104308068A22044060430C001C0204078010800139181A00";
    attribute INIT_05 of inst : label is "8618633180201400001C095800040404000082201630101486400228851440C6";
    attribute INIT_06 of inst : label is "C62104144070A6010B01964B05B2DB2DB2596CB24C904058600E02100106820D";
    attribute INIT_07 of inst : label is "08344061866188010000401C09420290CE2518380180500A0C30208084020414";
    attribute INIT_08 of inst : label is "02460672021415208A1142C003208260816001830842003004300A005081A631";
    attribute INIT_09 of inst : label is "086883088820988CC10016226001488C18010504254109020482015301411A8C";
    attribute INIT_0A of inst : label is "B4A1A4129C904209080498A24A491290C5182820140B000008423228CC086C66";
    attribute INIT_0B of inst : label is "208908202B9082242080A8100EB0ED8A533C900C18C82210540C2800E5530C34";
    attribute INIT_0C of inst : label is "C2502A808282333679B8173324C4A459CCCB4F25E8B24BD2C96A3993129249E4";
    attribute INIT_0D of inst : label is "C6A4932B20828901498CC9192148CC919214886221201838E621911111108024";
    attribute INIT_0E of inst : label is "492458060F008091244B58482001489199C8CC914B224E2E441C048A59265155";
    attribute INIT_0F of inst : label is "646244C638B9107008914B20926311811112622C52293324B255160B0106643B";
    attribute INIT_10 of inst : label is "334502488882CB8A201912200B96430C89319113246488C4444C919222188859";
    attribute INIT_11 of inst : label is "CB6630118460805139CAD9630749260E22838884922660824AC2719928188992";
    attribute INIT_12 of inst : label is "2002180002820AB0415628A679B81614E6D050249CB02220ACD644F3302C25AD";
    attribute INIT_13 of inst : label is "10842E01A23088605B8D0312A50000000000002D1442C99350000C8CC0842080";
    attribute INIT_14 of inst : label is "0914210842ADAB4C2112221086A144D44D810A2B50A22A26C005151124A92486";
    attribute INIT_15 of inst : label is "88C086081000C20B4B1126000084220000A4C0C1002004250834C04420388421";
    attribute INIT_16 of inst : label is "87CA9087070822300064800840CA11204114122200CB00040001201A20C210A2";
    attribute INIT_17 of inst : label is "B344A150C5000FE7FFF0B6A865490C99248E4515412294210D508942008924B2";
    attribute INIT_18 of inst : label is "00456A62504A252C0018A014AAA232818A848A9AA1552483692448AA042C4666";
    attribute INIT_19 of inst : label is "8CCD55E0332498066493045842A230088084088C20510140620C2142056851A2";
    attribute INIT_1A of inst : label is "1610C500431000C218A04310008040302012440400C1694021C7B14274E22225";
    attribute INIT_1B of inst : label is "619219004454400058000000378C0E00B01C04000209024300004A00D0900208";
    attribute INIT_1C of inst : label is "1342F750087420830104000034350350D020640C81041806C848A00000000430";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000102002889440100098029084210842";
    attribute INIT_1E of inst : label is "2D14882944402000100022006000000FFFFFFF0190201A8B29CE645AA69995A2";
    attribute INIT_1F of inst : label is "FFE41192F165B8809489964A382A000000000000000000000000000000026161";
    attribute INIT_20 of inst : label is "1588188558A0051800388D088CB2461161040832C97FAA281C0028C883122202";
    attribute INIT_21 of inst : label is "2882804F061483A28224338A1E20011041456BC080560E08CF039C00B110785C";
    attribute INIT_22 of inst : label is "A100E1800000013A30102020AA15854A08070880384AD9A42C0146DC48008245";
    attribute INIT_23 of inst : label is "000004000000001000000800400000000A80002AAA9430041C4B4192A82A1513";
    attribute INIT_24 of inst : label is "8218CF1080D0533A700080000000003F401FA00FD007E803F401FA0000000000";
    attribute INIT_25 of inst : label is "29652DCB7213080E411101884805BD36C4B180C2A74600E0800C482082349018";
    attribute INIT_26 of inst : label is "6E870B15869D111264000048C6A890800107C83000605901C003108B00029613";
    attribute INIT_27 of inst : label is "5444A852C25964A4D4880D4169D16D2D001C005106308053630582C1C25CD42A";
    attribute INIT_28 of inst : label is "0E8A2618800448C02656C0C07B0348004600110B00C0000020019D0800006C18";
    attribute INIT_29 of inst : label is "9809B5136A2C88845D45000401BA8A0009B440018A08A051A00C0003FF01812B";
    attribute INIT_2A of inst : label is "380480001369B6D9690CB802A80004C9B6D4DB45946000041406518000040A01";
    attribute INIT_2B of inst : label is "1500F64D7094A5455AD0BADB9810B60082243A20A93274CE2AE3218004EB2AD3";
    attribute INIT_2C of inst : label is "5555555555555EAAAAAAAAAAAAAAAFFFFFFFFFFFFFFFFE000000000000005555";
    attribute INIT_2D of inst : label is "0E0082963351210046006392AB10E22B14DA2649544420066C8D4849850201A2";
    attribute INIT_2E of inst : label is "5E458B984F2349911648BECD9F8A82CB99B2180599B8163222226222142512C0";
    attribute INIT_2F of inst : label is "4963324C91548322646D2D792597999169264C800992AAD111550091A490801A";
    attribute INIT_30 of inst : label is "6A959892A24092972097222262556920B447D459724CCC0B1A7264C926041323";
    attribute INIT_31 of inst : label is "225A204792216227440000000004C949913949272B2524CB2524CA49B5EA925A";
    attribute INIT_32 of inst : label is "82925100524B4B25E5DAC1085545509CE6605C4032223EA2CB926660588B55B2";
    attribute INIT_33 of inst : label is "5B36C046118D00F489F55415414E2444CF34E6605D0490512C059002AC00164A";
    attribute INIT_34 of inst : label is "0ACD6453A9CE6CF3702C1A1000040539080092252DA5711119CE799806B40A8A";
    attribute INIT_35 of inst : label is "0808CCC44444A201A5AD23246584C34B51004C888E933CCC0B313812A6F25254";
    attribute INIT_36 of inst : label is "A620192024D980E62CE399134D91974C5A49E0D9702B63828105B24B24B88020";
    attribute INIT_37 of inst : label is "3216089600101254818530005816A1840026464AF54E66E2A4996AD13C0008CC";
    attribute INIT_38 of inst : label is "9134900612F0E0011112022E4147E1B8052A4080C41060820C40508082220090";
    attribute INIT_39 of inst : label is "B1E0802100F02DA9226031B1B122D30060D80C222220038004088C4489054222";
    attribute INIT_3A of inst : label is "4A4A4A09494940004AC5A42C5A42C5A51162D203C808021B4A222222228A9600";
    attribute INIT_3B of inst : label is "F7FFFFFFFFBFFFFFFFFFFF7E37AFFFFFFDFFFFEFFFFBFFFFFFFFFFF015C3864A";
    attribute INIT_3C of inst : label is "0208AAAAAAAAAAAAABAEFFFFFFFDD75555555555555441000000000000000000";
    attribute INIT_3D of inst : label is "015554015F555000000000000015555555500002800005554055555500000000";
    attribute INIT_3E of inst : label is "5555555555555555555000AAFFFF5555FF755550000022AAAA200000155577FF";
    attribute INIT_3F of inst : label is "7F8000E03803C0383F87FFC1F9FFE30755540000000000000015555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
