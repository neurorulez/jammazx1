library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity berzerk_speech_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of berzerk_speech_rom is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"02",X"C0",X"02",X"E0",X"03",X"00",X"04",X"60",X"05",X"20",X"06",X"40",X"07",X"C0",X"09",X"00",
		X"0A",X"40",X"0B",X"80",X"0C",X"A0",X"0D",X"60",X"0D",X"80",X"0E",X"20",X"0F",X"80",X"11",X"40",
		X"12",X"00",X"12",X"20",X"12",X"40",X"12",X"60",X"12",X"80",X"12",X"A0",X"13",X"C1",X"17",X"C1",
		X"21",X"1E",X"21",X"7F",X"1B",X"58",X"1B",X"7D",X"25",X"1F",X"1C",X"49",X"27",X"5A",X"27",X"5A",
		X"2D",X"1F",X"1F",X"58",X"20",X"DE",X"2F",X"41",X"33",X"41",X"33",X"79",X"39",X"1F",X"37",X"58",
		X"38",X"DF",X"3B",X"51",X"3B",X"78",X"39",X"1F",X"39",X"1F",X"39",X"7F",X"3D",X"49",X"41",X"1C",
		X"41",X"1C",X"40",X"D8",X"28",X"59",X"28",X"78",X"39",X"1F",X"39",X"7F",X"27",X"59",X"29",X"59",
		X"2A",X"5B",X"2A",X"78",X"49",X"1F",X"49",X"7F",X"2B",X"59",X"2C",X"DE",X"4B",X"49",X"4B",X"7C",
		X"49",X"1F",X"4E",X"58",X"41",X"1D",X"41",X"1D",X"41",X"78",X"39",X"1F",X"39",X"7F",X"4F",X"D9",
		X"50",X"58",X"50",X"78",X"39",X"1F",X"39",X"7F",X"51",X"51",X"51",X"78",X"21",X"1E",X"21",X"7F",
		X"53",X"59",X"2C",X"DE",X"39",X"1F",X"54",X"59",X"41",X"1D",X"41",X"1D",X"41",X"78",X"39",X"1F",
		X"39",X"7F",X"55",X"52",X"57",X"49",X"5A",X"DA",X"39",X"1F",X"5B",X"58",X"41",X"1C",X"41",X"1C",
		X"41",X"6E",X"49",X"1F",X"49",X"7E",X"5C",X"51",X"5E",X"CA",X"61",X"5A",X"62",X"49",X"62",X"78",
		X"39",X"1F",X"39",X"7F",X"65",X"D2",X"67",X"C1",X"39",X"1F",X"6B",X"4D",X"6B",X"79",X"49",X"1F",
		X"6E",X"D1",X"70",X"59",X"41",X"1C",X"41",X"78",X"21",X"1E",X"21",X"7F",X"71",X"59",X"71",X"78",
		X"49",X"1F",X"49",X"7F",X"72",X"49",X"27",X"D9",X"75",X"59",X"75",X"78",X"39",X"1F",X"39",X"7F",
		X"27",X"59",X"29",X"59",X"2A",X"5B",X"2A",X"78",X"49",X"1F",X"49",X"7F",X"76",X"49",X"2D",X"1F",
		X"79",X"59",X"7A",X"D9",X"7B",X"41",X"27",X"59",X"27",X"78",X"39",X"1F",X"39",X"7F",X"7F",X"D8",
		X"7F",X"FE",X"7F",X"FC",X"7F",X"F8",X"7F",X"F0",X"7F",X"E0",X"7F",X"60",X"7F",X"E0",X"FF",X"FF",
		X"97",X"B0",X"3E",X"07",X"96",X"95",X"F8",X"2F",X"92",X"F4",X"2F",X"02",X"F0",X"78",X"F5",X"2F",
		X"5E",X"D0",X"BC",X"0B",X"87",X"83",X"F4",X"3F",X"D4",X"BC",X"1C",X"5F",X"50",X"BE",X"65",X"3F",
		X"76",X"98",X"5E",X"57",X"56",X"E5",X"75",X"7F",X"D4",X"B8",X"68",X"57",X"63",X"D4",X"B9",X"2F",
		X"96",X"79",X"66",X"17",X"67",X"95",X"AA",X"3B",X"98",X"E8",X"65",X"5A",X"96",X"A5",X"7A",X"6A",
		X"99",X"96",X"75",X"99",X"A9",X"85",X"67",X"AE",X"96",X"66",X"76",X"1D",X"9B",X"90",X"5E",X"BF",
		X"96",X"65",X"E8",X"5A",X"9E",X"80",X"77",X"BF",X"86",X"69",X"E5",X"6A",X"5A",X"90",X"6A",X"BF",
		X"59",X"E7",X"71",X"69",X"89",X"D4",X"AD",X"6F",X"5A",X"99",X"D8",X"66",X"63",X"A0",X"AC",X"6F",
		X"5A",X"99",X"D8",X"66",X"63",X"A0",X"7D",X"6F",X"27",X"99",X"D8",X"5D",X"8A",X"A0",X"AC",X"6F",
		X"99",X"96",X"66",X"66",X"62",X"66",X"7A",X"7A",X"99",X"98",X"99",X"99",X"89",X"99",X"AA",X"7A",
		X"2A",X"66",X"66",X"2A",X"56",X"55",X"EA",X"AB",X"5A",X"99",X"A1",X"7A",X"96",X"50",X"AE",X"AF",
		X"A5",X"56",X"B8",X"5E",X"5A",X"80",X"7D",X"EF",X"79",X"55",X"B9",X"9D",X"0F",X"D0",X"69",X"BF",
		X"77",X"17",X"A5",X"79",X"1B",X"85",X"99",X"AE",X"99",X"96",X"99",X"66",X"1E",X"96",X"66",X"7F",
		X"8A",X"85",X"E5",X"6A",X"1A",X"86",X"B5",X"2F",X"67",X"62",X"75",X"99",X"8E",X"82",X"F4",X"2F",
		X"8A",X"95",X"79",X"5E",X"1E",X"56",X"B1",X"2F",X"8A",X"95",X"79",X"5E",X"1E",X"56",X"B1",X"2F",
		X"99",X"8D",X"8D",X"8D",X"99",X"99",X"66",X"76",X"62",X"63",X"67",X"66",X"65",X"99",X"D9",X"99",
		X"99",X"89",X"66",X"76",X"99",X"99",X"89",X"99",X"99",X"9D",X"99",X"99",X"96",X"66",X"66",X"8D",
		X"66",X"67",X"66",X"65",X"99",X"D9",X"9C",X"99",X"99",X"98",X"D6",X"89",X"99",X"CC",X"A5",X"99",
		X"CA",X"66",X"23",X"29",X"A3",X"65",X"A2",X"67",X"28",X"D6",X"8C",X"C9",X"CA",X"5D",X"99",X"98",
		X"98",X"A6",X"26",X"97",X"35",X"CD",X"89",X"D8",X"A2",X"8D",X"73",X"28",X"D7",X"35",X"A6",X"28",
		X"9C",X"D7",X"29",X"73",X"29",X"73",X"28",X"CD",X"8C",X"9D",X"68",X"A3",X"32",X"98",X"A3",X"5C",
		X"75",X"9D",X"99",X"98",X"5E",X"95",X"D8",X"BF",X"66",X"75",X"67",X"76",X"26",X"76",X"28",X"7F",
		X"99",X"89",X"9A",X"A1",X"2B",X"82",X"61",X"FF",X"89",X"99",X"9E",X"66",X"58",X"98",X"67",X"AE",
		X"98",X"6A",X"87",X"E0",X"2B",X"55",X"62",X"BF",X"75",X"5A",X"AA",X"56",X"86",X"A8",X"07",X"FE",
		X"98",X"5A",X"A9",X"97",X"58",X"E5",X"0A",X"FE",X"96",X"29",X"E6",X"68",X"59",X"D8",X"0B",X"FD",
		X"8A",X"85",X"E8",X"5E",X"5A",X"82",X"F4",X"2F",X"96",X"A5",X"6A",X"1A",X"57",X"C1",X"F5",X"2F",
		X"98",X"A6",X"1E",X"59",X"C7",X"A0",X"F5",X"2F",X"98",X"A6",X"1E",X"59",X"C7",X"A0",X"F5",X"2F",
		X"8C",X"CD",X"75",X"A3",X"5C",X"D7",X"28",X"CD",X"73",X"5C",X"CA",X"33",X"28",X"D7",X"28",X"CC",
		X"A3",X"32",X"8C",X"A3",X"33",X"28",X"CC",X"CD",X"73",X"35",X"CC",X"A3",X"33",X"28",X"C9",X"A3",
		X"66",X"66",X"66",X"65",X"99",X"9D",X"E7",X"76",X"99",X"66",X"66",X"62",X"66",X"6A",X"77",X"6A",
		X"59",X"99",X"9E",X"57",X"96",X"79",X"99",X"AA",X"65",X"99",X"9D",X"99",X"99",X"E5",X"A8",X"7B",
		X"65",X"99",X"A6",X"5A",X"99",X"D5",X"E8",X"6E",X"26",X"A9",X"66",X"1A",X"A6",X"54",X"6B",X"AF",
		X"D4",X"5D",X"BE",X"05",X"9A",X"A5",X"27",X"AF",X"66",X"75",X"5F",X"86",X"52",X"F5",X"19",X"FF",
		X"66",X"65",X"6A",X"89",X"96",X"B5",X"69",X"D9",X"66",X"59",X"6A",X"63",X"66",X"A6",X"75",X"6B",
		X"98",X"68",X"7F",X"06",X"17",X"E5",X"2A",X"AF",X"56",X"AA",X"6A",X"07",X"D2",X"D0",X"79",X"FF",
		X"22",X"B9",X"75",X"5A",X"98",X"94",X"3F",X"3F",X"85",X"DE",X"A8",X"19",X"9E",X"94",X"3E",X"AF",
		X"1F",X"82",X"E4",X"7C",X"0B",X"A6",X"26",X"7F",X"3B",X"42",X"B5",X"1F",X"57",X"96",X"B1",X"2F",
		X"97",X"C0",X"BC",X"0B",X"D1",X"F4",X"B8",X"2F",X"8A",X"C0",X"FC",X"0B",X"C1",X"F4",X"B8",X"2F",
		X"97",X"A0",X"E8",X"5E",X"57",X"95",X"F4",X"3F",X"97",X"A0",X"E8",X"5E",X"57",X"95",X"F4",X"3F",
		X"8A",X"63",X"66",X"87",X"63",X"5A",X"59",X"CA",X"5A",X"5A",X"29",X"69",X"8A",X"29",X"5E",X"29",
		X"68",X"A5",X"A5",X"A6",X"66",X"66",X"66",X"66",X"62",X"66",X"63",X"67",X"26",X"69",X"96",X"89",
		X"1F",X"43",X"E0",X"BC",X"1F",X"5C",X"6E",X"0F",X"36",X"59",X"E1",X"A8",X"99",X"E4",X"BC",X"2B",
		X"59",X"9D",X"89",X"9D",X"99",X"D9",X"A9",X"9A",X"59",X"99",X"D6",X"69",X"9A",X"72",X"79",X"9A",
		X"99",X"86",X"76",X"98",X"6A",X"87",X"A4",X"7F",X"69",X"86",X"A5",X"59",X"AA",X"95",X"E5",X"6F",
		X"8A",X"58",X"98",X"59",X"EE",X"57",X"A5",X"AB",X"66",X"96",X"31",X"5A",X"7E",X"95",X"A6",X"7E",
		X"66",X"96",X"65",X"66",X"7A",X"66",X"98",X"AE",X"76",X"19",X"D9",X"8A",X"76",X"66",X"98",X"7F",
		X"8A",X"A5",X"62",X"26",X"6A",X"52",X"B8",X"AF",X"A6",X"66",X"21",X"A6",X"66",X"55",X"F8",X"6F",
		X"97",X"5A",X"5D",X"75",X"D8",X"D7",X"5C",X"A3",X"35",X"CA",X"33",X"28",X"CA",X"35",X"CA",X"33",
		X"5A",X"28",X"9C",X"A5",X"D6",X"97",X"32",X"8D",X"72",X"8A",X"35",X"D6",X"96",X"8A",X"28",X"A5",
		X"72",X"97",X"5C",X"A3",X"32",X"8C",X"A5",X"A2",X"8C",X"A3",X"28",X"A2",X"8D",X"73",X"35",X"CA",
		X"5A",X"29",X"75",X"A2",X"97",X"28",X"CD",X"73",X"28",X"A3",X"33",X"5D",X"75",X"A5",X"D7",X"5C",
		X"69",X"68",X"CC",X"A3",X"35",X"D6",X"96",X"8A",X"35",X"CA",X"27",X"28",X"D6",X"97",X"5C",X"CA",
		X"29",X"75",X"D7",X"33",X"5C",X"CA",X"28",X"CA",X"33",X"28",X"D7",X"5C",X"A5",X"D7",X"5D",X"73",
		X"8D",X"75",X"CA",X"32",X"8A",X"5D",X"75",X"D6",X"97",X"5A",X"29",X"73",X"28",X"A2",X"8A",X"5A",
		X"28",X"D7",X"33",X"5A",X"5D",X"75",X"D6",X"8A",X"5D",X"68",X"A2",X"8A",X"5D",X"73",X"35",X"D7",
		X"99",X"72",X"63",X"69",X"99",X"99",X"99",X"97",X"72",X"5A",X"66",X"59",X"99",X"98",X"A6",X"65",
		X"E2",X"97",X"66",X"5D",X"99",X"69",X"99",X"99",X"8A",X"66",X"59",X"99",X"9D",X"75",X"99",X"98",
		X"A5",X"A5",X"69",X"57",X"96",X"98",X"B8",X"2F",X"5B",X"91",X"E5",X"A5",X"2F",X"06",X"F4",X"3F",
		X"66",X"66",X"66",X"67",X"56",X"A2",X"B4",X"3F",X"69",X"59",X"99",X"D9",X"6A",X"67",X"95",X"7E",
		X"29",X"67",X"62",X"76",X"2A",X"63",X"A5",X"6E",X"65",X"99",X"99",X"D9",X"9E",X"59",X"E6",X"5D",
		X"95",X"A9",X"2B",X"43",X"F0",X"B1",X"B8",X"2F",X"95",X"B5",X"2B",X"46",X"E1",X"A5",X"B8",X"2B",
		X"67",X"72",X"29",X"98",X"86",X"A8",X"9C",X"AF",X"5E",X"65",X"9D",X"99",X"56",X"A8",X"99",X"AF",
		X"66",X"99",X"98",X"9D",X"8A",X"95",X"85",X"BF",X"1F",X"91",X"A1",X"BD",X"0B",X"D4",X"26",X"BF",
		X"96",X"76",X"76",X"27",X"19",X"95",X"A6",X"AF",X"5E",X"91",X"AA",X"7D",X"07",X"E0",X"59",X"FF",
		X"6A",X"16",X"66",X"F8",X"07",X"67",X"94",X"BF",X"96",X"69",X"A6",X"58",X"8D",X"87",X"E0",X"7F",
		X"9C",X"67",X"1A",X"5A",X"57",X"D4",X"F9",X"2B",X"78",X"69",X"66",X"5D",X"87",X"D4",X"F9",X"2B",
		X"99",X"89",X"99",X"87",X"96",X"76",X"A8",X"3F",X"A5",X"66",X"69",X"57",X"A1",X"A5",X"F8",X"2F",
		X"2F",X"03",X"83",X"F0",X"2B",X"96",X"E4",X"7F",X"99",X"66",X"66",X"71",X"7A",X"89",X"E0",X"AF",
		X"C6",X"55",X"7A",X"61",X"6B",X"C2",X"B5",X"3F",X"A1",X"98",X"6A",X"61",X"6B",X"95",X"E8",X"7F",
		X"A5",X"66",X"0B",X"D4",X"6A",X"AA",X"C0",X"BF",X"A4",X"3F",X"41",X"FC",X"1F",X"53",X"F0",X"6F",
		X"67",X"62",X"69",X"5A",X"C2",X"B0",X"B8",X"3B",X"67",X"61",X"AA",X"47",X"D1",X"F4",X"B8",X"3B",
		X"5B",X"81",X"B8",X"4B",X"C2",X"B0",X"B8",X"2F",X"9E",X"0A",X"D0",X"AE",X"07",X"D2",X"F0",X"7E",
		X"67",X"A1",X"7A",X"5C",X"0A",X"E2",X"75",X"6F",X"39",X"99",X"99",X"D8",X"57",X"A5",X"98",X"AF",
		X"98",X"99",X"99",X"99",X"99",X"E0",X"F8",X"2F",X"95",X"E8",X"6A",X"1E",X"1A",X"92",X"B4",X"2F",
		X"66",X"6A",X"98",X"66",X"1E",X"55",X"79",X"BF",X"76",X"16",X"B9",X"65",X"5E",X"D0",X"69",X"BF",
		X"6A",X"51",X"FA",X"26",X"0B",X"D0",X"66",X"BF",X"87",X"A0",X"AD",X"7A",X"02",X"F4",X"26",X"BF",
		X"96",X"76",X"68",X"99",X"85",X"E8",X"A8",X"3F",X"96",X"78",X"59",X"7A",X"17",X"A9",X"95",X"7F",
		X"A6",X"26",X"66",X"1A",X"85",X"E6",X"A5",X"3F",X"99",X"9D",X"5A",X"85",X"E2",X"71",X"B5",X"2F",
		X"A8",X"2E",X"0A",X"C1",X"B8",X"66",X"79",X"2B",X"A5",X"69",X"5E",X"57",X"63",X"95",X"B8",X"2F",
		X"66",X"63",X"78",X"62",X"6A",X"A1",X"98",X"7F",X"66",X"66",X"A5",X"5A",X"67",X"A1",X"75",X"7F",
		X"66",X"66",X"99",X"57",X"9E",X"95",X"75",X"7F",X"A5",X"59",X"E9",X"56",X"7A",X"A0",X"1E",X"BF",
		X"79",X"C4",X"7E",X"19",X"8E",X"E0",X"19",X"FF",X"67",X"A0",X"7A",X"69",X"4A",X"F0",X"17",X"BF",
		X"87",X"E0",X"5D",X"EA",X"07",X"F4",X"15",X"FF",X"96",X"79",X"86",X"A6",X"16",X"A5",X"66",X"7F",
		X"98",X"9D",X"5A",X"62",X"67",X"95",X"F5",X"2F",X"A1",X"79",X"66",X"67",X"1A",X"C1",X"F8",X"2E",
		X"A1",X"79",X"66",X"67",X"1A",X"C1",X"F8",X"3B",X"76",X"27",X"59",X"9A",X"56",X"D4",X"F8",X"2F",
		X"65",X"9D",X"89",X"9A",X"66",X"A5",X"E6",X"2A",X"59",X"D8",X"9D",X"8A",X"95",X"E9",X"9D",X"6A",
		X"79",X"58",X"7F",X"47",X"43",X"F4",X"69",X"6F",X"61",X"AD",X"5E",X"46",X"E6",X"60",X"2F",X"7F",
		X"39",X"9D",X"59",X"9E",X"A4",X"64",X"2F",X"7F",X"67",X"59",X"9A",X"76",X"61",X"58",X"6F",X"6F",
		X"67",X"5A",X"66",X"99",X"95",X"62",X"6A",X"AA",X"66",X"67",X"67",X"66",X"58",X"62",X"6A",X"AA",
		X"9A",X"56",X"69",X"57",X"99",X"96",X"B5",X"2F",X"8B",X"80",X"BC",X"0B",X"C1",X"F5",X"AC",X"2F",
		X"8A",X"C0",X"BC",X"0B",X"D1",X"F4",X"EC",X"3B",X"8A",X"C0",X"BC",X"0F",X"C1",X"F4",X"B8",X"2F",
		X"97",X"94",X"B8",X"2A",X"5A",X"92",X"F4",X"3F",X"97",X"94",X"B8",X"2A",X"5A",X"92",X"F4",X"3F",
		X"99",X"C2",X"E4",X"7A",X"57",X"95",X"F4",X"6E",X"96",X"A1",X"79",X"5A",X"87",X"95",X"F1",X"3F",
		X"C2",X"E0",X"7C",X"5A",X"5A",X"92",X"F4",X"3F",X"96",X"78",X"5E",X"57",X"87",X"95",X"B8",X"2F",
		X"98",X"A9",X"2B",X"06",X"E1",X"69",X"E8",X"2F",X"99",X"98",X"99",X"89",X"E2",X"67",X"78",X"3F",
		X"A1",X"AA",X"55",X"6A",X"56",X"97",X"A4",X"7F",X"67",X"57",X"A6",X"78",X"0B",X"D1",X"59",X"FF",
		X"5A",X"A6",X"65",X"5E",X"86",X"85",X"AA",X"AD",X"56",X"AA",X"75",X"5A",X"89",X"D0",X"7E",X"AF",
		X"85",X"E9",X"A8",X"5A",X"89",X"C4",X"6A",X"BF",X"85",X"AA",X"A8",X"4A",X"A2",X"94",X"2E",X"AF",
		X"85",X"A7",X"A9",X"56",X"5A",X"A4",X"5D",X"FF",X"89",X"96",X"AA",X"59",X"56",X"A1",X"9C",X"AE",
		X"A5",X"65",X"DE",X"26",X"5A",X"94",X"77",X"AE",X"A2",X"55",X"EA",X"1A",X"63",X"A0",X"69",X"AF",
		X"62",X"76",X"99",X"99",X"89",X"95",X"A9",X"EE",X"99",X"56",X"B9",X"1A",X"67",X"D0",X"69",X"FF",
		X"A5",X"56",X"B8",X"5A",X"5A",X"C0",X"79",X"FF",X"A1",X"95",X"BA",X"26",X"16",X"E4",X"1A",X"BF",
		X"76",X"65",X"AA",X"55",X"89",X"E1",X"79",X"7F",X"76",X"62",X"2A",X"56",X"5A",X"E1",X"66",X"7E",
		X"79",X"89",X"67",X"58",X"8A",X"A8",X"66",X"7E",X"99",X"98",X"9D",X"86",X"66",X"A5",X"79",X"AB",
		X"99",X"6A",X"26",X"17",X"66",X"A1",X"AA",X"6B",X"99",X"A5",X"66",X"26",X"99",X"95",X"EA",X"7A",
		X"99",X"66",X"99",X"66",X"6A",X"61",X"5A",X"AE",X"96",X"66",X"98",X"9D",X"6A",X"55",X"67",X"AF",
		X"66",X"76",X"65",X"99",X"67",X"95",X"9E",X"3F",X"99",X"69",X"96",X"36",X"1E",X"95",X"A9",X"7F",
		X"1F",X"86",X"A1",X"7D",X"07",X"A6",X"55",X"FF",X"66",X"5B",X"D0",X"BD",X"03",X"E1",X"E0",X"BF",
		X"39",X"2B",X"D0",X"BC",X"07",X"9A",X"D0",X"BF",X"2A",X"9E",X"43",X"F0",X"0F",X"C6",X"94",X"BF",
		X"67",X"98",X"79",X"89",X"56",X"B1",X"69",X"6F",X"67",X"57",X"A6",X"26",X"1A",X"A0",X"A9",X"7F",
		X"27",X"7A",X"55",X"96",X"7D",X"41",X"F7",X"BE",X"61",X"7F",X"1A",X"81",X"AD",X"45",X"A6",X"BF",
		X"66",X"39",X"6B",X"A0",X"1D",X"5B",X"C0",X"FF",X"A5",X"6A",X"86",X"65",X"9D",X"1B",X"D0",X"BF",
		X"66",X"A1",X"79",X"59",X"9D",X"4F",X"E0",X"7F",X"66",X"95",X"9D",X"86",X"A6",X"5A",X"B4",X"6F",
		X"66",X"62",X"68",X"6A",X"5A",X"A1",X"B8",X"2F",X"62",X"6A",X"55",X"DD",X"8A",X"67",X"A5",X"3F",
		X"96",X"66",X"76",X"59",X"D9",X"95",X"67",X"AE",X"C1",X"E1",X"BD",X"49",X"D7",X"94",X"3E",X"7F",
		X"D4",X"78",X"7F",X"07",X"92",X"B0",X"2E",X"6F",X"D4",X"75",X"AF",X"07",X"85",X"F0",X"2E",X"6F",
		X"6A",X"62",X"75",X"66",X"66",X"62",X"B4",X"3F",X"D0",X"FC",X"65",X"2F",X"02",X"E0",X"F8",X"3F",
		X"96",X"76",X"27",X"56",X"A5",X"A1",X"B8",X"2F",X"86",X"E4",X"3F",X"03",X"E0",X"B5",X"7D",X"2B",
		X"79",X"61",X"AD",X"0B",X"D0",X"BC",X"3C",X"2F",X"66",X"5A",X"62",X"69",X"99",X"A9",X"98",X"6F",
		X"66",X"59",X"99",X"9A",X"5A",X"A5",X"A9",X"6A",X"65",X"99",X"99",X"9A",X"66",X"99",X"A9",X"6A",
		X"96",X"69",X"65",X"9D",X"98",X"9E",X"95",X"EE",X"86",X"B8",X"0B",X"86",X"A5",X"3B",X"C0",X"BF",
		X"7C",X"1B",X"43",X"F4",X"1F",X"C2",X"E0",X"AF",X"7A",X"07",X"99",X"95",X"6B",X"95",X"A5",X"AF",
		X"79",X"66",X"15",X"F8",X"0F",X"C7",X"D0",X"BF",X"96",X"66",X"75",X"6A",X"85",X"AA",X"94",X"7F",
		X"D4",X"AE",X"42",X"A5",X"B4",X"2F",X"C4",X"3F",X"86",X"E8",X"47",X"95",X"F4",X"2F",X"C0",X"BF",
		X"8A",X"E0",X"69",X"66",X"94",X"7F",X"80",X"BF",X"6A",X"95",X"5A",X"62",X"95",X"6F",X"90",X"BF",
		X"66",X"62",X"66",X"66",X"76",X"76",X"69",X"DD",X"66",X"59",X"99",X"99",X"DD",X"96",X"79",X"DD",
		X"89",X"9D",X"85",X"9D",X"D9",X"99",X"9D",X"EA",X"99",X"99",X"D9",X"55",X"A9",X"9A",X"22",X"AE",
		X"82",X"F5",X"F4",X"1E",X"0B",X"91",X"B9",X"6F",X"72",X"B8",X"2C",X"0F",X"57",X"84",X"7F",X"2F",
		X"A6",X"65",X"69",X"5A",X"86",X"71",X"7E",X"3B",X"98",X"99",X"67",X"27",X"65",X"A6",X"2E",X"6A",
		X"99",X"A6",X"1A",X"17",X"98",X"A5",X"6E",X"6B",X"95",X"6B",X"9E",X"03",X"D1",X"F0",X"3E",X"7F",
		X"A4",X"3E",X"2F",X"02",X"87",X"B4",X"2E",X"2F",X"A4",X"3D",X"6F",X"46",X"52",X"F4",X"3A",X"3F",
		X"D4",X"E0",X"BE",X"1E",X"02",X"F0",X"69",X"AF",X"66",X"98",X"7A",X"66",X"47",X"A5",X"65",X"BF",
		X"65",X"9D",X"66",X"5A",X"96",X"A5",X"B8",X"6B",X"65",X"A6",X"27",X"1A",X"86",X"E1",X"B8",X"2F",
		X"A4",X"7D",X"47",X"8E",X"82",X"F5",X"78",X"3F",X"95",X"A5",X"7F",X"0A",X"02",X"FC",X"0E",X"AF",
		X"95",X"86",X"F9",X"55",X"56",X"F0",X"3E",X"6F",X"17",X"A3",X"F4",X"19",X"6A",X"A0",X"7D",X"7F",
		X"6A",X"99",X"C5",X"89",X"96",X"90",X"FD",X"AF",X"A6",X"58",X"99",X"9C",X"85",X"99",X"EE",X"7E",
		X"99",X"99",X"99",X"66",X"85",X"A8",X"E8",X"6F",X"A2",X"67",X"62",X"1E",X"81",X"F5",X"78",X"6F",
		X"76",X"59",X"99",X"9A",X"1A",X"C1",X"F8",X"2F",X"C2",X"B4",X"79",X"69",X"4F",X"82",X"F4",X"2F",
		X"A1",X"E8",X"2E",X"0B",X"47",X"C2",X"F4",X"2F",X"C4",X"BC",X"0F",X"83",X"D1",X"F0",X"BC",X"1F",
		X"B4",X"3E",X"0A",X"D0",X"F5",X"78",X"7D",X"1F",X"A4",X"AD",X"2A",X"1E",X"4A",X"D0",X"F5",X"2F",
		X"96",X"75",X"6A",X"1A",X"95",X"E2",X"A8",X"2F",X"A4",X"AD",X"0F",X"82",X"D6",X"A0",X"F8",X"2F",
		X"78",X"2E",X"0E",X"8A",X"57",X"D0",X"FC",X"2B",X"75",X"6A",X"57",X"67",X"56",X"D4",X"F8",X"3B",
		X"6A",X"55",X"E8",X"6A",X"55",X"6B",X"84",X"AF",X"99",X"96",X"76",X"18",X"9D",X"9E",X"85",X"FE",
		X"9A",X"9D",X"56",X"11",X"FA",X"19",X"A9",X"7F",X"1F",X"87",X"D0",X"A8",X"6A",X"80",X"AE",X"AF",
		X"57",X"E5",X"B0",X"2D",X"67",X"90",X"7E",X"AF",X"69",X"95",X"FC",X"0E",X"0B",X"C0",X"E6",X"BF",
		X"1B",X"D1",X"E4",X"BC",X"03",X"F4",X"7C",X"3F",X"C6",X"92",X"F0",X"2F",X"02",X"E1",X"F0",X"7F",
		X"99",X"A1",X"79",X"59",X"9D",X"87",X"B5",X"3F",X"98",X"9D",X"5A",X"62",X"69",X"99",X"B8",X"2F",
		X"57",X"A5",X"66",X"2A",X"96",X"99",X"A7",X"66",X"59",X"D9",X"66",X"66",X"A6",X"66",X"77",X"66",
		X"26",X"A5",X"69",X"5A",X"A6",X"66",X"6A",X"66",X"27",X"6A",X"62",X"19",X"E6",X"61",X"6A",X"AB",
		X"79",X"0B",X"DA",X"90",X"E9",X"A4",X"2A",X"BF",X"75",X"5E",X"5B",X"D0",X"E1",X"F0",X"2A",X"BF",
		X"79",X"1E",X"1F",X"C1",X"C2",X"F0",X"2E",X"7F",X"27",X"99",X"8A",X"A1",X"86",X"A5",X"66",X"7F",
		X"66",X"62",X"66",X"69",X"87",X"D5",X"B8",X"2F",X"27",X"98",X"5E",X"D9",X"07",X"E1",X"E1",X"BF",
		X"5E",X"84",X"7F",X"8A",X"41",X"F5",X"68",X"AF",X"E4",X"61",X"7E",X"9D",X"07",X"E0",X"7A",X"3F",
		X"E1",X"18",X"BE",X"1A",X"06",X"E0",X"A8",X"AF",X"9A",X"80",X"BE",X"79",X"07",X"A1",X"69",X"AF",
		X"9A",X"59",X"98",X"96",X"76",X"56",X"F4",X"3F",X"79",X"4B",X"D0",X"F4",X"AD",X"0B",X"E0",X"3F",
		X"3E",X"12",X"B4",X"2E",X"0B",X"83",X"F4",X"3F",X"8A",X"82",X"F0",X"3F",X"03",X"B4",X"AC",X"2F",
		X"D0",X"BC",X"2D",X"4B",X"C0",X"B8",X"A8",X"3F",X"29",X"8D",X"67",X"99",X"8A",X"A0",X"B8",X"2F",
		X"2A",X"25",X"9A",X"98",X"67",X"A1",X"E9",X"2F",X"66",X"62",X"66",X"67",X"66",X"79",X"99",X"9E",
		X"98",X"A6",X"26",X"97",X"35",X"CD",X"89",X"D8",X"A2",X"8D",X"73",X"28",X"D7",X"35",X"A6",X"28",
		X"9C",X"D7",X"29",X"73",X"29",X"73",X"28",X"CD",X"8C",X"9D",X"68",X"A3",X"32",X"98",X"A3",X"5C",
		X"73",X"59",X"9D",X"8A",X"86",X"69",X"66",X"98",X"9D",X"8A",X"35",X"D7",X"63",X"28",X"CA",X"65",
		X"A3",X"62",X"75",X"A3",X"29",X"68",X"A5",X"D7",X"35",X"CA",X"32",X"8A",X"29",X"8A",X"65",X"CA",
		X"69",X"8C",X"9A",X"5C",X"A3",X"63",X"5A",X"5D",X"73",X"5C",X"D7",X"32",X"8A",X"35",X"9A",X"29",
		X"8A",X"35",X"C9",X"A3",X"32",X"8A",X"36",X"28",X"D7",X"32",X"8C",X"A3",X"5C",X"D7",X"35",X"D7",
		X"66",X"77",X"59",X"66",X"72",X"61",X"7A",X"AE",X"C1",X"A9",X"EA",X"43",X"E0",X"B0",X"3E",X"3F",
		X"C5",X"D4",X"BE",X"1C",X"46",X"F4",X"2E",X"2F",X"D0",X"F9",X"A4",X"3F",X"02",X"E4",X"B8",X"3F",
		X"C4",X"F8",X"2B",X"42",X"F0",X"A5",X"F5",X"2F",X"99",X"67",X"17",X"98",X"9D",X"D5",X"F5",X"2F",
		X"66",X"66",X"56",X"99",X"D9",X"A5",X"A7",X"7A",X"5D",X"97",X"56",X"99",X"E5",X"A6",X"69",X"DD",
		X"67",X"99",X"85",X"96",X"A6",X"68",X"7A",X"3B",X"89",X"8A",X"A2",X"85",X"E5",X"A4",X"7A",X"7F",
		X"98",X"5E",X"8E",X"C0",X"F4",X"B4",X"2E",X"7F",X"C0",X"FC",X"68",X"2F",X"03",X"E0",X"B8",X"3F",
		X"75",X"A9",X"3D",X"0F",X"57",X"83",X"F4",X"3F",X"A1",X"A5",X"B4",X"7D",X"1F",X"42",X"F4",X"2F",
		X"A8",X"2E",X"1A",X"0E",X"D0",X"7F",X"43",X"F0",X"9E",X"4A",X"E0",X"1F",X"81",X"F4",X"EC",X"2F",
		X"3F",X"06",X"A8",X"0B",X"82",X"A5",X"F8",X"2F",X"9D",X"D8",X"2E",X"07",X"93",X"C3",X"F4",X"3F",
		X"2E",X"47",X"D0",X"B8",X"2D",X"6D",X"1F",X"C2",X"2E",X"0A",X"D0",X"EC",X"2A",X"2B",X"0B",X"C3",
		X"99",X"D1",X"F4",X"6D",X"2D",X"3E",X"0B",X"D0",X"3D",X"0F",X"82",X"B0",X"B4",X"F0",X"F8",X"3D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
