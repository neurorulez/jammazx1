-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu1 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFE2FFFFFFFFFFFFFFFFFFFFFDAFF4B4138A420B420B420B420B4C0";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0F";
    attribute INIT_02 of inst : label is "1882F8E2863A2B84E253844E4A700151431154312FC2E280AF68D28E20E03DBD";
    attribute INIT_03 of inst : label is "CA2E01BE9894F18D2FC6AD7760A5A317AD8ED3B6F03EF05FB450FFF8A5794E10";
    attribute INIT_04 of inst : label is "11A52AFC62EF760A5A317AF8ED3B6703E705FBE620D466EBFD82993F6E845378";
    attribute INIT_05 of inst : label is "239DBC10308000AE2478A5805823AE61466EBFD82993F6E845378CAFFFFFFFCA";
    attribute INIT_06 of inst : label is "A69540A1018825939565510D694173A103F4402AD50374049FE9DF21A3C64008";
    attribute INIT_07 of inst : label is "0B1B40000000092A9238AE0E13EA28E8AE0E13C0025147634D04C6420BD10874";
    attribute INIT_08 of inst : label is "5F3C371F39656142400009065722090653B1471041020612B0AD38138F88A3A1";
    attribute INIT_09 of inst : label is "20710400197CF0811CF16984472F8F501C38A431D7911541B948778154382464";
    attribute INIT_0A of inst : label is "E5958509000810400D1ED40C21803C4113CE319196066F3C1A9103F3CC3C3800";
    attribute INIT_0B of inst : label is "2071A945614A573A2B8E501D45F3C119430760385E608184AC28F8917CF0DC7C";
    attribute INIT_0C of inst : label is "C22A1253B4072BCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5A05A9328364";
    attribute INIT_0D of inst : label is "142405A03E220612B0AD0C21041803C43CF06AC40FCF30F0E01681C4100065F3";
    attribute INIT_0E of inst : label is "145397814844905A1384276964968D4945415A5CF3C904929845F3C371F39656";
    attribute INIT_0F of inst : label is "E14657340EA5AE23A83CE23A80C2E84CE4548E473C23417D146D4A15398F3CAA";
    attribute INIT_10 of inst : label is "04AF000884404E200F0138C1E0CA000A0ACA90C5899992F0C3C44F0F5A439590";
    attribute INIT_11 of inst : label is "A05A2EE894070589451939209901E831AE6338597CF04292A746BBCF27726D38";
    attribute INIT_12 of inst : label is "FFFFFFFFFEAF3C13CFFFFFFFFFFC84A9384D8840752D18F3CCD4221A5085412A";
    attribute INIT_13 of inst : label is "4FFFFCAC5432423B7E94000734FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF64293201947291A62B";
    attribute INIT_15 of inst : label is "A1105184734FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "D03000324640C040324FF7B40BE103D407D13CA7B02C40FE5EC0FD02F4074E53";
    attribute INIT_17 of inst : label is "555554B7E651D95F8A57B440FBD3B64AF964A902C0A3CF34240F01A6F53B41B1";
    attribute INIT_18 of inst : label is "1113FFFFFFFFFFFFFFFFFFF0000000000000000000000AECEE8AA4466AA62025";
    attribute INIT_19 of inst : label is "9E85DE15779550E053B1B226200E20060228040C0A2E2B9EA8EE658000111111";
    attribute INIT_1A of inst : label is "56A8E4FA97931279CBD2D33D0F390B666E6EEE65DD555D55C666AF9679DFA9C7";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFDFFDFFDFFDFFDFFDFFDFFDFFDFFDAA839391A7913FFFFFFF";
    attribute INIT_1C of inst : label is "77BA9747B3A8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF085B79FFFFFFFF";
    attribute INIT_1D of inst : label is "A0000000005A0000056AFFFFFFFFFFFFFFFF90E749D200EA150000FCE4FBFBA9";
    attribute INIT_1E of inst : label is "A80A80A8014000016969405AAAA02A02955015A556800002A000150150002A02";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0169400056AA0030000001680";
    attribute INIT_20 of inst : label is "41C40D80C94C850C49278154AEA65BFA67906F4D26E2D88D3030321032301030";
    attribute INIT_21 of inst : label is "F33F7FBF7FBF333FBF7FBF7FBF3F7F3B37BFC33233FF3C111C1F311D5D3C8508";
    attribute INIT_22 of inst : label is "46467DD9191D5F7447447D1D11D13C8A8C8CBBAB8C8CBC8CBC8BABCB9B8A89AB";
    attribute INIT_23 of inst : label is "111931DDDF1113CCECECCCFDFCFEFECCFCF232B2B2322A3232F272F2F22A3757";
    attribute INIT_24 of inst : label is "B3F3F333F333B3F3F333F333F3333C8A8A88B9B8A8AC8C8CBCBC8C8B9F11F1D3";
    attribute INIT_25 of inst : label is "EDFCFCCCFCCCFDFCFCFCCFCFCEDFF311D5D1D5D1D5D33C4757475747574CF333";
    attribute INIT_26 of inst : label is "30F030F0F0F0F0F0F0F030F030F030F030F0F0F0F0F0F0F0F3CCFDFCFCFCFCFC";
    attribute INIT_27 of inst : label is "7CE987610FE987610F24AC12F852D2F852D2F852D2F852FBA98BA98BA98BA9F0";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC8B8C9C9CBCBC8CBC8CBC8CBC8CB98F1476547655";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "D082D082D7450511FF0309744B09D79E4E9575BFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "0AFFA90638F14FAA418E3853CA3C18E30533F633D8DF60A50020B7539082D082";
    attribute INIT_30 of inst : label is "7D1B852E0C46E14F8F11B850E2E491A147A471B852E1124B1CE4463F500608E5";
    attribute INIT_31 of inst : label is "5E0C65BC95046A9D0A609FC444B909B3D87E0D6186853E1F71B850E2D46E1478";
    attribute INIT_32 of inst : label is "B8425D8409A0B288B5DBE8255555E63191A383FE5869058642E55555782E5555";
    attribute INIT_33 of inst : label is "C2D5C9505EA9D0A6BA2444525E0976809A0B288B5DBE82555551A86288B54D2E";
    attribute INIT_34 of inst : label is "6564EE3B4F0B472541BA990A5EA18A22D534BAE10898408A55A6666564DE8ED3";
    attribute INIT_35 of inst : label is "0000D98EEBB5010C040231648E040C0D0BE6618A22D534BAE10898408A55A666";
    attribute INIT_36 of inst : label is "FFFFFFFFFF73CCCD159E6F73CCDE2B389AB385681EF5EC1F1B9028BA987F1B20";
    attribute INIT_37 of inst : label is "1940AF29303C0757FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "CC064A4D2834AEB79A5443CD04A1111C4951147701B9511111C7171CA55AA612";
    attribute INIT_39 of inst : label is "5C39C571309C79F44388C1AA840B1E9256D19BCE21919110011D042413191B72";
    attribute INIT_3A of inst : label is "407051208393815B225250240B98209701EC55582356664ACBD6086340B0FDC7";
    attribute INIT_3B of inst : label is "9689162A0E56249BB44F06092342B9C84053E496D120014F9253B19AA630BE3D";
    attribute INIT_3C of inst : label is "AD4887862D01EA4BBA4B8B442F7274109B05A6613559E504D826664266BEE680";
    attribute INIT_3D of inst : label is "438056DB4904D04654104539D4D1027FB9C9FFFEF3D5302490152A4392938401";
    attribute INIT_3E of inst : label is "51043609999910A0486B2588BB443856B444B4BE3D44748DAF7A620E0F651400";
    attribute INIT_3F of inst : label is "903D242443E2B8574A91BB9198125BB7CADDDDDFB7CC65915401930E5622D0E2";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFC6FFFFFFFFFFFFFFFFFFFFFCEFF0A80007830F430F430F430F400";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAC6";
    attribute INIT_02 of inst : label is "06CD18F3C71F1F5279E37939812711AF90C4790C780E8690F78556996574235E";
    attribute INIT_03 of inst : label is "0D06F43DA3DAA638E24060A21878506A1A41D2C48128813A5719C638F92B8DF6";
    attribute INIT_04 of inst : label is "605F42240E0E21878506A1A41D2C40128013A553F0B81BE636C9F2383296F422";
    attribute INIT_05 of inst : label is "F061CDE2C06222704998F3C52C32F13F81BE636C9F2383296F4220DFFFFFFF5B";
    attribute INIT_06 of inst : label is "F0C550FF606CDEA350F57A08FCC4E2F7129788DC1ACB588824C6A011A695888E";
    attribute INIT_07 of inst : label is "24376222222226EFE21C7D4FE39B347C7D4F238006ACD0E555759D9C4E760412";
    attribute INIT_08 of inst : label is "277548AF7090808D80000F5154971F5158E71D75F45D43D0E0F949E3417433FE";
    attribute INIT_09 of inst : label is "35D453450C5DD6D57534BD2B3518867119F52E573D4ACD442B51DD4A6C541960";
    attribute INIT_0A of inst : label is "C2420236000D4534594B114D24100115ADD26F2F2E41A7750F85947750BD3400";
    attribute INIT_0B of inst : label is "168AD0A080858D531485711902775079D52CC124527750F4383C17409DD522BD";
    attribute INIT_0C of inst : label is "5B7F55014C4614DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4BD2F852F778";
    attribute INIT_0D of inst : label is "08D8007505DD43D0E0F94D24514100115DD43E9651DD42F4D001D7514D143177";
    attribute INIT_0E of inst : label is "5D234B412E6042056378B43431C7D08080808591775420015D0277548AF70908";
    attribute INIT_0F of inst : label is "B281BF7F14B0B6D74B1B6D74B2817A86285092977534C42B61BA81B637977566";
    attribute INIT_10 of inst : label is "B9A8400398EB5D9FC6AD767C52AEAAAEAE5EF5FF12222192A18E8EA920A44829";
    attribute INIT_11 of inst : label is "344D41215C462A422A8226626711A50E744C750D5DD581A1688189DD6896BAD1";
    attribute INIT_12 of inst : label is "FFFFFFFFFD2775F7DFFFFFFFFFF5985E340C04047012F9775810819297550816";
    attribute INIT_13 of inst : label is "5FFFF5B32987813C597D000E75FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF781856F43DE7A068D7";
    attribute INIT_15 of inst : label is "5F756045E75FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "990D40C69A643D00C697F1AC466711AC46763986611BC46619846F118C462363";
    attribute INIT_17 of inst : label is "00000100004400038F929B6520234D813BD81B1381A5DD48D64215B98E37D1E1";
    attribute INIT_18 of inst : label is "1113FFFFFFFFFFFFFFFFFFF00000000000000000000001102111003122221020";
    attribute INIT_19 of inst : label is "7070CF0C3152140083BA5053733DEEAD5C58595880C25D590A445508A0911111";
    attribute INIT_1A of inst : label is "000C63EC9803FEADC000006070A0B048C44C40C840C84C8C4400000000014731";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFF2AA7FF7FF7FF7FF7FF7FF7FF7FF7FF7FF3FE9498CCC0000000";
    attribute INIT_1C of inst : label is "BD2C9BF2FBD8CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF166440FFFFFFFF";
    attribute INIT_1D of inst : label is "05680000AA50002AA540FFFFFFFFFFFFFFFFFEA96504045515455100009E6EC9";
    attribute INIT_1E of inst : label is "01501501682A96A800002A0000054054000A80000016969405AA80A80AA94054";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA800296A0000557955AAA8015";
    attribute INIT_20 of inst : label is "551551151111111108510C1304C110CC11008004004832083311321021003200";
    attribute INIT_21 of inst : label is "F0400CCC0CCCB08CCC0CCC0CCF0C0044888BC20103CCFC000C0F0008CC355555";
    attribute INIT_22 of inst : label is "00111C44400CCB2213320C0884CCBC033C0C11113C3C1C0C1C0111C122330000";
    attribute INIT_23 of inst : label is "19DDF1D1D31597C03C33C3303C0101C222F0707070B08470B0B0F0B0B0847233";
    attribute INIT_24 of inst : label is "F03030F030F0F03030F030F030F33C2232233033222C3C3C3C3C1C100F1DB19B";
    attribute INIT_25 of inst : label is "003C3C1C3C1C003C3C0CC3C0C003F044C0040448488F300233023302330CF0F0";
    attribute INIT_26 of inst : label is "F1313131B131B131B131F131F131F131F1313131B131B131B3C1003C3C0C3C0C";
    attribute INIT_27 of inst : label is "3C444777722221111F26558845550845550845550845553012330122301123F1";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC746C3C3C3C3C3C3C3C3C3C3C3C333F2211110000";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "D0C3D0C3D7B62BA0B21405408D16A9D575A9C12FFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "05658794597F8120C5165BE878BA51657E0BBC10F053C05988B0526350C3D0C3";
    attribute INIT_30 of inst : label is "C6B84A2DB2AE3287686B84A1DA082BB28B4E8B84A1DFA0A63818C8BBD4D6343E";
    attribute INIT_31 of inst : label is "A37196CD061AE0E7108AAE088A92164092E4774CEECA0DB28B84A0DB2AE328F6";
    attribute INIT_32 of inst : label is "2443AE440C00F000DAF2513AAAAA3A065B80F09A98A71C2943FAAAAAB83FAAAA";
    attribute INIT_33 of inst : label is "83D3D061A20E710898C888BCAA0EB9C0C00F000DAF2513AAAAAB82B000D08E25";
    attribute INIT_34 of inst : label is "8A88260FC20F4F418698E710A20AC003423894910CE440CCEEC8888A882203F0";
    attribute INIT_35 of inst : label is "2000D88D649A01A0788101739238809D06578AC003423894910CE440CCEEC888";
    attribute INIT_36 of inst : label is "FFFFFFFFFC8CD159159D5919E6E62A6FB733CCCD115E2B7FC89E27F856AF805B";
    attribute INIT_37 of inst : label is "D6402962ED085593FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "7939B1A93417A03C2461819717EEEEE381869C98015186EEEE3A2824DAA00C53";
    attribute INIT_39 of inst : label is "742F35D101355B15D57705091C42165C849F2DD25F2F21E201D60A0818C636C4";
    attribute INIT_3A of inst : label is "C4605A386C544169CDD6B58D64D0D114012C5EBB20EAC943827FFB28C4281F02";
    attribute INIT_3B of inst : label is "6A8C005D49A230004D8E07DDEC452BD389CA32F8DA38EB28CB10665314D46219";
    attribute INIT_3C of inst : label is "593D868557118BD847D8545C594F9828240499BA31CD3A0AF088889092419752";
    attribute INIT_3D of inst : label is "C75041F90C208041580000063B622082E6063FF67F977520001007D8545CF881";
    attribute INIT_3E of inst : label is "9000BC22222B340043913131FB1C755485E824E239D8660C20CCA476436822D5";
    attribute INIT_3F of inst : label is "94C308DB8A33490CC90272207975923598F22225D7F509EAA84E607184C771D5";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFC7FF0F0338D01C781C581C781C58C0";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF768";
    attribute INIT_02 of inst : label is "AFA73E9A69A6A5E9CF99C6045328A384AB388AB3A0C569E86B4259E8966808ED";
    attribute INIT_03 of inst : label is "270FE8FF18741180F70CB45B5BC59314B2D3E948B390B3809D0A741E521C67CB";
    attribute INIT_04 of inst : label is "D8EF8770CF49B5BC59314B2D3E94833903380933402638FC1E032D9192389D8F";
    attribute INIT_05 of inst : label is "6BCF0AC378F33AE18E1E585A86196336638FC1E032D9192389D8F27FFFFFFF0F";
    attribute INIT_06 of inst : label is "6A4AA86CBAFA7159F2122D4214CE0953391F0E7BF84FB0C4938D0D3379EF0CCB";
    attribute INIT_07 of inst : label is "339FB3333333ACB94BA697A559159E9A97A559000544A39A6A9A3C48E4B94C38";
    attribute INIT_08 of inst : label is "D49224D7834343674000079B23A9A79B2349679A7A24A92A4A668299EB5E996C";
    attribute INIT_09 of inst : label is "1E7B6DBEA4924AE09ECA1B352AA06833A05ED8C72DCD488E8231C9C15C5EF470";
    attribute INIT_0A of inst : label is "0D0D0D9D0007B6DBE9A52CB2DB603A8B85238E9F99935492A688AF4928DE9C00";
    attribute INIT_0B of inst : label is "334D9353436B4799AC6B33A30D492E878F0CA1AC19292A4A929AB5C35248935E";
    attribute INIT_0C of inst : label is "2B970A5ACCE8AF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0D28688F4BB6";
    attribute INIT_0D of inst : label is "367404DEAD74A92A4A69B2DB6CB603A8924A9862BD24A37A701379EDB6FA9249";
    attribute INIT_0E of inst : label is "8E59E6C1948C71E7D9F0E38E9B6DB34343636F7A49271C3ACA0D49224D783434";
    attribute INIT_0F of inst : label is "416B58CBE0F2F24CCAA024CCAA022F00F41ACF6F9E388E8ABE1653219E649213";
    attribute INIT_10 of inst : label is "2726C00B280133262804CC5A7A0BFFCBCB4A332331111A1A0A3B641492472491";
    attribute INIT_11 of inst : label is "D0449314C8E835493509AD1AD23A3433D589DAA49249631AC46B3D248443342B";
    attribute INIT_12 of inst : label is "FFFFFFFFFCB492CBAFFFFFFFFFF0D6BD9CCF5CC07DFC664922CCD7616238CDF1";
    attribute INIT_13 of inst : label is "AFFFF0F5024A63B492BE000EBAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF63883E8FEEB58D63B";
    attribute INIT_15 of inst : label is "ECAA58C2EBAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "0A3B80FB6128EE00FB67FBD8E81A3A08E871924853A08E8D214E863A18E83F19";
    attribute INIT_17 of inst : label is "0000000000000001E521F12BC319DC531DC533391A792486728E21E4319F2A4A";
    attribute INIT_18 of inst : label is "3E97FFFFFFFFFFFFFFFFFFF00000000000000000000004554554554445555540";
    attribute INIT_19 of inst : label is "2330CF0C33F30000C33001E92925E5E5E5E5E5E63A39E55555555549CB543E94";
    attribute INIT_1A of inst : label is "000144D216A95556D7D94BFFFFFFFDDD99D9DD99DD99D9D99D5BE9759DD43230";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFF3FF3FF3FF3FF3FF3FF3FF3FF3FF3FF2AAEAAAA50FA40000000";
    attribute INIT_1C of inst : label is "711217511711FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF244000FFFFFFFF";
    attribute INIT_1D of inst : label is "0000AAAA5555AA95555500000000000000000000000009000000000000AAA921";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000030000000000";
    attribute INIT_20 of inst : label is "00C000C000C000C414541867110761D45411C618619054105555444477776666";
    attribute INIT_21 of inst : label is "E18885458546A285458545854424989ABABB82AA21F778CCF84C0CC888F000C0";
    attribute INIT_22 of inst : label is "66666D999995572221111CC88844785008888040888888888880400804049D9D";
    attribute INIT_23 of inst : label is "264662686A2A8B8D888D099298AA2A8AA2C182828282A8828282828282BBB555";
    attribute INIT_24 of inst : label is "226262226222226262226222622038D111515A19151898989898A8A2AE322234";
    attribute INIT_25 of inst : label is "2698982C98A026989820898A0269E088488844440003333222322232223CE322";
    attribute INIT_26 of inst : label is "22626262226222622262226222622262226262622262226233862698982C98A0";
    attribute INIT_27 of inst : label is "38AAA999999999999E333321032121032121032121032138888899999AAAAAE1";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFF0C55090909090909090909090909DDE2222222222";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "6071E0716E1C0ED43C13CFD0418D9566D7D4E2CFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "4E46FF3B5E674D7DDED795D37F75ED791D777A17E86FA8E7CCE8D919F071E071";
    attribute INIT_30 of inst : label is "354E458B7C538162DB14E058B5F494F166DB64EC59B2D2512E340867A0EB34E9";
    attribute INIT_31 of inst : label is "526309FF81253C533274D18445618D383F0792B4D3859B4E64E859B5E539162D";
    attribute INIT_32 of inst : label is "AC81D2C804A0428815E93835555525CC24F848126C6334C0B17555555C175555";
    attribute INIT_33 of inst : label is "31E6F81257C533277F8444485FC74B8C4AC428815E9383555554F3528810451F";
    attribute INIT_34 of inst : label is "4444DF87A0079BE0497C533257CD4A2041147EB2C7EC8C6F9944444444D7E1E8";
    attribute INIT_35 of inst : label is "5B20F6D7DF7C09DC70D332F14D30EC5E4C6F4D4A2041147EB207EC806F994444";
    attribute INIT_36 of inst : label is "FFFFFFFFFC000000000000000000000000001111111111112222222333330000";
    attribute INIT_37 of inst : label is "1DC0D3105E305D53FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "D63547725C3DB3C894124B16395999934049D97109804999993425142550C8E0";
    attribute INIT_39 of inst : label is "6A87C8A23128B2D9685CC4C4CCE83D340B3F9D23AE9F93C3097C0724972D5E8C";
    attribute INIT_3A of inst : label is "CE827C3CB326C9E774DF1AF6B72D716D091E4F4450F4C6E928265F1CCE8EB2E8";
    attribute INIT_3B of inst : label is "D3C70D34AB4F1C34DC64252B169BC3FF0CE0E864EC1C7383A1A6C02EC88E81A0";
    attribute INIT_3C of inst : label is "A31E4A49323A15E34DE34C98E1D7701C9326767C3CA8F80720C4444269CE2D2A";
    attribute INIT_3D of inst : label is "CDA25B5DC71C725BF030C3BCE1C1324C6D4CFFF5FF3B9A2C70976DE326F5F0C9";
    attribute INIT_3E of inst : label is "730CC8311113E0A248F9062767C8DAC848F50E81A0C68FCF18FBD4284DB30CAE";
    attribute INIT_3F of inst : label is "263226770CE8CE48A799D594E63A7CD23B2DDDD4899327D1544D5307589D336A";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFC9FF07B1247B38F338F338E338E080";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC951";
    attribute INIT_02 of inst : label is "47D13575D75F5C270D455A2A210962EDA2581A25BC8068A8F74E18A08E1A1C9D";
    attribute INIT_03 of inst : label is "150508FD44D0A044DDC41CE1F4613220DBA1C5C0335433776B022B157007153B";
    attribute INIT_04 of inst : label is "C45289DC49C61F4613220DBA1C5C0F354F377660C8511AF71E8134577334CF17";
    attribute INIT_05 of inst : label is "754A02EF247FF5708E5577D27E35F60D11AF71E8134577334CF1715FFFFFFF24";
    attribute INIT_06 of inst : label is "F7C028F3B47D1C4561F03885F44DD5D1356BBD1CAEFF3BFC3207CB9229EBBFFF";
    attribute INIT_07 of inst : label is "F2673FFFFFFF555E955D70978542557D709705400CEC2218638AC600D5108437";
    attribute INIT_08 of inst : label is "728E2CF181C1E1D1C00001BD0208E1BD0228E18668639705E5F3828554C5B6FE";
    attribute INIT_09 of inst : label is "0E18608E4E0A38E28639FE3D0554151354424CC4118F4C0DD331058300D95CD8";
    attribute INIT_0A of inst : label is "0707874700038608E09B018E38A00E1AECA0BF0D01A1028E4F382A28EBC64400";
    attribute INIT_0B of inst : label is "13CFD1D1E1D1C1A2541513568728E183CD4443440028E5C1797D4C61CA38B3C6";
    attribute INIT_0C of inst : label is "E3A829F544D554EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1467F3811B31";
    attribute INIT_0D of inst : label is "1D1C0C4E53139705E5F08E38618A00E18A393C20A8A3AF191031386182393828";
    attribute INIT_0E of inst : label is "9E0558806C075D59C57BF275F6DBE1C1C1D1D9CE28E5D7944A8728E2CF181C1E";
    attribute INIT_0F of inst : label is "90D1CCC4A343430F8E4430F8E47D3793F00148A39258CDD18A19213054628E04";
    attribute INIT_10 of inst : label is "0739C00027083E121120F849944555450545130130000454544E152830C30C30";
    attribute INIT_11 of inst : label is "5000BD0F4CD53E433EC3570573357C215800C27C0A391144501134A3900938F7";
    attribute INIT_12 of inst : label is "FFFFFFFFFC528E382FFFFFFFFFF2511C545DC45037DEC628EC85F1C0C0345FDD";
    attribute INIT_13 of inst : label is "EFFFF24F1A49114C2C4A00008EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB1138908CA08445114";
    attribute INIT_15 of inst : label is "5386445208EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_16 of inst : label is "42A18038A00A8E0038ABF34CD503354CD5105400A354CD50028D53354CD51C05";
    attribute INIT_17 of inst : label is "000000000000000157007B0AB2054621146211355628A38110A863503054E5E5";
    attribute INIT_18 of inst : label is "4003FFFFFFFFFFFFFFFFFFF0000000000000000000000CDDDCFFCFDDCFCDFFF0";
    attribute INIT_19 of inst : label is "13300C4030001454137552569696565656565656969654000000003A542A9555";
    attribute INIT_1A of inst : label is "000000C001555557C00000000000033FFFBB7777BBBB77333C00000000033133";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFF2AA3FF3FF3FF3FF3FF3FF3FF3FF3FF3FF55555550000000000";
    attribute INIT_1C of inst : label is "300003000300CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400000FFFFFFFF";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000002000000000000AAA800";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000030000000000";
    attribute INIT_20 of inst : label is "CC8CCC8CCC8CCC8208020832040110CC11008208108803081111111100000000";
    attribute INIT_21 of inst : label is "F122323232312232323232323323232212138888CCF33CDDFCDF3333333CCC8C";
    attribute INIT_22 of inst : label is "CCCCCF33333333CCCCCCCF333333384888888C8C48888888888C8CC8C8C88484";
    attribute INIT_23 of inst : label is "2222222222222384888488888888888888F23232323222323232323232223CCC";
    attribute INIT_24 of inst : label is "222222222222222222222222222338488C8C8888C88888888888888C8E122212";
    attribute INIT_25 of inst : label is "C88888848888C888888888888C88E3333333333333323CCCCCCCCCCCCCC8E122";
    attribute INIT_26 of inst : label is "2222222222222222222222222222222222222222222222221384C88888848888";
    attribute INIT_27 of inst : label is "BCCCCCCCCCCCCCCCCF33333332223332223332223332223CCCCCCCCCCCCCCCE1";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFC488C8C8C8C8C8C8C8C8C8C8C8C888F2BBBBBBBBB";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "CCE38CE38BBECFC87B3246B1CD476158B060407FFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "05B349340E3008D34D038C022428D038C022B4CFD33F445EFFF44A056CE3CCE3";
    attribute INIT_30 of inst : label is "B404C3421D0130D087004C3421D03070D0BE004C3423C0C6D51F372B533BCCAC";
    attribute INIT_31 of inst : label is "8103403F030CD0B130C34E3FFCF0472463E0914C01C3420F004C3422F0130D08";
    attribute INIT_32 of inst : label is "F8334B83CC3CE0DCD8101CB88888120D0344E459070130D423B88888073B8888";
    attribute INIT_33 of inst : label is "63C3F030CD0B130C2503FFC0058D2EF8C38E0DCD8101CB88888343D0DCD3C3CD";
    attribute INIT_34 of inst : label is "0200894D51CF0FC0C324B130CD0F43734F0F37E08FF838FECC400002008D1394";
    attribute INIT_35 of inst : label is "005BE3794F9E40C8FBF1A0833E3BC83CE798CF43734F0F37E0CFF83CFECC4000";
    attribute INIT_36 of inst : label is "FFFFFFFFFC000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "1780CD02CE2CE80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "4A0FC5F4E43813443C30C3C337C00000F0C34E3B4000C300000F1F74C88CCCD3";
    attribute INIT_39 of inst : label is "355100D02334130008C48CC0C4D52C2C81ED00A09F0D0EE7406E7F0C0217E7CF";
    attribute INIT_3A of inst : label is "4D502E4F720E40B1445F82C0B243934B400F04000C405097953F35004D554315";
    attribute INIT_3B of inst : label is "7451475095D1451D4415006ECF3921F39C5D37F1CE5D7174DFCE7103400D5054";
    attribute INIT_3C of inst : label is "4E33030353354062D462D40CDEBCF9FC3201DDCEF4CC8EFF1FC00000D749C825";
    attribute INIT_3D of inst : label is "4C2039445145103DBB1C7154BBEFF0CB27E4BFF04BA292451401F4620F6F39C0";
    attribute INIT_3E of inst : label is "E145C7700001D0301C5D3003434CC2800062195054415B1D084CC204C811441C";
    attribute INIT_3F of inst : label is "00310D1FBCB542CC55354E084659E0CF3414444440830E3E20C3F209C00D1309";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
