-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FCDA49A1B2060435CD735F28A0864247FFFB11167DF6806FFF118000673FB29B";
    attribute INIT_01 of inst : label is "34AB39933AE2B8F71B6694C80BA8D1FAC2469F82705EEAF000595C35EE2EBBDF";
    attribute INIT_02 of inst : label is "6A42A0B6110B3DC44D22D71CAD04A08DCFBA03C0131C4847218D2FFE777D7693";
    attribute INIT_03 of inst : label is "6DA147E984478604B1CF291708409B6B669A6B2CB7D9F4DADD102DB6FBA62840";
    attribute INIT_04 of inst : label is "FFC17FC16B3E7D977CFA66000227CB32F00EB0779A8487BCC97794D840203884";
    attribute INIT_05 of inst : label is "44A46B4B820120280292C240B4A52BD2A3FB1AD020E9AA14C9EC4E3679FFFFDF";
    attribute INIT_06 of inst : label is "085CFE599C27209112621F33995290B2B7DE779B24105168F2EDA530320524B1";
    attribute INIT_07 of inst : label is "671EA5F30F5EE8D706AF5F47FBB16EEC47467936BCE87ADE2AC8502E6D6AE7D7";
    attribute INIT_08 of inst : label is "AD89EA1B60F80E42A857D39389C6E13826302F6B56854904CCA700A5DE9A2185";
    attribute INIT_09 of inst : label is "6CFD49F18E38D97226FF5517554069112303449D27C9D3C108402A2C924924EA";
    attribute INIT_0A of inst : label is "BEDD319D3E9D319D3E9D21993C92E3A9DCE7393CD986D82FFA8B0504F6DDB635";
    attribute INIT_0B of inst : label is "6A639C7782062BD769191CFFCFA1A73EF3E9A17802502020EEA1EAFC001D311D";
    attribute INIT_0C of inst : label is "49BF7D54EC1F6258D4EB65091340EE247279A2A55686A838A10C0C08C1168C0B";
    attribute INIT_0D of inst : label is "43E7A9CA1FCEFFB6E9934A0900010616D0117E9CDF19D61EA34A4AD9D3D66007";
    attribute INIT_0E of inst : label is "82AAAAA00000AAAAA02C080114002C082100002C08310C149B92DB4A68A710F4";
    attribute INIT_0F of inst : label is "AAFD3CEB09DEEE3A9D460C4BD14005EAB4BB0D60A91D1014BD1AFD6DEDED4249";
    attribute INIT_10 of inst : label is "4A934DA46C5A3B0020AB27682B689800A25D57A8EAA3C29B0B1D8968D2AE2E9D";
    attribute INIT_11 of inst : label is "2480C0D6428A5CAD9A397ABAEBAE9AC88B6F4A002089249249A4014113493493";
    attribute INIT_12 of inst : label is "EC62893FE29260A9E808519A8061052A51AAFD1FBEEB4623E47CCF99E2BA59A1";
    attribute INIT_13 of inst : label is "A8BA8A28876498708445398F78124800000000004EAD0F5E75FC62D543814E93";
    attribute INIT_14 of inst : label is "3D34ABD30C65BD9E997DB35E4F9BEBB1A7346E62300252C2C2CF5AA05228A28B";
    attribute INIT_15 of inst : label is "882113A5411290BE318C4000F1884022237013878A00203BB406EC081BBB3DBD";
    attribute INIT_16 of inst : label is "7D0EA48E9F4CC3A29312BEE9C68E2E6F34D3F7BF269BE4D34FFE495FE69A4E79";
    attribute INIT_17 of inst : label is "A7F08F1A0C2166A77228FFB9C35BFDB7DB36095E96BB00AFF06D11A991ADF27A";
    attribute INIT_18 of inst : label is "79FE188CBD9D808C2D2206FB57DB7F7EDB10800815EC20C0A054B04094608022";
    attribute INIT_19 of inst : label is "14EB260462DB2A12000D5B2A195DB5640802CC5B580780A2BFF7ECBEDE63DD61";
    attribute INIT_1A of inst : label is "13082958EC25221AB33924920924920924924900920AEF520511AB8184E19889";
    attribute INIT_1B of inst : label is "45555C7A5A68261FE02D8A8060A2004083001020C00C100C404F174297FBBB4D";
    attribute INIT_1C of inst : label is "4104219D50B5FF5FC16B01A8491082400104015A6E80A0B70608998418540021";
    attribute INIT_1D of inst : label is "C4DBD209467F6D18AF9351EC02A10FD0B1E580928442017096D4BB3DDDC3540A";
    attribute INIT_1E of inst : label is "3C3A46BC8D0A95AB69371CC429B75057D4C30E737513C8EE85B9D529BC7ADB69";
    attribute INIT_1F of inst : label is "6E226D5AB89DB301F1E7CC8357188AB1CDDDBE0B67A9459D03D441361F2BFD74";
    attribute INIT_20 of inst : label is "96F2DA536C96522835A4A72FACD55555587FF4BC2CBF98F94AAA015262874A00";
    attribute INIT_21 of inst : label is "0C5EE95A2E84602082942F5979843B640E0DACAD65CCC30B4942BAD3576DAB36";
    attribute INIT_22 of inst : label is "D0F9A13500A87CA3947F87FFFAFFE12057151BD3D3A136405517FF2FDE9D2015";
    attribute INIT_23 of inst : label is "8B6D034E59B8C90AA833F3C50A00415B06091D27A85D0A1A094E4588510556E8";
    attribute INIT_24 of inst : label is "35555555555FFCFA80F5A162E5747293FDA692F2E9BF4ECA95FAC070D850C482";
    attribute INIT_25 of inst : label is "A86342EEEED4F7A200042509053C74A92BF8A49EDF44EADCEFF52751D6EB4E7A";
    attribute INIT_26 of inst : label is "0C9B60D9262FEFC2000B2FD60A71A74AE4E9499A5BA59B4A2306345AD28437A5";
    attribute INIT_27 of inst : label is "998685810458122599264892448160D8366C8B2188E209AA2E8B2289BA288B32";
    attribute INIT_28 of inst : label is "0801C13454013A2E1999A96EAA5DCED5C01BA48D5FA90298C5A068F2E926AA03";
    attribute INIT_29 of inst : label is "0D8173B374EDDD166864AAD2D4637DCCB2B5322FFC989C02E0B745BA2E198020";
    attribute INIT_2A of inst : label is "E6F245598F4C4835052E1609C44ED5D1EEBBA3E6AEBBA3D83611A1833666C0B6";
    attribute INIT_2B of inst : label is "460A928B3A44259CC5B4AA3EB0B7D5100158AC5632802090AC5625C0A43F9BC9";
    attribute INIT_2C of inst : label is "3C52B8B894BC04253694073410F5A5DC700272AA9FDD5AE9D5DAA0185A701797";
    attribute INIT_2D of inst : label is "944AAB51A8EFBCF4D2521A1B9FA583DA6B1824D574BC47B48D4A0A31138484F1";
    attribute INIT_2E of inst : label is "7C77F77464798448C4C4017B2F7B6F5C2224F93E4D767AFF5E6A1CAA01EF42E0";
    attribute INIT_2F of inst : label is "F0298A4B82F4390A03B4FF3F8ECC8515EE678766C0024E066C69B6D46E777F37";
    attribute INIT_30 of inst : label is "FD07FDFF7DFFF507F5DFF5DFFDFFFFFFFFFFF7D7F7DFF4DFFCFFFCFFFCFF0000";
    attribute INIT_31 of inst : label is "0F3CC36389C263091DD73F9E3FFF35F37FF3FFD3FFF7F7FFF7FFF5D7F5DFF5DF";
    attribute INIT_32 of inst : label is "1A3A91C7901E1E930210A116639E78EE8CF633B3D3113D38E8A79CCE3450A550";
    attribute INIT_33 of inst : label is "92B2564B6DDADD51CF6F2F6DB66639E76FF76D772F327AA4DFFF5755359A498F";
    attribute INIT_34 of inst : label is "043443002083231EAE4B288C23D8012057FCD8BD1800026D81E7CE9DB3566D95";
    attribute INIT_35 of inst : label is "0000A83CF3E040EBFFFFFFFE04385BF360000000000000000000014090803002";
    attribute INIT_36 of inst : label is "FFA8FF9FB54C600000205000894EC0000054219000000890C200000A04E88000";
    attribute INIT_37 of inst : label is "D974E4647419193D776A9391D3D351115158862511BC61D80BFFFF894327FFBF";
    attribute INIT_38 of inst : label is "E6F66F2F02368440429699BC029A0605E5E0400D20604A08206698000EBCEF5D";
    attribute INIT_39 of inst : label is "235042230B1BC8696D33E315C4A52B58ECC66C806A0F1704E5143968A9BC96D9";
    attribute INIT_3A of inst : label is "F2A70302B2928C100450A62C4C28020A267DDACE4133E564E3452D0008808800";
    attribute INIT_3B of inst : label is "DFBF793A87D24A4C44496D7D76C4D34457F6C5F137BD480A800B450015FB4A04";
    attribute INIT_3C of inst : label is "D54C3B4D707D9B56CD750AA1512E8B48EDDB759385DA242C40747C40466A1554";
    attribute INIT_3D of inst : label is "5692FDB35DA0E52DEE62C7696F7EC54E7E08854E7942AF3A4564D4BEEB97EC3A";
    attribute INIT_3E of inst : label is "A2C72158A46DD305E352D6ADBEB55C737AD67562E530D4B08243B2B319AD15CE";
    attribute INIT_3F of inst : label is "38447F060C031D61E0BC17F03661466200001010A3F22602176A8D0B212C1809";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C125925E871715040140400D12A08754800087881699CA0000068020E06F9629";
    attribute INIT_01 of inst : label is "4B828FD9802649612D89330187B1C4984BE001EFBDFF03C11119EC749D832DA4";
    attribute INIT_02 of inst : label is "6F4CF6F04892AA0499C1938D9F17AC0A82A05D892C762A0332C6090713CE8B64";
    attribute INIT_03 of inst : label is "10C8680FE3B033A86620667D9CDBC910502890116822D224928F092182D65459";
    attribute INIT_04 of inst : label is "0822894A298128C200512391EDBC199DF0105D4244DF6F8790D83333824A53CB";
    attribute INIT_05 of inst : label is "BD7AF8F87B53B754293BAECACE7BD48B8A06017B7A044F2A588C930C32001040";
    attribute INIT_06 of inst : label is "80EC0DDE3D1097426D8C60007BBE3C6D6CB7DDF21014451AC0A227EED7BC918F";
    attribute INIT_07 of inst : label is "4409F34A8499B15D889A348AA627C3B9F18A82F3A5AB7F32FE208304C0AF7E89";
    attribute INIT_08 of inst : label is "29EE876839E6F6258CC1E15FBA5A13F67EF3613D234A1F9D07E827E91328671C";
    attribute INIT_09 of inst : label is "8E02FFED659644978A1057659AE52DD2832570001880002239847AE492492459";
    attribute INIT_0A of inst : label is "5924CE665B24CE665B24DE66DB6826FA46318C40101A5FB81FF5C75A4DDB7779";
    attribute INIT_0B of inst : label is "8CE72CE19B206DEDDCF4B2452452B4114900AB1391D9B3AD64FC8FB49934CEE2";
    attribute INIT_0C of inst : label is "5468A1A82285A6280E92249180681B000B100C9526BABBABCE8C94B6AD723E5F";
    attribute INIT_0D of inst : label is "2C70FA0590030891265C3D925D234D2D1E7D42206050037061DCDD90A1C2A001";
    attribute INIT_0E of inst : label is "980000000000AAAAA0180D0010C0180D2000C0180D2008CDAEB54EC57BF34BD1";
    attribute INIT_0F of inst : label is "5F69D9093A215C8E11F957359AE9BACF6A38E19D5479EEA939ECA50D0D0DE6D5";
    attribute INIT_10 of inst : label is "D8012C82FAF1E60AC91D6FEF8E2E41E23364E9B45B2249D372424F5F5F4BCBC2";
    attribute INIT_11 of inst : label is "F6E8CB5AA3AE8512617FCA0802800A011D223C124ADB69BE9BE82495B6D37D37";
    attribute INIT_12 of inst : label is "0506CE1A05CC0758CF79CF39484A37B92A4400C08209A99812020000000CD0BB";
    attribute INIT_13 of inst : label is "C00C00006993A886109C99A3A581016DA0A090000DBDDC02948FFE00C508502B";
    attribute INIT_14 of inst : label is "0635D0636D7881A21A0434C8581936DCE9AE33664496CB7A5A576AE2D8000000";
    attribute INIT_15 of inst : label is "1871DABF084BDB58A52B5F778A52974CE4A22D4A55736F0AA683B85E0EE34686";
    attribute INIT_16 of inst : label is "40244904105131252454124A6936DCF08924111A8B2C026591B0256951248000";
    attribute INIT_17 of inst : label is "7A8E48A3112209BD0A4D0467141F2619488851B24A4D2B9245C578980C110430";
    attribute INIT_18 of inst : label is "DA88001580A3070CB4A63975CBA91E00022A15978E4A520D9F39021258EEA605";
    attribute INIT_19 of inst : label is "7D1D6F6DEE210B4F0007A10B57C4AF40AE583DE9465E4B0C1E10C45D46412797";
    attribute INIT_1A of inst : label is "82519DD95718F9EFCD482402410090490410402492410F7BF68CB4970B0E34F3";
    attribute INIT_1B of inst : label is "2001F894AED16F320E6427ADCBE9C4C9AF39226BCC3C7338CD8333E5A4CC891D";
    attribute INIT_1C of inst : label is "64BCEFE18F1001A1B62D26FC9A339986673333CC22319C433E725F92D7CA124A";
    attribute INIT_1D of inst : label is "10006DF31DC0EDA167BFEC04DBCCF04FB20B3668C67CB7BB38382812D2CEFA21";
    attribute INIT_1E of inst : label is "EA504D09DC1102BC35AD4A8E90857DF933CF310AAC8BB77F1265FD76090154AA";
    attribute INIT_1F of inst : label is "F1D4330162422EA0809442C820311BA82367FD314411A6099EADCCE10986BFE0";
    attribute INIT_20 of inst : label is "218C29DA4D005E2D61CAE8089860079FE01FEE27C00B8A25C3F9C42B667A3CDF";
    attribute INIT_21 of inst : label is "1CCC22CF1B28E42419DC902602FB85B7777080040109432963958C29B4D25E6B";
    attribute INIT_22 of inst : label is "B2B3B9402E01B40680C019FFE8FFF25D85D9C86DB7FA443B5C87EA834B7B5D83";
    attribute INIT_23 of inst : label is "9F9B5ED941A49DC3B7B33088FE1492132335E542F2165C8A855FF36083BFEA39";
    attribute INIT_24 of inst : label is "5980079FE01FE5F88A0FB1BB761C184048024823CFD9D0FE2C2BD77E0331CF50";
    attribute INIT_25 of inst : label is "1CB8ED1000703ECB4B6F8C422E42C4F5AD897CE800A0141C7F86B6B2E02D0326";
    attribute INIT_26 of inst : label is "090A0498A24FFE3DE00667DC553D997C86A23E2C208A098DFFBAC6D1D9899966";
    attribute INIT_27 of inst : label is "1006C90200902609924098A0098A4091340D9B6759D06DB30CDB348D2B6CDAA4";
    attribute INIT_28 of inst : label is "FFFD6ACEFADBADC3C601A322A8C903FE6C91C556C6406404C8B32C600242BEFA";
    attribute INIT_29 of inst : label is "E07A07FA4AADC785DA0F957E2AF7F769E5FF8519D58DE950B523E93D43C27FFB";
    attribute INIT_2A of inst : label is "B45A6CC1BC37BA6810B644A19F03F06A8DF0718F8FF0F18F81AC3CF8EDD03D23";
    attribute INIT_2B of inst : label is "E6195AC2460E73E0C8D38DB83EC83F2492F178BC579A493178BC43A616A29968";
    attribute INIT_2C of inst : label is "3E758B8BA3CB636A8206CB113437EFFD80030022C15118BA3D6AF3D435625D0C";
    attribute INIT_2D of inst : label is "9CAFFC2D36A498E009094140364FF79CCDE178489B8D9B6CCC8CC3563D6646F9";
    attribute INIT_2E of inst : label is "0AC1DE02D38E607063124F94719C310EF7800000007A04A0513020AF7D5626E2";
    attribute INIT_2F of inst : label is "CC97044908761FE0F12E7D136657475D7BAA78984BC46F612AB0DF009986B80E";
    attribute INIT_30 of inst : label is "55057DFF7DFFFD07F55FF5DFD5D5FFFFFD7FFFFFF7DFF5DFD4D5FCFFFCFF7867";
    attribute INIT_31 of inst : label is "E88200E86C1414DA02083FDF3FDF3FF717F3FFF3FD59FFFFF7FFF5FFF5DFF5DF";
    attribute INIT_32 of inst : label is "7863930CBB3284008848840C04228FFEAE37533893A1A0AD057003E0C6194579";
    attribute INIT_33 of inst : label is "81B03606D8CD77AD0F1E5E5BFD6D140FFF8001E1BE5B4F43E4A0232A1A40003C";
    attribute INIT_34 of inst : label is "820C908008500B2C8C23DB1B93E00A3047FC598CDA08A82EE8618005B036058D";
    attribute INIT_35 of inst : label is "00009414516D389000000002F68807F10079E781E0781E79E0781F3B5A860800";
    attribute INIT_36 of inst : label is "009C00404CE50000002D3800BCA58000005ED14000000BCA5400000BDA414000";
    attribute INIT_37 of inst : label is "4AF0B0B020B82C2CC732C2C2C080C0C482C9B3680C15094B800000B4A2800040";
    attribute INIT_38 of inst : label is "C909109CD37DB9AAD7B208D3F5BEAEA7878A4B5B6BFB5CC964E6916C9E9BD56A";
    attribute INIT_39 of inst : label is "949F64C325205AD373670627DC4CBD1A12D192C9B85837DCE9038FD78089B014";
    attribute INIT_3A of inst : label is "063026254ED91DD4C0A2511A20925967EE9FEB31CF740BEED4DF7A4A52A52A52";
    attribute INIT_3B of inst : label is "E24824CBBA1E707DCDF3838490531205F18250C3BEE8EC0A8009DAFB684DED9D";
    attribute INIT_3C of inst : label is "38A806424B1348F420DD58F2F3089E2BEE04004CA07BD290CAC280C8CA80E416";
    attribute INIT_3D of inst : label is "20A1C1283634191B8165C088DC09C970CBCD4970D6688BDF10471ED921D92AE0";
    attribute INIT_3E of inst : label is "911DB35903407DB7DA7B01D4501E00302039184002A0E050412111020802A565";
    attribute INIT_3F of inst : label is "720B28A11CC73434FBEF7F943022F0286265D452F1F0622B2D0AC54463B63CA1";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "8564964A88193901601807019120C394028089967B65C22EFF080040A00F0438";
    attribute INIT_01 of inst : label is "C9930C93A16018430C8970088220183282E105C738FE3299939174303D874D08";
    attribute INIT_02 of inst : label is "2F5EFCF88CEBE1C750DF3EC76AF33A6EE77B1AE00F6A320D21C327A4B21E1B24";
    attribute INIT_03 of inst : label is "4B68CDB27367B334FDE7659AC064F6DFECF64B6D925D66BFED2E25B2FF342D53";
    attribute INIT_04 of inst : label is "D7CC9C33409705012E0B1B19913DD88F0000194D9399257B29F7B1E3020A3EF2";
    attribute INIT_05 of inst : label is "9C73BC9C9EF3C3982A789262C63CE65B8EEC007872593BCDF1E8285FE62DAFD6";
    attribute INIT_06 of inst : label is "8072AD9E29949E7887733881C9ED657D703BEEF88550101F81F612EED19E77CD";
    attribute INIT_07 of inst : label is "E673569BB9C311C8CCB0E9CC088F1303C18EFB470F084504D44C5A8F8DCA0942";
    attribute INIT_08 of inst : label is "0442853C13F4F4E7CE15039FBB8E1382F082703E9F0F1E1DC76F732D0E18461E";
    attribute INIT_09 of inst : label is "178E6D6B5D75C0DB231FF93F99844E1043214842008200A2318650F49249245D";
    attribute INIT_0A of inst : label is "6DB36BDF6FB37B5F6FB36B5FEFFAA6FB918C6356788F4DB479D187962912445A";
    attribute INIT_0B of inst : label is "AEC1C839019C2E0AA5296C34D3039B0C30C00B131981838D0E71E70091236B5B";
    attribute INIT_0C of inst : label is "157D2DC0838C43CCB7EF424FA24123309399BA6DD8E4A9C1DA088464B964EB15";
    attribute INIT_0D of inst : label is "C840FB0292E21699871E70B4DA338E2DDCE0BE362B7007E013B899D64A5D0E44";
    attribute INIT_0E of inst : label is "0A00000AAAAAAAAAA0080002D8AF0BC032CCA708C0A2D8A9202404C55250F213";
    attribute INIT_0F of inst : label is "92A1E10AA7C022A609B19A335C8D19AC063FA3514B3588A6B58BF96969E9E0B1";
    attribute INIT_10 of inst : label is "9AD36EC672B1CF0A8A3BB7472D4E44C09380E8361D4C48E2E3D442340D0D0DD0";
    attribute INIT_11 of inst : label is "E720CA5304B32E64C12EC3430AA2A30B33B13A120A92492C92C8241524925925";
    attribute INIT_12 of inst : label is "AFCCEE2FD9C639D46C338E2C60AE83C38533E63CF3C794CF99F11E27C4FEA130";
    attribute INIT_13 of inst : label is "9FFDFFFFA113BCD6B4C8C1C4DDA92524800081200114B452F437BF15C61E5AB9";
    attribute INIT_14 of inst : label is "BC24CBCB2E672DDE59FE38C21B0804086C5958432CBF6242436552A7E7FFFFFF";
    attribute INIT_15 of inst : label is "9440D73BA111E30294E50A7339CE71EC46723B8B9E324C0DD603745C099B3CBC";
    attribute INIT_16 of inst : label is "7C4E2D8E5F5CC3A8B6563AE1A62AA31BADB6B225AFBEA2F7DA440776B5B6C328";
    attribute INIT_17 of inst : label is "25F4489A94434735C2E9456B77496F5C7C708516E38628EAD45D1CB45DB9F66D";
    attribute INIT_18 of inst : label is "D6CE7B9EC3BE220CA52028C2C619960C393999171866798E9D65B844616F2F89";
    attribute INIT_19 of inst : label is "ADDBB7250B152B0E0006952B174499A0A851A14C42D04A682651C824E4513F97";
    attribute INIT_1A of inst : label is "04649E545798E9CD47712090482482412082092492410129261AB0950A053843";
    attribute INIT_1B of inst : label is "89D8BC0D3CDA4841E8A4276599C944C9A831226A0E30622088C203E7B4387997";
    attribute INIT_1C of inst : label is "866B52C8DEBC2F99E7C622FC1B23190646322269E221984C30E3841C9768128A";
    attribute INIT_1D of inst : label is "9C48CE321BAB89E66864BC10E325E10EA189B664633997AB68E87D0E31DE9809";
    attribute INIT_1E of inst : label is "B20D4617118BC5ABCCFF7DC408002CAC220821FAE9A89BD59E40485E8959958B";
    attribute INIT_1F of inst : label is "0EAA3A13F384754030311A697418992C579FFF3173B86189CB3C88C403E33A96";
    attribute INIT_20 of inst : label is "646C959B4E0D1CAD09E6481FD9801FE0001FEB358DAB1C3CCB5D017C52E338DE";
    attribute INIT_21 of inst : label is "6A44838F09E0B0464BE4C04C19E619A767731818C3AD632153846C958D8EC2C5";
    attribute INIT_22 of inst : label is "3E1FC81564AB01DB3B7FE1FFEA14A499A48F2A6C6C48043373914A9B5122799C";
    attribute INIT_23 of inst : label is "C4965595089415E3C6BFE288D21410E29B31E05212135681322CC894E22AA51F";
    attribute INIT_24 of inst : label is "FE0019E0001FE5F86BA19DC387F8F1C0BEA24AA14FC7DE771DA17A1391C6A250";
    attribute INIT_25 of inst : label is "10AC28E4ECF4FEC9596EA94B6FA76850EE5130D47DD0139CFFD71BD3F4AB0177";
    attribute INIT_26 of inst : label is "4F13C4E91E0FFDC2020443F463BB1675F5363AC9AC92CDAC93D4B745451ADD47";
    attribute INIT_27 of inst : label is "390E830080300E0310E0308E4380E4301E4799C7F97C47B1E8721EC731CC7B3C";
    attribute INIT_28 of inst : label is "AD2DAA454A49B7CD5214BA286E84062A08D0D1DE4AE1461EA419388842C4ACFC";
    attribute INIT_29 of inst : label is "A1BA0DEE7FB69BA5B60B496D37BEF72F4DFABF4175C72950D524E925CDD26D99";
    attribute INIT_2A of inst : label is "140A6EE1B44A5EE904C610A0532129AA4963D40B4963541286AC253849B0DD24";
    attribute INIT_2B of inst : label is "250C52E5C52792B82C398C2D88C39A31C2AB54AAD518E1AB54AAC3C695605828";
    attribute INIT_2C of inst : label is "2A378FCFB38A336FA4965CB13F246AFD8002D001B499943B8092B3E5994D3467";
    attribute INIT_2D of inst : label is "0E015409048A2A6449494948676AC41A89B970BC39819C4846864B0777C262A8";
    attribute INIT_2E of inst : label is "0A00E7CACBCF4600068083FFAA002B10C7002C0B201552550BCD342B3E67C0A0";
    attribute INIT_2F of inst : label is "CF374E1B26FBBEE85BA6F13C6C660966EF7363300F4775700BB0DB5585D79C17";
    attribute INIT_30 of inst : label is "5505FDFFFDFF5505F557F5D7D5DDFD7FFF7FD7DDF7D7F657D4DDFCFFFCFF0418";
    attribute INIT_31 of inst : label is "F1E3808E2F1C1C5604103FDF3FDF377915F3FDD3FF51D7FFF7FFF55DF5D7F5D7";
    attribute INIT_32 of inst : label is "8B0C58715C9CCAA912192101120657285B9DCEAE3AEFEFCF7F5DE73A378C2159";
    attribute INIT_33 of inst : label is "4D6D2DA4884CF69F48D191DA4A58FE0B2605CCE85EC58533E39E93899EA20441";
    attribute INIT_34 of inst : label is "C688C887088823DF1B93E50BF8042C4757FDCC69CFDF5420DC94ECAD692D316B";
    attribute INIT_35 of inst : label is "0000C5C30C215870000000023588555D1F86187E1F87E1861F87E14852C60C00";
    attribute INIT_36 of inst : label is "00AD00200565C0000023580085270000005210C0000008D65C00000A426E4000";
    attribute INIT_37 of inst : label is "CEC00010837400043530000042404606024D124404D5C8E9E000008521C80000";
    attribute INIT_38 of inst : label is "64977F7471393B7E9F3A48D4072CB9A2829E34524A8A4C4266C0890C98D0C222";
    attribute INIT_39 of inst : label is "B6B6318329019ADA7A44DB36266DBD16A2B51673B878D526A5032DC5C8C139FB";
    attribute INIT_3A of inst : label is "E4BC2020EE5C2DE5F129139E14C2C967AAC09B1E8D560DF9FA518C4E56E72E53";
    attribute INIT_3B of inst : label is "818618C1799C72759CF68E8104030869A8F1FC73A35DF10A800991D1C634A19D";
    attribute INIT_3C of inst : label is "BC8E484DEBBC48AFCDA859BCADBAE5EE4828A28CC2A2C2808EC2808C8F2AC046";
    attribute INIT_3D of inst : label is "293317D36B65232B6AC309195B5F59D69FCC19D69F60A39E15165C43A88987C0";
    attribute INIT_3E of inst : label is "93DAB01012001C27DE7C05CFE03FAD1240EFD3522529E49467A2E94A910FEC66";
    attribute INIT_3F of inst : label is "D10020A308420D3271CE3F84264146427325E470B958A41A4AE0086761B61C30";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "84D249208DB8980060500601110203C182C4099769F44011509C0440801F20D8";
    attribute INIT_01 of inst : label is "24825B689D45114A32669168801D94A080E00E1EC3DFE1B97DC854283195592A";
    attribute INIT_02 of inst : label is "EEE4E8D360F0C443F84191C5E8A1DE23E5FF3F610D7B30060185B6F42A55F693";
    attribute INIT_03 of inst : label is "FB208FAF332E933CFD65279EA82CF6CFB6D6D96EDB7B34D2FF8DBEFBEDE66EB7";
    attribute INIT_04 of inst : label is "9A1C95F3795C3C27AAD83A41AC59494CC31C594DBF1D202939F690B908686E72";
    attribute INIT_05 of inst : label is "CC732829AF535788A1F19262EFD69451843411F172DBF3CEAF44BAD2DA2F347E";
    attribute INIT_06 of inst : label is "4863F0C2008FFDF882555CA068C8403C3C1966D8C37388C151E38B0A311CA499";
    attribute INIT_07 of inst : label is "0E9BDDD5CDAB96843D29DD7E6EEA509A88352757AC91A9D05DD4CB76AE731A2F";
    attribute INIT_08 of inst : label is "42C7B47D46FD49FF82FC17D4995F5E4B4EC764A6B17EBA3CB065ABE6BB7C56FC";
    attribute INIT_09 of inst : label is "C58A482F75557352A238FAFF2A836EB3048660280A1684B3B9E579E7B7FF6F9D";
    attribute INIT_0A of inst : label is "359D294F379D294F379D394FB7DF81395EF7BD7C78DE6E64D1933546B6AFEBB2";
    attribute INIT_0B of inst : label is "59E6ECDC94B60A1FA569355165939D565560813455D1E39C9B6D56C4F9FD29CB";
    attribute INIT_0C of inst : label is "0838890EE9001386F7EF1001AA4143A8A3DD3E68F17989CC7B0618EC1C3B715B";
    attribute INIT_0D of inst : label is "478D99C3CB8755D31F6CBEB3597F4D2CAB7A76142A50C4132A0828E288484877";
    attribute INIT_0E of inst : label is "9A00000AAAAAAAAAB46018F22C9E6098C22C916258F22C9B3D679DAE931F5135";
    attribute INIT_0F of inst : label is "1902D812B2002228C29B9433CFC839E7C60277790BBCFC86DCFB6B5FDBDFC4F6";
    attribute INIT_10 of inst : label is "0DF6F6C63065C7086133B4669797448696B5CD26D484EB645552C721485555D2";
    attribute INIT_11 of inst : label is "5561238E2D16053FC10F8327BCF9CD899BA1945868E506506500B1D0CB0CA08A";
    attribute INIT_12 of inst : label is "A8A50E2F3986193CA5B58E04602EB355B5672CE594585514A294728A59436174";
    attribute INIT_13 of inst : label is "8DB88A68832D9E79CF4AE4A4C83EDE5844B659614318C4F24A6E967E764C4AA1";
    attribute INIT_14 of inst : label is "4ECF54EDE53948A70E4C966ECF31CD2AE418522756FBE77F765FA6332A6CB6CB";
    attribute INIT_15 of inst : label is "9B7EAF8320D9AB66B5ED5BB7CA56947C51B2CDDC77F65E1DD2C267EB099DCECE";
    attribute INIT_16 of inst : label is "3FFB64BBCFCCFECD935DEFB5C74D36916CB3F3F56EBBE1F3CA6E2773ED964638";
    attribute INIT_17 of inst : label is "97854C1519D2C5506964210C40404B0C10E40265C086FB20994A69FCBB6CF64F";
    attribute INIT_18 of inst : label is "27DDD2FFD792461218E6FAFB945D25AA75FAF446BAB5FAAD1BEBF8366C3E1E81";
    attribute INIT_19 of inst : label is "64B3B5358F1835655F5C983562EC99E48D1EF3E8EB6F7DA5E1753DA2C92254FB";
    attribute INIT_1A of inst : label is "11751AEDFD66F1B26F295DB7FFFF7EFEFFF6DB7F6DF882B1CAF4D6DB3DBB35B7";
    attribute INIT_1B of inst : label is "933618E3F04B00E383E6F517ED75D0A56C3C295B2DB66BB0EDC4A13F9AACAD03";
    attribute INIT_1C of inst : label is "B6CA52DA2DE939982BFA85F8E96F39ADF6737ECD7780E0BFE95E9A3456CC58E8";
    attribute INIT_1D of inst : label is "F449C618372A76EE68410CB2DD54DB2D52CE0A7478B6DB41C09C78E011DF9C6B";
    attribute INIT_1E of inst : label is "E2BA9D79EA98E90C58B2BED43050C888871C79C776C0144CF66424069B49AD97";
    attribute INIT_1F of inst : label is "18CC6AD49D8D3550B8AD705C7C53BF4ED1B50334CD3ACB00AE19E8958EA62C9A";
    attribute INIT_20 of inst : label is "646C9DD7DF861FF941AD611CC01FFFFFFFE018298CA09F12C89D0D353569972D";
    attribute INIT_21 of inst : label is "F6C4A85008C0101751AED87C01A68F6A7D794C4E63C9848223C46C9D8DCEC6E7";
    attribute INIT_22 of inst : label is "C28C5D7FD7FEC593326001801B42180A84ABA39302001415B9FEB4C95EDD8AFE";
    attribute INIT_23 of inst : label is "50403000A1C4EA625E0E581CB210C2C5BAB4CC34E811120777333738C3128441";
    attribute INIT_24 of inst : label is "401FFFFFFFE0100718911DC2853560C16CA2478B088CCA8604980D2C11EF6941";
    attribute INIT_25 of inst : label is "1F9906F5577B05A52DA56718C7C77548CE342AAE14A052808FBF18715CC705D4";
    attribute INIT_26 of inst : label is "08900401326FD3FD1C0924C572174585D3B495ED1ED1E9A59FB5EEE0E0F99C7F";
    attribute INIT_27 of inst : label is "89228C1104C1120C9124C9924C010048300C832281605C2F2ECBF29C330CCB22";
    attribute INIT_28 of inst : label is "840EAA110D25D715D09C49EE52784188CAABA3FB6AE7FE7E6C0B178940D58EEC";
    attribute INIT_29 of inst : label is "A2BA18DAAE922BA524200380462480358C48D542032442E55508E84715508015";
    attribute INIT_2A of inst : label is "E773DC4C3A79C14D35DE50AC19260AAA535554A2535554A38AAC262803215D28";
    attribute INIT_2B of inst : label is "939D6FE5D3279394BAB0C57E84CA5D78E3D3E9F47ABC7153A9D464B1ADE397CB";
    attribute INIT_2C of inst : label is "D4F2D5D39962A4E47F9A9CB8EF77265CC032F3C4BF111839596637638C7D2463";
    attribute INIT_2D of inst : label is "E2E1110B85EFA63448C9C8C93563C7FAFDF3ACEAB0D3ECFE9E754D7EF20D8FD3";
    attribute INIT_2E of inst : label is "C1C2E7C1C3CF37FF368012001E001F104100681A0711F81C2FC25E63364DC552";
    attribute INIT_2F of inst : label is "CF1BC5D9E6419046D1866711E6C45A2CCAAD6EF22FF630232A68B2FF5587DD07";
    attribute INIT_30 of inst : label is "5D05FDFFFDFF5D05555D55DD5DF57F7F7D7F5FF557DD555D5E757E7F7E7F7E77";
    attribute INIT_31 of inst : label is "B2698206874C4D0E1DD71FDF1FFF1D755F797F797D755FFF57FF5575555D555D";
    attribute INIT_32 of inst : label is "A74D2A6B2FD84AA88000008008D7539D0783CB1E01E0EA67521D603B2BA5731B";
    attribute INIT_33 of inst : label is "2DA53587E0A4DC98329BDBDBFD2C474091AF3A788F88D922F399D2A9430A04E1";
    attribute INIT_34 of inst : label is "00840801040013E10BB8005EEEFC300742A83C103C0A2241748C58A3A835128D";
    attribute INIT_35 of inst : label is "555545122889080003748B7494B0500D678000000000001E0781E00A52408020";
    attribute INIT_36 of inst : label is "F005FDBFB028C37333090A7624289FFFFF929000000002428C33266252AE5555";
    attribute INIT_37 of inst : label is "C150D0D0D19034305D16034303014703434090241028C027B2AAAA242001F803";
    attribute INIT_38 of inst : label is "2DDE4DBC1D1812660C195000040060799983A4400606CE77D6FB65BE968F5FB1";
    attribute INIT_39 of inst : label is "D67596848E6348486CA0328A25E0DDA29714B879E9599FE5F80F0DC48A9013ED";
    attribute INIT_3A of inst : label is "905D0504E9ED87C3D03919A812DF6DBE6666F329A733CD9D9B1CE36B5F47F47A";
    attribute INIT_3B of inst : label is "238EBAD99AF6D2D0AADD08C30D2B4241714288A33F0CD72AAA6FB9B7F87D187C";
    attribute INIT_3C of inst : label is "920850EDF1B9488BDDEC09BC8D1B7157C238EBAD9AF9C981EDCB81EDFEFFB444";
    attribute INIT_3D of inst : label is "750B96D77AE540A9FB24AA054FD5B8FE7466F8FEEA37B569CDA59362CE6E6128";
    attribute INIT_3E of inst : label is "2B5EA3B9F23D55240E35C4891620182A488104287414AEA8440A43A9458804AC";
    attribute INIT_3F of inst : label is "5F0E380004A1252787B0F7F63170415B7B63C2D03808360808266C25717528A8";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "052592488399990842509715BB22D798D2D2C3E816492B2555840260824000E6";
    attribute INIT_01 of inst : label is "49841A4895775D03AD993165C0391C3E2D708594B28133D311DE935829171C0C";
    attribute INIT_02 of inst : label is "2EA4E4C1A8BB82849440128510412C6F92E8510DA853722DDB2091303059C96C";
    attribute INIT_03 of inst : label is "A0122A4A20A800AA02009024EAC904B04260269A2C149848B0A91900168177F3";
    attribute INIT_04 of inst : label is "28B2CA9A1049013192034B5560B02489015545412856DD4014004A06815D515A";
    attribute INIT_05 of inst : label is "694AB0B00A771B082575248AF3148423080815350B02856A528294C022825121";
    attribute INIT_06 of inst : label is "C01808B02900D90038A400F222ED6D2124924492D0A4D691B086C20A05580142";
    attribute INIT_07 of inst : label is "59C9DB4E64E99E2CB35934B26667DF99FDF18CD9E08B05D0DD8C1ADCA3090008";
    attribute INIT_08 of inst : label is "70C685604420042D40E15D07D75808E11CEB0A0D76DA121AA154AADD80204618";
    attribute INIT_09 of inst : label is "96B1B346BA6BA00DC0906264162184EA441CA9E2382E23B731EE50C2A5756E54";
    attribute INIT_0A of inst : label is "61B2085763B2085763B208D7E3FC3B170108423C50D80049052EE0FA00100440";
    attribute INIT_0B of inst : label is "20D522A550216AA4BDEDE38E38E318638E28CC8C7581C70C686906B2FDF21853";
    attribute INIT_0C of inst : label is "912080A83A10E4200E82E6CE102258192840AD19319D558CCD8852BD0F203044";
    attribute INIT_0D of inst : label is "1EC537B4990449069428AC361B66492A935A414824506910209190A261018461";
    attribute INIT_0E of inst : label is "5C0800A0800A0800AA228A12B8A722CAA2B4AC220AA2A4A37F6F95AE535EC7AF";
    attribute INIT_0F of inst : label is "1030E1B9310804A669807E34123D3A096800C8C7562123ABA125121296149400";
    attribute INIT_10 of inst : label is "94D34901F205881D45860194AC4CA1231820980F24484CC00018F7B06C0000D8";
    attribute INIT_11 of inst : label is "10410528290420DA10EE14220822AA05D04404154952C96CB6486A92E492496C";
    attribute INIT_12 of inst : label is "208FCE1A0D6C0D00CBB78C29488A771721AAF11EB8EA0623D4788F55EA320078";
    attribute INIT_13 of inst : label is "1A61A6DB16C532D294CCDA650929205964A48165B018EC85C686B415E60C8AF3";
    attribute INIT_14 of inst : label is "E053BE0CD39E627067A04D12A3227DE14DCF94144D9884343C3475530E9A6DB6";
    attribute INIT_15 of inst : label is "DB689A0A08610E5B7B9ECDFF37B9EDB5D4E3E718DCAF4C2205E080E38204E060";
    attribute INIT_16 of inst : label is "726905E91CD8AA4C167F24914575DC0284B7F62586BFE653DA4E4672B096C638";
    attribute INIT_17 of inst : label is "822542A33D9DEA310EE41631850D26584D509533620CA98A45A170801109C6F4";
    attribute INIT_18 of inst : label is "6590E7330654751053D5DA2810C06320666B6644D298D379524E62184ADF3F55";
    attribute INIT_19 of inst : label is "6AC600C9CCAC14C1CBE2AC14D0912241DF2F3982935C6B1F938E639214626192";
    attribute INIT_1A of inst : label is "0453B8D1002695214CA25121A4D34CA69344921A6D22703185A62D1219822432";
    attribute INIT_1B of inst : label is "311006E6349BD97A2CD811118444D7AF7EFDEBDFADF36EBEFD82226D76C1D055";
    attribute INIT_1C of inst : label is "3CB9CE30297120AC2B3114BA97671DEEE67B37910082203A5C323751F4961549";
    attribute INIT_1D of inst : label is "30028712600C8981402C805B927695A94B961A5C7AA49329454C200000002631";
    attribute INIT_1E of inst : label is "A0724CE941863C2720CDCF0892F2A88C235D732CECCEFC59B0A7664223039ECF";
    attribute INIT_1F of inst : label is "A089C8CE6E694440888C28743A2911EA8340C3348E130C008E2BB8928D264286";
    attribute INIT_20 of inst : label is "294528AC93699F4002A06D091FFFE00000000045480087A8C050C63147DE0769";
    attribute INIT_21 of inst : label is "38C6BA7C2808A4453B8E932113DDD58AF5F254D2A1116404FBA54528A894544A";
    attribute INIT_22 of inst : label is "63449D552EABB110A2007E000214A10AC9BDA3262449141558514AAD11226AB6";
    attribute INIT_23 of inst : label is "B016E5B1A0C0144010C440E8263B8E222BE5A65ECA50810CCCCCCCC2EB20A811";
    attribute INIT_24 of inst : label is "5FFFFE0000000007080E9DF2BD594D1000408C214011BA14280D09D8D5638864";
    attribute INIT_25 of inst : label is "4194A598000202C10925A508200FC644EF00EBA800E41420001F1EA9490C4144";
    attribute INIT_26 of inst : label is "600A0209802FFE32E0013B01E48508148A030500D00D004B4C614984041B4008";
    attribute INIT_27 of inst : label is "E03A428084812240900080A00000200908621884288872188229CA628CA229A0";
    attribute INIT_28 of inst : label is "BDB40B4779B783485A4E830760C7CF286A14184682C2542C8802253003515468";
    attribute INIT_29 of inst : label is "690B4528023691B1B68B076C0F9244208F26216156A76BB405A46D0148DA36D7";
    attribute INIT_2A of inst : label is "4B25102715108B6A18916097180B290B4112C69943124691A435151A4BB48D84";
    attribute INIT_2B of inst : label is "B5515D406C1ED2332A040BC05CDD2279A6211088693CD3E1108870618B992496";
    attribute INIT_2C of inst : label is "C92E4D097048849CB485DC09BC3E1AC38E20000500AAA5173CB55342AD06CAAB";
    attribute INIT_2D of inst : label is "40BD50AA55308B4810909190529A342681B38B2A840ECC01006442CE6B519124";
    attribute INIT_2E of inst : label is "E1E908E9E83040004112CE00000800C7FF06100400480301A0114255243A340B";
    attribute INIT_2F of inst : label is "322E8AAA3A8CA72AAA4AA62DA800520910060C843C2735219039DB548002A338";
    attribute INIT_30 of inst : label is "A60AF7FEF7FFA60AA6BAA7BAA7BAFEFEFEFEAFBAAFBAACBAACBAFCFE7C7E0C30";
    attribute INIT_31 of inst : label is "A0A2808A2D1414423BAE3FBE3FBE2EF2EEF2FEB2FEBEAFFEAFFEA6BAA6BAA6BA";
    attribute INIT_32 of inst : label is "62F3579EDA610107001801800E24D34A42B1500A90ADA00D0054012B8681D2A9";
    attribute INIT_33 of inst : label is "436C6C74980D48AA2636363248599D0BB70408130130255A2474786282F4B826";
    attribute INIT_34 of inst : label is "C00800810C0038005EAEFAF00104405757FD4CFD675FD63BA21B3709672C616B";
    attribute INIT_35 of inst : label is "9999B5BF5D75A9333044CC475AB80554782EA7A9EA7A9FE1F87E1FAD6AC00C10";
    attribute INIT_36 of inst : label is "3CD53DA7B6AD41B0E0F5AA5ED6AD0666666B5242AAAAAD6AD4E0E5ED6AC35999";
    attribute INIT_37 of inst : label is "5FF4F4E4E7B93939AF65D3939391D3D393DB775919F54A61D26666D6A4C79E4F";
    attribute INIT_38 of inst : label is "820422C068F921AC91217911B52488D0120D1B52588D9766C490C1D9DA049C22";
    attribute INIT_39 of inst : label is "9E99054414B430BEAA444C5799813040C606325DB17064588808029550396010";
    attribute INIT_3A of inst : label is "C4B49415284B5BE7EAA251E052924924FDC2237583EED383068E72CE76C76C77";
    attribute INIT_3B of inst : label is "6B2C306D0A34D4D088D454955441A4932B93088F2C09C4BB99ADBA156AEC9D1A";
    attribute INIT_3C of inst : label is "2026960049E41889924E407282211109D6B2C306122561298F63298DDC2AEAAD";
    attribute INIT_3D of inst : label is "0891BA44931650123517328091AB21288A49A1289A4D2A531151464229C9320D";
    attribute INIT_3E of inst : label is "8014AA0576DC65A198716910434820210D305A534328484400B1084298D3090B";
    attribute INIT_3F of inst : label is "574F6CB152D4BC72651CA042003AB02DBEF1E4EB555553A5ABC006505A3CAA85";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "0924924BCBDDDD2088621825D3A467D2CD8A978930814A68E903006101804997";
    attribute INIT_01 of inst : label is "49D66E4EE8862104248939B9AA73627B49E01995B2A1676555B89E5EF9CF4810";
    attribute INIT_02 of inst : label is "B58555C6CA9F9285A2EB56B1380B65DF0C84DC892E63BA7F138A9260C0228924";
    attribute INIT_03 of inst : label is "B6C12ED26CBA04B0630C1E78C8DBCD96982D120A4C024A4182490104248C4575";
    attribute INIT_04 of inst : label is "6C46F00B8C1983D8330687172D73076B4196655A6C524FE060D20C66424E634B";
    attribute INIT_05 of inst : label is "294AF6F20872936029792CDA63108507290919790AB6C52C8118E66DBB36D89B";
    attribute INIT_06 of inst : label is "0000CCD8BD2099433026519542FDF48980C611814AA02A99E39EAE1E455BD123";
    attribute INIT_07 of inst : label is "B125412A12D5590AAA1412A955468D51ACA94A0994495A2E343CBB10129B87B5";
    attribute INIT_08 of inst : label is "2BDE8A26C41116252593F0AC79A9801002961355764AD75CDBE6BA65D5865F5B";
    attribute INIT_09 of inst : label is "BE6493FCCBAEAAA4E157C2ACD32314A260242723C8C23086FB8576DEEB534472";
    attribute INIT_0A of inst : label is "0A90DEF088D0DEF40A90DE7088DA7D5981004010F169ECD725266A4A40200884";
    attribute INIT_0B of inst : label is "A5C518A31D2077E89CEDE30C30DBD8430C21A8CC77C58B6C605A15B99B30CEF4";
    attribute INIT_0C of inst : label is "50804002222200021E800000080000800004643B60BC19904488909585391240";
    attribute INIT_0D of inst : label is "506A5928BD41A26855A92416096ADB7CD24E9190A851511828D3F60300000051";
    attribute INIT_0E of inst : label is "1C080A8080A8080A8F03C05892020280589E000200589E05A0B44E84FAA15449";
    attribute INIT_0F of inst : label is "FBFBFD1CE84422B85B8CDAB8966D5C4B108211CD62A966B2A96510101012A51B";
    attribute INIT_10 of inst : label is "D1FEDA30FA099E1E49C65F64AEDC1B221520B85E05692ACE1E035371DC3838C3";
    attribute INIT_11 of inst : label is "92400908F94499DB02763CC61C7186219C9AA6364A7B7BB6BF7C6C94B6F36D3E";
    attribute INIT_12 of inst : label is "44D45FC145C04593893BCCB958D92B9D2DCEFDDF3EF2B73BF67EEF9DFBB78C32";
    attribute INIT_13 of inst : label is "600600410897D550844AD86AB34820012D208004AC7BC34F6F1BDD944FAEEBF4";
    attribute INIT_14 of inst : label is "034B9834D3181261A6034C428B64060A762830C4EDBCB9B9B9B5707388000410";
    attribute INIT_15 of inst : label is "3862BE9ED8C54A59214844EB921486B5E1830C28C4AEEC05148145F20514C383";
    attribute INIT_16 of inst : label is "6AE184415AD3205E10D6451659D7518406889A6E16C8885B25D496BDC0D10A61";
    attribute INIT_17 of inst : label is "B5044A077D1562B21C64C00020E0022882064B206414930405D368931109A685";
    attribute INIT_18 of inst : label is "822A2411689CA4809086A0118106815588292464B301552952C8063148E7AF25";
    attribute INIT_19 of inst : label is "D4C65E4D29468069A905468074A252A3EC482534224248320808030826AEAA92";
    attribute INIT_1A of inst : label is "8EC97CA3116C9527D5320349A64805269124349B20266EF78C816571E870AF0A";
    attribute INIT_1B of inst : label is "333224E737EAFE4459930181C060C881793270DA4C3872A6A8836CA59756069C";
    attribute INIT_1C of inst : label is "249CE732A91392C22A252494992F9B0D57762A2699CC63210282A89514A2364B";
    attribute INIT_1D of inst : label is "2810CE32EAB511B377B6815A966495A92392724D70A492AF7E78E60000003221";
    attribute INIT_1E of inst : label is "C0E2D80477951A6C83A1A49CB98052BB328A249244C9D80C8914C5410280180C";
    attribute INIT_1F of inst : label is "82EEDD250533A578100081C0E07B7FBF3D0043D960561897B84BB94910A40D6E";
    attribute INIT_20 of inst : label is "736E6DC59158BE048B3360387FFFFFFFFFFFE5653370C242A1F644390D4CA609";
    attribute INIT_21 of inst : label is "91E4624C4704EC6C97CB95302A8CB5AEF776B135872B40206BAF6E6DEDF6F6FB";
    attribute INIT_22 of inst : label is "B3E2115506AAB934268000000E7FE06AC8ACCE25B76862954C97EAA1F93B6AB2";
    attribute INIT_23 of inst : label is "9C1B56D2160B22D911B749A9263C93B467259552428E3C1EFCEDCFD5CF955399";
    attribute INIT_24 of inst : label is "7FFFFFFFFFFFEB0699615BC5CBDBC7069260126FD662CDBD8009C93189291E42";
    attribute INIT_25 of inst : label is "62B23849110908C1093263B9907744E2DEC79151CBC0B962104FDB9F2258190E";
    attribute INIT_26 of inst : label is "21984211864FEDCD0107614569CB333FA898A72632632619D83888E6622B3986";
    attribute INIT_27 of inst : label is "1106C9920098260902641886019064190661184191E6713C4F1B86A1386A1384";
    attribute INIT_28 of inst : label is "BCBF08672996E17043658D32E35C12D508345772728C88C91956662382211D79";
    attribute INIT_29 of inst : label is "6E18276BC27FE086DA4F2F7C9AD6CDB837EEC30DCF97E7F3841820E1304132D6";
    attribute INIT_2A of inst : label is "080531159D21086B11907024B041E618791C40CD791C40E1B80C961BFCD30C38";
    attribute INIT_2B of inst : label is "2C91505E0CCE54DA8AC86990E1E89022CA0502817011658502817A2BD9082010";
    attribute INIT_2C of inst : label is "01322F2B9A5A2DA56FC4EF853C9227208F01600519CAADD981F073CC59424F97";
    attribute INIT_2D of inst : label is "29E3AA2914A8DAEC02020202CCCC698D13FBCACAC86DFF002145624AB350D004";
    attribute INIT_2E of inst : label is "0C0D9C0C07CF53FF53364BFFADF78D69CD02A028080060180D0058072C9E2592";
    attribute INIT_2F of inst : label is "E0992421D0521C8681EA4611A419F2889CCE9DC0ACC7BDE54032DF543034B04C";
    attribute INIT_30 of inst : label is "F60FF7FFF7FFA60AA7BAA7BAF7DEFEFEFFFEAFBAAFBAAFBAF4DEFCFE7C7EFCFE";
    attribute INIT_31 of inst : label is "E49240E92C92124104301FBE3FDE2EFE36F27EB2FFD2AFFEAFFEA6BAA6BAA6BA";
    attribute INIT_32 of inst : label is "3671B38C99381D810210210217FFB74A42713849D499981CC0F309E48E4BC03B";
    attribute INIT_33 of inst : label is "754AA8AC823E6FC6C61E1E16DAFF3CAEFD8C1C9191190A972C763234AF46011E";
    attribute INIT_34 of inst : label is "810C008008002EFAF04104510140806047FCFDA0DB5FFC2581D931834568AA7A";
    attribute INIT_35 of inst : label is "1E1E943E8DE5296A6622AA2252B867F37E7FFE7F9FE7FFF99E6799294A810800";
    attribute INIT_36 of inst : label is "3F950FE1FCAD204BB12528BA94AFC969694A52D4C19CC94AD2B10BA94AF15E1E";
    attribute INIT_37 of inst : label is "0840404042501414A439010101034141410C421030E52AD5DA965A94A5AF9FFF";
    attribute INIT_38 of inst : label is "51010491DC7DA4ABDDA6CA1CB5F7AEBA3A2B897BEFFB177455D9E5CEB9749DB2";
    attribute INIT_39 of inst : label is "12092D20242ADCEFCB7786D64CD376301B80D2499272304D0A889297381FADA6";
    attribute INIT_3A of inst : label is "A6B286263C491CF5E4A657889D924925865C47B38CBA23E3C641081C64D44DC2";
    attribute INIT_3B of inst : label is "0F3CF30B072EB8B8AAB7E799658C37176D274DD3A445E7EBC3F9DC55214F4E5C";
    attribute INIT_3C of inst : label is "210000200DE48C89308D66F6876D301BC0F3CF3066680C4DAC0C4DACBDAAAF3C";
    attribute INIT_3D of inst : label is "00093A6C2334008AA647400455334D6B92DBCD6B9EDEE294170A285F3889AA1A";
    attribute INIT_3E of inst : label is "0998B391C2F02DAACB3951210A884009BA24200050000A000008000004A21000";
    attribute INIT_3F of inst : label is "9C042EA798E63C3AE57CA85401220118EA60F5F273F27A212800254E627F2C80";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "C6492494CDB8BA8561184790BD125989FFFA49325B6C312FFF1D0400673092B8";
    attribute INIT_01 of inst : label is "92C2975119725E6B89125A668119C42A34400D45A8A171BB33CA55882C05798C";
    attribute INIT_02 of inst : label is "E58C58F800E0C2C218E7DFC3C1631222E39302E4839971254D0325F6331BD248";
    attribute INIT_03 of inst : label is "596491257205D30CB8E3A1874F24365B2D965B6C96492596596C2496D9671D62";
    attribute INIT_04 of inst : label is "B7E86DF0E32668464CD072018518E986B249B88497292519196DD1D90F2B9CB0";
    attribute INIT_05 of inst : label is "86312C2D2B5ACB8CFCAED3215A5695B1D47424AEB04970C378CE5E32F1C96F84";
    attribute INIT_06 of inst : label is "0FFE79B2088E54B996F31F91BC4A4B1B158A228E5FF5554BA8F7802F781E6ED8";
    attribute INIT_07 of inst : label is "671764B38BC7799306264B05DDCF1E73C70C79269832FD0456C50802C8406387";
    attribute INIT_08 of inst : label is "2042859D40301CF7D64F178FFB8748090100369DDD2E561DCA6E232EDF1DCE1E";
    attribute INIT_09 of inst : label is "651E6D56BAEBB87B235F2813A980CE0D84F2D20EC3A0E00A779C50F45F0ABEDD";
    attribute INIT_0A of inst : label is "65B9738FE7F9738BE5F9738BE5F1EF8BB5AD29165C8712FEF8D3B3A73E9FA67A";
    attribute INIT_0B of inst : label is "D4F1CE39C98FA6B66A5A4F3CF3D3BBCF3CF481B431B1E30C9758C5CFFFF9738B";
    attribute INIT_0C of inst : label is "22113FF0E00DFFF8E44BFFFFE2F7FC23FFE111C08C4345C9321FCB4033604B2E";
    attribute INIT_0D of inst : label is "C3C57BE60DC76FDA050AB27D3CA7BEFDE9612E4F1796CC30620C2C44FFFFFF87";
    attribute INIT_0E of inst : label is "C31151111511115106328CFBB6CE328CFBB2CC320CFBB2DA514AB19A145C7025";
    attribute INIT_0F of inst : label is "B0B0E5F801D6EE0AC09B8476EDC23B768F16B638982EDC4C4ED2C84040C0B8E1";
    attribute INIT_10 of inst : label is "2A0006C661E5C32BBC71B73656064485D196AD164994C9612106090240C4C406";
    attribute INIT_11 of inst : label is "CB293CB764F32E64C12397010010010DD3B3B25BBF0504516104B77E4A2CA0C2";
    attribute INIT_12 of inst : label is "DDCC8E07F857B83C74B5AE0C2106C2C196BBD73A69AEDAEF4CEB9D33A6F4E122";
    attribute INIT_13 of inst : label is "CDBCDB2C9BADBDEB5AF9E69E7A69248329A4920CE308453EE377BF6B9EDC5E40";
    attribute INIT_14 of inst : label is "1E0441E104A1088F085E12BDD433CD29EE18527336DF6B4B4B4E8D1BE36DB2CB";
    attribute INIT_15 of inst : label is "D9E08B53A03163244210806344210A0EEB1F188F86664F1FFA63FC7D8FF11E1E";
    attribute INIT_16 of inst : label is "6E372DD79BC8E5C4B7EC1C79C70C32732DB6B9352FBEA0FFFFF40E7EA5F7C32C";
    attribute INIT_17 of inst : label is "03F006111D012754F8897B18E302D9443170800CC1A22861B018057CAA65B6CE";
    attribute INIT_18 of inst : label is "CC6E10DED9BA5A13CB5351C74E3D8FDCBBBCD006092C708C1824B80C665616D0";
    attribute INIT_19 of inst : label is "ADF1B7221330352C5EFAB035266EF9E0B8E4C26C692124F266F3D865ED63BBDA";
    attribute INIT_1A of inst : label is "0036161CDD2EC1947374D26D260941849829A6D34D2BE0108202133108007813";
    attribute INIT_1B of inst : label is "90002631F15C108DE0369111A4444A9528F2A54A3EF5EE619A46A2F7BB3D3D86";
    attribute INIT_1C of inst : label is "964A52D08C19CFB00267F1974BA77F1C4EBEE66CF6C0A024810F807C26685BBF";
    attribute INIT_1D of inst : label is "8C497DB83FF74ECC204906E8C136CE8C3969F1605232DAEF85CA3C000001885D";
    attribute INIT_1E of inst : label is "182403B398A88102D8973241082028AFA430CEFAEED8D8DDEF6C448E9E786934";
    attribute INIT_1F of inst : label is "5E221F18B98C13182031C060300819B8C5B9413B6110C38889988A2702C1F682";
    attribute INIT_20 of inst : label is "0C81902026EE9E54716C668FC000000000001A2D85A0BDB8CD1D0BBCF0E3B26C";
    attribute INIT_21 of inst : label is "4E692448199030836160CECC1BA25FC239BB585AD1D8C4E2CD60819010080804";
    attribute INIT_22 of inst : label is "91CACAAAFF57CE5BCB6000001856A480C40E094B4A949C01A3A56A324A54A0E8";
    attribute INIT_23 of inst : label is "4644A12C633198E5CCA660089257784392B2CCB3043306455665566AC3DAAC48";
    attribute INIT_24 of inst : label is "2000000000001F0600B0BCC1833171CD2CA249E1456FDC277FF859102584E349";
    attribute INIT_25 of inst : label is "C9E93A6800402BA5ADB2000477FFD51DE633904491DB7680D073BA57A5C335BE";
    attribute INIT_26 of inst : label is "40900401022FFFF01009A4904608E6A66134B1CD1CD1CD846C8C621D989E8761";
    attribute INIT_27 of inst : label is "8902081204882008020080A04882248020580623816248022088224812248902";
    attribute INIT_28 of inst : label is "4A6890D8864C10C406C4BB622EDC86AB900171DF1AA38A38E41911E8C48444FC";
    attribute INIT_29 of inst : label is "5090D12621A4890D25B09A82700367046035101B66E252AC48620310C406C988";
    attribute INIT_2A of inst : label is "A071BEED32D8CB6D2EC9901C012418808421012084210109420B4094912C4862";
    attribute INIT_2B of inst : label is "066C65619F258FBE6838D4A7C0B7C5B0C3D1F8DC62D86191F8DC63C31C4F8141";
    attribute INIT_2C of inst : label is "1C77DFDBBB3A25EF001A5C78B6710AA1C4033144CE20005BC34D1BE500FD22C0";
    attribute INIT_2D of inst : label is "8E615780C0678E5548484849A363C618CD7DF66878D3DCF79E944D367744C4D1";
    attribute INIT_2E of inst : label is "D8DB29D8D3FFC7FFC5EDB5FFC7FFE741CF58589627FF3BCDE6FF8CD1AE6998C9";
    attribute INIT_2F of inst : label is "8F05C25024310243D086150560EEC9E7E773C3300E5F75FB3060B2ABEC99E619";
    attribute INIT_30 of inst : label is "A60AF7FFF7FFF60FA6BAA7BAA79AFFFEFEFEF7DEAFBAACBAA49AFCFEFCFE0410";
    attribute INIT_31 of inst : label is "F2698206974C4D3E04303FBE3F9E37F226F2FED2FE92F7FEAFFEA7DEA6BAA6BA";
    attribute INIT_32 of inst : label is "C18E0C712EC6668C800000000000069C9F9FCF3E63E2E667331CF03A23AC668D";
    attribute INIT_33 of inst : label is "AC959393E995EEB571D1D1DD260AE763B7C1C69CD9CDDD613BCFD1DB0FAA36E1";
    attribute INIT_34 of inst : label is "0004004000000104510145051104000757FDDC69D80AAA61C6664E899C1381A4";
    attribute INIT_35 of inst : label is "1FE0E1D3FA38C0C04444CC478C38315C6BA8A6298A628A2F8BE2F9C630000400";
    attribute INIT_36 of inst : label is "3FE102604F0CCAABF178C155E30E803FC07181A7007F0E30CCF1555E30DE1FE0";
    attribute INIT_37 of inst : label is "4790D0D0D0243030481203030303434B434691243424C181B2A9AAE3034F9FFF";
    attribute INIT_38 of inst : label is "2592DB3E273012150858C8374841514FCFD4E4208405625BECEE3B299CD96259";
    attribute INIT_39 of inst : label is "5264B284F2D9CA58D8B0F04A20201D8830410975CD5D8FA0F28E0C60C8C21ACB";
    attribute INIT_3A of inst : label is "F15951398D6ECAC2DA190F8026CB6DB52EE192DEE9771949931001B9494C944A";
    attribute INIT_3B of inst : label is "11C71C9891CD373688B85CE28A3264D276FCDF3BF14FF3FEBEAA2B419790811D";
    attribute INIT_3C of inst : label is "84FFFF09794F6C16CB640D28181042C4711C71C9C0DC90939C90939F8F557AED";
    attribute INIT_3D of inst : label is "FFE26DB2D9CBF424DDF29FA126EED28CEEC6D28CFE36829644020C24A081E069";
    attribute INIT_3E of inst : label is "C2E6587C0101CF439CACCC1B66613E631984DFFFC7FFF8FFFFC3FFFFF1986FFF";
    attribute INIT_3F of inst : label is "410D1E136E5B9901515A2865F86DF86773A2C0CD1D5D12C487FF0C33AD12961F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "44000002C69090054150540094024901FFFA01125B6C102FFF11000167B0DB14";
    attribute INIT_01 of inst : label is "00C15799994A502A000019628128C0BA10C00C4508A06279115804A030063888";
    attribute INIT_02 of inst : label is "4508F8C80082264508A6CD06AB22200853B602C201092029040125F221134000";
    attribute INIT_03 of inst : label is "5B2053674005814494D31152454096DB6DB24964B6CB2CB64B6825B649228802";
    attribute INIT_04 of inst : label is "B7C52FC0C12E38025C7022010F20C523B3AEAA8D96A00018092589F80EAA9A84";
    attribute INIT_05 of inst : label is "021524252B4AAA44FAAA49454A52959252703AAA94596A1368C44A1259DB6F8D";
    attribute INIT_06 of inst : label is "88027124004E509556EA9F81B4494838301A6698400AAAC22055820D68126451";
    attribute INIT_07 of inst : label is "27326D9B994228B98E72598C888A9D22A6847B248C38B81406481002C84863A7";
    attribute INIT_08 of inst : label is "208480B5801018D654466289628D4889118214D8DE2C54314B0A220B4D15C432";
    attribute INIT_09 of inst : label is "649C2436BAEB9869615F2432B100C50107EA09280AB2AC8E251CC19530FDF3A4";
    attribute INIT_0A of inst : label is "2499739DA6D9739924997399A4D8DE4295AD6B14488D1296E8409AAD3F8FE229";
    attribute INIT_0B of inst : label is "D42184308106A41228484F3CF3D6934F3CE080A8313162189350454FF7E97399";
    attribute INIT_0C of inst : label is "00308009E0000001D4CB000026000060000300A14CA70529A017AC0822C0023E";
    attribute INIT_0D of inst : label is "4B8762E215C56F4A8408A2713AE2AAB171412D0C1700C410260424C20000004F";
    attribute INIT_0E of inst : label is "86104101041010410D6158020CAD6158020CAF61D8020CB3716EB51E460C5225";
    attribute INIT_0F of inst : label is "2090A7E821C62208C102002271001138846A8520082710046716C8C0C040A050";
    attribute INIT_10 of inst : label is "20000A442145012ABA6090745A080005D156B51A4192D99303000900404C0C00";
    attribute INIT_11 of inst : label is "8A89FA856A290A64800301010400430D5693E25AAEA104504114B57D4A08228A";
    attribute INIT_12 of inst : label is "C94C8C65E2D6223878A52800010A42A15699D73AE9AFDA675CE9BD33AEFC5122";
    attribute INIT_13 of inst : label is "4494492482BA25AB5AA8A75EF905DBFEC4164B6962108118A533196BD4C81600";
    attribute INIT_14 of inst : label is "0A0280A082910845044A0AAD5411C9288A30C6203FFD2929292ADC0B91249249";
    attribute INIT_15 of inst : label is "F1409158803152256B5AD42656B5AC84693F499CA22218155C0154F405508A0A";
    attribute INIT_16 of inst : label is "241264D28948C48193EC0821861866606492BB15669AA1DB6FF4046EACD34228";
    attribute INIT_17 of inst : label is "81700E1217092664F8C07B18C302DB4D3530014D89A62869B0590D78AA64924A";
    attribute INIT_18 of inst : label is "CC6610DA59284013A843D48324148ACC9BB5E004012C61881005B00C54341440";
    attribute INIT_19 of inst : label is "8160900719153438931C15342C2A50A0A8D5E324293126BA22694920A9C4BB5A";
    attribute INIT_1A of inst : label is "00521508990A81153656990090D26C12434D1008699EE0210400231018816806";
    attribute INIT_1B of inst : label is "00002510E114808DF01290132404839718A0E5C638E14E218AC4C4D62D353480";
    attribute INIT_1C of inst : label is "552108408808CE1182E3E99542E25514CCEAE22455064104912A8454A4205AAF";
    attribute INIT_1D of inst : label is "842128E84237C72AA00000E882368E881570F1405222DACEACE015FFEE21105D";
    attribute INIT_1E of inst : label is "1806439289008122D8B236C408A000A7A638EE788A984891640C040814547138";
    attribute INIT_1F of inst : label is "5E22551899843100202180402018111045B840130112CB8089B0886702C9CC04";
    attribute INIT_20 of inst : label is "44E89D2002A61A54604C46075FFFFFFFFFFFF01A0C8F35988D440BBAA043E268";
    attribute INIT_21 of inst : label is "04642048008000852150AEC819804BE66BE9484A40D487E30744E89D1D0E8E87";
    attribute INIT_22 of inst : label is "888AABEAFD574E4B4960000018420000C20D294B4A901001D1A420214A54A0E0";
    attribute INIT_23 of inst : label is "A24020042110888528888088025574C102A30C308001020FFEEDDFFB86000444";
    attribute INIT_24 of inst : label is "3FFFFFFFFFFFFB0208B195810A7060A125E828C4066F14310018110005004141";
    attribute INIT_25 of inst : label is "59A13A2000400BA52DA2108477FFD54CAC33914CB54062BC9076904E20880599";
    attribute INIT_26 of inst : label is "60882608824E322EEEECE44442A8EEB26092E0A48A48A4886C0C601195980561";
    attribute INIT_27 of inst : label is "8080E89A0681A0280A228020681A0681E0389A2080A2283A2E83A2E82A2E8A80";
    attribute INIT_28 of inst : label is "290980144520300C00C40A62029C84818011708D4A818918401028A440040072";
    attribute INIT_29 of inst : label is "098010806000180000200A805000010C2004300A022242A4C02601304C02A404";
    attribute INIT_2A of inst : label is "E0F0A22C22D8C3572FA8311C101641900C0380320C038018260029820000C006";
    attribute INIT_2B of inst : label is "420075011E142D2E6968588EC833DFB0C3F1F8FC47D861B1F8FC4242102783C1";
    attribute INIT_2C of inst : label is "3C4456522E322109001C5868A15108214B1130274E200042C35C0B9402B09400";
    attribute INIT_2D of inst : label is "8860030180E7863C2000040181634208456FD6292853D8FE8A544E366444C4F1";
    attribute INIT_2E of inst : label is "C8CA21C0CBFF0FFF0DA005FF87FFA7418E4058160401384C26400CC0A9214040";
    attribute INIT_2F of inst : label is "908F20E8C832008160383E0FA2AAD452AD538320085D21C33060B2ABEC194611";
    attribute INIT_30 of inst : label is "A60AF7FFF7FFA60AF6DFF7DFA79BFEFFFEFFA79BF7DFF7DFA49BFCFFFCFFF4DE";
    attribute INIT_31 of inst : label is "CB0C0300D84061A8379E3FDF3F9F26FFE7F3FF93FE9FA7FFF7FFF69BF7DFF7DF";
    attribute INIT_32 of inst : label is "000810413016078080080000021045B4941A0D10710306083040C10064286607";
    attribute INIT_33 of inst : label is "A1943217E898A0147B0303076E42F06102C0468050051829194F16114DAE0081";
    attribute INIT_34 of inst : label is "4000000000000145051105550514000042A838103CA000600066CF88943200AC";
    attribute INIT_35 of inst : label is "E00081FE0FE000D3BBBB33BA00383801745141D0741D1450741D070000000400";
    attribute INIT_36 of inst : label is "C080F01E040C05540EA002EA800E0A8015400187FFFFF800C00EAAA800D89FFF";
    attribute INIT_37 of inst : label is "0440C0C0C1D030305407030303034B434341D074347401810155558003406000";
    attribute INIT_38 of inst : label is "24B2597A26100104084AC0140041404F4F44D2800405225B4C2CB3688449A2DD";
    attribute INIT_39 of inst : label is "5050A207EA19C2141030EA0C1470249800C0094545C55A94528C042058400ADB";
    attribute INIT_3A of inst : label is "7165E928A76A868288100D9816AB6DB588A330CE7C45D11021108529C984984A";
    attribute INIT_3B of inst : label is "81A61A1981E9A3A288AACE424828404176FD977AD376AAAAAAAAB14157900031";
    attribute INIT_3C of inst : label is "80000019794D0C36C92404A4350826CA380A20A148FC080A9800029A9955D045";
    attribute INIT_3D of inst : label is "0026EDB249A002685DA3801342EFCB4C6D884B4C6442808644020C24A000E028";
    attribute INIT_3E of inst : label is "264254EA41D1490312AAC40D46208027188440000C0001800006000013882000";
    attribute INIT_3F of inst : label is "D50D1E0324491B151142282404E404E732A280440404324000009C11241B4500";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
