-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu2 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu2 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "4654BD72E82D544810A1C62B22A2A0DDDD169646A5529A4601C512864ED8457F";
    attribute INIT_01 of inst : label is "8894A388B606259D2E822A4AE0D85E4229285764E55594C074B44A9938644616";
    attribute INIT_02 of inst : label is "8C2E1E8EC562F83EFD74210AF04AB165391B48410A206A982BB90B558929F0B6";
    attribute INIT_03 of inst : label is "842516934DCA4927611B64924A4D36046832AF46EECEEFD9D734AB06B8036BB1";
    attribute INIT_04 of inst : label is "A64F3CE24E2C02C3F246B0F24A42F587649272934DC940BE55506F9F542BE415";
    attribute INIT_05 of inst : label is "3AA0A9900B9853453FFFFBFFFFFFFFFFFFFFFFFFFFFFF6947B5447A5527A6953";
    attribute INIT_06 of inst : label is "2E408AA308C5061142F17608C1A92AF65239594A05A2A92AC65209194A351902";
    attribute INIT_07 of inst : label is "3958E08A140B2B5881670441A57A99C110699D4B454A5642846A866722A14E8A";
    attribute INIT_08 of inst : label is "FFFFFFFFFF99C78D54205BBD50215BB154E1D78846062695514464B5D8A42825";
    attribute INIT_09 of inst : label is "6D610098B4B402581029E9B5B462B87A472A026D610098B484025810C6BFFFFF";
    attribute INIT_0A of inst : label is "049EC9624B90155038530519D2F02E5A348F34018D28E1E9B58462BB7A442A02";
    attribute INIT_0B of inst : label is "B35AD39290AB9C406098207C4B12969C9D6C01AD608063A1253018254C061095";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5A04";
    attribute INIT_0D of inst : label is "0820BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "20281F325ABF1365AFD12FC4E979FCC895AC0CA96AC0C9979D15A8FD340FD600";
    attribute INIT_0F of inst : label is "C2B8E8B58B06BFA400001929EBDE71018260819F13E5AB5820281942FA609A58";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFF5726D9321610BD9CBA66F44B10998C17082080653B9094224D";
    attribute INIT_11 of inst : label is "2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "91007B503D4901069010B5590103D480F1790B1490D5641D5E600001062C7A44";
    attribute INIT_13 of inst : label is "6A1A05D22A8BC88B87D10181970249303DE64D8DE9F84DC7CA51585190007564";
    attribute INIT_14 of inst : label is "091A02440906660121118867CEA665AD05AD34168681BC4EA1A07D20A8681344";
    attribute INIT_15 of inst : label is "06918842E8D04A0000000000000000519694D694907EA45B01851CADDA040911";
    attribute INIT_16 of inst : label is "9D0DB4B959D2C031802E02C10A1041BAFFFFFF1BCD04104106C1B91D020BF6C4";
    attribute INIT_17 of inst : label is "57284124D5C5484524D1C0635B80B5C3541B01D0F4B778D0EE143DADDC1541B0";
    attribute INIT_18 of inst : label is "8D92A44A686B6706041FFFFFFFFFFFFFFFFC97945394518450A4924D5C613493";
    attribute INIT_19 of inst : label is "935C4AE39407F3C12B62AC09B72AC262B4EC885F3BCF01A5C7495A4794A47D48";
    attribute INIT_1A of inst : label is "02F9042C006E4A5552F5C89E5DCB966C9C89E5DC9966E9C8925C8519090906D6";
    attribute INIT_1B of inst : label is "334B2B752B5D39B2B5DB1F04AC0000000000026400009B0B52DAC144004F56B0";
    attribute INIT_1C of inst : label is "875D2C407AD5C59E2258F3CEDDDB1E6C9D4C12C9DD49DA39B276AC776C79B2B5";
    attribute INIT_1D of inst : label is "5FB678B6BD9B2C0A72A455DD110406E9B96E1CC844C2778D2BA416A4D24EB00F";
    attribute INIT_1E of inst : label is "8F3CE4F7896BD91985314E7462941DAD13AD41CC5BFA97F273C5BFA9749F06FC";
    attribute INIT_1F of inst : label is "E92B2763F64441C6614C539901219D0005195602BAC1E1E107C22146C9D34189";
    attribute INIT_20 of inst : label is "35A515851C85539B264C78E4FFFFFFFFFFF6218D91519D56144C588E65EA6280";
    attribute INIT_21 of inst : label is "E0D40764914EE29407F465613FFFFFFFFFFFD3A6466200006600A323B6E2FDC5";
    attribute INIT_22 of inst : label is "0ECCCCCD413C198FE2D40748AD01CE570196F1AE59CBE1D40757019631EE1BC7";
    attribute INIT_23 of inst : label is "823C0A42361B828B88AB71A68222292A8BE84174222291AA1A2BD3C403600350";
    attribute INIT_24 of inst : label is "C2241E2241D28A41E2241C2241D28A41D2241E2241C28A41E2241D2241C28AC4";
    attribute INIT_25 of inst : label is "3255866A1975CA1998FF64F13D024D907089074890789A41D2241C2241E28A41";
    attribute INIT_26 of inst : label is "4238099DC3A6D8D915066A4C0E2800004E54EC816792C829CC6B200019B20424";
    attribute INIT_27 of inst : label is "14104D2411804395785501CA7D89046C86953923EABA8D0A8AD8879DEB051BE6";
    attribute INIT_28 of inst : label is "4042BD8141C181C101814140C909D074C06D0822FB0743FFFFFFFFFFFF64D141";
    attribute INIT_29 of inst : label is "395176644B346789515C7BBAD9A524A128AD24A914E1FE407040606060706040";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF68B1C118";
    attribute INIT_2B of inst : label is "90A684A3FFA8AE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "38B66A4A9F8D0DF0D3E713C43436351DC3E1D74B101FA4C5C898D0F434F46753";
    attribute INIT_2D of inst : label is "CE31750144C9259999AEA038FEE534A94965217545ACCD852154A6D116B03699";
    attribute INIT_2E of inst : label is "992EE0F832910C52148D2A14A3482EAB0BAA6629B98A1A63F6118456D61096FB";
    attribute INIT_2F of inst : label is "5495274AA529D20BEAC2DA998E6E6186983D846115B68427CE31750944C9A599";
    attribute INIT_30 of inst : label is "6585F096504D485E648965742721391E5321D539152A95555D66664B53B0B04F";
    attribute INIT_31 of inst : label is "242A85149C56A0961411426850314053D014D14F9543692A2D99992C4E0916CE";
    attribute INIT_32 of inst : label is "000000000000095019715644CF569999D5A27E999966683D75999925A50A6149";
    attribute INIT_33 of inst : label is "ACBD00E428642421DC91800000000142DD8E8E29503318016A045104149B9000";
    attribute INIT_34 of inst : label is "01E98160A95594959A3481249A9A942B9451385321DA5144014F43507900CA3C";
    attribute INIT_35 of inst : label is "9775E97019548093A85857880230308FEC37CE15299992E6DD5DB82D68000000";
    attribute INIT_36 of inst : label is "1A55D4822320C23DEA455232BAD56752088D8318FBA4EB2CE0696B6A4702625A";
    attribute INIT_37 of inst : label is "CFFFFFFFFEAEB89A59F562A705E7A959232BAD255D48A23E0C027A5592027AB0";
    attribute INIT_38 of inst : label is "482640728CE0844200D55568394A28BE3D4078B53A520E6668259590C5F64EB2";
    attribute INIT_39 of inst : label is "5048DE53A69F3CEA549D1857ADB34A1819AFD0BA6C0BBA2501C1625176614A4E";
    attribute INIT_3A of inst : label is "64A4060999989300000048C9D3B7EFFA74EDBBC9F8904CAE3940751151D1AD89";
    attribute INIT_3B of inst : label is "D845CA14661614A45AFA9C502F8F501E99AABA98003250159843921229CC6848";
    attribute INIT_3C of inst : label is "122240181509C360A6E667911BD1DA069F612868000038000235235A35988B15";
    attribute INIT_3D of inst : label is "441E598A514A910A91CAD18A114A910586A2940760A86501D985C61409C01418";
    attribute INIT_3E of inst : label is "6E5104112C96B59A5440910E4429106529D03FCF1809A4226528442A472B4529";
    attribute INIT_3F of inst : label is "C8A7E67E6D13BD9AD101C21129484123AF65D53584E4644441949269A495C988";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C9E80F087306AB8010478001034341AAAA38A08AB4E4D28C119B604E8DD88508";
    attribute INIT_01 of inst : label is "212201B2DC427723280EE1FC69B5A0883E3A9EA82A7A728462CD81BA368E8EE9";
    attribute INIT_02 of inst : label is "754F168932E4E759FD48FE2520554178C2048C812300533844840DAA4236807E";
    attribute INIT_03 of inst : label is "C5E34EC30C340000EDB5430C0D34C147F4134A009E924AEA4C7FC459601D108C";
    attribute INIT_04 of inst : label is "55B7758227994010F781043A2CC4AB1D40001DC30C37136055C4D81F71360552";
    attribute INIT_05 of inst : label is "D42C4723565F2DBE32CB27FFFFFFFFFFFFFFFFFFFFFFFB8D68135681C7683763";
    attribute INIT_06 of inst : label is "0735CD1449975A65C43FA81DDD403C48D43D6350012F403C48D40DE35031721E";
    attribute INIT_07 of inst : label is "3E48F0CF1F5061790A3828915952CE0A2456155B5EA9F9E48F9AAE9C43531300";
    attribute INIT_08 of inst : label is "FFFFFFFFFF69388D79E058BD79E058B175A2C5989C7D7950A38B98DA5FE81431";
    attribute INIT_09 of inst : label is "2C6C753881A1D4F164153081A1E4390A1E43D42C6875388191D4F164C57FFFFF";
    attribute INIT_0A of inst : label is "48524EBA5F601C445A446C540D45758D06565DC5D56995308191E43A0A1D43D4";
    attribute INIT_0B of inst : label is "DDA3906FF444E080582E14508DEADCD0693211552DBDC6A57740160910052824";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5D48";
    attribute INIT_0D of inst : label is "FE1E5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "1515147585C44718503A0911E615111F627001E624001C6261EA6E09E8E093B2";
    attribute INIT_0F of inst : label is "D0641F890E056598B88811461653820160B8515447D8500E151517138838450E";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFF5B7D064EA4E4E06DD4192E82E2146014BE38E054CCB5A8949B";
    attribute INIT_11 of inst : label is "5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "CE205665014652566525457652501440C146585565055951517000029871061B";
    attribute INIT_13 of inst : label is "2866053E4A14710754620A015B410600301A83CDE435522BDC28202060007057";
    attribute INIT_14 of inst : label is "E866B08882056A92322203D80D0D7A60C260001619810B1E866043C4A19814F5";
    attribute INIT_15 of inst : label is "45578F8915D045000000000000000035E983C98000409749DDEE40092606C222";
    attribute INIT_16 of inst : label is "171F4250256F2E3162393291FB000025FFFFFF4B5E000000020D25BD0B44D700";
    attribute INIT_17 of inst : label is "3D6B0C33CF17BE0C2383D0431E4CA4845C6A1171037D2535695C40174845E6A1";
    attribute INIT_18 of inst : label is "13A1614E091A2C7C7C7FFFFFFFFFFFFFFFFE82B1C7A1F791E690C234F9A0200C";
    attribute INIT_19 of inst : label is "857505215C46775015C4FD00DD4FD011583D6C5425DD6076DC06F7DC547DCD07";
    attribute INIT_1A of inst : label is "9606C0BD0270054BA096DE4DA2DE41A2ADE4DA2DC41A0ADE41A28C4F7F7F4611";
    attribute INIT_1B of inst : label is "42BF7214320D46F720D0DF4050000000000001F70000AF6CE63BDF80A650AEF6";
    attribute INIT_1C of inst : label is "827A0BC46F42832D754F775951AF51BDF810EFDF850F8F46F7E3C346BD46F720";
    attribute INIT_1D of inst : label is "8F2FDFEBEF3EFAF83F2ECFB690689761D8769F5F5F1CBD505E989889052BE108";
    attribute INIT_1E of inst : label is "9775BA0FDAAC262BCA41498F8D62720D72022886FEEC9BE85B6FEEC9B3EDB6F2";
    attribute INIT_1F of inst : label is "57AF5D8EF7889A29F2905266DE690F77740F4BC3D219F431B0ACDB15BDAFDE37";
    attribute INIT_20 of inst : label is "8242820224EAA263BC0EFC63FFFFFFFFFFF59639EE22709F2A5053499BAC8D0C";
    attribute INIT_21 of inst : label is "209C46608101215C4604B9467FFFFFFFFFFFD27A9E8D555543C0613E5FD57D12";
    attribute INIT_22 of inst : label is "22000003C540174E209C466C13118D4801424F43750E209C464801420F43750E";
    attribute INIT_23 of inst : label is "22A132130DA5410F8C11C73F200001400E319FC6000014040438F41622C623C6";
    attribute INIT_24 of inst : label is "8C8518C8508C18528C8518C8508C18528C8518C8508C18528C8518C8508C284D";
    attribute INIT_25 of inst : label is "13AA7DB9E60B9AD67909272764569514A3214632142338528C8518C8508C1852";
    attribute INIT_26 of inst : label is "8BC1166F35791B1EC61B958002C400001993306CC82F06820C5C180002C14608";
    attribute INIT_27 of inst : label is "00800000010551508827118DB38C1012817635BC23D7FB13F392F083710C0596";
    attribute INIT_28 of inst : label is "F6E793D7DB9F9317DB9F13975B5FD16B03560E1A284447FFFFFFFFFFFF60C20C";
    attribute INIT_29 of inst : label is "EAF084C5C214E985BEBC6265D52561A5692165A171D554C5F6F7E4D5F6E7E4F5";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF75CF5606";
    attribute INIT_2B of inst : label is "58009197FF389D7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "16CC9E0F685F2A29F192A3AA4D5C6C4F82209E82F1198273D0B5F28E7C625A63";
    attribute INIT_2D of inst : label is "168FA919C84F5A22227A64A0672CA0F52C74B51EB0B35F04B912C77A02CE7CFB";
    attribute INIT_2E of inst : label is "22BA6460A98A282E0A8EAB6053ABC4A1F1606C8F0B270581AAA228AEAE2B7409";
    attribute INIT_2F of inst : label is "0B82A3AAE814EAF1287C581B23C2C9C160AAA88A2BA88ADD168FA915C84F9A22";
    attribute INIT_30 of inst : label is "7430627C81092C223A8EE0BD7EC716AACAAA9CAB151CEAAABFC88886234B8286";
    attribute INIT_31 of inst : label is "26631B4C9F0809806DB16631B6414C2199ED7086708A1614B32222198DB9C185";
    attribute INIT_32 of inst : label is "0000000000000319B090966907EE2222BE1493222209C50A9A222208599806D3";
    attribute INIT_33 of inst : label is "382710BF481D4010F50040000000038107C1A3252B831623C748621912641000";
    attribute INIT_34 of inst : label is "0355C0213CC068CCCD404CCCC5C9D815A87E2454A62EA1F89153F6C42B108B28";
    attribute INIT_35 of inst : label is "0A25A84016179ABEAC754C39BE50A9C6B962A460922221AA3F29C034E4000000";
    attribute INIT_36 of inst : label is "16C5F398E572A619A878DE5BAA1736CE63958A986888D649A54959697C7EC42F";
    attribute INIT_37 of inst : label is "9FFFFFFFFDABA90B1094BC281286A18DE5AAA1DCDB398E532AC26A185E6BEAC0";
    attribute INIT_38 of inst : label is "9899C4638040C8A2842AAA8501FF102239C467C6354D4088A41A6A642F948D64";
    attribute INIT_39 of inst : label is "6181319CFB077551A8A2045859CC8ADA7AD3916571104857118A908A808AB089";
    attribute INIT_3A of inst : label is "08C04582666E60000000D812766F26089D9BC9B10158045205C466EE6A68A350";
    attribute INIT_3B of inst : label is "22A9C8089B29285AD24071F1088E711895C08182D6F4B1095C082F01820C5C06";
    attribute INIT_3C of inst : label is "9D42F6399E6B9BF4D71998AAE0916605533614BC0000390001826C2A027F1848";
    attribute INIT_3D of inst : label is "9C7E2356E75E2756A71E2716E71EA71E81E35C462058D7119317178C67DAFD8A";
    attribute INIT_3E of inst : label is "559A000094E80E501451614185061418D13109DD5C55B35C8E5B9E7A9D589C7B";
    attribute INIT_3F of inst : label is "6D895DE5E8DC65A227118136053F88D8D978023AAF215888C4236606A26F9B39";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "D4A4D20E212557081CE4062928E0A2111104D26F6810E35C3A0794EF677C4187";
    attribute INIT_01 of inst : label is "3893BBEC08EF03D293E71C8BA7A8524E39BE4A46FD29780E886E53BD9E4A63F4";
    attribute INIT_02 of inst : label is "24A123EB50EE0492FFF07C39C25B72F6F94D0C413A226B8AE9990155898D3CDF";
    attribute INIT_03 of inst : label is "487BAB30C37CC30DBE658C30CECB1E079437EC46FE32AC18C8C9E69F881D79D4";
    attribute INIT_04 of inst : label is "EF14922B9CF282EFEA63B8DB008E0235CC30DF30C37D67CCA959F32F567CC958";
    attribute INIT_05 of inst : label is "2E53E3D638BDC71C3CF3CBFFFFFFFFFFFFFFFFFFFFFFF1EEFCFD3FCC8FFCF319";
    attribute INIT_06 of inst : label is "252342AAB6223D988C95471E21EC8454AE3DD2BB0991EC8474AE0D52BB39BD11";
    attribute INIT_07 of inst : label is "84961961223E7F330D353441A495CD4D106926978A44C48D5F495F48C8E2378A";
    attribute INIT_08 of inst : label is "FFFFFFFFFF6F454533524A7523924B792391E4B448FCF6B09044F4157DD63A52";
    attribute INIT_09 of inst : label is "9F9F23CB7F7C8F23A82B7C7C7CBEC7D7CBEC8F9F9F23CB7F7C8F23A8C6BFFFFF";
    attribute INIT_0A of inst : label is "8411415238D097B847B84CE8D7B867577EA8A62AE59E8B7C7C7CBEC7D7CBEC8F";
    attribute INIT_0B of inst : label is "155D2BD7788384426C9C204C41C18F64D33401A792408C8E7B901B26E4261C9B";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF484";
    attribute INIT_0D of inst : label is "4F279FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "214C1BAB533B86B533ED42E18D4CEE1BD6CC01BD6CC01BD4CF72C733707333D3";
    attribute INIT_0F of inst : label is "34ED3972E4268470CCCC924CE8761109B27081BB8635373C214C123924F09B3C";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFF8AB4D31C88E46E2AD34DF50C324CC9DC71C726C5F64709892";
    attribute INIT_11 of inst : label is "AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "CC3258EE725EE2E6EE2E326EE2E725C0327EE327EE897B8C9FF00002A89A7E29";
    attribute INIT_13 of inst : label is "DBAC24C8C6E3277DADC10D89B8B75D700DF703418DDAC935E8D4D0DAD0027D7D";
    attribute INIT_14 of inst : label is "39ACD244C926E2A1011288B4EB93E2CB3ECF2C9EEB013231BAC24C8E6EB01323";
    attribute INIT_15 of inst : label is "06BE4F0DE5E25B0000000000000000BB8B2CBB3CB24D3D85488CFCA36C274911";
    attribute INIT_16 of inst : label is "22323AD99F877339B3323301BF30C3AEFFFFFF4D280C30C30CC18FE24E4CFF4C";
    attribute INIT_17 of inst : label is "CBE7C73CF23D1FC73CF6F2639C8CCC9889C6622339D922231888CEB249888C66";
    attribute INIT_18 of inst : label is "A3DAE2C3C7C7C8CCCCDFFFFFFFFFFFFFFFFC4F7C8E7CBE7CBC6C71CF2F531C30";
    attribute INIT_19 of inst : label is "89DE6B1ACCE84923AFAE620BF8E621EAF062B813AD24BAEE235D2DE325DE3E5E";
    attribute INIT_1A of inst : label is "113C1CE2009CEBCF941E22D34E23DF4D622D34E23DF4F622D74E9CC7878788DF";
    attribute INIT_1B of inst : label is "3208A599259A3C8A59A33E8EB4000000000002840000C8B781E6225CD58F398B";
    attribute INIT_1C of inst : label is "503940CE89AB02D68BCD492277C88F22864C82286648663C8A198CDF223C8A59";
    attribute INIT_1D of inst : label is "0E80511411410519768154457F90CA328CA32232323449CE38F0F484E3925340";
    attribute INIT_1E of inst : label is "649234FABD171C1205306B5F639233C83233288554D217D657554D21755D4430";
    attribute INIT_1F of inst : label is "BBFF8960FF704134C14C1AD95C1AF2333CA4A5699912AA16C8363A3A1F863D8E";
    attribute INIT_20 of inst : label is "4D0D4D0D14055AD3856D7144FFFFFFFFFFFC6183D9C1324C148C18EB67FD638E";
    attribute INIT_21 of inst : label is "1A0CE8CCB1EB1ACCE83E93BEBFFFFFFFFFFFFAE44F635555C3CEF100C96A7F0D";
    attribute INIT_22 of inst : label is "058888888C4C97E41A0CE8FAB33A27F109910B305CE41A0CE8F109910B307CE4";
    attribute INIT_23 of inst : label is "FF936D304851EF81427A8DCDF2222C8AC0FBAA4B2222C8AA9E03FBAC02CC02CC";
    attribute INIT_24 of inst : label is "0EF290EF290ECF290EF290EF290ECF290EF290EF290ECF290EF290EF290ECFB3";
    attribute INIT_25 of inst : label is "10558B462D32312D233119F904CBE7CA43BCA43BCA4397290EF290EF290ECF29";
    attribute INIT_26 of inst : label is "0EB21DD231F6FCFD4127674C010C0000327178B4C4938B094E6E2C0009E20724";
    attribute INIT_27 of inst : label is "0C30C30C738BA6F144523A2B7EC30E7EE7219FB7BB5FD23B5B32D343951E9C2E";
    attribute INIT_28 of inst : label is "DEDE72B3B3B37737F7F7FB3A37B7F0E1426C0C2CC30787FFFFFFFFFFFFCC30C3";
    attribute INIT_29 of inst : label is "7522488890A6B469AD268ACAF212271223522352236BFCBCECECEDDDFDFDFEEE";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD2D5E58D";
    attribute INIT_2B of inst : label is "FC8C4C8FFFBEB6BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "AF7473A68332A0132A31D90CCCCCCCF210140E5033A169C2F8232A18CA893919";
    attribute INIT_2D of inst : label is "2D0947520840B51111E5DA8E8ECA4A6B949E524E4452328E527949291148CA72";
    attribute INIT_2E of inst : label is "1125FA8E8CCDA0190445CF5AE171346D8D17A709F9C2A77A2E511461A9D23CC7";
    attribute INIT_2F of inst : label is "06411173D6B85C4D1B6345E9C27E70A9DE8B9445186B748F2D09475E0840F511";
    attribute INIT_30 of inst : label is "DD2A4ACF73A394511445114CCC8DADE4A41E4A438BA4D5555344446899DCD368";
    attribute INIT_31 of inst : label is "8B718CAA2224ADC632E8B318CB38989A3C722268E2689DAEDD1111A367FFA92B";
    attribute INIT_32 of inst : label is "0000000000000B2326724CEDE4B311113190521111252C395511112677DC6326";
    attribute INIT_33 of inst : label is "92823A08D4D8E6B3279AC00000000263326BCDAF8CD39B30C60411241AD32000";
    attribute INIT_34 of inst : label is "016B412FB4EAF04EA3348F286F63D638702DAC135515C0B7A04E8DCE8E3A29A2";
    attribute INIT_35 of inst : label is "E083CC909BBB205F382FAFB2FC9280A8E4F9D8FA71111A3F3E83D8043C000000";
    attribute INIT_36 of inst : label is "98AE7B2EC92A01A3CC8EEC92B322B9ECBB2468068ED673AAE88484848CC8CF86";
    attribute INIT_37 of inst : label is "AFFFFFFFFD3FFAE12E3A17FF383F32EEC91B320AE7B2AC92A043F32EEC827390";
    attribute INIT_38 of inst : label is "46B48E80CC70047504D555643D887E81908E8BB19EC50C4465B1D1D0F91D673A";
    attribute INIT_39 of inst : label is "124DC375F784926A7011AC13A3D70CCE3D8FD8CAF764C5323A0D524D424D626B";
    attribute INIT_3A of inst : label is "24CC06C95DD1D3000000EC1C397CF3370E5FFCC131B042B1AC8E8811551842F8";
    attribute INIT_3B of inst : label is "9342BC36341416B7616F3333A06423A36BCC4C4CBC9D23A4BCCC9332C94E6CCB";
    attribute INIT_3C of inst : label is "DAE09FB7EDFB7EDC2F7774CD53AA2C66B7F5AE1800002200024D14D18D323834";
    attribute INIT_3D of inst : label is "48D952311231523512351239923992376BD9C8E85AD6723A37333FCEF37F37D7";
    attribute INIT_3E of inst : label is "A67C0C32B417DC2F7CE9D3A74E9D3A767BE38124BFE87DA148C648C448D448D4";
    attribute INIT_3F of inst : label is "18700D70BE538751123A23794F1F0E77A1F441164C6B6445CC99D1AD1ADA3363";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "60C0F10F1F76239C4672CF0E75730644440CF0C1E032C3C7354108471535C008";
    attribute INIT_01 of inst : label is "3C33C370CCCD3141540D10DC3F3430CFFC250F00943C174D57C4211C550F0950";
    attribute INIT_02 of inst : label is "06930251F06D17ACFEB9CEF4B039208C308793C43F701CCCE3764D884357274D";
    attribute INIT_03 of inst : label is "C0D3855D75D471C4C4330410534D1503DC7E51FD1B3F514E4CC704BD7331D17C";
    attribute INIT_04 of inst : label is "5BB28EC970D5806209111A890CCD5332871C755D75D5EE483C7B920F1EE48147";
    attribute INIT_05 of inst : label is "374371403763EFBE3BEFB7FFFFFFFFFFFFFFFFFFFFFFF14E344C3344CC344105";
    attribute INIT_06 of inst : label is "75034DC090A33438CF32103023706FB0FC7883F04003706F90FC40C3F07C1434";
    attribute INIT_07 of inst : label is "6C01B6DB00305113CF0F3DC01C2003CF70070B030D0040CC040C070CF6573CC3";
    attribute INIT_08 of inst : label is "FFFFFFFFFF66CF0013C00F3C33C00F3C3307F0C3CCC4CD2070DCDCD8A31115B0";
    attribute INIT_09 of inst : label is "0D01030C04040C331BD2C00404CC00404CC00C0D01030C04040C3319F13FFFFF";
    attribute INIT_0A of inst : label is "9C004E1333740128C328C4D4B128CDF128238258218A0AC00404CC00404CC00C";
    attribute INIT_0B of inst : label is "DC85D57C1972EFD00C305009CDE1C55E7E0C401A8200CCCD02B4430CAD00FC32";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA09C";
    attribute INIT_0D of inst : label is "43576FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "53F40281F9228C1F123C84A307F48A337C480337F480337E4AF8872EF972E0D7";
    attribute INIT_0F of inst : label is "3E7A1C0055013839CDFC00E493AFBF4030C140228C1F121053F40F3540417510";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFA38DC720C00D5D4E379C8721E70E480BC75F7008F33C390BF3";
    attribute INIT_11 of inst : label is "9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "0E70278620C46C6E46C620E46C620C4020C4620D4603D18839800000A28EE4E0";
    attribute INIT_13 of inst : label is "00880080D02203E42BE7CF002385C7200B1F914014828B3C68747874701037DB";
    attribute INIT_14 of inst : label is "3288D0FFC300B8673CC1FC9C95F5B8893485D408220820300881080C02204203";
    attribute INIT_15 of inst : label is "006FB39C93C03900000000000000003AE224D217500B5B404044F83EC80343FF";
    attribute INIT_16 of inst : label is "0331266366ECF37C3F4DCFC0341C7165FFFFFF74EE471C71C48046F9FFC4F8C5";
    attribute INIT_17 of inst : label is "4DF1755453BBB17554537007C373F8180CC0603326460E33038CC9918180CC06";
    attribute INIT_18 of inst : label is "A1C44E8C40404CC4C4CFFFFFFFFFFFFFFFFF2614EE14DF14DF17564537C9D592";
    attribute INIT_19 of inst : label is "3A86D50544D528E147CC86F13CC86C5479C63C0244A3B478E2D714620D462CD4";
    attribute INIT_1A of inst : label is "312E07C6FD0A518DC868E179C8E175C80E179C8E175C80E179C8C4C1818180B5";
    attribute INIT_1B of inst : label is "2F818233C2382E18238220851C000000000000300000E1B2E1F86107CD0BBE1B";
    attribute INIT_1C of inst : label is "211C844D52C67340898328EDAEE18B8618CBE0618CF18B2E1862C8BB862E1823";
    attribute INIT_1D of inst : label is "0C000000000000003000000020BBC0D0340D003030340589D37BD0C09D64A384";
    attribute INIT_1E of inst : label is "628ECDBC9C020E73432011C4117EEEBBEEEEEBB000C003C003000C00300C0030";
    attribute INIT_1F of inst : label is "14D08D11F8F9C33C50C804773E1441AAA85C1B57E03429F0C7751335F2EC9044";
    attribute INIT_20 of inst : label is "0787478774F8847F000C3000FFFFFFFFFFF9F04638E710C50D080451DCD01131";
    attribute INIT_21 of inst : label is "0644D5875E590644D529B512BFFFFFFFFFFFE4510711AAAAB01275324509BE07";
    attribute INIT_22 of inst : label is "40999998CCC80E590644D5BD913559BB40200033F4990644D5BB40200033E499";
    attribute INIT_23 of inst : label is "11630033440195CF0D9FCC051FFFF3830C8CAFC1FFFF383767320868474C474C";
    attribute INIT_24 of inst : label is "434E6434E64334E6434E6434E64334E6434E6434E64334E6434E6434E6432483";
    attribute INIT_25 of inst : label is "138809C027233027332E070838186A3990D3990D3990C0E6434E6434E64334E6";
    attribute INIT_26 of inst : label is "BF0A1441E18D24A3C30CDD08000400003DE3C974503097C3DF025C00C325030C";
    attribute INIT_27 of inst : label is "C71C71C71E082F63C0F33555F341C5915930568C54D83334D46233015AC465DB";
    attribute INIT_28 of inst : label is "4C4C13717171717131313130357520BBD00EF05CB2000FFFFFFFFFFFFF871C71";
    attribute INIT_29 of inst : label is "5430C0C06150F01430355671E000330033003300330A54DC5C5C5C5C4C4C4C4C";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF823C6444";
    attribute INIT_2B of inst : label is "6F0404CFFF1590BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "443C0D7F17314563144E855CC4C4C4C1A108472113540703F333144CC5174205";
    attribute INIT_2D of inst : label is "2CC21230354CD8000010391511C597F26C29B0C40C203139B0E6C23CF080C411";
    attribute INIT_2E of inst : label is "00101915104F44FC3C03044750C0445011183C440F11D9C47F0C8330FC001800";
    attribute INIT_2F of inst : label is "3F0F00C111D430111404460F1103C476711FC320CC3F00042CC21230354CD800";
    attribute INIT_30 of inst : label is "AB01944503766CF02C0B03C4C40C471859018591824CE22201C00011057273D1";
    attribute INIT_31 of inst : label is "80D2E0BE000C334F82F8052E08780034610230D130D167470F00004715170651";
    attribute INIT_32 of inst : label is "0000000000000103198D98A1E445000018301100000F24261800000D9E34F82F";
    attribute INIT_33 of inst : label is "7953354CC04CCD51333540000000011113951E66ECF7C3F4733C3F0C06720000";
    attribute INIT_34 of inst : label is "0086BF3F08477B84DD2F710F999D1114393044020400E4C0A008CC4D53355B65";
    attribute INIT_35 of inst : label is "1D76343403002444DF3344020091145108C62CF19000044D1D76313414000000";
    attribute INIT_36 of inst : label is "00C0102009145146340C00914D030040902451451241558E3800000004C04C7F";
    attribute INIT_37 of inst : label is "EFFFFFFFFD934E1F01C5F50F3748D0C00914D00C0102009145498D0C00910DF4";
    attribute INIT_38 of inst : label is "C15CCD53C944F3004CA2220C20DC119064CD50B0558F08001F984840B4E81558";
    attribute INIT_39 of inst : label is "30CC85EF0CC28E9DF94044024E3F98361CCBC5718CEF43D3354F90CFB0CFB0D5";
    attribute INIT_3A of inst : label is "0F0501C3F44172000000143EC611CD2BB18433402363B19064CD5E3300C80330";
    attribute INIT_3B of inst : label is "B3F0361D5E0E0D1FC001131364193354C20C0C0C2C0E33D9605C3015C3DF0057";
    attribute INIT_3C of inst : label is "41CCDD1745D1745CD8D111E042FC48E06F44457C0000060001C70C70C710341C";
    attribute INIT_3D of inst : label is "0CC00330C3300330433003308330833019064CD50641933561313845D1751741";
    attribute INIT_3E of inst : label is "49EEC71594E04504F9267499D267499D9EF344A3A0E400900CC20CC10CC00CC3";
    attribute INIT_3F of inst : label is "CC3BC49CC5823A40033561108633BD92DE8CCF0F05D61FFC4C36706706733103";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
