-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "63B7C1BBFD90FF6F3A2FE7AECCAE37BA095FD3C08A3EBB948F77D345FAA5BAFF";
    attribute INIT_01 of inst : label is "8D651C393A37FFBCB2CB80C85E379789E04598E621EF31BD18D9C783BBE2A095";
    attribute INIT_02 of inst : label is "56E2EDE2C97E1ECB77FEE3F1F1F8F8FC7C7E3ED22488EBC7379E3D4235267B58";
    attribute INIT_03 of inst : label is "C4F6369C6B4FF9AE8D2E66B8FCE3ADD7B73CEE908A6C89679B78EF1AFAEF36BD";
    attribute INIT_04 of inst : label is "A876A5FF51FCA3A9BB3FA94C4C748F1AB427A7F175AECF7974BA3EC5B0EF039E";
    attribute INIT_05 of inst : label is "B9B6679FC7FB27739F1FC8AE3B329764E2D200FCE31CCBA4CE979D1DF8D643B3";
    attribute INIT_06 of inst : label is "3D16186B95C6FDB778C96DB25F6F26FABFEFDF6FEE5FFB449D7F67F93FA7F8E7";
    attribute INIT_07 of inst : label is "7AEFAD7E6FCBC1F07BD4FDDA7E6BD71CD096CE06677779CF582325FE7F9FE277";
    attribute INIT_08 of inst : label is "5817F5AAEBEAA2FF52D57E6FEA5AAFE2EBD6AB925B648F1FA46BE2C4E27ED3F7";
    attribute INIT_09 of inst : label is "FDF3D9B19F86EDDE6FDB2BF5399BD6F6B2F9345E6B45FE37F9F917F2D6ABEFEA";
    attribute INIT_0A of inst : label is "FFDFFFFBB9B99B9BB99B98FF37DFE4F1FA8B06FDF179ED265FA2A8001FE3FFFA";
    attribute INIT_0B of inst : label is "7CF7D9B3F6977DE79E7FEEDF7FEFBFF9FFB64FF1C73EBFFEBEBB5FDEF5439F9D";
    attribute INIT_0C of inst : label is "EDBEDBEDBEFFFDBFDFFDFFDBFDBFDFEFFEDFEFF76FEF5BBEF3EF3DF76FBFFFDF";
    attribute INIT_0D of inst : label is "FDF7FF7FF7DFFDF6FFEFBFFBFFBFFFEFFFFBFFFEFF367F4DADB6DB7FDBEDBEDB";
    attribute INIT_0E of inst : label is "FCDBB7DB537F6FECDF4D8FFFFBF68B6F766DFF76EDB7DFFD5E2DDB3FDFFFD2DF";
    attribute INIT_0F of inst : label is "9B3EFBBFFE66DDF7FFCCD66DFAFF77D6FEEFBFEFF7F7EEDDFFDDB6DEB2D6FDDA";
    attribute INIT_10 of inst : label is "BD6D3F7BBEE3ADFBDFEFBFFEFDFEEFFFDEFDBF7F7FFFFEFBF7FF7CE34FBB7E7F";
    attribute INIT_11 of inst : label is "BA6872B1D44B3712EB19FD566BECF65B2B17B632CD17B9FFDEBE7BFD5EFBF698";
    attribute INIT_12 of inst : label is "F9899B1F3A9F7DBFFC056A5A94A4ED9FFF8F2ADCEF22E863A1AD0DE8FAFA19D1";
    attribute INIT_13 of inst : label is "C4BFFCCDCBF1DAAE008E9FDFD9C6987DF7C0BF679FD7CEF2D6FA7B3F9FEFF7F3";
    attribute INIT_14 of inst : label is "ECBF97B8BFC4310C6316E97CDFAFE7B7C9CF2F9FF3973E3E3CFDC47FF639CD7E";
    attribute INIT_15 of inst : label is "B79F7BDECFE5F2B1FC4BFE461894BA5E7A49E4885FE6F9BFDFCEFCCFF0F1EC57";
    attribute INIT_16 of inst : label is "8DD8F9B43EE3B8B177B3FDDF702C5BEFF7F265B32E4A700E8B5989B3A7EE9158";
    attribute INIT_17 of inst : label is "CD75D43EA3ACDC5DE8FF57E828DB3A7EE9158B79F7BDECF65B2B17CE4E88EEBA";
    attribute INIT_18 of inst : label is "C1C0E042B7FAB41DFFBC63C9F8FF1BFF765CBBDE56595C4CF77DEFE733B94832";
    attribute INIT_19 of inst : label is "955E7A4DEF68B396C22D1511FCBFF5E9EAA89F23DF7DB337390BC1D07C0F8FC2";
    attribute INIT_1A of inst : label is "8B561682012B3A8BB70859973A8476775DC6573736750A301681DECCF12B4938";
    attribute INIT_1B of inst : label is "9F2BDC672ABA4AD8CDA6B0EB8D617F0D442038CB2BA67D5329D38B60E85198DE";
    attribute INIT_1C of inst : label is "7EE6DD3E75D6ECB7B756481EDE3CC7F6F94BECBFF2EA033CF95EA8D9CAAE94CD";
    attribute INIT_1D of inst : label is "A5618000BEB7FD553AD3C8629B6C8E0C8D686B6CB741ABF5D97029C59D3FA32D";
    attribute INIT_1E of inst : label is "3D8700EA1DD9FC7231C3A3AA88AF086A8751A102701028BA65D8DFF5EFC8CD74";
    attribute INIT_1F of inst : label is "FA1F8E7523EA755AEAF6A435C8F9CB9C86721371EBA010F29F136D0CE42465C1";
    attribute INIT_20 of inst : label is "C8E2BB0B6E0E16315209C8D7677E26A395E4CA1251B4DFC23F952D11F511EDB0";
    attribute INIT_21 of inst : label is "5505C85DA3288A18D763C6571840B54518908EA2617C3D21DBB0F2A422EA2617";
    attribute INIT_22 of inst : label is "FFDFFDFFDDEDAD6EB5BF2BAFEAABA08ACBD52DE59BE69EC49C6DCA908CA29751";
    attribute INIT_23 of inst : label is "0DEF5A3FFF7AFEEAC7DEFBE677B2B6B9CF7CABFFABDEB5BB9DB19BDF957D67FF";
    attribute INIT_24 of inst : label is "9D23D98B636E409EC5BB7319BFFDFFFFFFBEFCF71C71E78FBEEBAEDFF7AF7AE7";
    attribute INIT_25 of inst : label is "DB5AF8BF6EEEDF9ACA53BEAE07EC41FE759779F79EBAEBBEFABD2B0C71CC9571";
    attribute INIT_26 of inst : label is "44A2E2E5FBEDFBBD7FFE2AB8C462313F89327393818B17E489D2719116247FDB";
    attribute INIT_27 of inst : label is "7E63978FFFC04C96306A462F9FAC27FB623A68C34CE6A6ADD7BA777D9CA63ACD";
    attribute INIT_28 of inst : label is "E386F0BCA31FE638DFFA9B60505383523A2EA61343FF1817434C8782C28A77FF";
    attribute INIT_29 of inst : label is "E9D95B77D5578A2E8A377C517DDD45BFDFFF75555C0300C105010550541505BA";
    attribute INIT_2A of inst : label is "FBFEFFFFFFFFEFFEFFEFFEFFFBFFFFFFFBFFBFEFEAA02D5FFFFAAAE8A8B0F0FF";
    attribute INIT_2B of inst : label is "444C50F25E27DD0EF617D85EA7882320AF926FFBFEFBBEEEFBBEEFBBEFFBFFBF";
    attribute INIT_2C of inst : label is "1117DF68B8844C2E20BA9133C43D1197275D5F772ED450827515517546875800";
    attribute INIT_2D of inst : label is "DB22DA64782DA07BA69E0B463523066932398DA351694B479E18C68BAB71D2A6";
    attribute INIT_2E of inst : label is "FF0C3B80A8855CFF8375C6D4B9AFF6605F6154FD8462EC91068CA07EBB7ABDBE";
    attribute INIT_2F of inst : label is "DB857FF57D575DF311600103B6D248A00192FC99208808FC0446AC17B2841DCF";
    attribute INIT_30 of inst : label is "C9D313EC4558BA566F134E5B2AD92AFCC7E26111E15924FA6BE470A9C15DE2D5";
    attribute INIT_31 of inst : label is "455E4CD190F508A5321D6274CD7D72469594223457798F793B88EF25B8A6F334";
    attribute INIT_32 of inst : label is "104235A4AF70C913215C99990842B96670C94464808944653718BE423EB81572";
    attribute INIT_33 of inst : label is "3842410138913193133541D8996C84E8527CC7929284601293028BC0C14C2151";
    attribute INIT_34 of inst : label is "7A0478886489468A391617043C8808111E888818081289148048488929A6BDD2";
    attribute INIT_35 of inst : label is "EECD408F4894E08B5889D6C9844C8AC6AE23401209F9AD15FE108422A415C9CC";
    attribute INIT_36 of inst : label is "1A533412CB2A0A710FB4EEE3D3D6767656DEFE7E5C55757D5DD5D5DDFAEEEEEE";
    attribute INIT_37 of inst : label is "228CE6E4E94CE6572B8774A76E44125156A727BAA83D92C503E73A298F184D1E";
    attribute INIT_38 of inst : label is "7D39BF044C09826B2976A4FA73315C41F36521306C4C130124D992B12851A6C9";
    attribute INIT_39 of inst : label is "5AD9DD475E1D7875F0BDF32E3FF5E7F4B64179FF6C8B933403EBC4CFDF97E72A";
    attribute INIT_3A of inst : label is "F7C371C638E18CECB81CEB5B9DCD06B177AF1265E565EC575A5E3DC2A27F47AC";
    attribute INIT_3B of inst : label is "6DFE05E902F7FFC09C3AB1BC743A4A5B31E45EEA82C6FEE2261442F17DE8D9B9";
    attribute INIT_3C of inst : label is "8F54443FFEFFDF7FBEBAFD7D5D7FAFBEFF5DD7FFC5D65D5DFEF6FEF6FE2A823E";
    attribute INIT_3D of inst : label is "70E82DE9E4B83A1BFBFBF5FF557FBEFDF7DFFBBBABBFDF5DFAFF75EB38EAB8E3";
    attribute INIT_3E of inst : label is "E5A379C37F597B26A31B79EFE6FF272F5CFEEA6DF8EFBC9DD71F55E1CCE718E6";
    attribute INIT_3F of inst : label is "8FE13DE5C7ABBC1D5B32FB150D963597914132F5D8BAF0FFD89EA49D3D873E17";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0B72D80C8DB4FF69B9EFE8CADBBEDBBA309EB2CBBEDD0A54B06B932DDCA1362E";
    attribute INIT_01 of inst : label is "B1B623C47F0FFDB4B6DEDBD0EE1EB3DEC8F79DC3EC48F7273B03EF1A3BAFED8E";
    attribute INIT_02 of inst : label is "E876E4EC6B96CF9996E73F7BBF9DCFDEEFE772DB348DC4299CDC43CEC7B0DBDB";
    attribute INIT_03 of inst : label is "E4FF204E6C7E119FB986641AFDEBCCBD34706390C7685131DA1B27BC1B27B025";
    attribute INIT_04 of inst : label is "9B76E3E91390D3554FF8ED676F7783081DA43F1820CC85F190DF3132DAEB809F";
    attribute INIT_05 of inst : label is "E606A53676DF31897CFDBEFED96D96E6FBDA66047FFE1BE6DC981F9D9D9E7809";
    attribute INIT_06 of inst : label is "0F3C6FC2001475B268CB64925F006E99EE7E3B19EEDFFB4DEC28180660580221";
    attribute INIT_07 of inst : label is "6EC9CF726E4B54EB183E650013D3D77E594486DAB127F8CD6B253A0180600B13";
    attribute INIT_08 of inst : label is "CE974CD9908492E4D66CC52E9ACD99D2F133606934DA2F5E202B9E07A67C403B";
    attribute INIT_09 of inst : label is "1B5E8B51F044E9E76CBA3369B95BD988BBF61A5A72A5A297E31F9726B366D11A";
    attribute INIT_0A of inst : label is "DDFDFFFDFDDDFDDFFFDDDE4AB780FCD69FEFD6F16F79973E6055F7D7C1406AAC";
    attribute INIT_0B of inst : label is "FFFFF8C14033FFFFFEFBEFFFFFFFFEFBEFB58A0184502000002C50000041DDDF";
    attribute INIT_0C of inst : label is "7DFFDBFDF6DF7DFEFF6FFEFFEDFEFF7FF6FFEDB18200197DF7DFFFFFDF7DF7DF";
    attribute INIT_0D of inst : label is "7FFFDFFFF7DFFDF6FFEFBFFBEFBFFBEFFEFBFFBEFF1820881EFFEFFFFBFDF6DF";
    attribute INIT_0E of inst : label is "8122C80400000040609208005480000020A0001832481110000464102140007F";
    attribute INIT_0F of inst : label is "8C5102C0002B064840046832402018000AB00022038004160016490820200883";
    attribute INIT_10 of inst : label is "005E40204802320160100088120081042812001EFFEFFFFB58A8084400138002";
    attribute INIT_11 of inst : label is "207F0080FBC2027080C0030F2F3C361F1F9DB40976D03FA951002C0005641920";
    attribute INIT_12 of inst : label is "F9B962829042131D266D6B5AD6A4428BCFCF10673F787F01FC0FE07F001FC0FE";
    attribute INIT_13 of inst : label is "030FFC30400C0881FF70003185CBF92D6B9D1D468FFE5333FCC63B1D86C7E3B1";
    attribute INIT_14 of inst : label is "8507EC877E3DEF7BDEE880C68EBB25CD44CBDA873B972E373B0403C105C73042";
    attribute INIT_15 of inst : label is "098B348EC361F1F9C6DBA36F7B843E17D60DFE7DA0818D1D876C76CFD1F94499";
    attribute INIT_16 of inst : label is "70A01483C81E0827020C103188D784C763B30CBB6EFE7BD37B59FEFB6DEDB98F";
    attribute INIT_17 of inst : label is "041C83C81E0809C083040C6F7BEFB6DEDB98F098B348EC361F1F9C6EDE608390";
    attribute INIT_18 of inst : label is "3C1E1E3E07FE03F0011F0100770407E3218D089FC618A6A2E9F9C763F0D87CEC";
    attribute INIT_19 of inst : label is "DF277E6DEFE5BB365CECB7371766A6B20A468D2344DD9FCEC1F0FC1F0FCF703C";
    attribute INIT_1A of inst : label is "E073C0F0781E3FACC3EF79B3739E0A3BC68E3BA6377D7A739F7A6CCDF36E799C";
    attribute INIT_1B of inst : label is "5E6DDDC7F9BF477B8F3E06087C0C209FCEF6DE7D0F336FF10F876E21F9BBDEDC";
    attribute INIT_1C of inst : label is "3D0F9BC20FEF83007FB207C09008BC201E490F0210176F1AF76ECC71FE6F87E9";
    attribute INIT_1D of inst : label is "587F10857F78FDF7CA6783F6FFFF7FCEDE70EFBFDFCFCDD29ED39A040C1F9AC3";
    attribute INIT_1E of inst : label is "B7999AFE79F9FE6733532CF30F38766FA587534F369EED87EFBE8577BECEB7AF";
    attribute INIT_1F of inst : label is "83BEEF7C6B352622DAF175B1C48ECB9E921A70D9115B7E71DFFBBDDEE7BE77CF";
    attribute INIT_20 of inst : label is "DDC53D4B434E9ECFF469D1DF41981E3335E87E2B1976DFD5249EB196E596E9D4";
    attribute INIT_21 of inst : label is "F73BD06CB5CCBEE32B2BC2F764AD9FDF3BD3B633E97D564939A49FE86D633E97";
    attribute INIT_22 of inst : label is "EF1EF1EF1CE1AD68B5BDFEAAFFFEF156816739E7315D5ED888788D185ECFFF67";
    attribute INIT_23 of inst : label is "0D6B5A3DEF7BBFBA8F9FFFCEF7A6F7B3FFFFFFFEC3FF37B3BD3393FFFFD7E7BD";
    attribute INIT_24 of inst : label is "CF33CDDB3B6665FDECD821B93FFDFFFFFFBEFCF79E79E7AE38E38E1EF78F78E7";
    attribute INIT_25 of inst : label is "9E1A9B7B02AABFB673BD6E01E0659FFE9E99EB9EB869A61A61CC31857D6EF5F1";
    attribute INIT_26 of inst : label is "7CB6F6E7FBFFB6BDEBE2C46DE6F379BFC3B3799B2CC996E99A3039981460F89C";
    attribute INIT_27 of inst : label is "EFEF8D3B8FCCDDB431E523122FF8A779EE3E6DCE6CFEE7BDD3BAF77D9EB2BEBD";
    attribute INIT_28 of inst : label is "4D2EF6D1CC4862BF9D537B98E3338F2C3B8ED30F23EA7336ECFF9DD261B07FFB";
    attribute INIT_29 of inst : label is "AAAAABAAEAABAAAFFFFFFFFFFFFFFFFEABEBFFFFFFFFFFFAABFEAFFAAFFEAAA0";
    attribute INIT_2A of inst : label is "FFFFFFEAAEAAFFFFFFEAAEAAEBFBFFBFEBFEBFAFFFFFFFFFFFFFFFFFFFFAFAFE";
    attribute INIT_2B of inst : label is "CEDF766992CF90CA22D75C778DDA762E04B1AFBFEEEBFAEAFEBEAFEBEBFEFFFF";
    attribute INIT_2C of inst : label is "F331EB26F3BCDFBCEE1EF37F65379E5F473DFE7F4FC657CCCDB3DC3DEEF7D3E3";
    attribute INIT_2D of inst : label is "59E24B6EF31C2CF9E2DF6F67F73004F9B776F64937BD409993BCFEE1EDCDF3E0";
    attribute INIT_2E of inst : label is "BF3BD77D7998AFFFB2B7F39C9B57F7EA5F4C66FFDA52DC333615A4EDEB3B3CB6";
    attribute INIT_2F of inst : label is "FE577DD77DDD7BBA99F24993B6D2499659927C993F7F54EBEABB372AFEE37CDB";
    attribute INIT_30 of inst : label is "FDFBDBFB6ADEFEFF7FDBFB77FDFFB7DEEBFB7FDBBDB6D6FF7FFEFEDF7DBBFBF9";
    attribute INIT_31 of inst : label is "7EFFEEFEDEDFEF7EDBDFFB5FEEFFFB9EFBFFBCF7EFFDDFB5ADEDF6B7DEDF7BDD";
    attribute INIT_32 of inst : label is "DF3FBFF3DFBEEFBFB99FDD7DCCCF7CF77DEDDEF79ABDDEF6FBDD6F79BFF6FFFF";
    attribute INIT_33 of inst : label is "7B7B7ADDBDBDAEFBDD7EE7DEDF7EDDEF7F3BEFFB67F6C97B67BB7FF6FBAEF5F5";
    attribute INIT_34 of inst : label is "FF76FEED36EDD7EFEEBF5F76BAEF327BD6EDF7DFF77BADDB25ED6DED29F777DB";
    attribute INIT_35 of inst : label is "FFFD9FDF6EDDEEDCF5EF59CFDFDEF399FF6BF2CF7DFDFF9FFE7BFFFB99FB9DEE";
    attribute INIT_36 of inst : label is "7B7B779ECB6E649BD9DADE7BFBEF6FEFEBFBFBFBFFEFEFEFEBFBFBF3EBFEAAAB";
    attribute INIT_37 of inst : label is "C7EAF6FCF87C3E1B1FDBFCE3AF6F7299011805DC2F3D92CFCE47BF69CF136F3A";
    attribute INIT_38 of inst : label is "79FBD9737CFBDE63F9B6BCF3F7B71F98737F3DF3CDDEF3653999D3516F7F3CC9";
    attribute INIT_39 of inst : label is "82041FD9F767DD9F74B584F97BF9D2F7BE7A74B124B99B7F5B8846F3CF9907BE";
    attribute INIT_3A of inst : label is "2D4F7CE7BE678EF0B179F0CF87E9C00F0082701B031C09A0C630083A9D083F81";
    attribute INIT_3B of inst : label is "6B2C04D702162C59EDFB35BD863E6E733DE46EEA506254F66CE4DB7DFDFC71BC";
    attribute INIT_3C of inst : label is "04FEBF880400802410002020000204100200000080000000080000080157D584";
    attribute INIT_3D of inst : label is "CC0FE40814774E56000009040000000000088000000408200004000000000000";
    attribute INIT_3E of inst : label is "2118780C1207001880C207E818911820438603890E883F05046014043398EE31";
    attribute INIT_3F of inst : label is "AE03B421EFAE94DF9BFEC1225C9221DB9F010E04432083844388238104611070";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "3E43A5B73D7969BF6B280F00092D1C03BE801E4B65240D244F4C43D9FA9936D8";
    attribute INIT_01 of inst : label is "477D88288E349242C8B06E373135FCB0595C7626D3CB692D74FEB131C0798E33";
    attribute INIT_02 of inst : label is "D4D98F537EED9A75ECFDEFAFDF97CFEBF5E5F32CD9763EC375950CD51CEFA7D5";
    attribute INIT_03 of inst : label is "890C6FDA4ADF7226323BBDE50214B6F641479F6CC65EE1D997F6CD6BF4CD4FFB";
    attribute INIT_04 of inst : label is "6C8DB9BD5FF7F1B7AC7EE033B9CD9D1AD1CB6FD9763B2FFFD7D1FEDD93550F21";
    attribute INIT_05 of inst : label is "79B97FDBFA5B6FEB7EBF26452BF79BED8EF4CDFF9084FD6D6EB7D4D397BEC796";
    attribute INIT_06 of inst : label is "C9E89FF2270DEEDA086FD9B25F1F91E7F99F84E569A40112722E23F82703F9F9";
    attribute INIT_07 of inst : label is "C566A5FF7FEE008951E3FAF26D0C210474092D645975619AD40324FE3F0FE597";
    attribute INIT_08 of inst : label is "7ED4A70F3F7C3A9A63879BA94C70F33A9E9C3FEDA6DA685124024FDFCAC497EE";
    attribute INIT_09 of inst : label is "AB4EB0101FDDB3E5A231BECE246A2722EE4FC755C47558D41674D4D31C3C304C";
    attribute INIT_0A of inst : label is "45F75F711911311117701915D47FA2036EE6DA8C1B425B66DF7786363EDA8806";
    attribute INIT_0B of inst : label is "B7FBEB27B632EDB6DFFDF7BBF9F7DF6FF7D366756E7EAFBFAA3B17DE93439F0C";
    attribute INIT_0C of inst : label is "B6CB64B6DB6C924924924924924924925B49A49A552AB9F6DB4FFEFBFDFEF3EF";
    attribute INIT_0D of inst : label is "FFF7FFF5DF5D77D6EFBEBBEFFFFEFFFFBDF7CF7DF3A5523D1925B6C924B6DB6D";
    attribute INIT_0E of inst : label is "FFF9BDFBB91F5E7997690F4D9FE7FB8BBCE9F724E9B7E7FE10859237DFFDD55F";
    attribute INIT_0F of inst : label is "B216BBBBD22C9D77FC44D66FFE2F37F2BE6FA5AAF7F5E7996FCF7ED3E6D2BCF0";
    attribute INIT_10 of inst : label is "97F1ADDF239FED7ADFCDB6DECDF4ECFF5ECDBD7B6BB7DF7DA577BC6345BB5C2F";
    attribute INIT_11 of inst : label is "AF681ED2F02FDE8BEB0C383DCA377F9FCBBF0DB699148DBDACD5F2D7F6B2B6D2";
    attribute INIT_12 of inst : label is "BA669F675FBA6D69F16C025AC4054D761DD513DB32A7F81DA14D0DF8921E13D1";
    attribute INIT_13 of inst : label is "5CBFFECDFD33CBAE1903A81B98F1DE643C855015FAD0C6DFBDDBB3CBEDD66D3C";
    attribute INIT_14 of inst : label is "603F14C0BE4539CE5296BC69B4F4FD67FDFA8FFD67AF5EFF6CEF5C7BDE010A77";
    attribute INIT_15 of inst : label is "3674FBBCF6F97CBAF3EC74B186BBEBF7FBFF058A46CCD369B34D7CFFFCFBFCDD";
    attribute INIT_16 of inst : label is "09C59AFC0EC1BFA85BB0DD9BB28C9B5EED37F36EC986F256792234393864F89B";
    attribute INIT_17 of inst : label is "BCBEF80D014F7A16D0368695D30393864F89B3674FBB5F6F93CBA731E98FEFDF";
    attribute INIT_18 of inst : label is "43416182FFFEF80F77BC1DCBF834E3B4A6FFDF4672480C0C85B45A7FBDFE6DB3";
    attribute INIT_19 of inst : label is "76DBC6D554534E7252626769B8FC0DCC15B1E75EB7DE39352701C350BC3F0500";
    attribute INIT_1A of inst : label is "0FD31FCB016FE9BB6D31C6497B0D37B6CCD796DAEDC08DB4284AC457B7B99961";
    attribute INIT_1B of inst : label is "725B6A7C55E9F3D4BAC6F9EE8DF13C64DB9BB40BC9DDDB83C978B28633676BD3";
    attribute INIT_1C of inst : label is "E32F943B75F7ECD8B7DF682EB34D83BB18FBFC8A9A6EB0C396DBC4DF157AE7B6";
    attribute INIT_1D of inst : label is "240CD8C06C8211234B271249820109821111DA4121890B253142808FE5701634";
    attribute INIT_1E of inst : label is "5D9586A66B6F012C9E138B99A5116777AC972E1AA4A3D83E4931308000C64010";
    attribute INIT_1F of inst : label is "F8614609EFF77CD99A87B1E605E49036A27A5F09E5ADCC92A6D52EBB6CE41189";
    attribute INIT_20 of inst : label is "19E10C5A1F54B4B690EA82B607860ED2B50E120369C3D0113EB6A6947494EAC5";
    attribute INIT_21 of inst : label is "A323C2596F742C24858A18B45E60725932D72ED38F411349D38DFFA149CD38F4";
    attribute INIT_22 of inst : label is "EFDEFDFFDFFD39EED4B40000400141879C2739A72E80CC16B1491B369E837744";
    attribute INIT_23 of inst : label is "CDEFFF35AD68A8A10FCF7FEFBDF7D7B9DAD000148BDFBFFBDEBFFBDE002AA7FD";
    attribute INIT_24 of inst : label is "1B67A33FFDBECF72216120C2C5B64924927D24FFFDFFDFCFFBFFBFDFFFEFFEFF";
    attribute INIT_25 of inst : label is "0ABBFCFFF4006BC2C801DFA1932E21FC708F697492EA8E3AEBA396214B5B9370";
    attribute INIT_26 of inst : label is "CC6BDF6D0082041A0C1911130984C2601CFD2FB1BA7CF54F719969B6B9E26509";
    attribute INIT_27 of inst : label is "998C3265211B4CE484522479B17F5C8353EAFF92FFA5A760000000003660A784";
    attribute INIT_28 of inst : label is "9A70291F5B5FD0A7E00C7A2D2CAC368E9924B9E27080C6164906B2913C138120";
    attribute INIT_29 of inst : label is "516905EE3BEC4D339E4EE0410CC33CCEDBFC788DDB3044140004444EEEEFEE9B";
    attribute INIT_2A of inst : label is "FAAAAA6AAFFFEAAEAAEAAFFFEAABFDFFFEA5FF2FFEB5695AFAFBAE13131EFEF4";
    attribute INIT_2B of inst : label is "FA90AC8A8C385C40C0B404313E6098886FBD707FDF03F0F5FD7F0FC3F7FDFDFF";
    attribute INIT_2C of inst : label is "3A26006B330E90CCC2A0BA52618594530E5B4157009A44CA4964B541359B5720";
    attribute INIT_2D of inst : label is "CFE7FE5305A3C3176F91B8FD6CE8115B598CA51DDF40DC6AFC6FADAA89F695A4";
    attribute INIT_2E of inst : label is "033800001B17020042811303B9080812D009B10F52643CB22B2ECB1BB060A07C";
    attribute INIT_2F of inst : label is "8E855DA0255F61963360019001325B205B92FC800AAA8B80018025A1A1BDDDC8";
    attribute INIT_30 of inst : label is "CE9C5EEE31289077CB1E234B4E0A3A7CB1A3A58C50C1679D4567B86941D1206B";
    attribute INIT_31 of inst : label is "C74CAB198D4406AD31A101C46F0C02631D41031870296B49EB862D3C886ADA20";
    attribute INIT_32 of inst : label is "02D2501860643010A63CE3113333AA17A28F2120654E210343C61A4E669B191B";
    attribute INIT_33 of inst : label is "86E3C570D241C50A388730F070E8627C07D0F15B89C356D98941810886DC3A5B";
    attribute INIT_34 of inst : label is "17C31987A98728813D15A7C74180CD9CE986085A889C530C5B669A46B7E1A5E1";
    attribute INIT_35 of inst : label is "008E68E1D862BAED5641A42962203CE4AE954DB38349B060EF9C0000E69C3E43";
    attribute INIT_36 of inst : label is "8DADE9D02DB691DCE616AEFFDB3F37BE343D757CF67F7DFCDE7F5DFCC0000000";
    attribute INIT_37 of inst : label is "7D75AB2BAE5F2F97CB74E5B9B1B9CDAC0080B31253A07BFB9A7C7EF62854B9C6";
    attribute INIT_38 of inst : label is "CB4E96D3A4B09234F27F6B969D2CA5999E9E4E92C68491F74E8F6615F989647A";
    attribute INIT_39 of inst : label is "43CBE59D2894AA52AAC2FC8FEC050F040E9D43CEF6CE7692646F99AA8531F975";
    attribute INIT_3A of inst : label is "BF90D5BD4AC87B2F97C5A6FBE4B614707DB683E59DE6EA434B934CC2A2BF87BE";
    attribute INIT_3B of inst : label is "87D0401E2041D3196DD6E6A178AAF697E10DEF4A4879A9ECD9B96E775F38D76B";
    attribute INIT_3C of inst : label is "FFEAEBF7DBFB5FFFBEBBD1D65D5FFFAEEC7754A3551FDD75B5FDDDF5DFD775FB";
    attribute INIT_3D of inst : label is "415FFF6A29A15BF3EBBAFDD7577BBEF9E7DFF2BB3BBF777DF2FF1BCEBFF33FFF";
    attribute INIT_3E of inst : label is "F5A7F1E373501A47CB3F1023079FC4FB7C74DA7B886FA0ACB786D36042100401";
    attribute INIT_3F of inst : label is "A80127FC589821B493687E68D8A2EE6630E73375C876CCF57C6DB82B440DD99F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "716AF4912D69DAE77CEBE3EAFFE7B3BAAC1F57F1EF986097CAD2691023ADC648";
    attribute INIT_01 of inst : label is "EF28F7D3CE55B6D3CDA3B6BF89D57AB4F16D633AFA957C555EAED7736267EDB1";
    attribute INIT_02 of inst : label is "F24912F1F6278AEDA2FEF3F5F1FAFCFD7C7EBFB7FDFED35D6EAAF4C7BD4B93DB";
    attribute INIT_03 of inst : label is "27913B163ACD0B0EBB1D57DD8E769F5BFF9EFBFFBEFC11FFBF9E45695E456589";
    attribute INIT_04 of inst : label is "ECCDBDD88FE6FBBEEE7EE3ED18FF9B0BC8FB6FC93E7DEF7C1A158C91A038A6F2";
    attribute INIT_05 of inst : label is "D71FFC7DEFBF6E221A996AFFBAFA8FEDB4EE1927B18DBEEDE7A275F37A5EDA0F";
    attribute INIT_06 of inst : label is "FEE6E30891DFF3FB6DCB6DB6DF15D077A4CD1EFF85EDB71A09EB1FFFD858077F";
    attribute INIT_07 of inst : label is "275294D5DA390A02E1B42A1024D41309BDFFFDB6FFDD6BDF9E92BFFFC0601FFD";
    attribute INIT_08 of inst : label is "B475DAB754BFAEADBD5BA4EBB7AB754EB76ADEFFEFBFCB7FA12C4C51EA32ADA2";
    attribute INIT_09 of inst : label is "5DF2A499C659D3BCAC92F7732BAAF74BE6D6A1D2C81D3275FA8C756DEADD1D56";
    attribute INIT_0A of inst : label is "99BBB9BDDDFFFFDDFDFDDD4A55AAAAD7EACF0ABDF75F274E8A5DF7D7ED757FF1";
    attribute INIT_0B of inst : label is "FDFFDD2ADC7EFBEFBF7FFE9E7BEFBFFFFFFE5DA2FFADBFFFFFF2DFFBFE49DBF9";
    attribute INIT_0C of inst : label is "FDFFDBFDFEFFEDFEFFEFFEFFEDFEFFEFFFFBFDFA55BEBFFFF7DF3FF76FBFF7DF";
    attribute INIT_0D of inst : label is "7DF7DF7DF7DF7DF7FFEFFFFBFFFEFFFFBFFFEFFFFBE5DA2FFEDBEFFFDBFDFEDF";
    attribute INIT_0E of inst : label is "6EDF27F9FFFFFFFE966DC6FFFEE3FFFFFFDFEFE54DB46EEFFDFEDBAFD0BFFFDF";
    attribute INIT_0F of inst : label is "D2EEF72FEBF4B9B47F7EC749F9F7E4EFFF4AFFF7F97FFFF936F9B6ABDFFFFFFC";
    attribute INIT_10 of inst : label is "37D1BC57A3FEDDEC9FEAFF97ED7B7EF7B7ED5FFBFBFFBEFB245A9FCFFFB57FFF";
    attribute INIT_11 of inst : label is "080730200BC0097008C9964466BFA3F1FA2BAD60DD828E3F0CFFB2F7FCBA64DF";
    attribute INIT_12 of inst : label is "AB6EF994A6EAA5F8896719C6719C55AE2FCD7C48BF7B17601CA0E88720C1D80F";
    attribute INIT_13 of inst : label is "03100238A92D000FC07E0B66A8A75454BC7AA3EBF12F6A5D63EBD1E8F57A3F1F";
    attribute INIT_14 of inst : label is "935F7B37C1B8D635AD7C2199FC6BBAD87175F0F0B56EDDCE579943A641CEF50C";
    attribute INIT_15 of inst : label is "52AFD9FC7A3F1FA2A1F64CF796BF6B8B0FACD8F1F26333F82A89A8BFCCF23C7C";
    attribute INIT_16 of inst : label is "FC7CA52FF45F1017151E48E65BF5A97EBF16D36499A835AA99F3003310EE4BEB";
    attribute INIT_17 of inst : label is "014137F29EA025C52B9159D2B843310EE4BEB52AFD9FD7A3F1FA2A19F5E04426";
    attribute INIT_18 of inst : label is "BD5E3E78500053F1760360000F930FCEEA74E9071EFFE5E441587E3D5EAFC15D";
    attribute INIT_19 of inst : label is "B7CABEDCDFFB615306EF6748D8CC42AC7C77FD7C396BAAAFE8FA3D4F13C0FFBE";
    attribute INIT_1A of inst : label is "6504CA30783BEA191D5AD642769FD7D1D557F1EAE88785B427354E9FF7FABB65";
    attribute INIT_1B of inst : label is "26F0EE7D26CBFE1CB958570070AC48E5D12DA18BFAEBB193F8B85AB63A76F1F5";
    attribute INIT_1C of inst : label is "EEF7FCD02A38473648E007C44A703D06C7026321C0F2DAE13787D75F49B0FD7A";
    attribute INIT_1D of inst : label is "66EC8C217D69FF552A6BDEFB2499FB598AF5F3DB4DD35AFDF7143AAEB2307F96";
    attribute INIT_1E of inst : label is "D7A5B1AE7FBFFDFEFF41F3EFFB7EB8EB02A8163AF961F222A297F5ED6CDEB4A3";
    attribute INIT_1F of inst : label is "79DFCE6DB2B842DEAEB6C1F7C0799FBF047E9769F4F69DBEEE5DCF7FED46CCD5";
    attribute INIT_20 of inst : label is "CAF7BF076FCE0F3372DC4AE377DEFAF51D61FEAD7AF557C61F0E6FADBD8DEDB0";
    attribute INIT_21 of inst : label is "37490AD7C93D6998AFA7D27591123FDF3C39C2F5E55C67E0D9B064E5F02F5E55";
    attribute INIT_22 of inst : label is "FF1FF9FF1DE1BDECBDFFFEEBAAABE082FBEF7FBD7D443CE7DDBDD7BFC9399E9D";
    attribute INIT_23 of inst : label is "2DEF5ABFFF7BFBFB8F1EF78E7386B5A3DEF7FEEEE3FF37B3BD3393FFFFDDF7FD";
    attribute INIT_24 of inst : label is "6F6EF73EFFDEC6965313E9DB5FFDFFFFFFBEFCF79E79E78E38E38E1EFF8FF8EF";
    attribute INIT_25 of inst : label is "6BF874FEFFAEFB5A894AFD3731EB7703F79F79F79EFBEFAEBAFB8EFCF659B623";
    attribute INIT_26 of inst : label is "906FBFAD6DB4D27ADC0BD55BFDFEFF7FFFDBFFB75AEDDEF734E99EB4E993BE62";
    attribute INIT_27 of inst : label is "27EDB56B5FFAAAFDB5F8EFD2CF32ED37FBEADBD2FBA717EDDDBB377DD6EE782D";
    attribute INIT_28 of inst : label is "591E6FBB599CFEFBAD55FF8FEF3BAFD7E2B8CB6E4BAAD6AF4A0EB09F6D757B6D";
    attribute INIT_29 of inst : label is "5757F788D75F555C20B00EFBF88FFDFC03C3BFFFFFFFFFFBBEEEEBBEBBAEEB61";
    attribute INIT_2A of inst : label is "FFFFFFEAAEAAFFFFFFEAAEAAEBFBFFBFEBFEBFAFE00A82A0803FFFC080B0F0FD";
    attribute INIT_2B of inst : label is "7921F9B6B537EAEF7EFF5C65B4E88CD265F4F57FDF57F5F5FD7F5FD7F7FDFFFF";
    attribute INIT_2C of inst : label is "1C43CF3537C7254DF3EB9C913DF7BB5D2FCE7FD76F5EBCBBFF7DE7D77F2E5BAE";
    attribute INIT_2D of inst : label is "77EFBED916EA7397EFB2DAFD79F939FB7C85AD5A1267B515C5FFAF3EB82B832B";
    attribute INIT_2E of inst : label is "B11FD1015BA6A2003D7C6DB655580105D753FC7DB42FF8B74F4BF383F3A609DD";
    attribute INIT_2F of inst : label is "73F0A228A22A0CCA99600192925249B24992FC9935FF7D680A396ECA6CDE9AAB";
    attribute INIT_30 of inst : label is "5E553C09E23AEEDD413CC0719CB87223B0AF003CA7933F88DB4F41C9238C2302";
    attribute INIT_31 of inst : label is "DE015AB4FF2F1F378FF6A70D9A13532BB8A0395DE49360C3ED3E3B795BC3B68D";
    attribute INIT_32 of inst : label is "1887FDEFC2F1B8AF353FC3C9AA67078D045F7776A99E777E2B346C7685D533A4";
    attribute INIT_33 of inst : label is "24CFA4A3CACF8BD6A1BE52B9FB83CA707A83A297080E14870DC734B5A90A722B";
    attribute INIT_34 of inst : label is "328E399EC99E2B0CC27D278E418F85382D1D7F35253CD338521C9ABFB31D0847";
    attribute INIT_35 of inst : label is "14FD23C0D9E611C0022F7A2F4966C428F0B4E927FF876D5E63397FFBC2386B7A";
    attribute INIT_36 of inst : label is "8DCDF8C4F7AE9A3E32808F77E7C357C3776B7FEBDFCADEC2F6E2F6EAF0141414";
    attribute INIT_37 of inst : label is "3CB529030F57A3F5FAB6653F13F6DD2C000FD0227189EFD1D2D97ABE226EF4C6";
    attribute INIT_38 of inst : label is "9A269AC58C2186D42A6BC3344D3C61FAAC8546307B0C36BB47B6343BF29DC5BA";
    attribute INIT_39 of inst : label is "900665D17605D8176343C9E430088CD1368D23FA97BDE695262DF9ABD7A5D979";
    attribute INIT_3A of inst : label is "1FF3D5FD6AFDD9A77A9EEFE7FD7AC4DF5709703EA27845F59C2A71FD7F133815";
    attribute INIT_3B of inst : label is "8AAC48CB247FAFF4DDBEF6FE6AEADE96EB3D0D47145D95E8C7DF2472563B574B";
    attribute INIT_3C of inst : label is "FF05012579AF35FEBDF7DF7FDBFFBB6DFDDF7FFB7DF7F7FFDFFFF7F7FE080A5F";
    attribute INIT_3D of inst : label is "6CE002A19FAEAB8BBFEFD7FFEFCB7EF75FBFEEB7EF7F76FBEEEFFDBBEFFEEFBE";
    attribute INIT_3E of inst : label is "101D084D04073B1A60E847C75A2C3D1517E049A466239F18916E02A318C2B08C";
    attribute INIT_3F of inst : label is "1DB3327F57BA9575E799E5FD379C5EEFEF401EA09B92537A2B94039C31602A6C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "7A7924FBBF7988DDFB5FF5453441219AB9CD97B241184F7D46D6F9C9F7EE33DA";
    attribute INIT_01 of inst : label is "4F3CE7C19A74924B6D33B6BF9B756EB4792D736E1A7B49EDE42E767359E6E9A5";
    attribute INIT_02 of inst : label is "FEC9B2912E619AACE4FBDF97EFCBF3E5F9F2FDBFEDBFF4DB6DACDD493DEB335A";
    attribute INIT_03 of inst : label is "67B32FCC50DE6B3A277D55F7BBDEBAFCCA9CF1B73672A1BD9C86CD6946CD65B8";
    attribute INIT_04 of inst : label is "64DDBEE6B3937B3D89FA8CAF39CD1A159FF66F514C79C7FD9AD0F36ED9F447F6";
    attribute INIT_05 of inst : label is "E80DBDFFBFE569C93CB76A1131AF3AAD96E4BD455EF625AD3DB165E6CFCAC265";
    attribute INIT_06 of inst : label is "E7E51F576D0F9F6B09890924801693D5EB5EBABEEDC0966C9A208000B88005BC";
    attribute INIT_07 of inst : label is "4F36B47F8FF25FF19CA1FCF1FE17F5F7F4A01BB43EE9435ED49284003F0017EF";
    attribute INIT_08 of inst : label is "E8EF1E5D7C1C1DE1EF2EB1DE3DE5D71DFC79777B7DBEBFEE12DDB43748762D66";
    attribute INIT_09 of inst : label is "EDFBDB7BFADAF5ED9C3EDF737AE7F1606647BFBED2FBE5EFE2C9EF0F7975F43D";
    attribute INIT_0A of inst : label is "DFDDDFFFDDDFFFDDFDFFFF10CFEDAE2C5E8519F48CFF356AC655F7D7E853BFFC";
    attribute INIT_0B of inst : label is "FEFFFD2A5C527BEFBFFFFFBEFBEFBFFDFFFB74A6CE9FF976775BBEF5FF27DFFF";
    attribute INIT_0C of inst : label is "EFFEFFEFFEFFFFBFDF7DFFDBFFBFDF6DF7DFEFF247FF8B3DF7DFFFFFDF7DF7DF";
    attribute INIT_0D of inst : label is "FDFFFF7DF7FF7DFFFBEFFEFBEFFFFBFFFEFFFFBFFF64FF9BBFDFEFFEDFEFFEFF";
    attribute INIT_0E of inst : label is "F79BB4BA3890FEF9DB698F49D3D4D61F7C3B7F76E937F578BE8C937CDF77A8FF";
    attribute INIT_0F of inst : label is "9B56F9BFDD66DDF6BFACD66FFA7F37DDFEEDF563F3FFEF8DA4CD26FCCDA9FFF2";
    attribute INIT_10 of inst : label is "09FDAF7D3FA77977D2CD48DFC9D7FCBD5FC9F5DEFFEFBFFBE5CA3F67EFBF6FF7";
    attribute INIT_11 of inst : label is "FAF8918DF4122A049C3A357FCA9F9FEBF1F7AD4F265B7FCFFEF5DBCCF6F3E4F3";
    attribute INIT_12 of inst : label is "5B6F9B4F16A8EDF7AD2F7ADEF5AC9DAEE746CFDB98237883A21D1068443A26F0";
    attribute INIT_13 of inst : label is "E47FFF8063213DCA0702C8D73AB6D63A9E7D2344EF7FA6DEDF5BCBE7F3FD7EFE";
    attribute INIT_14 of inst : label is "00579688BF0621884313EB5DFBC87D8FFDFB5FE595BD7ADDEC057041340100C2";
    attribute INIT_15 of inst : label is "76AAE6FAFDFEBF1F552EEEFED6BD6B967FA5668C5B9ABBF7AD4DD4DB95AFF00D";
    attribute INIT_16 of inst : label is "80D6F0DC48200C60A2037057624D3B797EF5B366D3AA75D6AAB35CA9DD873778";
    attribute INIT_17 of inst : label is "461CB4486018A82884DC35D6A18A9DD87377876AAE6FAFDFEBF1F55B2D918396";
    attribute INIT_18 of inst : label is "016001076FFF6C01577C833678DC1BEECEF9F36D0CB39D9CAEFEFDFEFF5FBFF1";
    attribute INIT_19 of inst : label is "B4D98AD15B9A426745AF4549E237AD7701E7FB7EF5FB9AAF3300C1700C2F0540";
    attribute INIT_1A of inst : label is "96FB2DC686E6EA9B5D5AD7414496F3CB5293CF7EECD695D4AFBAC61BD6FBCA69";
    attribute INIT_1B of inst : label is "F399B25D2762FDC4B9E769580ED22564512DB289E76BB911E7E95AA66A4DA9A7";
    attribute INIT_1C of inst : label is "A14A930AD5D78011B756D8119EDAC0A2386F2C46B546DAEF9CCD3BD749DAF3DF";
    attribute INIT_1D of inst : label is "1E9B14A6FC21FF576A5AAC3192028951386E990920511A2C70B4E1ABE55FE463";
    attribute INIT_1E of inst : label is "76A0A32A47C7829F4FB2D0FEFEEBD7C7A728063BC9E39A1C1C31601EF210872C";
    attribute INIT_1F of inst : label is "90208410CB1F3485F1FBF42DEC9290BB960E8CF9ECC6D596BFD7EF6D6D6A885D";
    attribute INIT_20 of inst : label is "E6B3864D41C8990E6138443550C0EAA7A3F780915383BFE3239B6D395D190064";
    attribute INIT_21 of inst : label is "954345D36B29CF2901DAB5AF85D21D9724F242A60CFE3DE902A49EC2112A70EF";
    attribute INIT_22 of inst : label is "FF9FF9FF9DE9BDECBDFED415000051867B5EF3CE7C19F7E39AB9AF4F99339F98";
    attribute INIT_23 of inst : label is "4D6B7B3DEFFD45104F9FFFCEF7A6F7B3FFFB541463FF37B3BD3393FF6AA807FF";
    attribute INIT_24 of inst : label is "6D6B3675F6BEC9944CB325FFFFFDFFFFFFBEFCFF9E79E7AE38E38E1EF7CF7CE7";
    attribute INIT_25 of inst : label is "63C3D6FAA154717C4C41FD1039C770017D35597514594514513ADC2153512352";
    attribute INIT_26 of inst : label is "D4CD6D6D009200CB1FF191A78BC5E2FF16ED94B75A66EEF331DEB5B77EF5F36B";
    attribute INIT_27 of inst : label is "8EEBA0615FFB3349C698884FB17F6C9693EBFF53FFA1924CCD99333CDC40A8A8";
    attribute INIT_28 of inst : label is "18782D7B784250F93006D7D78E4C34DBEABAFC752880C689A2CAB54D0C658900";
    attribute INIT_29 of inst : label is "AAAAABFFFFFFFFFFFFFFFFAEBFFEAABEABEBBFFFFFFFFFD054141051505415FB";
    attribute INIT_2A of inst : label is "FFFFFFEAAEAAFFFFFFEAAEAAEBFAABAAABFEABAAFFFFFFFFFFFAAAEAAABFFFFE";
    attribute INIT_2B of inst : label is "F924CDA62D981C45D0AFA00419F926256AA0EFBFEEEBFAEAFEBEAFEBEBFEFFFF";
    attribute INIT_2C of inst : label is "3C47FFA5A64F256991E93C960C5F3A1D10D360954154E931A20D33D259AD52AC";
    attribute INIT_2D of inst : label is "6EAB76913EEA5B36ADA6DAFD4D694FAB68939C0CD7EA40AD5C7FA99E93FB5289";
    attribute INIT_2E of inst : label is "0C2807FE8AA20EFF8BF93BB24607F763BFF35C0DA64C14514D4B532FFBDCB5ED";
    attribute INIT_2F of inst : label is "7D62A0A2A0AA05F499F659B3F7D6599249B27D9B20020303F58260A1A41AD230";
    attribute INIT_30 of inst : label is "FFFFFEDFFFFFFFFFD7FEFFFDFFBFFFF7FF7FFFFEFFFFFFBFFF7FFFFFFFFEFFFF";
    attribute INIT_31 of inst : label is "FFFFFFFFFFDBFFEFFFFEFFFFFFFEDFFBFFEFFFDFFDBFFBFFFFFF7FFFFFFBFFFF";
    attribute INIT_32 of inst : label is "FFFFEFFBFDFFFFFDFFFFF7EFFFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFFBFF7FEF";
    attribute INIT_33 of inst : label is "EFFFFFFFF7EFFFFFEFFFFF77FFBFFB7BFFBFFBFFFFFFDFFFFFFFF77FFFEFFEFE";
    attribute INIT_34 of inst : label is "BFBFBF7FFB7FFB7FFFBFEFFFDF7FFFFEFF7F7FFFFFFFF6FFFFFFB7FFFFFFFFFF";
    attribute INIT_35 of inst : label is "01FFFFFBB7FFBFFDFF7FFDFFFBF7FFFDFDFDFFFFF777FFFFBBFF7BDFFFFFFF7F";
    attribute INIT_36 of inst : label is "C4E4CC5AFCD280CE369FFCEFEFCFCB5BDFC7C3D3F7E7E3F3F7E7E3FBDD540154";
    attribute INIT_37 of inst : label is "1CBDAFA38F9FCFC3E1B645BE3AF6DF6DFDEA2E4558B5FDB95BDD4EDF2D7EF5EE";
    attribute INIT_38 of inst : label is "CF3E86C5CA7D0DF62B4D639E7D0C7577BEC56729BFE86FB7633F3659DAD561FB";
    attribute INIT_39 of inst : label is "2EA2B51143E50F943FE72BEFFFF55FE6BAC6573EFB7D76D536B57DAD5AB65D61";
    attribute INIT_3A of inst : label is "BFFFD4FD6AF959AEDAC1CDBFF1DF2F40B5C20C05C96518416B5ED842A00907DA";
    attribute INIT_3B of inst : label is "84046E40372800BD8526477E2CCBFADFEA7D6FAD873D81ACDFDF66F37F69D76B";
    attribute INIT_3C of inst : label is "F614403AFE5ACBE00A69BA3AB416569A0AB88D42F1ADEE6E0F676F6F64A880D5";
    attribute INIT_3D of inst : label is "325FEE3C6F8F5BB974D3A30673F6882A094CD46852ACED3454868952DF954F7D";
    attribute INIT_3E of inst : label is "3965767192C89E82D42A883282930671E41D6A290939A04ED5075A33CEF718EF";
    attribute INIT_3F of inst : label is "FF6B1EBA51196B356C5313785D165663605BC00EC43AE49DE80EA44B8E171C99";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "9E65B8BF80B04C89104C00351155D0CE5BE7F3E77D413655508D06F9B2B5A8FC";
    attribute INIT_01 of inst : label is "51BE1032A53E5B277B6A5B49753B657A37B6AEA7D41FEA7E9505C72A0C9FFF5B";
    attribute INIT_02 of inst : label is "6CFBC8DC5FF5DD9B7CD9CCDA6E2D13369B8B44DA2681CFE787C72FB546F1EEBD";
    attribute INIT_03 of inst : label is "F2BFC01214EC1BF713800803C10F41918A3D26031712F805C417EEF415EED87D";
    attribute INIT_04 of inst : label is "17EF6601494083D704B074BBFDEEE1539960760A4CDD89C3098315FFF9068057";
    attribute INIT_05 of inst : label is "8150A22D1082B1025858BDDD70CE0CD6DB15AE004AD226D723782A2B0E0D6540";
    attribute INIT_06 of inst : label is "305A19D26A44D8038FABE2DB6F20F598982C2B0A8E765E5EF3C0000D00300826";
    attribute INIT_07 of inst : label is "C72D7F6D2DA6008748067D98FB02ADD682A000CD040EB426F5BE80037FC02041";
    attribute INIT_08 of inst : label is "07460021004948C00010888C000211A8C000800984D20C41A250344D5894005D";
    attribute INIT_09 of inst : label is "FEA9425C60A811A681588349B2A31905916C09182C9185461E0E460000841200";
    attribute INIT_0A of inst : label is "DE6C55F31BB9BDFDD9CB928146015D2E05D2E8C2846092DDE0A8F3CBC20BFF7E";
    attribute INIT_0B of inst : label is "BFDB6923F627FFFFBF6DB6DF6DA6DB7FB6D76CA4E73679E7F5BB74FDE851B111";
    attribute INIT_0C of inst : label is "92592D925B6C924B6DB6CB64B24B6DB6C924925F7DBEED7FFFFFB6DB4FB4DB6D";
    attribute INIT_0D of inst : label is "B6CB2CBEFBEEBAEA6DB61965F7DF75D75F7DF75D7576DACB996CB6C96D925B25";
    attribute INIT_0E of inst : label is "BFB5B5FA9836F66F93DF5BDFCFCF60FCB7BBB3A569B6F4DA3826DAB7DBF74F6D";
    attribute INIT_0F of inst : label is "B23E9BBCF9248D77A774946FE68A77D94EEDD120B3FE76D96FDD36F1E8BDEEDC";
    attribute INIT_10 of inst : label is "4BEDA7FF3FBBDDAB97E805D2ED6D2ED6D2ED5B1DF7DEBBEFE5FFA5E5E73F5F3B";
    attribute INIT_11 of inst : label is "657E2CECD8668AD9D1048D968B9CC2451440921FBF54900D36F59BCE36F324B1";
    attribute INIT_12 of inst : label is "019C165655067F2606FE9DAF2FEBCEDBB2B512FF9A857E5BB98FCAEE259F86DC";
    attribute INIT_13 of inst : label is "38DFFC2AD8D2AD942A8946409F9B71518F47BAA488E68FF23B7E45329944A4D3";
    attribute INIT_14 of inst : label is "054604D83E4729CE728195069360267C414CB8844E8D1A6CA0A734696E318C53";
    attribute INIT_15 of inst : label is "3FD8049349A4D1450737030E3900763BC60B440C029A0D264882C10D82648F31";
    attribute INIT_16 of inst : label is "02911AE05D435D2DA7505AC081AE9FC924C217BFFCDF4A7F369CFA54CCF3B99F";
    attribute INIT_17 of inst : label is "147EA85E038A2B69E017102F37A54CCF3B99F3FD8049048A4514407D3205D7D5";
    attribute INIT_18 of inst : label is "6B35B5471FFB1D5B335E5B86F016DB41674897F3A75C4E4F8EDF49A25148B2C1";
    attribute INIT_19 of inst : label is "4AFE0D792BD6DE606ED6FEDAAED55F7F9FE698370469AFC22BA9EB3ADEAF8A2A";
    attribute INIT_1A of inst : label is "11FA238D50C757F78EEF2BD0D9FB3A6DBB3A4D213BE6E22F9F4FE369680E17F0";
    attribute INIT_1B of inst : label is "69550BEAEB5E45B74F071C9C8E3AA13BB556D8F520106CFD228E651B9EEE76BC";
    attribute INIT_1C of inst : label is "3081DA0327F6D62C3FDBA2A4B118C4259CE91E571C8D6D574EB8C4FABAD58A48";
    attribute INIT_1D of inst : label is "1F063FAEA63300FE97E547DDCB260CBFFDF0DF65B2ED9E26D8AB27C991C01C66";
    attribute INIT_1E of inst : label is "115BEBD7E5E58192C9A5CCF38F3C2A734980C55426AA5DCF0978C80630478628";
    attribute INIT_1F of inst : label is "0220729A46204C65E8C086741011EC49C785688018DB3E490DA1B1F3979FBBFE";
    attribute INIT_20 of inst : label is "06C9C297E0ED2CC7FA65A9BFE80137B35980D652D948980A47D9D59B63BF7CA9";
    attribute INIT_21 of inst : label is "FEB2E8F377EC5FC213534566618C9EFFD3493FB392609E7235F10FF44DDB2926";
    attribute INIT_22 of inst : label is "FFBFFBFFBFFF7FFFBFFFFEAB955533DC84A30863109136085437CF98D75FFEEB";
    attribute INIT_23 of inst : label is "DFFF7B7FFDEFEFB57FBF7FDFBFFBDFFFEFFFFC4407FF7FF7FF7FF7FFFFAAAFFF";
    attribute INIT_24 of inst : label is "F2B8BEC68A996BA13EE2C03917F7EDBEFA4FFFFFDF7DF7FFBEFBEFFFFFDFFDFF";
    attribute INIT_25 of inst : label is "BE209132095535309A9F0400304AB9FC151D41561EF3EF3AE3AC3B4A60377BBF";
    attribute INIT_26 of inst : label is "FFD1B517B2DB644DD000CCC190C86430232288580D932601CE208E58645090B4";
    attribute INIT_27 of inst : label is "DF7D5A11B00CE764295C209421B0B6D8D57D24F425DDDB5AAF556AAAC3553116";
    attribute INIT_28 of inst : label is "046CB620E41045311A0B8358E3E24EE4374FD71BFA5023B8585F58F4E3104DB2";
    attribute INIT_29 of inst : label is "B0ED1127C25E21D825E05EAFE05CA7EC37C408D8DE3705DFFFFFFFF555555540";
    attribute INIT_2A of inst : label is "CFFEAAAAA3FF3FF2AA2AA3FF2AAFFEBFFFFABDFF71101004C46ABF82177AFFFF";
    attribute INIT_2B of inst : label is "54C82EDB2F5810951506ADB1481ABEF40A69AFBFFEEBFFEAFFFEAFFFEBFFFEFF";
    attribute INIT_2C of inst : label is "5390A4165114CFB445BDD32E1E5FDD3FA27BE0EAB0B62ABC9AE7BB6B85F3F975";
    attribute INIT_2D of inst : label is "A45833FF4B345DCC5CF96D0EEE0282958FA46233EDF460003F91DDDB5DCCF976";
    attribute INIT_2E of inst : label is "03FC23C2B5D91754C0CBB5B9A62293B8982D738BEC930F2BB05B55C88FCF67A7";
    attribute INIT_2F of inst : label is "3000352BD28DD12000F25AB64816C9B6C892FC9B6AA2881014807C2536836920";
    attribute INIT_30 of inst : label is "35B898557BEE4B1D9D981E2757853CAA6BB9EF1ADDF5F6961BBABCF398E393C4";
    attribute INIT_31 of inst : label is "6B98038B5AC5CDEC4B4033964BCDF196EE5E34A6B849DA198AED63349EF892D6";
    attribute INIT_32 of inst : label is "9D7F0305FC48AB5118C9F4A0C49FC125ABC58CD7127C8CF7D71F0E6179C0DBEA";
    attribute INIT_33 of inst : label is "C3194A09B5B4C030CF7F859CD41AF1AA707139E1E667C971E033C3887365FCDD";
    attribute INIT_34 of inst : label is "8067AECD16CD94CC03D9CE6396CC3A7E804E0096527B2D9F25C72DAC0157D363";
    attribute INIT_35 of inst : label is "AA65D5796CD94C79F12D4F8A72DEE39F516AF2CF019D4E9FA8FE042B9D6E9CEF";
    attribute INIT_36 of inst : label is "E1686AB376CDA335FFF0DC5D713DFC7DFEFFBE3D3E3DBE7DFE7DFE7DAAAAAAAA";
    attribute INIT_37 of inst : label is "CF8B5D7179A4DA4914493BE65E0F380155B39EC45566E997F72FE58C59C70F75";
    attribute INIT_38 of inst : label is "A6EF57F07DFFAA651EED514DDEEEAF99F7A3D1F7CCFD530EF89AED5C973ED4D7";
    attribute INIT_39 of inst : label is "23282AA8A1428D0A17530368300318CCF5A8C637D3302FAEEF102FD4B9EE0E90";
    attribute INIT_3A of inst : label is "2629F90EF4961FD18AA0D8249A4811414ADAD5A1ADB64B1363511A0280D883C7";
    attribute INIT_3B of inst : label is "B2404816242840A3F2C12A3180552DE17EB0CD001A4FC89F6CC6C101BA94E9F4";
    attribute INIT_3C of inst : label is "F64444FBDE7ECF48DA6AFF1ED47626BA8ADCCFEBD72DEEEEBF575F5F6D777704";
    attribute INIT_3D of inst : label is "F19FF4C94259FE25F7DFBABDD1728B3AFB4DDF2A5AACD534F58A9F5ABFA74F7D";
    attribute INIT_3E of inst : label is "6B51FAA89A8929B3998EA9E593DD956674EC533B4C2ABC0CA5CA90C3DE7B5BFF";
    attribute INIT_3F of inst : label is "CA001823BDDD4BFBD6CD8111B5D7C2AB698B19AECA74D4664ECD34B32ECB9A86";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "E4F9609DC0DD25C1E0177F7524C32845CD63EF2EE33E9930EF88C512A69C9002";
    attribute INIT_01 of inst : label is "CF6977DC91824B274DA025EDAA82E277A70BE750B80418104EC61CB7840C5161";
    attribute INIT_02 of inst : label is "B41D30322483013A895004864A4325018280C02C9923B11C0A2AF1233C41822A";
    attribute INIT_03 of inst : label is "53628E21B989CB118F63318DA63663004BDEA56E1DC7D60F710C00C60E00E602";
    attribute INIT_04 of inst : label is "C4D9289C55444E681227108C50CC60C75848C4F61A7B33082D249932DD96106C";
    attribute INIT_05 of inst : label is "98032EC00C00E214D342D12B84916D9C47B3180D3109A49DB667B2F62B21C010";
    attribute INIT_06 of inst : label is "444B8FC20025584F9FA649B24FE09B1E4069CBE8C7D6DE4DDB7127F9A0A7FC28";
    attribute INIT_07 of inst : label is "9F92C6819034D57D19C926B9B7204A891EBB722B1898D6758ED9C5FE7F9FF189";
    attribute INIT_08 of inst : label is "216B93648C1B6D7929B240972536488D6E4D9000000815AE8251B840FD981008";
    attribute INIT_09 of inst : label is "5FF7CCAAAF6D9212DC0ECDBE5AB5E0804C25A1AE991AF54BE91B6BC94D920825";
    attribute INIT_0A of inst : label is "200222064CE44664664000006BC0172C91912D7E90BE00C19F0AA80280155D59";
    attribute INIT_0B of inst : label is "0000052AFFDC00100504100000004104104A557EFBED1B6DFFF2CDBFFC02C840";
    attribute INIT_0C of inst : label is "249249249248024124124124124124100024020A55FF6E800002000020020000";
    attribute INIT_0D of inst : label is "020800800000000000000000510514414510514414A55FEFF000001249249249";
    attribute INIT_0E of inst : label is "6C9525B3FFFFFFBF964976DB7AFFFFFFDF5B6FA54925FFFFFFFB92ED97FFFFA0";
    attribute INIT_0F of inst : label is "52ACB52F7FDCA925FFFB95C93FDEE5BFFD4BFFD5B8DFFBF96DB924BFFFFFFF7C";
    attribute INIT_10 of inst : label is "FFA90D5B2F7D596F96CBFF76C93F6CB7D6C97FE006484000E5DFEFBB7FAE5BFD";
    attribute INIT_11 of inst : label is "207C0080FC420210800004B301CD02814262BB9B76F6B016EC37F29FFA92E497";
    attribute INIT_12 of inst : label is "2A57830310850152C395EF7BCC52206F6326AB02C9207C01F00F807C001F00F8";
    attribute INIT_13 of inst : label is "000FFC00400008823F80004043FE3F81087F82A8B86E38161122A142A050AA55";
    attribute INIT_14 of inst : label is "0DFA9488BE45294A52908103A9502C16D2586DBE0CE9D3C0F404044106010042";
    attribute INIT_15 of inst : label is "8069A8AB55A8D427BBB6C19DE5B146D262C6668C40820752E1B713703F072BA8";
    attribute INIT_16 of inst : label is "80C018844822082102001041877040552A57F26CD3318FF8C6772366B31A8542";
    attribute INIT_17 of inst : label is "041C84482208084080041070EE3E6B33A85428069A8A255A894273BBB7808390";
    attribute INIT_18 of inst : label is "0000004607FE0410011C010078040803903060088001F1F01258D4A8542A0310";
    attribute INIT_19 of inst : label is "2DC3C1D83B326CE6161E4CE8866D505774D2A95CC80FC4FF0100C0100C0F8000";
    attribute INIT_1A of inst : label is "807300C00023C4700C94BE46C26242812172A5DDE9918F8E60FF1B7A4C99E66B";
    attribute INIT_1B of inst : label is "A5322679EC47D58C7AE600088C0021323B8944355288E22D527D95DB671437A3";
    attribute INIT_1C of inst : label is "13046C0217F78000BFD208009008C42018490C02102117C929812A1E7B13A377";
    attribute INIT_1D of inst : label is "8D00F39A9235EE9DC494FC17096704330CCB312D9338B118298ECEC3EDB5F0D7";
    attribute INIT_1E of inst : label is "E8767519D7D7825F2FA8BA420AAE1C48524FB6F9DD73337B4548208C61A18C70";
    attribute INIT_1F of inst : label is "4600949784109994695E8C1EFA577CFA59C9CE84165CA7AEF17EDAA19C719827";
    attribute INIT_20 of inst : label is "718AC5A1E92B4BAA6FD43E65FC856BC852BF8D54E4292D7A924A6E494369941A";
    attribute INIT_21 of inst : label is "0CE23F8AC4B2492601D5952BD61B09E7EEA8E3C954B7A8348CF246DF383C954B";
    attribute INIT_22 of inst : label is "10E10E31631252154A02011015545E3A4294B5D4982233F54FB6F5E811B318D8";
    attribute INIT_23 of inst : label is "9290A4420080FCA4107298B14E492A44810001548C21CC7CC7CC7CC700088842";
    attribute INIT_24 of inst : label is "30EC63268691C1D76CB77876E1260000004C0100A08228B1C70C31A008310B10";
    attribute INIT_25 of inst : label is "2EAD1D23ED557DD514A61707A35261FF0A6AEF2EF124964B6CC3DC7ABEBB8E1E";
    attribute INIT_26 of inst : label is "8369A91C92C96DE76805BBBE9F4FA7FF364CC4767B264BBF3789C674CD933264";
    attribute INIT_27 of inst : label is "44D360E0DEFA77128CB314E3C0862A4CBBCFFE32DF133AE22C45088269ED5E73";
    attribute INIT_28 of inst : label is "3A999CD33A245D5C302685619E1C75980E414C708841CE99B411726B8E8904B2";
    attribute INIT_29 of inst : label is "427AB1AA030C861030CDD3AE8881C780400449999A205505111015410444411E";
    attribute INIT_2A of inst : label is "100000400555400400400555540401000007418040357D5F00FBEF2BEBD00004";
    attribute INIT_2B of inst : label is "BBB69D1C91802195DD4BA38CF33A776401C5DAC031A80A1A0281F03C1C030100";
    attribute INIT_2C of inst : label is "AE66B5D168EBB27A3AEF2ECCB72B4FA9FD86208DF1392933365965DE7B08F8DE";
    attribute INIT_2D of inst : label is "B41D2693A4EE392C19A49FF89979FF0769D6F2F010C6B7E0415F132EF2C22A5B";
    attribute INIT_2E of inst : label is "4CE40082A67403020979ADE0CE0041992BBB8388A5172388E1E73930178403CB";
    attribute INIT_2F of inst : label is "6017D50A8020BA6C661FB7FD6DBFFECFFFFF4FEFDDD55E801446EA801250B674";
    attribute INIT_30 of inst : label is "148758C450F1DCDDC112CBE0F5703590A103A11801BA0683586A10D52124C763";
    attribute INIT_31 of inst : label is "5EAD6BB5186A0C768313C3D9E89E572922A47B49EFB94AB9A78C3034D0D56A89";
    attribute INIT_32 of inst : label is "38C7ECF3578088BCF53BB243AA775E95A4C9330EA95D3306B85246F8BBFE3F97";
    attribute INIT_33 of inst : label is "8EE375B19249CADAA09EEB20D2ECAA5CED53319B5A8754DB5CC37D3CA9AE6A72";
    attribute INIT_34 of inst : label is "1B47090CA9096B9CD8ADA1C5411FCD3C5B8F7755AD3A521AD36E920DBB455D53";
    attribute INIT_35 of inst : label is "FF3B63E190C23AACDC1FB1E72925CCE17695E9A777396C4AA9357BD7662BE30B";
    attribute INIT_36 of inst : label is "9FDF9CC164998F2CE0E160F0D44262CAEAC363CBE94068406AE3CBC38BFFFFFF";
    attribute INIT_37 of inst : label is "39B39D331A150A85422A8B2A139CAE357EEA6F563982C9B33218C9C7A0CC1CC9";
    attribute INIT_38 of inst : label is "96746881B182313CEE5CC32CC899A6541E9DC6C6A71189B8C64F4EAF98E2E266";
    attribute INIT_39 of inst : label is "020833629D8A7E29FA6F72A094002DC079CC0B78D340E489E6C03D302070E889";
    attribute INIT_3A of inst : label is "00B19A38E51ED39C68804620A877001100821005050408414A500842A2084780";
    attribute INIT_3B of inst : label is "D5020C3D062902A2326E9A5F75E7F997C76D9528E079039C916D2D86AA460F44";
    attribute INIT_3C of inst : label is "FFBFFABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDD7501";
    attribute INIT_3D of inst : label is "D00FE408234FE2E5BFFFDFFFFFEFFFF7FFFFEFFFFFFFFFFFEFFFFFBFFFFFFFFF";
    attribute INIT_3E of inst : label is "2100780012010000800201E8009100204086020908883C050400140CA5A94A72";
    attribute INIT_3F of inst : label is "A6D6882B71716B265EA7B9DFA6596A2571010204402080844088208104011010";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "4BEAA8BF85B6FFE939FF78DFFF5D5BFE78BE32EF5D5D505470CF2C5005A5DABC";
    attribute INIT_01 of inst : label is "5BBA67C4AFBFFFFFFF6EDB91FCBEF7FFC3F73F97DC6BEBAFB50767BA3F9FEFAF";
    attribute INIT_02 of inst : label is "ECFFD4DC6FD5DF99D77FFFF3FFD9EFFCFFF67A9226CDE6FB89EDDFDD6FD17FDF";
    attribute INIT_03 of inst : label is "EC7F604E55FE97DF77C4CC13D9CFCCBDBEF563DADBB8C936EE17AFFC17AFF835";
    attribute INIT_04 of inst : label is "2FEFF5E2ABD0DA5D5DF9EDFFBDFF83089DF4FF3824DDC5F1A8F260049661188F";
    attribute INIT_05 of inst : label is "E604B57B7F6F7199FDFDFEDD79AF9AEEFB993A066F7B2DEF6EB82F2ADEDEF809";
    attribute INIT_06 of inst : label is "BF7D60000016F5B6FB4B6DB6DF00BC91EE7E7A1FACDFFD57DFA0180640580237";
    attribute INIT_07 of inst : label is "777FFE7F4FEB9E85A01B36BDFFC3977BDBF6DCD9A7EBEFECE5FDFA0180600A7F";
    attribute INIT_08 of inst : label is "CDDF5CD991DFDBE5DE6CCFBEBBCD99FBF173604DB4933DFE6B7603C79A7C287F";
    attribute INIT_09 of inst : label is "BB5E87F6F04AF5F7BDFEB33BFFEFF99CFFFE7B7BF7B7A7DFE71CDF2EF366DBBB";
    attribute INIT_0A of inst : label is "DDDFFFFDDFFFFDFFFFFDFEEFDF81F9FE0FDFBBF3EDFFB77EE055F7D7C3CEEAAF";
    attribute INIT_0B of inst : label is "7DF7D5BBDFDFFFFFFFFFFFFFFFFFFFFFFFEF7FBFFBFFFFFFFFFBFFFFFCD9FFFF";
    attribute INIT_0C of inst : label is "6FFEFFEFF7FF6FFEDBEDBEDFEFFEDBFFF6DB7FEF7FBFFFFFFFFF7DF7FFFFFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFBFFFEFFFFBEFFEFBFFBEFFEFAF7FBFFFFDF6DF7DFEFF7FF";
    attribute INIT_0E of inst : label is "FEDDB7FFFFFFFFBEDF24DFFFFBFFFFFFDFFFFDF7E497FFFFFFFBDBFFDFFFFFFF";
    attribute INIT_0F of inst : label is "5BBEFDBF7FD6ECB7FFFAD76DBF7FB7FFFDEFFFDFFDFFFBFDFFFDB6FFDFDFF77D";
    attribute INIT_10 of inst : label is "FFAD9F7FBF7D6CFECDAFFF5FADBDFAFBFFADEFFEFBEFBEFEF7FBFFBFFFED3FFF";
    attribute INIT_11 of inst : label is "000300000380006000C003BFAFBEB77BAFD5A4404431BDE6FE7BFBFFEAFBF6DF";
    attribute INIT_12 of inst : label is "D93C608080435FBD346D6A52D6A56E9BAFDF9BF7BEF803000C0060030000C006";
    attribute INIT_13 of inst : label is "03000030000C0001C0700038DFDF7B3FFDBD6D56CFFFF5BBFE9F5BADDEEB77BA";
    attribute INIT_14 of inst : label is "A8C768074038C6318C6800E4DEBB35CD65EBDAC5FD9F3E5FAB00038001C63000";
    attribute INIT_15 of inst : label is "BD9A54DEEB77BAFD4F6F326E73847F37570D9871A001C9BDCBEEBEEFD9FDC499";
    attribute INIT_16 of inst : label is "70200403801C0006000C00390CDFDEEF77B21FFFB5FE5FD5FA3FDFF36EEDBDDF";
    attribute INIT_17 of inst : label is "000003801C00018003000E4775FF36EEDBDDFBD9A54DEEB77BAFD4FD6C600000";
    attribute INIT_18 of inst : label is "3C1E1E38000003E000030000070007F237DFBEF7A71DBFBEFFBF6F77FBDDEEAC";
    attribute INIT_19 of inst : label is "DEF67EF5FFDEDBD12AEFDF7F940954A48AA6D53704DD9FCEC0F03C0F03C0703C";
    attribute INIT_1A of inst : label is "6000C03078167FBEEFEF73FEFBBF7B5BDEBF7BB27FECF2378DFABDFFF7FF3AF6";
    attribute INIT_1B of inst : label is "6ED5DBCFFBDF6FF79F980600700C00BEDFF6EF6DBD3337F5BDCE6E6BBBEDEBEE";
    attribute INIT_1C of inst : label is "3D0F3BC008080300402007C0000038000600030000176E7376AEEEF3FEF7DEEC";
    attribute INIT_1D of inst : label is "DD7F1087FFDCEFF7C877ADFDFFBF7FD77F7ADFBFFFDEF5CEDED79644082A0226";
    attribute INIT_1E of inst : label is "9FBB2F7CE9E9FF2793F31C738FBA7677E7CF5F7F6FFCDFC7EBBECF7BDFEE3BCF";
    attribute INIT_1F of inst : label is "83BEDEFAAB3D27A7FFD9F7FCFC9EFFDC3092F0D9125B7FD7CFF9F9EF6FBEBBDF";
    attribute INIT_20 of inst : label is "7DEF78CE121D9DCFB57BD5BE19387EB87FBBF77B5CDFFD7F242C5DCBE58BC38C";
    attribute INIT_21 of inst : label is "F77FD5AE75AE5D637A7FEFDFEC9FCEDB77F776B9BFF7F759370C9F6ADF6B9BFF";
    attribute INIT_22 of inst : label is "FF9FF9FF9DE9BDECBDFF2AAAAAABE116C777BDF7B3FF6FF9AA9AA5483D77CFBB";
    attribute INIT_23 of inst : label is "4DEF7B3FFFFEFEFA8F9FFFCEF7A6F7B3FFFCAAAB83FF37B3BD3393FF957FE7FF";
    attribute INIT_24 of inst : label is "FF7FBEFDFFBEEBDFF6BFA9BD9FFDFFFFFFBEFCFFDF7DF7EEBAEBAE9FFFCFFCEF";
    attribute INIT_25 of inst : label is "DF5E9B7B1BFFBFBA7FDD7E3040A7FE00FF1FF1FF1E71C71E79C8B5DFFDF77BF6";
    attribute INIT_26 of inst : label is "FDDF7F6EFBFFBF5EEBE7FFC9F4FA7D3FE7FBFDBE7FFFFEBBFA5AFFBD5ABDFADE";
    attribute INIT_27 of inst : label is "FFEFAFFFCEFEEEA6BDDC73926FFAA7FFD67E4DDE4DFDFF5FFBFF7FFFF75FFEFE";
    attribute INIT_28 of inst : label is "7DBEFE93DC484FFFAFFDFF9DE7EBEEFE3B8EFF3F7FFFFFFBE8FFBDD1E7397EFF";
    attribute INIT_29 of inst : label is "AAAAABAAEAABAAAEAABAAEAABAAEAABEABEBBAAAAEABAAFAAAABFFFAAAABFFFA";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAEAAABAFAFE";
    attribute INIT_2B of inst : label is "DFFA6BEFCB4F915F3FFFFCFF54D8FAFC0519BFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "F7F9F9A6FB7DFFBEDE7D77FBB593DEAF56FBFEBF5FD73BB5FAEFBCFAEDF787CD";
    attribute INIT_2D of inst : label is "FFEF7FB7DB78155FEFEB6E6FEFB7EBFBFBE4672648009CF19BBDFDE7D5CDE7C9";
    attribute INIT_2E of inst : label is "F773FF7FFBB9FFFDFFBBFFEDFDF7BFFBFBDF77FFAE47D97776F79D4DEFBD3FF7";
    attribute INIT_2F of inst : label is "0435F7DF5D7DF3FE99F24993B6D2491249927C9935D5FEFFFEFDD73FDEE37FEF";
    attribute INIT_30 of inst : label is "004A820200100800408040012011004002003000801040300340000100080001";
    attribute INIT_31 of inst : label is "000200C80010002000080042C010808400440021008804002100020400083004";
    attribute INIT_32 of inst : label is "00003184011008000014100800000860500144600000446012000A0202101842";
    attribute INIT_33 of inst : label is "18400040008004401120488010680420100000000300810001100A4001100118";
    attribute INIT_34 of inst : label is "0600140124004402001053002800000090001082000288000000408129402100";
    attribute INIT_35 of inst : label is "FF0400064004C002080012480640004284230000182801000C009420800018C0";
    attribute INIT_36 of inst : label is "BB7B6B1FFDAEED9FFDDBDE7EFEEFEFEFEFEFEFEFEBFBFBFBFBFBFBFBCAABFFFF";
    attribute INIT_37 of inst : label is "CFEF7B7D7D7EFF7FAFDDFD75B76F78D17CFEB576163FFF57D64BDFACCFFF6652";
    attribute INIT_38 of inst : label is "BAFFD5FB7EFFDF6DFABA5D75FFAF2FDD75BF5DFB6DFEFB6559DAD5F6B77F5ECA";
    attribute INIT_39 of inst : label is "80042FBBE66F99BE67DB86E97BF9FEF7FEB27FB5FFB92FBF6F384BFBDFAF0BB6";
    attribute INIT_3A of inst : label is "2F4FFDCFFE673FF0F4B9F1FFDEECC00E0000601A021801A0842000381D003801";
    attribute INIT_3B of inst : label is "FB7F18F28C3E7CF9EDF76FFF835E6EF37EA47FCD264FFFFBECE49BFDFFBEB3FC";
    attribute INIT_3C of inst : label is "55ABFFAAB556AAD55555AAAAAAAD55555AAAAD56AAAAAAAAAAAAAAAAAB557F84";
    attribute INIT_3D of inst : label is "EC00000014B7575B5555AAAAAAD5556AAAAAD555555AAAAAD556AB5555555555";
    attribute INIT_3E of inst : label is "0018000C0006001800C00600180018000300018006000300006000077BDAD7BD";
    attribute INIT_3F of inst : label is "3C93FC32FFDFDFFFD5F94126FCB2D2EBEE000C00030003000300030000600060";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
