-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GAL_FIR is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GAL_FIR is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "B49F904476A3E9B9F97709E4423FC0B3C059765C5D9075B7D8340D8699240FE0";
    attribute INIT_01 of inst : label is "B3982EBF45D4DCC8D327B46D00AE2E0BBA280206C1A39D9C8BDC3A1017DF0FD2";
    attribute INIT_02 of inst : label is "83E261BA7033AD1EBAB7E1E7F9C1AA28D082C334ACE0361F375F494CA48250D7";
    attribute INIT_03 of inst : label is "177FF2F46153EDAD517F1E782C29184B6093317AFC5699E23D4B5C8016A578CD";
    attribute INIT_04 of inst : label is "EBD3F3F0FB1B04ADB7EB5D381B79DCD4DF6F5EDC594C5F142BEAF8D93CD356C2";
    attribute INIT_05 of inst : label is "E003D10B7526FEEAAFC13D6C25CD9DAB78CA36FC7828E64CC9DF0AB6B3CD27D6";
    attribute INIT_06 of inst : label is "5BF4378C229A8F914D522AB42C7B72E3ACAD87EC45EBBB4DD2DE1DBB1EF28A63";
    attribute INIT_07 of inst : label is "547321F99B74C941149FC667F4A88BB52CDCF9418DCF2D5868FC816E825BE5AF";
    attribute INIT_08 of inst : label is "23E5082436702A32F9E613E7D602C16E8D8655FA560E9C31576B72DF6EFAAF65";
    attribute INIT_09 of inst : label is "5A780FF894C7FE42B170E7A365E5B891B27CB95DDBF7DD08DDD9BA95AB88B903";
    attribute INIT_0A of inst : label is "772A3B7A5ADB389A6846CFD111F10717E225EACD6628D6E6DB966C504F92569A";
    attribute INIT_0B of inst : label is "2B2A5B4B51AB2DC741FA214218C6A99DBD888EB3F1AF367883B3EC7A648DB8F6";
    attribute INIT_0C of inst : label is "E4A598CE4617BDFD20F1D0932552A5B74E5E263AC5491406D63862A2DDEAACA9";
    attribute INIT_0D of inst : label is "E6085A0442B7926326D52E7B98354BEA8691C45979D00120D597477E788916CA";
    attribute INIT_0E of inst : label is "FE20582C16BD0834FBCC65372B90CFF9F7F4C71F29E541EE96079C1F4F0C3CC2";
    attribute INIT_0F of inst : label is "0A3AD70AE3E31C989DD19C803BD816D54760D35695830B179C094C1E9554147D";
    attribute INIT_10 of inst : label is "9388D9014AFBEAB97AFA96CBB77C197ECAA4C0BCD7C2B4838C2846C300D40E7D";
    attribute INIT_11 of inst : label is "96532749F87EAC7E0BC57455684CEE3FF10D899106D9296D6884AA0D253BAB28";
    attribute INIT_12 of inst : label is "789D99C009E3BDA221EF247AB653E2F87B6AA211AD60DD61E624D693FB7F7CC4";
    attribute INIT_13 of inst : label is "EACD1F3960BF0947768A724E4883C53B61084A2E4FB653C866E19FCCCD30539A";
    attribute INIT_14 of inst : label is "A68EC4571B9FC6B75F36991993820A9498120A8617164983B1C04A5B7E0BC70C";
    attribute INIT_15 of inst : label is "A1BD22CFEE3C118FF2787485E08102A060BBFB76715C1981675837446B60F06E";
    attribute INIT_16 of inst : label is "E2AF9EF9398394E66218C4D9A8AC57F2FCCCD61F9017CCEFE6B68ED623F9D396";
    attribute INIT_17 of inst : label is "FAC01577435ADA8AF1F50D4041FFDFA10F1761336E957F1A3369B752DB6F7FD3";
    attribute INIT_18 of inst : label is "AC9BD155183D5F93D065596C9620CC659A88F7DDE5FED7068D4546D35F3186F8";
    attribute INIT_19 of inst : label is "88E5546B6CC405484A055D103C9900F79DFE6F781A66D8CF29CBBB370CBE3772";
    attribute INIT_1A of inst : label is "FCFEFBA7868828BB223577E86E8EA29D98E283A4A795AED095EAA5D7A0D0E5E8";
    attribute INIT_1B of inst : label is "0D291B5C786708F35701EB807D25FFE9C06E5BB38A4E9E365C2416E6C66C2662";
    attribute INIT_1C of inst : label is "F2F7FE9E1245442568C27C58EC56B968E9932CE611BF0D38E1ED384437DF1A83";
    attribute INIT_1D of inst : label is "3B8518C3C8F4F4E575514F80B44791BD5F5C116CEE11278AED318AE68C7720D6";
    attribute INIT_1E of inst : label is "EA4DC7E9F12E6A21EDB6C9D7A0784E10FB401A7E52DA3BCBFEFE9FE9CEA40C73";
    attribute INIT_1F of inst : label is "E59EC0B37735C70A1A5D7D66D6A592F1DFE9C45944613AEAF3A002FDC1FB84C0";
    attribute INIT_20 of inst : label is "FFB978477B3F9E072D702DFB7F4C33C99DF91F1053A71E7C171A9D71A190BBDD";
    attribute INIT_21 of inst : label is "BD756E0820CC67243D2EBCAF5D120BB57F32D8116B13786F07ABD3179B31D6EB";
    attribute INIT_22 of inst : label is "AA2F35A3D3CFC619E648CA7F53820B433054636F4660407F110748261E9482EF";
    attribute INIT_23 of inst : label is "371D56769E7C1B61FD58B80805775BD1B57E04AADF71B0C17D16878CF145D050";
    attribute INIT_24 of inst : label is "6BBAB2332D41A4579B74E059075D99EF933AD2AA479662846B766554555AE5FF";
    attribute INIT_25 of inst : label is "D6D3FD340740C6A1B83120A959275EB4E8B8442729AEA4B4A35F5F94E6BEAF99";
    attribute INIT_26 of inst : label is "BF7F1F8E7A25B8DF822D8932315B09BEE9B4BB6E5F94B06EC2038C9B311307CA";
    attribute INIT_27 of inst : label is "FF9E589A39131C843B17CFA79F6DBBDE0B7ACB86A4F79DB117F538D5E1EBC238";
    attribute INIT_28 of inst : label is "2B4A74480964D593F0745EB157CA37973C9B75FD67A294096AF327C8D510375D";
    attribute INIT_29 of inst : label is "3DDB5449F1721BB3EBCA2213EA311632653594CFF913C9BB3BED9E9CC64B7A98";
    attribute INIT_2A of inst : label is "1F15D24A81940C9FF29F6032092C43A1F08C849764B5773EF961CA2D5CA4AB59";
    attribute INIT_2B of inst : label is "8ECB188C15E69C4BF0ADA30E83AFA0749412DDBA283D51932E70DE3F1C83FC1C";
    attribute INIT_2C of inst : label is "D936F6E82A6FC47BB852B16A706215C1B12F682C17D2B67C7C241E7D6B69AACE";
    attribute INIT_2D of inst : label is "E36D61AA9524299145A87458CF938CA9C48A94C378A87067BA7EA3B0C8920DBF";
    attribute INIT_2E of inst : label is "257279DB8A2E01A0BD52D2D074E748B48BA652DF3D7023FCBB1F6C3B76BB239F";
    attribute INIT_2F of inst : label is "6D6A791CEB99C7472579BEF261959CBDDFA696ADC80457E97CD21DC431928A7A";
    attribute INIT_30 of inst : label is "3291BBAD7497E8E7C1DED0F6813D1CADA39DCA67A005EF0A07C7D043381F103B";
    attribute INIT_31 of inst : label is "D129D9EEC377619D59F796914F6A1A0A1A1A379E27B2B36D37A95F98F9EAA832";
    attribute INIT_32 of inst : label is "3A1609C6B5838C8F9B5DAE30BDACC3EDB946AE5D0A178C16F93E519B5DB207A7";
    attribute INIT_33 of inst : label is "2C862D633FA12FA34739E46894CF79B798184163CB76B0175278F5985EDCECC1";
    attribute INIT_34 of inst : label is "E069855595036F0BC562ECCF7B1D50601285CC9F3C94F8917576F739BC592631";
    attribute INIT_35 of inst : label is "57EC02577D4DC4C33C5C373271C3D42E3C18B8B401CFCF5751F37FF1C2575C34";
    attribute INIT_36 of inst : label is "D091619310341013722E371C4FC9115F5103B01D73EC66DC43834DFAED4C1001";
    attribute INIT_37 of inst : label is "F1F4BD0047B364012CC163B3463B0395ED440C434FB46F30940749B0DC4F8395";
    attribute INIT_38 of inst : label is "DB99A2C009028B04334024CF8F4746402BE1050380B940CE21904046B9E3065D";
    attribute INIT_39 of inst : label is "7079030A1C0D7D7EA7D107345F439DC1312BE4A0EBD1DCD0DC032ADADAB01C70";
    attribute INIT_3A of inst : label is "A807AC5E9C5A8A1D3725F5AD7A4C4A73D1DDF1761DF9E9FAA77A04118A67D00E";
    attribute INIT_3B of inst : label is "A7B7A7A2564A7AA47A7A61074D41DCD3D794C5F50F9F892970DFE7C474370E9E";
    attribute INIT_3C of inst : label is "A8E5795AF5C25094E9F985E56B7A7C40E9E886840E93DC43D4EFB7A0EA9FEAB7";
    attribute INIT_3D of inst : label is "45485AF1940AB03B3E156503BEC840948439494EF102507B322165029FEAAD42";
    attribute INIT_3E of inst : label is "9BA576E3945662194E5252E7641B8190220269E26106E799880AA788BAB80F89";
    attribute INIT_3F of inst : label is "0BBF6E88B8980EC88586B6B2EFCB9B86B06BF9BA26B76B923982E99B809B06BF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1DFDDCAD17FD2D44AEE05E81B180C6E1B43C12682B82DBC331EFDE800A038C4B";
    attribute INIT_01 of inst : label is "71C912FDA4D347533C6ABB383EB040A062CA54BB19EE82B17AA9B6ED7E22B497";
    attribute INIT_02 of inst : label is "AD2DF7C78F042CCEB29512BC4B12568AD6D33BB3ABA0AD82996EA9FC813F8F97";
    attribute INIT_03 of inst : label is "E13615354BDDB76AD8C98185367EE2930A248D19DDEBC7710F2CD2E470F728C1";
    attribute INIT_04 of inst : label is "9FBF1C9F3E81F58FD066148E375E4FBA7B42C263150EC8686D1D5F240739E60A";
    attribute INIT_05 of inst : label is "20BECF269B4C9FA6C486D4D6CA4892F2A89841C2B896AED676C33DE016C3B216";
    attribute INIT_06 of inst : label is "F3A7E4FEABA5CBF9C2D6F5E834A8FC3C887C4990E5A005104022A20503EABCD4";
    attribute INIT_07 of inst : label is "FEE5E763042B739AF7A37E5C099392C321282478AF83035910C08BB9EA75515C";
    attribute INIT_08 of inst : label is "92FAB62711E9DA8EAA9E073E6A2B0EF07963A3C7C0F0B2039568100703824B2B";
    attribute INIT_09 of inst : label is "8E48ADE1880AA3CAC5DB70A1653409DDD2AA806F7824249D347E960B339E1E89";
    attribute INIT_0A of inst : label is "D1220E11D0158BF9FACCA83119B08F191A45C81E670DCB5547B1D150CB943A88";
    attribute INIT_0B of inst : label is "646320E90EE1D94B9254AC193212767A8F1A7B6CFA4F142B936DA3682800FFF8";
    attribute INIT_0C of inst : label is "5A511874E3B576B2739E59DBA8AA9BB238A8EBDD2D1733BC6726D5CD55A05A64";
    attribute INIT_0D of inst : label is "CF4DBB259E3E8B1D0ECB8FEA5D66BCD09A31C439184E49B651A2D3581FABDD5E";
    attribute INIT_0E of inst : label is "6661F62738B2A4CED12AAEC57D579698248F907E8F2F4D948DBE850F3562F464";
    attribute INIT_0F of inst : label is "0B58EFD2D9D049C1979EC1D3FD503BB7962634401D43AC54092F65C4EC25CC21";
    attribute INIT_10 of inst : label is "A6A49C20D7C6EA2764F8BF064951F220732415DAB4D0F81914FEE958E3A8FD1B";
    attribute INIT_11 of inst : label is "0C336943351979046B1BD28B05D21C2ACCE0082DFFA9A4B30B2DA54D137B016F";
    attribute INIT_12 of inst : label is "4D52ED6A68F9F5946C89E1D99E412FEFAB2AFC051AF42C7D3E2C9C068225DF43";
    attribute INIT_13 of inst : label is "A7154E3B95DB025BAD9F5F7DF4BCC8DE806B5305D969CD8272F7ADFF785AA210";
    attribute INIT_14 of inst : label is "C58E8515A606C713C228A4E0198C9D3CDA743163D394D8D15FC5A812EB11C2E6";
    attribute INIT_15 of inst : label is "ED4648DBD8460832B38F427B0A51D9BE30CE7FE2905583DD1D48E5D705D85B1C";
    attribute INIT_16 of inst : label is "B85514A835B2792DB3277CF09519E3A02774E831126830836F905A564FE8E12A";
    attribute INIT_17 of inst : label is "A2D50D666EE7BA7E6B7DDF12E44537B6179D57BECB5CEFFFD3950B37CF017483";
    attribute INIT_18 of inst : label is "3BADE1289DAD1D25B46E4704A01803CDC270F2386652F496122C7C31D9881CE2";
    attribute INIT_19 of inst : label is "A2DFF1F8AD28BFE39D113432F3D994EAB333FE5001EE68719470F658249DB733";
    attribute INIT_1A of inst : label is "BAE28709E094176EF77E42C103E8F50077BD0807D1EEFE8F94C175596F7E1021";
    attribute INIT_1B of inst : label is "2C07DCFA903C0212112C827B1EE70FFE9ED93EF3B2E42C407D556BD3821801E8";
    attribute INIT_1C of inst : label is "7D9265D0A863B0DFA5E8697C67635338F5B8762303D01A0372618633A7CFF8F4";
    attribute INIT_1D of inst : label is "9BD0D862EBD00C376C805BBC6C2B6EF03CF6E9A9C8624A033873C96C7D3E7951";
    attribute INIT_1E of inst : label is "8767CC1DF48F8E7D3330E16311C901F4566DC598D851369DA18DBF0363CEA438";
    attribute INIT_1F of inst : label is "4A2349A4055BDE7A780C0239FE5E3378F757C4A83D1A8E647E3DD15A68F35BBF";
    attribute INIT_20 of inst : label is "E4E38DC5282F0F955A0B8D2F8746250CD822D927C00A8150F0B6B7925B277405";
    attribute INIT_21 of inst : label is "E37C10CE0FFE85443A3DBE34DF1F200DEB234F36178849FBA12D32E06F843799";
    attribute INIT_22 of inst : label is "BF37F3CF89F053020D11F0FA3E90CEE0C9A002622F388008E06B763D186F4A30";
    attribute INIT_23 of inst : label is "0F73BF080AF9D80CDFC15C1F8FF7C3FBF732FCEC404748A9F33C5307BD0849D8";
    attribute INIT_24 of inst : label is "C8C5330F73E3331CCCC3DFB2730AA8C8F370A53DCD201584F7C0AC84FE5321AA";
    attribute INIT_25 of inst : label is "3A2DCE4EE4ED4C603C0D30C301BC09CDD78931B77DC9CAC8F00FA9980EBC5316";
    attribute INIT_26 of inst : label is "923E5BD3C30C36393D63C0C0C0E7E33F0F1CF63F288057A22BD0C3ACCF41CF75";
    attribute INIT_27 of inst : label is "3E4E439036763D3D6C7C0CF81A5A59497C3366925DB9393F496618625F0D8360";
    attribute INIT_28 of inst : label is "F9A697EA9F7DFD393760DB97C7366C6033696608669791DCDBC6C76060F5E0A9";
    attribute INIT_29 of inst : label is "90B4E1C45A3EA59A4CA8970D99FF88460D8619CB153DFD2CF4A5A7D6D361A4D9";
    attribute INIT_2A of inst : label is "660AA5E5C970EBA5697573A2E0DA515CEBE885A8DA8FD2D299709249CB5A89F7";
    attribute INIT_2B of inst : label is "FAE1150B887384844B3578616A3A884E1959E28D9FD38618612EEDF4ABE2DD9C";
    attribute INIT_2C of inst : label is "18B5757213572E311C2BB8B55215B8484AD68E5C21C2D3573B8BA132A5A84D68";
    attribute INIT_2D of inst : label is "CAAE0BB3B8B8545B0AEE3562D5CAA2CEE22CE2E112CE1215A3B4CB56E2D56AB5";
    attribute INIT_2E of inst : label is "5B3B844C6D518B8B86EE487A15552B3B96AE2ED107B0B912A384D21135A38B57";
    attribute INIT_2F of inst : label is "B4B4B4878C78D55B5B1E31AB96D6C792CD2CEE345605B3796AE88C62B2B12113";
    attribute INIT_30 of inst : label is "6CD6DE34B5B37AE3492D2078D61BBAE1BB8C7921E596C6D6D696AF2E0606D631";
    attribute INIT_31 of inst : label is "BBC78792C1E3492186DE49258C6D235B5B5B1E1BAC6C6D2C1E348C6C78787849";
    attribute INIT_32 of inst : label is "37C1F484B483484B1B1B37F5B1B4837878492D21F3BF48492C1B124861B1F4B4";
    attribute INIT_33 of inst : label is "F7C7CD234B7C1B7DF06CC7DF1F1E31E31807C1231B34B5F31231B487D38D2CD6";
    attribute INIT_34 of inst : label is "87DF1F1F1F124B06C7C79F1B37CC7C7D7DF493CC6C7C081F31E4B3486C484861";
    attribute INIT_35 of inst : label is "F30804F3793CD3D203CD234F7CC79302481F31E4C48080F31F0230B484F34834";
    attribute INIT_36 of inst : label is "C7C7C7C7C1F4C04F34F0F7CD3C3C07DE4C120C4863087CDF121F48C2087C1301";
    attribute INIT_37 of inst : label is "3CC30F01330F7D34C3C1F0231F02003CC3D30D303C21F0F1F1331F03CD3C303C";
    attribute INIT_38 of inst : label is "3C3DF0301F4C30C1F7C07C083C30C7C07F0C1F4C300F01F0C7C1301F0F0F07CC";
    attribute INIT_39 of inst : label is "F00F0030C31F0F30F30C1F7D3C303CD303020C0CC20C3C0CC31F7C3C3C3C030C";
    attribute INIT_3A of inst : label is "C300F0C3C0C3DF030F7CC30F30C0C0F30CC3C330C3C3C3CF0F0F4C07C0F30C00";
    attribute INIT_3B of inst : label is "F0F0F0F03030F0F00F0F0300C0C03C30F30C0C3C03C3C0C30C3CF30C0C0F03C3";
    attribute INIT_3C of inst : label is "3CC330C3C3C0300C3C3C0CC30F30F0C03C3C0C0C03C0F0C30C3CF0F03C3CF0F0";
    attribute INIT_3D of inst : label is "C0C0C3C30C00F00F0F030300F3C0C00C0C30C0C3C300300F030303003CF0F0C0";
    attribute INIT_3E of inst : label is "C3C330F30C0C3030CC3030F30C03C03003003CC30300F30C0C00F30C3C3C03C0";
    attribute INIT_3F of inst : label is "03CF0F0C3C0C03C0C0C0F0F0F3C3C3C0F00F3C3C30F30F0330C0F0C3C00F00F3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "9C94FAA821FD8AFD03A33E1F878008C3F8ED27784BE2C1EF791BEC8883690D3A";
    attribute INIT_01 of inst : label is "04B10012EF411260DE30E41C644FB18F09E8C7D1AAE0F2DA8798CF3E1EE0FD2A";
    attribute INIT_02 of inst : label is "8459E4170438245B332BC32087FC444D5FB2DE3EECD2345387DFF1E24DC786C5";
    attribute INIT_03 of inst : label is "48B853EBF59E0433239BF1669FF9C44A8011303CF7B81314C7B9051CC33C20BF";
    attribute INIT_04 of inst : label is "8D4878765AB497BF70BB911E564421FADF9C47BD387016642641B812CD578BA5";
    attribute INIT_05 of inst : label is "3A3EEC426C7B88CC923B34BB32BE446A9398314E862CF7C601704592116530FB";
    attribute INIT_06 of inst : label is "E512609DA3CC003AC01A3CD1511201B621E2B8F1C7C42FF5F6051B2F1ABC2EE4";
    attribute INIT_07 of inst : label is "F0DB8525CD39F33700FA0968010D5A0DDE37B884885AC4454607090915BBB380";
    attribute INIT_08 of inst : label is "BA56428C1E82BDF19B08D4A79E528DBF31360ABF0D3B6552D3D5B15E9B0D7444";
    attribute INIT_09 of inst : label is "562C26D2015E2E7A84684341AB6A6164DA181D490CC78F349631361E0A68316A";
    attribute INIT_0A of inst : label is "B43680E8E037D4B0ADFD0D5EF40E8174C436700C7EEE066E59368965DFCF3596";
    attribute INIT_0B of inst : label is "2C162C1C0193C6990684B556BE286E8F9CB072867E19C8539D05807B00D1F7CE";
    attribute INIT_0C of inst : label is "573AACABFD7154FA5F589634E6988084CCE303B34F7DC1F0D5F77759E50835F8";
    attribute INIT_0D of inst : label is "C561590A08A3B67FA0849BC348C478AD445B5EEC08B2739FA4F77B261FA50D61";
    attribute INIT_0E of inst : label is "222428D83DA8888F3738FDCB5F378C0926BABC1008CF2890D445FC562A36DCDD";
    attribute INIT_0F of inst : label is "0D43EB98A876C3C98BFD2B27F69B38E6317E2BBDFF7162A3C1E7762215437B2A";
    attribute INIT_10 of inst : label is "FAC9FCE14875C54FC0EA839D95336CBDC2215A1F6E7B4DF717FF3D92A3F664F8";
    attribute INIT_11 of inst : label is "FF925705EDC0EC94D808F9D39DD84FC3272C047F8239C5B30E7C5D0500F543C3";
    attribute INIT_12 of inst : label is "E725CB0393CE76E8993C6963F30C0595360F2F4C2BFC19A648673C00B7170E67";
    attribute INIT_13 of inst : label is "4096A593639FAC0A41BC359E4F0E46FC13360FA933F1863C0E1B088E6310F91C";
    attribute INIT_14 of inst : label is "8736FAC79570663A8C796391CDF393666203A3879C993269A56A5893CD30893D";
    attribute INIT_15 of inst : label is "823D18514848437DA1A0C59B934DA450C36265921E4F47B76DE48787EF3EB1A4";
    attribute INIT_16 of inst : label is "072867D52A8A2A2AC2A158A8AFAE0F79752127FA94872EDF8168609F44D85A24";
    attribute INIT_17 of inst : label is "61C8B24852D5DCA61D585618AF72498BB572A09BAEAE0B7435EFB548CABA0ABD";
    attribute INIT_18 of inst : label is "579E15E8521C872BA82795555E0AFAD742AEBAEEC92AC92726E8A255D5D592DF";
    attribute INIT_19 of inst : label is "A286AE1EC5BBAC7B272E5E09F57EE2D3A95C772B2EB55C92A86E1D55927ED09F";
    attribute INIT_1A of inst : label is "7D112FB879785447D134B06CB9146E0BA45CACB87876D44D1842A0916AB6EEFB";
    attribute INIT_1B of inst : label is "AA21EC6ABA1E0ACAEB54EE1B91AB8DD1EC5492B46B4B06CB92EE5AD5C5BE2055";
    attribute INIT_1C of inst : label is "F7AB4BD2AEB1BAD11B1B1E34B1B05486DB4B06F4AE48BB5B4E3BABB87BE415A0";
    attribute INIT_1D of inst : label is "2F18D23AD5EBEB34BD288DB61BADE1A168DE1B4BD21FAF5B1B3AAE34B1B786D6";
    attribute INIT_1E of inst : label is "1B1BD21E09278DE1E06CD21E121EBD2C1B1B1878D21231BDEAD2F084B3787AE1";
    attribute INIT_1F of inst : label is "492348DF121EDE4E37D3C1E79E1E34B60B1B186C4B06CDE49E31B06C6D2F1B7B";
    attribute INIT_20 of inst : label is "E1E31B186D20F0861B06CD2F1B7D21F1B7C78D231F06C184B06DB6D21E06F192";
    attribute INIT_21 of inst : label is "B3781F1B1E0B7C7C792DEC6CDE1E07CDE0231E37D2C18DE6DF4B34B06F1F378D";
    attribute INIT_22 of inst : label is "0E30E3083DB7D212487DE48230848C3CDF7C1237DE31F048C7DE37C3CD209234";
    attribute INIT_23 of inst : label is "CC230B7D3C2CDF1FC2C7C31B1BC2D2C2C20208C3C1F37C09E7C3C6182C7D3CDF";
    attribute INIT_24 of inst : label is "3CDF37CC230F37C08C0FC20F37C083DFC27C0F3080F07CD3C2C7C3C1B0F37CC3";
    attribute INIT_25 of inst : label is "30F083CC3CC3DF34F0C0F00F07F0C08C3C3DF7C2083C3C3C3D3F083D3C2DF37C";
    attribute INIT_26 of inst : label is "0F33CCF30F030F30F0F30C0C0CC20F33C3C3F0F3C3C1F30F7F0CDF083C303F0F";
    attribute INIT_27 of inst : label is "33CC330C0F0F0F0F0F30C3F0C3C3C3DF0F30F0F7C3F0F0F3DF0F7DF7C3CC330C";
    attribute INIT_28 of inst : label is "CF0F0F3C3CF3CF30F0F03CF30F0F0F0330F0F0C30F0F0C3C3CF30F0C0C3CC30F";
    attribute INIT_29 of inst : label is "0C3CC30C0F33C3C3CC3C0F03C3F3C0C0CC30C3C3C30FCF0F3C3C3CF0F30C3CC3";
    attribute INIT_2A of inst : label is "0F03C3C3C0F03CF0F0F0F0F0F03C303CCF3C0C3CC3CCF0F0F0F030C3C3C3C3CF";
    attribute INIT_2B of inst : label is "CFC30303C0F30C0C0F30F0C30F33C0CC30C3C3CC3CF30C30C30FCF3C3CF0FC3C";
    attribute INIT_2C of inst : label is "30F0F0F0330F0F303C0F3C3C3030F0C0C3C3CC3C03C0F30F33C3C330F0F0CC3C";
    attribute INIT_2D of inst : label is "C3CF03F33C3C0C0F03CF30C3C3C3C3CCF03CC3C303CC3030F33CC3C3C3C30F3C";
    attribute INIT_2E of inst : label is "0F33C0CC3C30C3C3C3CF0C3C30C30F33C3CF0FC303F03C30F30CC30330F30F0F";
    attribute INIT_2F of inst : label is "F0F0F0C3CC3CC30F0F0F30F3C3C3C3C3CC3CCF30C300F33C3CF0CC30F0F03033";
    attribute INIT_30 of inst : label is "3CC3CF30F0F33CF30C3C303CC30F3CF0F3CC3C30F0C3C3C3C3C3CF0F0303C330";
    attribute INIT_31 of inst : label is "F3C3C3C3C0F30C30C3CF0C30CC3C330F0F0F0F0F3C3C3C3C0F30CC3C3C3C3C0C";
    attribute INIT_32 of inst : label is "33C0F0C0F0C30C0F0F0F33F0F0F0C33C3C0C3C30F33F0C0C3C0F030C30F0F0F0";
    attribute INIT_33 of inst : label is "F3C3CC330F3C0F3CF03CC3CF0F0F30F30C03C0330F30F0F30330F0C3C3CC3CC3";
    attribute INIT_34 of inst : label is "C3CF0F0F0F030F03C3C3CF0F33CC3C3C3CF0C3CC3C3C0C0F30F0F30C3C0C0C30";
    attribute INIT_35 of inst : label is "F30C00F33C3CC3C303CC330F3CC3C3030C0F30F0C0C0C0F30F0330F0C0F30C30";
    attribute INIT_36 of inst : label is "C3C3C3C3C0F0C00F30F0F3CC3C3C03CF0C030C0C330C3CCF030F0CC30C3C0300";
    attribute INIT_37 of inst : label is "3CC30F00330F3C30C3C0F0330F03003CC3C30C303C30F0F0F0330F03CC3C303C";
    attribute INIT_38 of inst : label is "3C3CF0300F0C30C0F3C03C0C3C30C3C03F0C0F0C300F00F0C3C0300F0F0F03CC";
    attribute INIT_39 of inst : label is "F00F0030C30F0F30F30C0F3C3C303CC303030C0CC30C3C0CC30F3C3C3C3C030C";
    attribute INIT_3A of inst : label is "C300F0C3C0C3CF030F3CC30F30C0C0F30CC3C330C3C3C3CF0F0F0C03C0F30C00";
    attribute INIT_3B of inst : label is "F0F0F0F03030F0F00F0F0300C0C03C30F30C0C3C03C3C0C30C3CF30C0C0F03C3";
    attribute INIT_3C of inst : label is "3CC330C3C3C0300C3C3C0CC30F30F0C03C3C0C0C03C0F0C30C3CF0F03C3CF0F0";
    attribute INIT_3D of inst : label is "C0C0C3C30C00F00F0F030300F3C0C00C0C30C0C3C300300F030303003CF0F0C0";
    attribute INIT_3E of inst : label is "C3C330F30C0C3030CC3030F30C03C03003003CC30300F30C0C00F30C3C3C03C0";
    attribute INIT_3F of inst : label is "03CF0F0C3C0C03C0C0C0F0F0F3C3C3C0F00F3C3C30F30F0330C0F0C3C00F00F3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "297568A2D7475686D689D35A2C6B96785B16CA86B16C75A1C75A175B5A89E2D6";
    attribute INIT_01 of inst : label is "D6A5B6D5A1B5B5CB289E1B578B568B569CA2786CA31E1A8A3875749A568B46CA";
    attribute INIT_02 of inst : label is "39758E5A978B5D74A68A368B5A4D6D6A34CA34D292A5A96D38691B1CD7569696";
    attribute INIT_03 of inst : label is "A387968A1CA35DA29C74A5D72892A5DA5B978B8728696D5E38696D7578D38E29";
    attribute INIT_04 of inst : label is "5729C9C9A31D7291CB4A2D74DA5B5D292935D692C78E5D7368E5C797575CA28D";
    attribute INIT_05 of inst : label is "A3592978D392A2A29D5CA5A4D71A5DA28D72CB2A29D34D2CB5CB3696D75CD74A";
    attribute INIT_06 of inst : label is "2975CB28A875B389A6CA875797975E4D75A59A1E29978C97297974E4E292D28D";
    attribute INIT_07 of inst : label is "968A5A9A2A5995D5CE26972A6CE35CB28A8A275A9A5C7979797697697598C9A7";
    attribute INIT_08 of inst : label is "8A35A99A666992968CA99A632669A29299CCD964B5A28D793935CDA4D6757369";
    attribute INIT_09 of inst : label is "A5CA6966A9A6598A5B5769A68CA35D6999A5D7366972A28DA5CA98E4E6638D72";
    attribute INIT_0A of inst : label is "96CA3A2A2A995D668A25D69963A2A68D769999E358A29CA2A5CA369728728D69";
    attribute INIT_0B of inst : label is "CA75CA976A665CA69A39973658DA59963299CA3658D97368CA9A3A59A75D6259";
    attribute INIT_0C of inst : label is "5CA63299265CD74A3599A5CA65A35E5D728D7628D8A5735A5A58CA359A69A659";
    attribute INIT_0D of inst : label is "9A5D72A975CA28D2975D71A5A96A6599A759A28A75CA68A269662968E4A5D69A";
    attribute INIT_0E of inst : label is "DA5DA5A38A2A36995CA34A59A1CA35D75C9963979A34D976975D63696968A5A2";
    attribute INIT_0F of inst : label is "B57928A5A5A65D36964A68A64A35CA28D75968A2928DA59CA7289A5D75B59968";
    attribute INIT_10 of inst : label is "1A29935D75A5A5D65B1A5A59A5D68A6575D76968A28A5A28DA18A575A595CA65";
    attribute INIT_11 of inst : label is "58A6969D65768A67576995A65A29D65A5A65E758A68A368A695A5A75E695DA5A";
    attribute INIT_12 of inst : label is "2969969A5A568A29A5A5A5A5969A75A5A5D65969D61A69696A5A59B695D69696";
    attribute INIT_13 of inst : label is "A6A5A5A65A595A759D65A5A296969A25DA5A68A5A5969A5A696969A2969D65D7";
    attribute INIT_14 of inst : label is "A5A595A65A69A5A59A5A5A5D6965A5A5A69A5CA65A5A6969696969A659A69A59";
    attribute INIT_15 of inst : label is "9A65A9A69A6A6A596969A695A66969A69A5A5A5A96997595A569A5A596596696";
    attribute INIT_16 of inst : label is "A696A569A5A5A5A59A5A96969656995A5A69A595A6A5A595A696A6966996A5A6";
    attribute INIT_17 of inst : label is "696A5A69A65A56969696A5A9965A69695A5A5A959656995A66595A696965A959";
    attribute INIT_18 of inst : label is "A5966996A696A5A596A59A69A5A965696A59596569A569A5A65A5A696969A659";
    attribute INIT_19 of inst : label is "696965A569965695A5A5A5A95A565A59969695A5A596969A5A65A5A69A565A95";
    attribute INIT_1A of inst : label is "569A95969696A6A5699A5A96969A65A96696969696965A669A6A5A9A65965959";
    attribute INIT_1B of inst : label is "969A569659A5A96965A665A59A59665A569A695A65A5A9696965A5696A569A9A";
    attribute INIT_1C of inst : label is "5965A569965A5969A5A5A59A5A5A9A6965A5A95A65A695A5A599659695669A5A";
    attribute INIT_1D of inst : label is "95A669996659659A569A6659A5965A5A9665A5A569A595A5A599659A5A596969";
    attribute INIT_1E of inst : label is "A5A569A5A699665A5A9669A5A9A59696A5A5A69669A99A5659695A6A5996965A";
    attribute INIT_1F of inst : label is "A699A665A9A565A599696A5965A59A59A5A5A696A5A9665A659A5A969695A595";
    attribute INIT_20 of inst : label is "5A59A5A6969A5A69A5A96695A5969A5A59696699A5A96A6A5A965969A5A95A69";
    attribute INIT_21 of inst : label is "5996A5A5A5A596969696569665A5A9665A99A599696A665965A59A5A95A59966";
    attribute INIT_22 of inst : label is "A59A59A6965969A9A6965A699A6A66966596A999659A5AA669659969669A699A";
    attribute INIT_23 of inst : label is "6699A596969665A5696969A5A569696969A9A6696A5996A6596969A696969665";
    attribute INIT_24 of inst : label is "9665996699A5996A66A569A5996A69656996A59A6A5A96696969696A5A599669";
    attribute INIT_25 of inst : label is "9A5A69669669659A5A6A5AA5A95A6A6696965969A69696969695A69696965996";
    attribute INIT_26 of inst : label is "A5996659A5A9A59A5A59A6A6A669A59969695A59696A59A595A665A6969A95A5";
    attribute INIT_27 of inst : label is "996699A6A5A5A5A5A59A695A69696965A59A5A59695A5A5965A59659696699A6";
    attribute INIT_28 of inst : label is "65A5A5969659659A5A5A9659A5A5A5A99A5A5A69A5A5A6969659A5A6A69669A5";
    attribute INIT_29 of inst : label is "A69669A6A59969696696A5A969596A6A669A696969A565A59696965A59A69669";
    attribute INIT_2A of inst : label is "A5A969696A5A965A5A5A5A5A5A969A966596A69669665A5A5A5A9A6969696965";
    attribute INIT_2B of inst : label is "6569A9A96A59A6A6A59A5A69A5996A669A6969669659A69A69A56596965A5696";
    attribute INIT_2C of inst : label is "9A5A5A5A99A5A59A96A596969A9A5A6A69696696A96A59A59969699A5A5A6696";
    attribute INIT_2D of inst : label is "6965A9599696A6A5A9659A69696969665A966969A9669A9A599669696969A596";
    attribute INIT_2E of inst : label is "A5996A66969A69696965A6969A69A5996965A569A95A969A59A669A99A59A5A5";
    attribute INIT_2F of inst : label is "5A5A5A69669669A5A5A59A59696969696696659A69AA5996965A669A5A5A9A99";
    attribute INIT_30 of inst : label is "9669659A5A599659A6969A9669A5965A5966969A5A696969696965A5A9A9699A";
    attribute INIT_31 of inst : label is "596969696A59A69A6965A69A669699A5A5A5A5A596969696A59A6696969696A6";
    attribute INIT_32 of inst : label is "996A5A6A5A69A6A5A5A5995A5A5A699696A6969A5995A6A696A5A9A69A5A5A5A";
    attribute INIT_33 of inst : label is "59696699A596A5965A966965A5A59A59A6A96A99A59A5A59A99A5A6969669669";
    attribute INIT_34 of inst : label is "6965A5A5A5A9A5A9696965A599669696965A69669696A6A59A5A59A696A6A69A";
    attribute INIT_35 of inst : label is "59A6AA5996966969A96699A5966969A9A6A59A5A6A6A6A59A5A99A5A6A59A69A";
    attribute INIT_36 of inst : label is "696969696A5A6AA59A5A59669696A965A6A9A6A699A69665A9A5A669A696A9AA";
    attribute INIT_37 of inst : label is "9669A5AA99A5969A696A5A99A5A9AA966969A69A969A5A5A5A99A5A966969A96";
    attribute INIT_38 of inst : label is "96965A9AA5A69A6A596A96A6969A696A95A6A5A69AA5AA5A696A9AA5A5A5A966";
    attribute INIT_39 of inst : label is "5AA5AA9A69A5A59A59A6A596969A9669A9A9A6A669A696A669A596969696A9A6";
    attribute INIT_3A of inst : label is "69AA5A696A6965A9A59669A59A6A6A59A669699A69696965A5A5A6A96A59A6AA";
    attribute INIT_3B of inst : label is "5A5A5A5A9A9A5A5AA5A5A9AA6A6A969A59A6A696A9696A69A69659A6A6A5A969";
    attribute INIT_3C of inst : label is "96699A69696A9AA69696A669A59A5A6A9696A6A6A96A5A69A6965A5A96965A5A";
    attribute INIT_3D of inst : label is "6A6A6969A6AA5AA5A5A9A9AA596A6AA6A69A6A6969AA9AA5A9A9A9AA965A5A6A";
    attribute INIT_3E of inst : label is "69699A59A6A69A9A669A9A59A6A96A9AA9AA9669A9AA59A6A6AA59A69696A96A";
    attribute INIT_3F of inst : label is "A965A5A696A6A96A6A6A5A5A5969696A5AA596969A59A5A99A6A5A696AA5AA59";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
