-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "813864D36D435B69E9B9A490D4F50A404088AA9A42498AC9282FFB807AE11162";
    attribute INIT_01 of inst : label is "20481A048120481A04831BA7A61C3C1FFAFF3FF8FF23931F69A69A569A69A049";
    attribute INIT_02 of inst : label is "C74CA2DFF62483A7A639E2E59659C80A14080082EE4D3273CA49C92048120681";
    attribute INIT_03 of inst : label is "403D813E433D0380EC03F60CFF204481F808484848024920C925122804464221";
    attribute INIT_04 of inst : label is "B3488EA40282A80120080120080126648532428C010101008A3E2E5401BC0701";
    attribute INIT_05 of inst : label is "F33A89084484220200264A530484FF775664A532529829008890844100848484";
    attribute INIT_06 of inst : label is "B0058548161400051208890444005850140C29402A2401120088000050585280";
    attribute INIT_07 of inst : label is "E2DC2F80D856FF88F421101025101058356E181200D820A611B822E5A2480480";
    attribute INIT_08 of inst : label is "D02880C8099999202A66666808D999920AA66664808975D00000A1E499400000";
    attribute INIT_09 of inst : label is "0EFE9C962DC2FD20A44881002000881020148D225A6078445111F00000000000";
    attribute INIT_0A of inst : label is "810000148D22FF8EF48291200400000200548D228D6978D44444F00000000000";
    attribute INIT_0B of inst : label is "C8284A80DC80808B7742F9480480FFE0FFCEFF48291220548D22FFCEFD20A448";
    attribute INIT_0C of inst : label is "C2FF41C7CD264583458A5013430C4C2903453B10040054820042190445194E20";
    attribute INIT_0D of inst : label is "8B548E54C2C4959682C34A568005FBE84800000DFBF1325544A164641570C201";
    attribute INIT_0E of inst : label is "FFEEE23AFFC9D282E6755555554AAABFF5555A641C822E840595632CA0881110";
    attribute INIT_0F of inst : label is "6003880C808080604CFDFF47FF8C04A9180101284300222042180514098E7598";
    attribute INIT_10 of inst : label is "D02880C8099999202A66666808D999920AA66664808975D00000A1E499400000";
    attribute INIT_11 of inst : label is "0EFE9C962DC2FD20A44881002000881020148D225A6078445111F00000000000";
    attribute INIT_12 of inst : label is "810000148D22FF8EF48291200400000200548D228D6978D44444F00000000000";
    attribute INIT_13 of inst : label is "C8284A80DC80808B7742F9480480FFE0FFCEFF48291220548D22FFCEFD20A448";
    attribute INIT_14 of inst : label is "C2FF41C7CD264583458A5013430C4C2903453B10040054820042190445194E20";
    attribute INIT_15 of inst : label is "8B548E54C2C4959682C34A568005FBE84800000DFBF1325544A164641570C201";
    attribute INIT_16 of inst : label is "FFEEE23AFFC9D282E6755555554AAABFF5555A641C822E840595632CA0881110";
    attribute INIT_17 of inst : label is "6003880C808080604CFDFF47FF8C04A9180101284300222042180514098E7598";
    attribute INIT_18 of inst : label is "D02880C8099999202A66666808D999920AA66664808975D00000A1E499400000";
    attribute INIT_19 of inst : label is "0EFE9C962DC2FD20A44881002000881020148D225A6078445111F00000000000";
    attribute INIT_1A of inst : label is "810000148D22FF8EF48291200400000200548D228D6978D44444F00000000000";
    attribute INIT_1B of inst : label is "C8284A80DC80808B7742F9480480FFE0FFCEFF48291220548D22FFCEFD20A448";
    attribute INIT_1C of inst : label is "C2FF41C7CD264583458A5013430C4C2903453B10040054820042190445194E20";
    attribute INIT_1D of inst : label is "8B548E54C2C4959682C34A568005FBE84800000DFBF1325544A164641570C201";
    attribute INIT_1E of inst : label is "FFEEE23AFFC9D282E6755555554AAABFF5555A641C822E840595632CA0881110";
    attribute INIT_1F of inst : label is "6003880C808080604CFDFF47FF8C04A9180101284300222042180514098E7598";
    attribute INIT_20 of inst : label is "D02880C8099999202A66666808D999920AA66664808975D00000A1E499400000";
    attribute INIT_21 of inst : label is "0EFE9C962DC2FD20A44881002000881020148D225A6078445111F00000000000";
    attribute INIT_22 of inst : label is "810000148D22FF8EF48291200400000200548D228D6978D44444F00000000000";
    attribute INIT_23 of inst : label is "C8284A80DC80808B7742F9480480FFE0FFCEFF48291220548D22FFCEFD20A448";
    attribute INIT_24 of inst : label is "C2FF41C7CD264583458A5013430C4C2903453B10040054820042190445194E20";
    attribute INIT_25 of inst : label is "8B548E54C2C4959682C34A568005FBE84800000DFBF1325544A164641570C201";
    attribute INIT_26 of inst : label is "FFEEE23AFFC9D282E6755555554AAABFF5555A641C822E840595632CA0881110";
    attribute INIT_27 of inst : label is "6003880C808080604CFDFF47FF8C04A9180101284300222042180514098E7598";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "F817412CB6B98C9636C6D96D451150035410F5796D689F8CBD9AA8FB93199D6D";
    attribute INIT_01 of inst : label is "4B32C4B12CCB32C4B128F305055272555455555C551ADE1E420820E020820A00";
    attribute INIT_02 of inst : label is "BB577B75565B6F0507D04DA49249E85B6B64AD260932B59AA249ECCB32CCB12C";
    attribute INIT_03 of inst : label is "530B8A6B328D27CC4731AC21FD1A2293FABABABABDB49249FFEE697EE0BD3028";
    attribute INIT_04 of inst : label is "7D3337EC94545E4BFA7E4BFA7E4BFD9B5ECDAF6302CACAC9F3FF4760B81EE398";
    attribute INIT_05 of inst : label is "C45F66D3B369D9B4ECC895E44969F88BF19B5ECDAF66D783322539164B6B6B6B";
    attribute INIT_06 of inst : label is "F49E8FD16A3FD24ACDB766DBB309E8F926F47FA4B59B7ECDBF66DFB3A9E8FD49";
    attribute INIT_07 of inst : label is "C7EE7F49E8FDFF33F43B5BF59B49B4CEA7277F7EEE4AEE7DCC9D04540F6DB249";
    attribute INIT_08 of inst : label is "D08DA9D49AAAA8036E2AAA00FB8AAA883672AAA20D9CCBCA0220DF934FC00000";
    attribute INIT_09 of inst : label is "994A11CC76E5F00700ED79834E6057894E201805AFDC13C02008F00000000000";
    attribute INIT_0A of inst : label is "F9836E601805FF77C11C23B6E60DF9816E2118456B97C9C80200F00000000000";
    attribute INIT_0B of inst : label is "EA6DA7A98D49A91EABE7F96DB249FFC0FF77FC11C23B6E611845FF77F00700ED";
    attribute INIT_0C of inst : label is "47FF48F2C08366910D188C850D20D4B0D88D29726A86D4945A52544CD8333C49";
    attribute INIT_0D of inst : label is "64CC95CD96A7373AC4729B9CE34242470903C0520252D94CC9B191D87FDA8B28";
    attribute INIT_0E of inst : label is "FFEDD55FFFF30E5A03D99999998CCCD559999FBE7D7FF6622373251B9F937A8D";
    attribute INIT_0F of inst : label is "2909DA9D49A9AB6CF774FF4EFF1109A95BB24268552D0CAE42A96C30401CEDB9";
    attribute INIT_10 of inst : label is "D08DA9D49AAAA8036E2AAA00FB8AAA883672AAA20D9CCBCA0220DF934FC00000";
    attribute INIT_11 of inst : label is "994A11CC76E5F00700ED79834E6057894E201805AFDC13C02008F00000000000";
    attribute INIT_12 of inst : label is "F9836E601805FF77C11C23B6E60DF9816E2118456B97C9C80200F00000000000";
    attribute INIT_13 of inst : label is "EA6DA7A98D49A91EABE7F96DB249FFC0FF77FC11C23B6E611845FF77F00700ED";
    attribute INIT_14 of inst : label is "47FF48F2C08366910D188C850D20D4B0D88D29726A86D4945A52544CD8333C49";
    attribute INIT_15 of inst : label is "64CC95CD96A7373AC4729B9CE34242470903C0520252D94CC9B191D87FDA8B28";
    attribute INIT_16 of inst : label is "FFEDD55FFFF30E5A03D99999998CCCD559999FBE7D7FF6622373251B9F937A8D";
    attribute INIT_17 of inst : label is "2909DA9D49A9AB6CF774FF4EFF1109A95BB24268552D0CAE42A96C30401CEDB9";
    attribute INIT_18 of inst : label is "D08DA9D49AAAA8036E2AAA00FB8AAA883672AAA20D9CCBCA0220DF934FC00000";
    attribute INIT_19 of inst : label is "994A11CC76E5F00700ED79834E6057894E201805AFDC13C02008F00000000000";
    attribute INIT_1A of inst : label is "F9836E601805FF77C11C23B6E60DF9816E2118456B97C9C80200F00000000000";
    attribute INIT_1B of inst : label is "EA6DA7A98D49A91EABE7F96DB249FFC0FF77FC11C23B6E611845FF77F00700ED";
    attribute INIT_1C of inst : label is "47FF48F2C08366910D188C850D20D4B0D88D29726A86D4945A52544CD8333C49";
    attribute INIT_1D of inst : label is "64CC95CD96A7373AC4729B9CE34242470903C0520252D94CC9B191D87FDA8B28";
    attribute INIT_1E of inst : label is "FFEDD55FFFF30E5A03D99999998CCCD559999FBE7D7FF6622373251B9F937A8D";
    attribute INIT_1F of inst : label is "2909DA9D49A9AB6CF774FF4EFF1109A95BB24268552D0CAE42A96C30401CEDB9";
    attribute INIT_20 of inst : label is "D08DA9D49AAAA8036E2AAA00FB8AAA883672AAA20D9CCBCA0220DF934FC00000";
    attribute INIT_21 of inst : label is "994A11CC76E5F00700ED79834E6057894E201805AFDC13C02008F00000000000";
    attribute INIT_22 of inst : label is "F9836E601805FF77C11C23B6E60DF9816E2118456B97C9C80200F00000000000";
    attribute INIT_23 of inst : label is "EA6DA7A98D49A91EABE7F96DB249FFC0FF77FC11C23B6E611845FF77F00700ED";
    attribute INIT_24 of inst : label is "47FF48F2C08366910D188C850D20D4B0D88D29726A86D4945A52544CD8333C49";
    attribute INIT_25 of inst : label is "64CC95CD96A7373AC4729B9CE34242470903C0520252D94CC9B191D87FDA8B28";
    attribute INIT_26 of inst : label is "FFEDD55FFFF30E5A03D99999998CCCD559999FBE7D7FF6622373251B9F937A8D";
    attribute INIT_27 of inst : label is "2909DA9D49A9AB6CF774FF4EFF1109A95BB24268552D0CAE42A96C30401CEDB9";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "F897536DB694A5B616C6C96C0D43540AFC0E77C12D188E8EFFAAA8935E341409";
    attribute INIT_01 of inst : label is "1A5695A5691A4691A46A518D8FD353555C55555C550A10BE1A69A6A1A69A7A04";
    attribute INIT_02 of inst : label is "AC97B5B982124B8D8D50833CF3CFC01249248002225BA62A87FFC11A5691A469";
    attribute INIT_03 of inst : label is "43085051B88C220C6831A341E85E231180A0A0A0AA492492FFFA08F4607A3168";
    attribute INIT_04 of inst : label is "B864CFF88E1E1566939566939566955266A9334A02A2A2888600506B38B0E018";
    attribute INIT_05 of inst : label is "DBBF5498AA4C55262A95276A8ACAFA67FD5266A933549982A549CAA28ACACACA";
    attribute INIT_06 of inst : label is "00890780741F9002A9315498AA08D07900E83F20055262A9315498AAC8D07E40";
    attribute INIT_07 of inst : label is "C39E3008D078FF08E00B40B40B40B41C804E7B1F6098E63EC13900E523000000";
    attribute INIT_08 of inst : label is "80A908C400EEE801623BBA00588EEE801623BBA00588E1422022B3E278C00000";
    attribute INIT_09 of inst : label is "3213183435E1F12124211C00470015C04704892164BED7420008F00000000000";
    attribute INIT_0A of inst : label is "1C0047058961FF0FC484908570011C0047048921201912C00202F00000000000";
    attribute INIT_0B of inst : label is "E2206348D840080C47E3FC000000FFC0FF0FFC584B0847058961FF0FF1612C21";
    attribute INIT_0C of inst : label is "03FF04AAC23799AA4730CC0553014C6CF0845B10112D51C01457024645055CD0";
    attribute INIT_0D of inst : label is "2588048C202666D8C1C8B35ADDA2888C408C0062C88051488331C4202A924B18";
    attribute INIT_0E of inst : label is "FFE2DBBFFFE1D6B250FE1E1E1E0F0F199E1E030528AE54430223011118070C8E";
    attribute INIT_0F of inst : label is "080B118C401808816EF5FF16FF225AAA0AA096A88309492244184840C2022038";
    attribute INIT_10 of inst : label is "80A908C400EEE801623BBA00588EEE801623BBA00588E1422022B3E278C00000";
    attribute INIT_11 of inst : label is "3213183435E1F12124211C00470015C04704892164BED7420008F00000000000";
    attribute INIT_12 of inst : label is "1C0047058961FF0FC484908570011C0047048921201912C00202F00000000000";
    attribute INIT_13 of inst : label is "E2206348D840080C47E3FC000000FFC0FF0FFC584B0847058961FF0FF1612C21";
    attribute INIT_14 of inst : label is "03FF04AAC23799AA4730CC0553014C6CF0845B10112D51C01457024645055CD0";
    attribute INIT_15 of inst : label is "2588048C202666D8C1C8B35ADDA2888C408C0062C88051488331C4202A924B18";
    attribute INIT_16 of inst : label is "FFE2DBBFFFE1D6B250FE1E1E1E0F0F199E1E030528AE54430223011118070C8E";
    attribute INIT_17 of inst : label is "080B118C401808816EF5FF16FF225AAA0AA096A88309492244184840C2022038";
    attribute INIT_18 of inst : label is "80A908C400EEE801623BBA00588EEE801623BBA00588E1422022B3E278C00000";
    attribute INIT_19 of inst : label is "3213183435E1F12124211C00470015C04704892164BED7420008F00000000000";
    attribute INIT_1A of inst : label is "1C0047058961FF0FC484908570011C0047048921201912C00202F00000000000";
    attribute INIT_1B of inst : label is "E2206348D840080C47E3FC000000FFC0FF0FFC584B0847058961FF0FF1612C21";
    attribute INIT_1C of inst : label is "03FF04AAC23799AA4730CC0553014C6CF0845B10112D51C01457024645055CD0";
    attribute INIT_1D of inst : label is "2588048C202666D8C1C8B35ADDA2888C408C0062C88051488331C4202A924B18";
    attribute INIT_1E of inst : label is "FFE2DBBFFFE1D6B250FE1E1E1E0F0F199E1E030528AE54430223011118070C8E";
    attribute INIT_1F of inst : label is "080B118C401808816EF5FF16FF225AAA0AA096A88309492244184840C2022038";
    attribute INIT_20 of inst : label is "80A908C400EEE801623BBA00588EEE801623BBA00588E1422022B3E278C00000";
    attribute INIT_21 of inst : label is "3213183435E1F12124211C00470015C04704892164BED7420008F00000000000";
    attribute INIT_22 of inst : label is "1C0047058961FF0FC484908570011C0047048921201912C00202F00000000000";
    attribute INIT_23 of inst : label is "E2206348D840080C47E3FC000000FFC0FF0FFC584B0847058961FF0FF1612C21";
    attribute INIT_24 of inst : label is "03FF04AAC23799AA4730CC0553014C6CF0845B10112D51C01457024645055CD0";
    attribute INIT_25 of inst : label is "2588048C202666D8C1C8B35ADDA2888C408C0062C88051488331C4202A924B18";
    attribute INIT_26 of inst : label is "FFE2DBBFFFE1D6B250FE1E1E1E0F0F199E1E030528AE54430223011118070C8E";
    attribute INIT_27 of inst : label is "080B118C401808816EF5FF16FF225AAA0AA096A88309492244184840C2022038";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0AA4029B68A52369ED3934D1581640228C0E70536314CFE6C75FF8BD93D0C041";
    attribute INIT_01 of inst : label is "4250942509024090240AB0AAAAD59592A52A42A52A08DDAE0924922892492815";
    attribute INIT_02 of inst : label is "E1790ADE03524AAAAAD000D96596C14008001249604B1622CDB6C14250942509";
    attribute INIT_03 of inst : label is "021C7840D80806984B6173E1E86E0023A0B0B0B0BA492492B6DA081040082140";
    attribute INIT_04 of inst : label is "7F1AA6E212121556D2B546D2B556D55AD6AD6B4B0AC2C2E17AD090C810324130";
    attribute INIT_05 of inst : label is "E21B5691AB48D5A46AD5AC6AEB4BFC436D5AD6AD6B56B582B5695ABAEB4B4B4B";
    attribute INIT_06 of inst : label is "4115AD8846B60342AD235691AB211ADC30AD6D06855A56AD2B5695AB615ADB0D";
    attribute INIT_07 of inst : label is "F31D30811ADAFFABE00908908908909102488D20A4950A41492204A12B0C30C3";
    attribute INIT_08 of inst : label is "A02631B0D31110462684441189A1110462684441189A07C5C594CD830DC00000";
    attribute INIT_09 of inst : label is "99C913C731F1F92925210C80432014C84324A9291BC700C90E26F00000000000";
    attribute INIT_0A of inst : label is "0C804324A929FF8FE4A4948432010C804324A929EBA7C9C11110F00000000000";
    attribute INIT_0B of inst : label is "C06023519B0D31CD17D3F8451451FFE0FF8FFE4A49484324A929FF8FF9292521";
    attribute INIT_0C of inst : label is "D6FEAD0942AF11B66B361E84D3A1EEB5C0A85377555D8AAB44AAAC2C91467CDD";
    attribute INIT_0D of inst : label is "FA8DDE91E5BDA554B716D2B6A3170A15BD71C2874A1B76B6ED2D1AD7777405A0";
    attribute INIT_0E of inst : label is "FFC1E03BFFD9AB0C9C5FE01FE00FF01E1FE011BDFC75AF6C7BA477DD25DA3128";
    attribute INIT_0F of inst : label is "410242190D212B0980F3FE92FFAABB14A9BAAEC52BA80D44A95D427402DCC9CD";
    attribute INIT_10 of inst : label is "A02631B0D31110462684441189A1110462684441189A07C5C594CD830DC00000";
    attribute INIT_11 of inst : label is "99C913C731F1F92925210C80432014C84324A9291BC700C90E26F00000000000";
    attribute INIT_12 of inst : label is "0C804324A929FF8FE4A4948432010C804324A929EBA7C9C11110F00000000000";
    attribute INIT_13 of inst : label is "C06023519B0D31CD17D3F8451451FFE0FF8FFE4A49484324A929FF8FF9292521";
    attribute INIT_14 of inst : label is "D6FEAD0942AF11B66B361E84D3A1EEB5C0A85377555D8AAB44AAAC2C91467CDD";
    attribute INIT_15 of inst : label is "FA8DDE91E5BDA554B716D2B6A3170A15BD71C2874A1B76B6ED2D1AD7777405A0";
    attribute INIT_16 of inst : label is "FFC1E03BFFD9AB0C9C5FE01FE00FF01E1FE011BDFC75AF6C7BA477DD25DA3128";
    attribute INIT_17 of inst : label is "410242190D212B0980F3FE92FFAABB14A9BAAEC52BA80D44A95D427402DCC9CD";
    attribute INIT_18 of inst : label is "A02631B0D31110462684441189A1110462684441189A07C5C594CD830DC00000";
    attribute INIT_19 of inst : label is "99C913C731F1F92925210C80432014C84324A9291BC700C90E26F00000000000";
    attribute INIT_1A of inst : label is "0C804324A929FF8FE4A4948432010C804324A929EBA7C9C11110F00000000000";
    attribute INIT_1B of inst : label is "C06023519B0D31CD17D3F8451451FFE0FF8FFE4A49484324A929FF8FF9292521";
    attribute INIT_1C of inst : label is "D6FEAD0942AF11B66B361E84D3A1EEB5C0A85377555D8AAB44AAAC2C91467CDD";
    attribute INIT_1D of inst : label is "FA8DDE91E5BDA554B716D2B6A3170A15BD71C2874A1B76B6ED2D1AD7777405A0";
    attribute INIT_1E of inst : label is "FFC1E03BFFD9AB0C9C5FE01FE00FF01E1FE011BDFC75AF6C7BA477DD25DA3128";
    attribute INIT_1F of inst : label is "410242190D212B0980F3FE92FFAABB14A9BAAEC52BA80D44A95D427402DCC9CD";
    attribute INIT_20 of inst : label is "A02631B0D31110462684441189A1110462684441189A07C5C594CD830DC00000";
    attribute INIT_21 of inst : label is "99C913C731F1F92925210C80432014C84324A9291BC700C90E26F00000000000";
    attribute INIT_22 of inst : label is "0C804324A929FF8FE4A4948432010C804324A929EBA7C9C11110F00000000000";
    attribute INIT_23 of inst : label is "C06023519B0D31CD17D3F8451451FFE0FF8FFE4A49484324A929FF8FF9292521";
    attribute INIT_24 of inst : label is "D6FEAD0942AF11B66B361E84D3A1EEB5C0A85377555D8AAB44AAAC2C91467CDD";
    attribute INIT_25 of inst : label is "FA8DDE91E5BDA554B716D2B6A3170A15BD71C2874A1B76B6ED2D1AD7777405A0";
    attribute INIT_26 of inst : label is "FFC1E03BFFD9AB0C9C5FE01FE00FF01E1FE011BDFC75AF6C7BA477DD25DA3128";
    attribute INIT_27 of inst : label is "410242190D212B0980F3FE92FFAABB14A9BAAEC52BA80D44A95D427402DCC9CD";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "DEFE85F6DFBDEEDFDBFFEFBF7E9F68724E29C196904C5CB9896BFB6E5220E815";
    attribute INIT_01 of inst : label is "82A1A86A1AC6B0AC2B0B957776E6E6E7FF7FE7FF7F3C64DE8514517051451CE7";
    attribute INIT_02 of inst : label is "AB8F1640017FFD7776E10DB5D75DD145ABFFE4B1E6898623BEDBC282A1A82A0A";
    attribute INIT_03 of inst : label is "0602BB1472024488002088ECE2388002A0F0F0F0F7FFFFFF6DBE29B050DA29B0";
    attribute INIT_04 of inst : label is "10508B6010505F47FA1F57FA1F57FBFF47FFA3EF03C3C3C15352B29910444110";
    attribute INIT_05 of inst : label is "CAAFFFD4FFEA7FF53FFFF57FCF4FF845E3FF57FFABFFD587FFFD4FF3CF4F4F4F";
    attribute INIT_06 of inst : label is "0011EC8157B2034BFFA1FFD0FF011EC8228F650697FF53FFA9FFD4FF411ECA0D";
    attribute INIT_07 of inst : label is "D75774115EC8FF3BE8189989989989852682E76CED05DED9D8024C200F659659";
    attribute INIT_08 of inst : label is "80005120D49999860D2666618349999860D2666618348CC090C16E8799D68698";
    attribute INIT_09 of inst : label is "1A1851C97575F24D49AD5D834760D1DB4769324D72D71ED90A62F74715DD1C56";
    attribute INIT_0A of inst : label is "1D835769324DFF0BC93526B4760D5D834769324D27834B429899F5ECEED7B3BB";
    attribute INIT_0B of inst : label is "D44DED41000D415D55B7F82CB2CBFFC0FF2BFC93526B5769324DFF0BF24D49AD";
    attribute INIT_0C of inst : label is "76FE2F9B8E8A5504AE3E8E9C84A43280C3AA21237FCF8E274E389929082E10FD";
    attribute INIT_0D of inst : label is "C889D091A4B56514B512B2949CC250159D8FC302101A4290EB292AD7608701A0";
    attribute INIT_0E of inst : label is "FFC2C22FFFF91C6E139FFFE00015554015555A79AC7E10747324749921D6354A";
    attribute INIT_0F of inst : label is "510025120D414B4FAABAFE80FF7F9F1C909BE7C724A023CA3925011C0E5BAB15";
    attribute INIT_10 of inst : label is "80005120D49999860D2666618349999860D2666618348CC090C16E8799D68698";
    attribute INIT_11 of inst : label is "1A1851C97575F24D49AD5D834760D1DB4769324D72D71ED90A62F74715DD1C56";
    attribute INIT_12 of inst : label is "1D835769324DFF0BC93526B4760D5D834769324D27834B429899F5ECEED7B3BB";
    attribute INIT_13 of inst : label is "D44DED41000D415D55B7F82CB2CBFFC0FF2BFC93526B5769324DFF0BF24D49AD";
    attribute INIT_14 of inst : label is "76FE2F9B8E8A5504AE3E8E9C84A43280C3AA21237FCF8E274E389929082E10FD";
    attribute INIT_15 of inst : label is "C889D091A4B56514B512B2949CC250159D8FC302101A4290EB292AD7608701A0";
    attribute INIT_16 of inst : label is "FFC2C22FFFF91C6E139FFFE00015554015555A79AC7E10747324749921D6354A";
    attribute INIT_17 of inst : label is "510025120D414B4FAABAFE80FF7F9F1C909BE7C724A023CA3925011C0E5BAB15";
    attribute INIT_18 of inst : label is "80005120D49999860D2666618349999860D2666618348CC090C16E8799D68698";
    attribute INIT_19 of inst : label is "1A1851C97575F24D49AD5D834760D1DB4769324D72D71ED90A62F74715DD1C56";
    attribute INIT_1A of inst : label is "1D835769324DFF0BC93526B4760D5D834769324D27834B429899F5ECEED7B3BB";
    attribute INIT_1B of inst : label is "D44DED41000D415D55B7F82CB2CBFFC0FF2BFC93526B5769324DFF0BF24D49AD";
    attribute INIT_1C of inst : label is "76FE2F9B8E8A5504AE3E8E9C84A43280C3AA21237FCF8E274E389929082E10FD";
    attribute INIT_1D of inst : label is "C889D091A4B56514B512B2949CC250159D8FC302101A4290EB292AD7608701A0";
    attribute INIT_1E of inst : label is "FFC2C22FFFF91C6E139FFFE00015554015555A79AC7E10747324749921D6354A";
    attribute INIT_1F of inst : label is "510025120D414B4FAABAFE80FF7F9F1C909BE7C724A023CA3925011C0E5BAB15";
    attribute INIT_20 of inst : label is "80005120D49999860D2666618349999860D2666618348CC090C16E8799D68698";
    attribute INIT_21 of inst : label is "1A1851C97575F24D49AD5D834760D1DB4769324D72D71ED90A62F74715DD1C56";
    attribute INIT_22 of inst : label is "1D835769324DFF0BC93526B4760D5D834769324D27834B429899F5ECEED7B3BB";
    attribute INIT_23 of inst : label is "D44DED41000D415D55B7F82CB2CBFFC0FF2BFC93526B5769324DFF0BF24D49AD";
    attribute INIT_24 of inst : label is "76FE2F9B8E8A5504AE3E8E9C84A43280C3AA21237FCF8E274E389929082E10FD";
    attribute INIT_25 of inst : label is "C889D091A4B56514B512B2949CC250159D8FC302101A4290EB292AD7608701A0";
    attribute INIT_26 of inst : label is "FFC2C22FFFF91C6E139FFFE00015554015555A79AC7E10747324749921D6354A";
    attribute INIT_27 of inst : label is "510025120D414B4FAABAFE80FF7F9F1C909BE7C724A023CA3925011C0E5BAB15";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "8B9465249256949212424924CC33C2AAC4AFD1D7B119DFABCB9AA85EFF30A815";
    attribute INIT_01 of inst : label is "6698A6298A6699A6699875DDDC4B4B5D55D55D54D509F4BE0000002C0000088C";
    attribute INIT_02 of inst : label is "E37F83F5434B2FDDDC584BBCF3CFD155A9A6DB6E0012C4C0A7FFC26299A6699A";
    attribute INIT_03 of inst : label is "0AA8B015513094AA80AA22C0EAA84D4A80B090B0932D92CBDF6BAB155588AB71";
    attribute INIT_04 of inst : label is "57322220D55553425A1752CA13425CCB46ECA3290252D24DCF4088CC55015555";
    attribute INIT_05 of inst : label is "C88832D4BB2A4CB52EDD9566490BF80108CB56ECAB32D583B7654992CB090B09";
    attribute INIT_06 of inst : label is "0254AC0542B01B6A65A17650990D0AC1AAA56036D4CB42ECA132D0BB4D0AC26D";
    attribute INIT_07 of inst : label is "D74570250AC0FF3BF01F99F99F99F9C517A08961264502C04E8A2F00CD659659";
    attribute INIT_08 of inst : label is "C0D94D66D4888A66EEE22299BBB888A66EEE22299BBBC2E00008DAA14B6F5BC5";
    attribute INIT_09 of inst : label is "9CCE36D97855F48D91ADCD837360D8DB63723C8D69EC31408080F66F5119BD45";
    attribute INIT_0A of inst : label is "8D8373723C8DFF42D33666B7360D8D8363733CCD198AD9602000FBD4566F5159";
    attribute INIT_0B of inst : label is "F344A58D046D4D5F3115FC2CB2CBFFC0FF62FD33666B63733CCDFF62F48D91AD";
    attribute INIT_0C of inst : label is "56FF2C8ED1DADD9DAF58AEA70BA0CEC2CC6E18235CD5BC2B46F0AA2A4C23055D";
    attribute INIT_0D of inst : label is "DCABD4BBADBB2BCD759695AD4062B8F9BD03D402F8FA57BAE95ACEF75552ABA1";
    attribute INIT_0E of inst : label is "FFC6D988FFDB145FEB5FFFE00019999559999ED05D0E077EFB2EF5D97DD3B9EC";
    attribute INIT_0F of inst : label is "8D0D94D46D4D4BCDE634FF0DFF39AB78A01AEA5E2BA444F8F15D223013528A0D";
    attribute INIT_10 of inst : label is "C0D94D66D4888A66EEE22299BBB888A66EEE22299BBBC2E00008DAA14B6F5BC5";
    attribute INIT_11 of inst : label is "9CCE36D97855F48D91ADCD837360D8DB63723C8D69EC31408080F66F5119BD45";
    attribute INIT_12 of inst : label is "8D8373723C8DFF42D33666B7360D8D8363733CCD198AD9602000FBD4566F5159";
    attribute INIT_13 of inst : label is "F344A58D046D4D5F3115FC2CB2CBFFC0FF62FD33666B63733CCDFF62F48D91AD";
    attribute INIT_14 of inst : label is "56FF2C8ED1DADD9DAF58AEA70BA0CEC2CC6E18235CD5BC2B46F0AA2A4C23055D";
    attribute INIT_15 of inst : label is "DCABD4BBADBB2BCD759695AD4062B8F9BD03D402F8FA57BAE95ACEF75552ABA1";
    attribute INIT_16 of inst : label is "FFC6D988FFDB145FEB5FFFE00019999559999ED05D0E077EFB2EF5D97DD3B9EC";
    attribute INIT_17 of inst : label is "8D0D94D46D4D4BCDE634FF0DFF39AB78A01AEA5E2BA444F8F15D223013528A0D";
    attribute INIT_18 of inst : label is "C0D94D66D4888A66EEE22299BBB888A66EEE22299BBBC2E00008DAA14B6F5BC5";
    attribute INIT_19 of inst : label is "9CCE36D97855F48D91ADCD837360D8DB63723C8D69EC31408080F66F5119BD45";
    attribute INIT_1A of inst : label is "8D8373723C8DFF42D33666B7360D8D8363733CCD198AD9602000FBD4566F5159";
    attribute INIT_1B of inst : label is "F344A58D046D4D5F3115FC2CB2CBFFC0FF62FD33666B63733CCDFF62F48D91AD";
    attribute INIT_1C of inst : label is "56FF2C8ED1DADD9DAF58AEA70BA0CEC2CC6E18235CD5BC2B46F0AA2A4C23055D";
    attribute INIT_1D of inst : label is "DCABD4BBADBB2BCD759695AD4062B8F9BD03D402F8FA57BAE95ACEF75552ABA1";
    attribute INIT_1E of inst : label is "FFC6D988FFDB145FEB5FFFE00019999559999ED05D0E077EFB2EF5D97DD3B9EC";
    attribute INIT_1F of inst : label is "8D0D94D46D4D4BCDE634FF0DFF39AB78A01AEA5E2BA444F8F15D223013528A0D";
    attribute INIT_20 of inst : label is "C0D94D66D4888A66EEE22299BBB888A66EEE22299BBBC2E00008DAA14B6F5BC5";
    attribute INIT_21 of inst : label is "9CCE36D97855F48D91ADCD837360D8DB63723C8D69EC31408080F66F5119BD45";
    attribute INIT_22 of inst : label is "8D8373723C8DFF42D33666B7360D8D8363733CCD198AD9602000FBD4566F5159";
    attribute INIT_23 of inst : label is "F344A58D046D4D5F3115FC2CB2CBFFC0FF62FD33666B63733CCDFF62F48D91AD";
    attribute INIT_24 of inst : label is "56FF2C8ED1DADD9DAF58AEA70BA0CEC2CC6E18235CD5BC2B46F0AA2A4C23055D";
    attribute INIT_25 of inst : label is "DCABD4BBADBB2BCD759695AD4062B8F9BD03D402F8FA57BAE95ACEF75552ABA1";
    attribute INIT_26 of inst : label is "FFC6D988FFDB145FEB5FFFE00019999559999ED05D0E077EFB2EF5D97DD3B9EC";
    attribute INIT_27 of inst : label is "8D0D94D46D4D4BCDE634FF0DFF39AB78A01AEA5E2BA444F8F15D223013528A0D";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "949890000108400000000003449188234231001C906C496D8D96A89635AB2130";
    attribute INIT_01 of inst : label is "84701C060180701C0600B35556A4A4B55A55A55A5554EB9ED861865186187024";
    attribute INIT_02 of inst : label is "43A271198534995556A282E49249C91C834D34D2A25B36A0E249D980601C4711";
    attribute INIT_03 of inst : label is "1194C41D84CB12464919D110E6433189B2E2C2C2EC9B6D264DA4844232211924";
    attribute INIT_04 of inst : label is "A10B362FC707081B30DC0BB0DC0BA3340F1207840B1B1BBC059B73388C36308C";
    attribute INIT_05 of inst : label is "ECD8CD06C4836261B9B360F9AE2EFC8B0F341F120F8987866CD82E6BAE2C2C2E";
    attribute INIT_06 of inst : label is "2446A41C1A90D9219A0D8906C42C2A45983521B243341B120D8986E66C2A4364";
    attribute INIT_07 of inst : label is "F26D06C46A43FFC4E469669669669616C84B2D95B1925B2B6325919370924924";
    attribute INIT_08 of inst : label is "B06D2CB643AAA889332AAA324CEAAA889332AAA324CE1F600800A7118762888A";
    attribute INIT_09 of inst : label is "BAFA8F9726D0FB706E102A040A8102A40A8DC370D7C202608000F02208808822";
    attribute INIT_0A of inst : label is "2A041A8CC330FFB6EDC1B840A8102A040A8DC37062247AE00020F88220220880";
    attribute INIT_0B of inst : label is "DB32106C9B642CC88B10F9924924FFE0FFB6FECC19841A8CC330FF96FB306610";
    attribute INIT_0C of inst : label is "D2FEE49A868E664664180E0C66825A10C1A1B39936460C8308320A25A18C4874";
    attribute INIT_0D of inst : label is "4E08CA18C013836C7260418C403608528C71D80648592398E418B34B2AA20D86";
    attribute INIT_0E of inst : label is "FFCBECD8FFD6A7205E1FFFE0001E1E199E1E10E3DCDC0A763386329C32C853C9";
    attribute INIT_0F of inst : label is "6C06D2CB642C2C731171FE60FFEC8C18084923860690534A3034829006C66894";
    attribute INIT_10 of inst : label is "B06D2CB643AAA889332AAA324CEAAA889332AAA324CE1F600800A7118762888A";
    attribute INIT_11 of inst : label is "BAFA8F9726D0FB706E102A040A8102A40A8DC370D7C202608000F02208808822";
    attribute INIT_12 of inst : label is "2A041A8CC330FFB6EDC1B840A8102A040A8DC37062247AE00020F88220220880";
    attribute INIT_13 of inst : label is "DB32106C9B642CC88B10F9924924FFE0FFB6FECC19841A8CC330FF96FB306610";
    attribute INIT_14 of inst : label is "D2FEE49A868E664664180E0C66825A10C1A1B39936460C8308320A25A18C4874";
    attribute INIT_15 of inst : label is "4E08CA18C013836C7260418C403608528C71D80648592398E418B34B2AA20D86";
    attribute INIT_16 of inst : label is "FFCBECD8FFD6A7205E1FFFE0001E1E199E1E10E3DCDC0A763386329C32C853C9";
    attribute INIT_17 of inst : label is "6C06D2CB642C2C731171FE60FFEC8C18084923860690534A3034829006C66894";
    attribute INIT_18 of inst : label is "B06D2CB643AAA889332AAA324CEAAA889332AAA324CE1F600800A7118762888A";
    attribute INIT_19 of inst : label is "BAFA8F9726D0FB706E102A040A8102A40A8DC370D7C202608000F02208808822";
    attribute INIT_1A of inst : label is "2A041A8CC330FFB6EDC1B840A8102A040A8DC37062247AE00020F88220220880";
    attribute INIT_1B of inst : label is "DB32106C9B642CC88B10F9924924FFE0FFB6FECC19841A8CC330FF96FB306610";
    attribute INIT_1C of inst : label is "D2FEE49A868E664664180E0C66825A10C1A1B39936460C8308320A25A18C4874";
    attribute INIT_1D of inst : label is "4E08CA18C013836C7260418C403608528C71D80648592398E418B34B2AA20D86";
    attribute INIT_1E of inst : label is "FFCBECD8FFD6A7205E1FFFE0001E1E199E1E10E3DCDC0A763386329C32C853C9";
    attribute INIT_1F of inst : label is "6C06D2CB642C2C731171FE60FFEC8C18084923860690534A3034829006C66894";
    attribute INIT_20 of inst : label is "B06D2CB643AAA889332AAA324CEAAA889332AAA324CE1F600800A7118762888A";
    attribute INIT_21 of inst : label is "BAFA8F9726D0FB706E102A040A8102A40A8DC370D7C202608000F02208808822";
    attribute INIT_22 of inst : label is "2A041A8CC330FFB6EDC1B840A8102A040A8DC37062247AE00020F88220220880";
    attribute INIT_23 of inst : label is "DB32106C9B642CC88B10F9924924FFE0FFB6FECC19841A8CC330FF96FB306610";
    attribute INIT_24 of inst : label is "D2FEE49A868E664664180E0C66825A10C1A1B39936460C8308320A25A18C4874";
    attribute INIT_25 of inst : label is "4E08CA18C013836C7260418C403608528C71D80648592398E418B34B2AA20D86";
    attribute INIT_26 of inst : label is "FFCBECD8FFD6A7205E1FFFE0001E1E199E1E10E3DCDC0A763386329C32C853C9";
    attribute INIT_27 of inst : label is "6C06D2CB642C2C731171FE60FFEC8C18084923860690534A3034829006C66894";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "128840000080200000000001401080210018000800208BE000CEA84A0AB90120";
    attribute INIT_01 of inst : label is "405110451100501005003600029494800800800900523F8E4820824082083094";
    attribute INIT_02 of inst : label is "B21BF63E06000A00028213420820D8080192D92EA2C91220E000C90441140401";
    attribute INIT_03 of inst : label is "181CE019C00B82E04B81F380ECE001C196A686868A412002A000004300218100";
    attribute INIT_04 of inst : label is "3A0B36268606041A80D01A00D01A04001E000F000A0A0A2842CB93C8C07701C0";
    attribute INIT_05 of inst : label is "ECD8000680034021A89121E8AA6AFD9B0C000E000700838224482A2AAA282828";
    attribute INIT_06 of inst : label is "6E0684381A10F000000D000680386847101420A000000A00050082A228284140";
    attribute INIT_07 of inst : label is "E26C06E06843FF80EC004004004004330059A504A1B34A094166009320000000";
    attribute INIT_08 of inst : label is "B06D28B403222050028888040082220100208881400A81C00000C1B208D57575";
    attribute INIT_09 of inst : label is "1183120626C0FB20640068001A0006801A0C8B20109F04C00000FDD5F77757DD";
    attribute INIT_0A of inst : label is "28001A0D8B60FFB6EC819001A00068001A0C8B20A0C780C00000F57DDDD5F777";
    attribute INIT_0B of inst : label is "DA2000689B4028899B00F9000000FFE0FF96FED81B000A0D8B60FF96FB606C00";
    attribute INIT_0C of inst : label is "C2FEC400428E33A6C118080453014C30800352440105140404501001D1544450";
    attribute INIT_0D of inst : label is "8E090E1944968678C2324318C01458071071C004180133188431999C00321E00";
    attribute INIT_0E of inst : label is "FFCBECD8FFF99A04995FFFE0001FE01E1FE0030328650E5652864394330863C9";
    attribute INIT_0F of inst : label is "6806D28B402828213371FE50FFA008281020020A0308081A5018425002865088";
    attribute INIT_10 of inst : label is "B06D28B403222050028888040082220100208881400A81C00000C1B208D57575";
    attribute INIT_11 of inst : label is "1183120626C0FB20640068001A0006801A0C8B20109F04C00000FDD5F77757DD";
    attribute INIT_12 of inst : label is "28001A0D8B60FFB6EC819001A00068001A0C8B20A0C780C00000F57DDDD5F777";
    attribute INIT_13 of inst : label is "DA2000689B4028899B00F9000000FFE0FF96FED81B000A0D8B60FF96FB606C00";
    attribute INIT_14 of inst : label is "C2FEC400428E33A6C118080453014C30800352440105140404501001D1544450";
    attribute INIT_15 of inst : label is "8E090E1944968678C2324318C01458071071C004180133188431999C00321E00";
    attribute INIT_16 of inst : label is "FFCBECD8FFF99A04995FFFE0001FE01E1FE0030328650E5652864394330863C9";
    attribute INIT_17 of inst : label is "6806D28B402828213371FE50FFA008281020020A0308081A5018425002865088";
    attribute INIT_18 of inst : label is "B06D28B403222050028888040082220100208881400A81C00000C1B208D57575";
    attribute INIT_19 of inst : label is "1183120626C0FB20640068001A0006801A0C8B20109F04C00000FDD5F77757DD";
    attribute INIT_1A of inst : label is "28001A0D8B60FFB6EC819001A00068001A0C8B20A0C780C00000F57DDDD5F777";
    attribute INIT_1B of inst : label is "DA2000689B4028899B00F9000000FFE0FF96FED81B000A0D8B60FF96FB606C00";
    attribute INIT_1C of inst : label is "C2FEC400428E33A6C118080453014C30800352440105140404501001D1544450";
    attribute INIT_1D of inst : label is "8E090E1944968678C2324318C01458071071C004180133188431999C00321E00";
    attribute INIT_1E of inst : label is "FFCBECD8FFF99A04995FFFE0001FE01E1FE0030328650E5652864394330863C9";
    attribute INIT_1F of inst : label is "6806D28B402828213371FE50FFA008281020020A0308081A5018425002865088";
    attribute INIT_20 of inst : label is "B06D28B403222050028888040082220100208881400A81C00000C1B208D57575";
    attribute INIT_21 of inst : label is "1183120626C0FB20640068001A0006801A0C8B20109F04C00000FDD5F77757DD";
    attribute INIT_22 of inst : label is "28001A0D8B60FFB6EC819001A00068001A0C8B20A0C780C00000F57DDDD5F777";
    attribute INIT_23 of inst : label is "DA2000689B4028899B00F9000000FFE0FF96FED81B000A0D8B60FF96FB606C00";
    attribute INIT_24 of inst : label is "C2FEC400428E33A6C118080453014C30800352440105140404501001D1544450";
    attribute INIT_25 of inst : label is "8E090E1944968678C2324318C01458071071C004180133188431999C00321E00";
    attribute INIT_26 of inst : label is "FFCBECD8FFF99A04995FFFE0001FE01E1FE0030328650E5652864394330863C9";
    attribute INIT_27 of inst : label is "6806D28B402828213371FE50FFA008281020020A0308081A5018425002865088";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
