-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "001503FFA80000005400FCC0082B0000001503FFA80000005400FCC000000000";
    attribute INIT_01 of inst : label is "019906D1B940000047201364002900000090003C1C00000000404D10012B0000";
    attribute INIT_02 of inst : label is "FD000000FD000000000000000B7E000024D402676DC0002014600E8106B20000";
    attribute INIT_03 of inst : label is "FFFFFFFF0BFF000BFFE0E000000300000000003FFE0000000000FFE0FD00FFFD";
    attribute INIT_04 of inst : label is "00000BFFC00000000000FC00003F0000000003FFF00000000000FF0000000000";
    attribute INIT_05 of inst : label is "4FF1FFFF4FF0FFF000040FFC00BD00200A803C2A7E00080002A0A83C00BF0000";
    attribute INIT_06 of inst : label is "03C0F57CF03C15E0F028157C7D543F80F0287D5005F8B5780F000F8070B42D60";
    attribute INIT_07 of inst : label is "FFFFFF00FFFF00FF0FF10FFF000003C015540000014000007800B578F50C2578";
    attribute INIT_08 of inst : label is "F0B455E0003C557C00F055F0783C2D7CA0B4B5E0F03CB57CF57C2DE0D743B55E";
    attribute INIT_09 of inst : label is "F03CB578FD3CF0BCF13CF8BC00F000F02F7C783CF828F0000F005F50F03CF03C";
    attribute INIT_0A of inst : label is "7DF4F03C1FD0F03CF03CF03C0F005F50F0282D782F7CB57C07D00000157CB57C";
    attribute INIT_0B of inst : label is "000000000000000001E000B0FFFEEEEE0B400E0001F8FD540F00F0F0BDF8F8BC";
    attribute INIT_0C of inst : label is "00EF0000000000B7E80000005780BD50FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "02400000001E030600000000AA8000200009000001BA0E7A00000000D8008D00";
    attribute INIT_0E of inst : label is "001F1FFF7FFF7FFF02FF0002FFFFFFFFFF808000F400FFF4FFFFEEEEFFFFEEEE";
    attribute INIT_0F of inst : label is "FFFEFFFEBFFEBFFE7FFF6EEE0BFD00097FFF7FFFFFFFFFFF7FFE7FFEFFFEFFFE";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFF0000FFFF000000000000C0030000C00025587FFD96960000A800";
    attribute INIT_11 of inst : label is "007F7FFF007F0000007F0000000000003FFF2AAA3FFF3FFFFFFCAAA8FFFCFFFC";
    attribute INIT_12 of inst : label is "FFFF0AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFF0FFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFF3FFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFA0FFFFFFFF";
    attribute INIT_14 of inst : label is "FFFCFFFCFFFFFFFF3FFF2AAA3FFF3FFFFFFFBFFFFFFFFFFFFFFFAAAAFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFBFFEFFFFFFFF3FFC3FFC3FFF3FFFFFFFFFFFFFFFFFFEFFFCFFFCFFFCAAA8";
    attribute INIT_16 of inst : label is "0FFF00A3000700FFFFF0CA00D000FF00003F000B03FF0A7FFC00E000FFC0FDA0";
    attribute INIT_17 of inst : label is "3FFB000005FC5FFFFA0000000000FFDD00AF0000000077FFEFFC00003F50FFF5";
    attribute INIT_18 of inst : label is "3FFF2AAA3FFF3FFFFFFCAAA8FFFCFFFC3FFF2AAA3FFF3FFFFFFCAAA8FFFCFFFC";
    attribute INIT_19 of inst : label is "3FD52AAA3FFF3FCCD5FCAAA8FFFCCDFC3FFF2AAA3FFF3FFFFFFCAAA8FFFCFFFC";
    attribute INIT_1A of inst : label is "CFD7D555C0FFC0FF77F35557FF03FF03FE00FC0000BF003FF3FFFFD5FFCF57FF";
    attribute INIT_1B of inst : label is "C000D555C150EFFD0E03555705432FF3C000D555CFFFCBEF00035557FFB3FBE3";
    attribute INIT_1C of inst : label is "CE6ED555C000C3666C03555700FB6503C000D555C555CFF4000355575553FF83";
    attribute INIT_1D of inst : label is "C2FFD555C7F4CFFFFFF355570063F403C0AAD555C550CF5F800355570003FA03";
    attribute INIT_1E of inst : label is "FCFFFCFF03C057FF3F3FFFFFFCFCFFFF03C0FFD5FAAFFFFF0BFF000B00000FFF";
    attribute INIT_1F of inst : label is "0000FFFFFFFFFFFFF400FFF4BFFFBBBBFFFFBBBBFFFDBBB900005555FF3FFF3F";
    attribute INIT_20 of inst : label is "000003FF0550002A0000FFC00550A80000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "003F0BFF05550000FC00FFE055500000003F0BFF05500000FC00FFE005500000";
    attribute INIT_22 of inst : label is "007F01FF05540000FD00FF401550000000BF0FFF05550000FE00FFF055500000";
    attribute INIT_23 of inst : label is "07FF02FF01FC003FFFD0FF803F40FC000FBF00FF0154002AFEF0FF001540A800";
    attribute INIT_24 of inst : label is "0A90807FF3F5003F4FDDFF007FF4FC00004103FF055000FF3F80ABC0FF3CF000";
    attribute INIT_25 of inst : label is "3F9A00FF0055003FA6F4FFE01BF0FC00038403FF0AA0003F12FCFA901540FC00";
    attribute INIT_26 of inst : label is "2BFF00FF0055003FFFF8FFE03FD0FC002BFF0BFF0BFC003FFFE0FD341540FC00";
    attribute INIT_27 of inst : label is "F3E1E0FF53FF000301B8FFFCF810FFC02FFF05FF0154003FFFF8FF501540FC00";
    attribute INIT_28 of inst : label is "0BC409FF0105000013E0FF60504000003FD0FF833FFF00000000F028F02FFFF0";
    attribute INIT_29 of inst : label is "0A5A0C87007A0000FE80FFF06FD000000D980FD700BF0000D7B0FFD0D0000000";
    attribute INIT_2A of inst : label is "0000000A000000000800000000000000000000BC0000000000003E0000000000";
    attribute INIT_2B of inst : label is "3FD0FF833FFF00000000FAA8F02F00000000000000000000B000A00000000000";
    attribute INIT_2C of inst : label is "3FFF3FFF00002AAAFFFCFFFC0000AAA83FFF3FFF15552AAAFFFCFFFC5554AAA8";
    attribute INIT_2D of inst : label is "3FFF000000002AAAFFFC00000000AAA83FFF155500002AAAFFFC55540000AAA8";
    attribute INIT_2E of inst : label is "0000000000002AAA000000000000AAA81555000000002AAA555400000000AAA8";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "00AF0FBF00FF0002FA00FEF0FF008000003F0A7F03FF000BFC00FDA0FFC0E000";
    attribute INIT_31 of inst : label is "0FFE1FFF007F0000FC00FF74300000003FFB5FFF05FC0000FA00FFDD00000000";
    attribute INIT_32 of inst : label is "03000000000002FD00C0000000007F80023F00FF003F000BFC80FF00FC00E000";
    attribute INIT_33 of inst : label is "0000000000000000007F000B05540000EAFFFFFF00000000FA00FFDD14000000";
    attribute INIT_34 of inst : label is "2FFF3FFF0FFD0AAEE3C0FFE05FD0A800FB0F0FFF2DFF0FEFFA70FFF8FD5EFA00";
    attribute INIT_35 of inst : label is "07F3FFFF1FDFFEAFF3F8FFD7FFF4FA2F2FFF3FFF2D5F0ABFA9C05FE8FFDEE800";
    attribute INIT_36 of inst : label is "0BFF0FFF2DFF0FEFFFF05FF8FD5EFA002FCFD7FF1FFF28AFCFD0FFFFF7F4FA28";
    attribute INIT_37 of inst : label is "2FFF5FFF2D5F0ABFFFC0FFE0FFDEE8002FFF35FF0FFD0ABFFFC0FFE05FD0E800";
    attribute INIT_38 of inst : label is "2FF75FFF1FDF28AFF7F8FD7FFFF4FA282FDFFD7F1FFFF8AFDFF8FFF5F7F4FA2F";
    attribute INIT_39 of inst : label is "0BFF05573FFE0ABF8000FE00FFF8FEA00004017F0555000F13C0FFFFFFCFFF00";
    attribute INIT_3A of inst : label is "0C330C33014100000CD00CC050400000AFFF0057BFFF0ABF0000FE00FFF8FEA0";
    attribute INIT_3B of inst : label is "007F001F0B80BD30FD00F40002E00C7EE0FE00AA00010030BF0BAA0040000C00";
    attribute INIT_3C of inst : label is "000008F0800000000000FC0840307000F8FE001F5E000024BF2FF40000B50C00";
    attribute INIT_3D of inst : label is "30000001000000000004FE80000028002800003F800000000000FF0000347000";
    attribute INIT_3E of inst : label is "00140005000000000000403000401C0000000002000000000000FE0004000700";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000002A2033300000000A2A0333000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "000001FFFF8000000000FB4002FF025E000001FFFF8000000000FB4000000000";
    attribute INIT_01 of inst : label is "000000FCF2C002E00000FE0000C600100000002FE680090000003A0002FF045E";
    attribute INIT_02 of inst : label is "D000FFD0D0000000D000000000D4008A000003F7041000300400FB40025C06A8";
    attribute INIT_03 of inst : label is "FFFFFFFFBFFF00BFFFFEFE00000F0000000000FFFF80A0000000FFF0D000FFD0";
    attribute INIT_04 of inst : label is "00000FFFF00000000000FF0000FF000A00000FFFFC0080000000FFC000000000";
    attribute INIT_05 of inst : label is "FFFF8FF2FFF08FF00BBF177D205F003811500007F5082C000544D00002FF000A";
    attribute INIT_06 of inst : label is "01401E0015502ABC1550B55414003C7815502F8055547E8055500F000540F03C";
    attribute INIT_07 of inst : label is "FFFFFF00FFFF00FF0FFF0FF20000006000002AA8000002800550FAB415501AF4";
    attribute INIT_08 of inst : label is "5540A83C00142ABC55502AF00554F03C1540003C15547ABC5014F03C7AADEB83";
    attribute INIT_09 of inst : label is "1550F03C5014FBFC5014FFFC555000F0541407BC1550F00055500F005014FABC";
    attribute INIT_0A of inst : label is "1010FBBC0100F8BC1550F03C05000F0015502AB45414F83C00000BE00014F03C";
    attribute INIT_0B of inst : label is "000000000000000000100B40FFFEFFFE040001E055541F8005003AC050141FD0";
    attribute INIT_0C of inst : label is "03B700170000005FE78050000000DD00FFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0D of inst : label is "022002A8000001E0000000000000554002DD017A00000D669000AA0000005980";
    attribute INIT_0E of inst : label is "000101FF7FFF7FFF2FFF002F7777FFFFFFF8F8004000FF40FFFFFFFF7777FFFF";
    attribute INIT_0F of inst : label is "7776FFFEBFFEBFFE77777FFFBFFD00BD77777FFFFFFFFFFF77767FFEFFFEFFFE";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFF0000FFFF00001554BAAE160490030140C00300005400";
    attribute INIT_11 of inst : label is "000707FF000707FF00070000000700003FFF3FFF15553FFFFFFCFFFC5554FFFC";
    attribute INIT_12 of inst : label is "FFFFFFFF05FFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFCFFFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFF0FFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF50FFFF";
    attribute INIT_14 of inst : label is "FFFCFFFC7FFFFFFF3FFF3FFF3FFF3FFFFFFFFFFF5555FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFF7FFDFFFF3FFC3FFC15553FFFFFFDFFFFFFFFFFFF5554FFFCFFFCFFFC";
    attribute INIT_16 of inst : label is "05BF03FF0007003FFE50FFC0D000FC0000FF000B00530FFFFF00E000C500FFF0";
    attribute INIT_17 of inst : label is "AFFF0AFC00003FF7FFEE00000000F500BBFF00000000005FFFFA3FA00000DFFC";
    attribute INIT_18 of inst : label is "3FFF3FFF15553FFFFFFCFFFC5554FFFC3FFF3FFF15553FFFFFFCFFFC5554FFFC";
    attribute INIT_19 of inst : label is "3FCC3FFF15553FEAD4FCFFFC5554EAFC3FFF3FFF15553FFFFFFCFFFC5554FFFC";
    attribute INIT_1A of inst : label is "C5D6CBFEEAAAC0FF9B53BFE3AAABFF03FFEAFC00ABFF003FF3FFF4AFCFCFFA1F";
    attribute INIT_1B of inst : label is "C2AAC000EAAAFFFF0FA3AF03AAABFDD7C08AC000EAAACFFFA2030003AAABFFF3";
    attribute INIT_1C of inst : label is "CE67C277EAAAC05E6703A003AABFC603CBFEC000EAAACFCB80030003AAABFF43";
    attribute INIT_1D of inst : label is "C3FFC02AEAAACFFFFF43FFE3AAAF4003CBFFC000EAAACFB5F8030003AAAB7F03";
    attribute INIT_1E of inst : label is "FC55FCFF03EA03D5BF3F7F2AFCFEA8FDABC057C0FFFFFFFFBFFF00BF00000000";
    attribute INIT_1F of inst : label is "00000000FFFFFFFF4000FF409DDDBFFFDDDDFFFFDDDDFFFD00000000553FFF3F";
    attribute INIT_20 of inst : label is "00BF0FFF2FC000BFFE00FFF003F8FE0000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "02FF0FFF2FC00000FF80FFF003F8000002FF0FFF2FC00000FF80FFF003F80000";
    attribute INIT_22 of inst : label is "0FFF02FF2FF0003FFFF0FF800FF8FC0000BF0AFF2FC0002AFE00FFA003F8A800";
    attribute INIT_23 of inst : label is "00FF03F803F40F7FFF002FC03FC0FDF005FF03FF2FF000BFFF50FFC00FF8FE00";
    attribute INIT_24 of inst : label is "0FFEF3FF00000077BF40FFFC0150DDAA007A0BFFBFC001DF5FF0FFC0153C7400";
    attribute INIT_25 of inst : label is "01FA03FF00BF0A7DAFC0FFF0C1407DF82FFB0FFF15500A5DE5FCFFF0FF8075A0";
    attribute INIT_26 of inst : label is "1DFF03FF00BF007FFFFC7FF0C500FD003FFF07FF0FD0007FFFFCFE80FF80FD00";
    attribute INIT_27 of inst : label is "53FAF3FF0000E007AFFCF5FC0000DF703FFF03FF0BFC007FFFFCFFC03FE0FD00";
    attribute INIT_28 of inst : label is "0C3B0F3F00000035EC30FCF000005C0000027FFF0FFF0001A000F08FFC5D5554";
    attribute INIT_29 of inst : label is "0C4B05A5000000B5FFF0FD4000009FE0001B07EB000002D0EBF0FF000000FE00";
    attribute INIT_2A of inst : label is "00000015000000003C0000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "00027FFF0FFF0000A000FFFEFC5D000000000000000000005000700000000000";
    attribute INIT_2C of inst : label is "3FFF155500003FFFFFFC55540000FFFC3FFF3FFF00003FFFFFFCFFFC0000FFFC";
    attribute INIT_2D of inst : label is "1555000000003FFF555400000000FFFC3FFF000000003FFFFFFC00000000FFFC";
    attribute INIT_2E of inst : label is "000000000000155500000000000055540000000000003FFF000000000000FFFC";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "05FF07FF00010007FF50FFD04000D00000FF0FFF0053000BFF00FFF0C500E000";
    attribute INIT_31 of inst : label is "2FFF0FFD000000BFFFB8FC0000003000AFFF3FF700000AFCFFEEF50000000000";
    attribute INIT_32 of inst : label is "00000000000003D000000000000007C001FF00FF00BF000BFF40FF00FE00E000";
    attribute INIT_33 of inst : label is "0000000000000000000700BF00000AA8FFFFD5FF00000000FFEEF50000002800";
    attribute INIT_34 of inst : label is "3FF01FFF07BE07FFFBC0FFFCAD00DF007FFF07FF1EAD01FFFFB0FFFF1EADD7C0";
    attribute INIT_35 of inst : label is "ABFD7FFF0FC03FE77FFEFFE90150DBF43FFF1FFF1EAD07FFFEC0AFFD1EADDF00";
    attribute INIT_36 of inst : label is "0FFF07FF1EAD01FFFEF0AFFF1EADFFC0BFFD6BFF0540FFE77FEAFFFD03F0DBFF";
    attribute INIT_37 of inst : label is "BFFF0FFF1EAD07FFFBC0FFFC1EADFF003FFF1AFF07BE07FFFCC0FFFCAD00FF00";
    attribute INIT_38 of inst : label is "BFFD2FFF0FC0FFFF7FFEFEBD0150FFFFBFFD7EBF05401FFF7FFEFFF803F0FFF4";
    attribute INIT_39 of inst : label is "3FFF0BE3FFFF02FFFE00FFE0FFF4440003EE0BFF2FF0001DAFF8FFFD3D6DF740";
    attribute INIT_3A of inst : label is "0C330C33000002800CC00CC00000A0801FFF0BEA7FFF02FFFE00BFE0FFF44400";
    attribute INIT_3B of inst : label is "0005000105E050BD500040000B507E057C05001F9FA0003E103DF4000AF6BC00";
    attribute INIT_3C of inst : label is "000001471A0000000000F430004001200005B8070000203E1000D02E0000BC08";
    attribute INIT_3D of inst : label is "50020000002A0000000001C0A4000480502F00047A0000008000000800400120";
    attribute INIT_3E of inst : label is "000B00000000000AFA0000D000000048016A0000000A000000005F00A9000012";
    attribute INIT_3F of inst : label is "00000000000000000000000000000000033301510000000033B0515000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "3FEA3C0057FCAAA8ABFC033C3FD42AAA3FEA3C0057FCAAA8ABFC033C00000000";
    attribute INIT_01 of inst : label is "04D403240E000020035020700026000004940093B10000000440F1183FD42AAA";
    attribute INIT_02 of inst : label is "FD000000FD0000000000000000A1600233790050AA10400AE9806E89076D0000";
    attribute INIT_03 of inst : label is "FFFFFFFF0BFF000BFFE0E00000000002029000002000000000000000FD00FFFD";
    attribute INIT_04 of inst : label is "0000000000008000068000000002000200060000000000008000000000000000";
    attribute INIT_05 of inst : label is "F00F0000F00000001FF805543FFB0002057F03FFEFFC8000FD50FFC000080000";
    attribute INIT_06 of inst : label is "03C0F57CF03C15E0F028157C7D543F80F0287D5005F8B5780F000F8070B42D60";
    attribute INIT_07 of inst : label is "FFFFFFFFFFFFFFFF000F0000000003C015540000014000007800B578F50C2578";
    attribute INIT_08 of inst : label is "F0B455E0003C557C00F055F0783C2D7CA0B4B5E0F03CB57CF57C2DE0D743B55E";
    attribute INIT_09 of inst : label is "F03CB578FD3CF0BCF13CF8BC00F000F02F7C783CF828F0000F005F50F03CF03C";
    attribute INIT_0A of inst : label is "7DF4F03C1FD0F03CF03CF03C0F005F50F0282D782F7CB57CF82FFFFF157CB57C";
    attribute INIT_0B of inst : label is "FFF0FFF00FFF0FFF01E000B0FFFFFFFF0B400E0001F8FD540F00F0F0BDF8F8BC";
    attribute INIT_0C of inst : label is "00EE0000000000BFFA00000057C0FF50FD05FFFFFFA0F0C0487FFFFF0AFF000F";
    attribute INIT_0D of inst : label is "00B80000001F03FF00000000FF00FFC0000000000045018500000000250072C0";
    attribute INIT_0E of inst : label is "007F7FFFFFFFFFFF0BFF000BFFFFFFFFFFE0E000FD00FFFDFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF2FFF002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFF0000FFFF00000000000000000BE0C02E255842819696F7E0A800";
    attribute INIT_11 of inst : label is "007F7FFF007F0000007F00000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000F5000000000000000000000000000000F000000000000000000F00000000";
    attribute INIT_13 of inst : label is "00000000C0000000000000000003000000000000000000000000005F00000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000255800380000300025582C000000000000000006000C0000000000000000";
    attribute INIT_17 of inst : label is "C0002400C000200000A00000000000200A00000000000800000300080003AA98";
    attribute INIT_18 of inst : label is "02A2000000000333A2A000000000206002A2000000000333A2A0000000003320";
    attribute INIT_19 of inst : label is "002A0000000000332A0000000000320002A2000000000333A200000000003300";
    attribute INIT_1A of inst : label is "0FFF0000005500FFFFF000005500FF00F1FFF3FFFF4FFFCF0FFF002AFFF0A800";
    attribute INIT_1B of inst : label is "0000000006A42FFD0F4000001A902FE0003000000FFF0BEF0C000000FEB0FBE0";
    attribute INIT_1C of inst : label is "0C0A0000000003000C00000000F801000AA0000000000FFF000000000000AA80";
    attribute INIT_1D of inst : label is "02FA000007C00FFF7F5000000060400000AA000005550CAF8000000055503F00";
    attribute INIT_1E of inst : label is "CFFFFFFF0F000AAA0FF0AAAA0FF0AAAA00F0AAA00FF00000000003F403FC0FFF";
    attribute INIT_1F of inst : label is "00000000FFFF0000F400FFF4BFFFBBBBFFFFBBBBFFFDBBB900005555FFF3FFFF";
    attribute INIT_20 of inst : label is "000000000FD0002A0000000007F0A80000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "001520000FD500005400000857F000000015000017F000005400000007F40000";
    attribute INIT_22 of inst : label is "28D5000007F40000572800001FD0000000AA00000FD50000AA00000057F00000";
    attribute INIT_23 of inst : label is "000002FF010028150000FF8000405428004000AA03F4002A0100AA001FC0A800";
    attribute INIT_24 of inst : label is "0E6F002A0FF50015B00FAA007D40540001BE3F000FD00055C0005500FFC05000";
    attribute INIT_25 of inst : label is "286F00FF007F0015F93CFFE0140054003C7B02AA01540015ED00AFD0BD405400";
    attribute INIT_26 of inst : label is "00003CAA007F00150000AAB000D0540004000AAA000C00150000AAF0BD405400";
    attribute INIT_27 of inst : label is "0FE600FE07FF0001FE400000C550554000003CAA03F400150000AA3C1FC05400";
    attribute INIT_28 of inst : label is "003B00A000510000EC000A00510000000002FF803FC00000BC0002000FD05550";
    attribute INIT_29 of inst : label is "00A5037C000500003FD00FF000000000026F002A000000002A00FFA030000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000FF803FC00000BC000AA80FD0000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "00BE001F00000000BE00F4000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "1D10000C0601000004740000009000000000000C000600000000000000000000";
    attribute INIT_31 of inst : label is "30000000160000000280008003800200C0002000C000200000A0002000000000";
    attribute INIT_32 of inst : label is "008025000000000002000058000000000C00000C00060B8000300000000002E0";
    attribute INIT_33 of inst : label is "00000000000300081400000050000000000000000000000000A400206A9D0000";
    attribute INIT_34 of inst : label is "000C0064082F002EFDC00000FE008000F9F300102E000280FDF00000AFFE0000";
    attribute INIT_35 of inst : label is "2CCF50002FE02E00CF00002900080000000F00682FFE0000F7C0A0A8007E0000";
    attribute INIT_36 of inst : label is "000300182E000280FD70A0002FFE000000F3682A20150000F32800050BF80000";
    attribute INIT_37 of inst : label is "000FE0002FFE0000F5C00000002E0000000F0E00082F0000F5C00000FE000000";
    attribute INIT_38 of inst : label is "00CBE0002FE00000CB00028C0008000000E3328020000000E300000B0BF80000";
    attribute INIT_39 of inst : label is "0002007F3FFF0ABFF400AA00FFF8FEA0201B000007F50005EC000000FFF05500";
    attribute INIT_3A of inst : label is "0C330C33014100000CD00CC0504000000002007FBFFF0ABF7680AA00FFF8FEA0";
    attribute INIT_3B of inst : label is "FFF02FFF747D028B0FFFFFF87D1DE2801FF53FFF1FFFBF8B5FF4FFFCFFF4E2FE";
    attribute INIT_3C of inst : label is "BFFF77F07FFF00AFFF800380BFC08A0007F5FFFF017F2FCB5FD0FFFFFD40E3F8";
    attribute INIT_3D of inst : label is "0FFF3FFF17FF00AAFFD00140FD008000D7FF3FC02FFF0ABFFF800000FFC08A00";
    attribute INIT_3E of inst : label is "2FEB3FFF07FF02AFFFE0BFC0FD00E2800FFF2FFD1FFF00ABFFF80140F000F8A0";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000002A2033300000000A2A0333000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "15553E00007CFFFC555404BC3D003FE115553E00007CFFFC555404BC00000000";
    attribute INIT_01 of inst : label is "0400022FBD20006000007D80063B0018000000121980090000006E003D003FE1";
    attribute INIT_02 of inst : label is "D000FFD0D0000000D00000000DF3093408508C9816C001C4000685B0009D0210";
    attribute INIT_03 of inst : label is "FFFFFFFFBFFF00BFFFFEFE0000000000014000009000400000000000D000FFD0";
    attribute INIT_04 of inst : label is "0000000000000000014000000001000100010000800000004000000000000000";
    attribute INIT_05 of inst : label is "0000F00F0000F00000401DD51FF22FC700043FFF8FF4D3F81000FFFC00060001";
    attribute INIT_06 of inst : label is "01401E0015502ABC1550B55414003C7815502F8055547E8055500F000540F03C";
    attribute INIT_07 of inst : label is "FFFFFFFFFFFFFFFF0000000F0000006000002AA8000002800550FAB415501AF4";
    attribute INIT_08 of inst : label is "5540A83C00142ABC55502AF00554F03C1540003C15547ABC5014F03C7AADEB83";
    attribute INIT_09 of inst : label is "1550F03C5014FBFC5014FFFC555000F0541407BC1550F00055500F005014FABC";
    attribute INIT_0A of inst : label is "1010FBBC0100F8BC1550F03C05000F0015502AB45414F83CFFFFF41F0014F03C";
    attribute INIT_0B of inst : label is "FFF0FFF00FFF0FFF00100B40FFFFFFFF040001E055541F8005003AC050141FD0";
    attribute INIT_0C of inst : label is "03FF00000000005FFFA000000000FD00F001FFFFFFFFFC10500FFFFFFFFF003F";
    attribute INIT_0D of inst : label is "03FF0000000001FFA00000000000F54000220000000002996E0000000000A640";
    attribute INIT_0E of inst : label is "000707FFFFFFFFFFBFFF00BFFFFFFFFFFFFEFE00D000FFD0FFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFF02FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFF0000FFFF000000001FF4167B90033FFCC003307FFE00";
    attribute INIT_11 of inst : label is "000707FF000707FF000700000007000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "00000000FA00000000000000000000000000C000000000000000000300000000";
    attribute INIT_13 of inst : label is "00000000F000000000000000000F000000000000000000000000000000AF0000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "00000001000000003000600000000000000000341AA4000C00001C001AA40000";
    attribute INIT_17 of inst : label is "1955C0001800C000001000000000005004000000000005000024000300040003";
    attribute INIT_18 of inst : label is "0332000000000151B310000000005150033300000000015132B0000000005150";
    attribute INIT_19 of inst : label is "00330000000000152B0000000000150003330000000001513340000000005100";
    attribute INIT_1A of inst : label is "00FF0BF0000000FFFF000FE00000FF00FE15F3FF54BFFFCF0FFF0BFFFFF0FFE0";
    attribute INIT_1B of inst : label is "02FE000200003FFF0F80AF800000F77400BA000900000FFFA60060000000FF70";
    attribute INIT_1C of inst : label is "0C0502550000005A0300A000001486000FF80000000001FF000000000000FFF0";
    attribute INIT_1D of inst : label is "03FF022A00000FF4F400FFE0000406000BFF000000000EF7D00000000000EA00";
    attribute INIT_1E of inst : label is "FFFFCFFF0F000F000FF00FFF0FF0FFF000F000F00FF000000000034003FC03FC";
    attribute INIT_1F of inst : label is "00000000FFFFFFFF4000FF409DDDBFFFDDDDFFFFDDDDFFFD00000000FFFFFFF3";
    attribute INIT_20 of inst : label is "00000AFF000000AA0000FFA00000AA0000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "00550ABF000000005500FEA00000000000550AFF000000005500FFA000000000";
    attribute INIT_22 of inst : label is "000002FF000000150000FF800000540028400AAA0000002A0128AAA00000A800";
    attribute INIT_23 of inst : label is "000003F8000000D500002FC000005700000003FF000028AA0000FFC00000AA28";
    attribute INIT_24 of inst : label is "00150BFF00000F5D400FFFC00000750028550BFF00000175AA00FFC01540D400";
    attribute INIT_25 of inst : label is "3C0503FF000000D7503CFD500000D7003C050FFF000000F75AA0FFF00000DF00";
    attribute INIT_26 of inst : label is "3C0003FF000000D5000055F000005700000007FF000000D500A0FFC000005700";
    attribute INIT_27 of inst : label is "07F90FFF0000000550000AA0000075D0280017FF000000D50028FFD400005700";
    attribute INIT_28 of inst : label is "03C500FF0000000A53C0FF000000A0002A037FC00FC00001F0000F7003A05554";
    attribute INIT_29 of inst : label is "03BC005A0000000A0FF03FE00000000003F4003F0000002A3F00FF0000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "3F827FC00FC00000F0000AAA03A0000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "00FF000100000000FF0040000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "000C00060150082800000000054028200000000C1AA40034000000001AA41C00";
    attribute INIT_31 of inst : label is "029530000000290050400140010007401955C0001000C0000010005000000000";
    attribute INIT_32 of inst : label is "034000000000000001C0000000000000060C000C000309340090000000001C60";
    attribute INIT_33 of inst : label is "0000000000040003000028000000A000A955000000000000501000580000956E";
    attribute INIT_34 of inst : label is "000F000007FF037F7EE00000FD00EA007C0D00001FFD0100FEF800005FFDAA00";
    attribute INIT_35 of inst : label is "947F00001FD03FBFFD0A00140554FE34000700011FFD0342FBE055FD1FFDAA00";
    attribute INIT_36 of inst : label is "000100051FFD0100FFB850001FFDAA80A07F157F1550B8BFFD16400007F4FE2E";
    attribute INIT_37 of inst : label is "AA0750001FFD0342FEC000001FFDAA000A87050007FF0342FBE00000FD00AA00";
    attribute INIT_38 of inst : label is "A07F50001FD0B8BFFD0801540554FE2E207F154015501CBFFD0A000507F4FE34";
    attribute INIT_39 of inst : label is "002F0BFFFFFF0024FE00FFE0FFF4BA00FF050BFF000000175000AA803D505D40";
    attribute INIT_3A of inst : label is "0C330C33000002800CC00CC00000A08000AF0BFF7FFF0024FEF0FFE0FFF4BA00";
    attribute INIT_3B of inst : label is "7FFBFFFF0010AFEBEFFDFFFF0400EBFA03FBFFFF005DFFE3AFC0FFFF7500CBFF";
    attribute INIT_3C of inst : label is "FFFFBEBA05500FFFFE000BC05500FFC0BFFB07FF0000DFE3EFFEFFD00000CBF7";
    attribute INIT_3D of inst : label is "0BFF3FFF00150BFFFFD0FE004000FBE00FD03FFB0550BFFF7D00FFC00500FFC0";
    attribute INIT_3E of inst : label is "3FFD3FFF000007FD0540FF000000FFF002173FFF00550BFFFFD0A0004000FFFC";
    attribute INIT_3F of inst : label is "00000000000000000000000000000000033301510000000033B0515000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
