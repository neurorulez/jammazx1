-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA5555AAAA5555AAAA557BB3F9ABBCB6496F58ABC5BE53ABAB5353A9AB";
    attribute INIT_01 of inst : label is "529A950417AD6B6B0D251E0145336F4E9A7BECFA785ECD9D244BB9AF75B4DAE3";
    attribute INIT_02 of inst : label is "8F2EB3B67CBF6749F63CBF6749B63C924C01102004A477FF3DFEC965901A0406";
    attribute INIT_03 of inst : label is "0E10E9E126D72218044935C80681126D722180468A124D722282EB3B67C9AC6D";
    attribute INIT_04 of inst : label is "9261BBDE95CAD6232B430ED372C9FB9E800302086819EAA56E1E90E1B87A4393";
    attribute INIT_05 of inst : label is "0CC30C300330C30C3ACBD65DA466C9892766C98926E240516598B26C68015CD1";
    attribute INIT_06 of inst : label is "073940739439C2F23AF7C9B3D67FDC7A1D1CF64F05DC9773900F5DB05C4DBCE0";
    attribute INIT_07 of inst : label is "C963FE42BEEB12E8153DC93409BB8DCC5753435E9DC9209DC97EDDCE71D0E71A";
    attribute INIT_08 of inst : label is "18A3D03CA76FBEC427204C4D6496A422128072188004AC28139924D14AB1A0C5";
    attribute INIT_09 of inst : label is "C15DEE944A75A043A6FDBF5CDFBFE91A0920CD3A504AA4A894A1248287FC4012";
    attribute INIT_0A of inst : label is "3A47C1C8592F48DFFF7F74092DF01F41F01B6225AA65B34C2AB5048AAD806242";
    attribute INIT_0B of inst : label is "66EC859A1217340801DD5434BC3D70444474966988ECE01FA05028284500BC2A";
    attribute INIT_0C of inst : label is "8088160282960AFFFF76B5B0641973637FCFC36E63FE0632DC6E7E3F1CB66D9B";
    attribute INIT_0D of inst : label is "8FDF6DAAC3414D61B4B0CDB815BC32B656F0CAEEB1FF319BE0785C0E0703806F";
    attribute INIT_0E of inst : label is "F66B39DD1653B4A30BA4BACBBCBACB24902945EFFBCD7D35BCDED37BC97D2010";
    attribute INIT_0F of inst : label is "FF602DFF64EA69B6D27DF9F7FD963B710670A97264B49CB776B3DD273A5339AD";
    attribute INIT_10 of inst : label is "48AA08D1157C83D35D296A6DE7D80290D10558A0A885527907A6A7F7F0FFFE7F";
    attribute INIT_11 of inst : label is "ABEDDB90B52AB7E9BD00042E588CAFDB4A1B6942E173B7C5BE9B27A2050BC000";
    attribute INIT_12 of inst : label is "D0550DFB77FD411BC101A00622A2F6F51159E9015281FD8B6EFFFB16FDFD54A0";
    attribute INIT_13 of inst : label is "410073A69E74D2D06D4B580800256ABED11ADA215A217EE15EE152D484FFE67B";
    attribute INIT_14 of inst : label is "E62A9A492005AC398E638080BFD6E79CDFBA351A8C01E59E5B47983EB20C5EEB";
    attribute INIT_15 of inst : label is "0000D49C001B3AE800065660000062080004B7300002C180000055800CF5B92C";
    attribute INIT_16 of inst : label is "000F4230000FB0640001CF800000A40400155050000FDAFC000AC4D400101AC8";
    attribute INIT_17 of inst : label is "54A50412855A168A28A28A28A2882B4A4000A300000136E00006B75000082308";
    attribute INIT_18 of inst : label is "8BCF5DEEF4C49637F55F150C48987A709B9C6849E18A2811A55295114A515129";
    attribute INIT_19 of inst : label is "FC5AEDA7BB739CE7057FDEF7BC17FFCD4454D33D377A01EC20816A5AD05107FF";
    attribute INIT_1A of inst : label is "02801B8229E2A8AF390E3490A5DF6337320FE08B09E7C11613CD90793F230A3F";
    attribute INIT_1B of inst : label is "4994694E090D553899D3093244C10B970C78A881418E0A3C48C2E183869B14F0";
    attribute INIT_1C of inst : label is "88E7044E549648CE19E324CB25560248E14C98C23D09D988865A95D5A651C8E1";
    attribute INIT_1D of inst : label is "26173920E92B913BB7C57EA84093930B576901C35BCEF780000003423148533C";
    attribute INIT_1E of inst : label is "7CB1E64E80013334D9B40F2F1F11CF2A8F1F11CAF6778145310F40E89EAA502F";
    attribute INIT_1F of inst : label is "1E94E6CFB67F9F3B4F55A7AF3B4F55A7AB75BD994FCE3754024EC8FC385EF6B5";
    attribute INIT_20 of inst : label is "9ADE7DD9F7FEEDFE697F32DB0C9B7DC17CBAEB2405327064D5DFACC12F850000";
    attribute INIT_21 of inst : label is "065E7843CF2A5019F7EFDFBF3FFEFD0FAFDDBE496F7FD9E6B6EEDF37BDF9F3EF";
    attribute INIT_22 of inst : label is "00014B2E005214F9820000016C41D72B08164E6B059098026C4F013B4684ACB3";
    attribute INIT_23 of inst : label is "38E38EE38E389C71C75588AACFD9711559EB2E22AB3E75C20220220092888020";
    attribute INIT_24 of inst : label is "987663BAC168630C4C55D86EB01A18C3315DA6E31D0CCC776BAAAA0071C71C8E";
    attribute INIT_25 of inst : label is "134D6CECE1BEAF73D8113964C4214040CC333858210C98AB2099808108462B24";
    attribute INIT_26 of inst : label is "F7B595047AC200C323F5883B906CC8331F70EAA9265844CB00C51A79392EEEF1";
    attribute INIT_27 of inst : label is "F74A6A13B17DC129B084F3A2A94554A137F2DCAA26FF5E8F68FEAF53F9424E91";
    attribute INIT_28 of inst : label is "4A372215BAADBD1268F856F51EFB5150058004D903C9206D023840884179F267";
    attribute INIT_29 of inst : label is "11BBBBB2AAAAAAAA000BCE15BB7251BE910ADFF45937CD2372215BF68935E8FE";
    attribute INIT_2A of inst : label is "EE7B1AC7B9EC290A6398A4298E6290A2198202826C5F7049412B3028F0144111";
    attribute INIT_2B of inst : label is "154D04AD8142A4FB16DED08B05A96B41442AEF7DBCF57E69A69AB1AC7B9EC6B1";
    attribute INIT_2C of inst : label is "4AC73EB208A8A8CBF815337118929494CA35A267ABC8FDD733D8410297F8BCCD";
    attribute INIT_2D of inst : label is "415106395919961179CE0A32C902AC6C6C48B02B336A5A8519971EEFB6F8A970";
    attribute INIT_2E of inst : label is "860160A0A0A04DC15E9FA559C4624494F4D94914A8D20511173644E40865290A";
    attribute INIT_2F of inst : label is "800086DBAA000004056DBB71AC6B1AC6A28732C22E2C3161D3E74D7EF5D7EF5E";
    attribute INIT_30 of inst : label is "9DE77EF15BE8B9E2BFB66E4E4AE78AAFFB6FD67EFA8880ADE05316E23542A54C";
    attribute INIT_31 of inst : label is "1040ADBB7DB55F9165F068E7C458C3F87C50142B6FEE7F63FBD424A750895707";
    attribute INIT_32 of inst : label is "1580276FB7DBD294B6C12911001015A960ADBEE2F0569261A26F021072A21518";
    attribute INIT_33 of inst : label is "99690D25A4349610C2F1004050108094EE7E299FB4FC167742415EF31F202424";
    attribute INIT_34 of inst : label is "6252280310620C498B7F3F7F3E5EA0F0F0F0F1AE80000200675D136AA9A77799";
    attribute INIT_35 of inst : label is "59F4F7CEF73BBA6B8AFBEC397E9B60F9A71FE931C2020A2D3FF99BA73ED25260";
    attribute INIT_36 of inst : label is "5B9DFB9FA4DB564FAF4C67CD9D689BDF4FE7A739FDAEB36B3663F59F59F4FD9F";
    attribute INIT_37 of inst : label is "FBE96EBA54BAF4846CCF56EEA3ABCF4B3695F776FDF4DDDD999DD44B7482CB9B";
    attribute INIT_38 of inst : label is "01ED56EEEC51A7FEBC113D2CC77413E18CFFEE6F9BF768C77B89AD8FDFDFBE65";
    attribute INIT_39 of inst : label is "2333768DE6F379BBDE6F379BBDD1EBE9E8772B5D759741DBA0DF5414BAA0BB14";
    attribute INIT_3A of inst : label is "9310211BDFC9846EDF2019BF242A19B3C58541190CEA1C4B70E25B8400882732";
    attribute INIT_3B of inst : label is "4B28ED615D6B35A5EB8F0B823118ED73E1FAE2D094C4A4013309084C42441312";
    attribute INIT_3C of inst : label is "B8FDF90141DDC640798D8219F4D900B7E119B7102A0EFC42F3F92235910BAC44";
    attribute INIT_3D of inst : label is "D196F03B67F9FFFAD19C231C72F5F43319A5759727A513BCF47796F7AE0ED6B6";
    attribute INIT_3E of inst : label is "86C91C0059852CC315D6910C1AFBEF224CA3654AEB59911DE5BDE18BA6B6B005";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA555586030D9238F1";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA5555AABA5555AAAA5549F00CC0482101B02F5F66C053ADAD5351A9A3";
    attribute INIT_01 of inst : label is "5B72DA62DDE2B90756949445F246009364A489EF8F9BA106926E561CA6DC0971";
    attribute INIT_02 of inst : label is "D6C158CB1BACB4BA8B438CB0388B0BEDBF5EBBDF78B7D4AA542A879372E371BD";
    attribute INIT_03 of inst : label is "6AD5420A59379B7575B65DE6DDDD65B37997775BB96DB779ACBE95ACB5B2D6B2";
    attribute INIT_04 of inst : label is "74DA011B3993DB58CF65B3719BAD2908ED9812E5B6CC1132993B39C8ECECE722";
    attribute INIT_05 of inst : label is "60E79E799839E79E4D302882CB4B969E5A4B969E580F4976B3766E9B0B657BB3";
    attribute INIT_06 of inst : label is "0001C000080006F5EFD994C379B35312E954DD4DE1F806E02D88A33141E64226";
    attribute INIT_07 of inst : label is "400D092E4C8431AB2CD84208B8AF3979B5856B30AC8030AC803253800170002E";
    attribute INIT_08 of inst : label is "F9A50B05AB22F30A759329CE820CB6453BB35AC959DF5694A00240522DBFF20F";
    attribute INIT_09 of inst : label is "1E34C0636DCA4D260C2E1C93098B1160B4B7DE91092F366B294B89252FFC94DA";
    attribute INIT_0A of inst : label is "C9682D06E0B53DE58B16C9E4B922D26D26D20D394B3064068B17635ED0B5B037";
    attribute INIT_0B of inst : label is "23006E02A1B8C9F6DEB2E707C3438729C05D000024B90560578EFB182372B086";
    attribute INIT_0C of inst : label is "3A514A446ECCC719324DAC20601A0ECA5C9CA149CAE502A1B349E4722DC2308C";
    attribute INIT_0D of inst : label is "BE45E64B2E263392411B46AD5A724AC369C92B756572AF3C4E8B6DD6EB75BA71";
    attribute INIT_0E of inst : label is "D03C6002676F722DE7FA77A7F27727F219F7D952903E20EE1BF06EE93F26B3ED";
    attribute INIT_0F of inst : label is "FF8D627688FAA68A660508953B48CE31B4766CAC283B05D19BC721F643E1B238";
    attribute INIT_10 of inst : label is "26915D262E42349C314611C44E61CBF719DFC3ACB145EC0469386FF3F9FFFE3F";
    attribute INIT_11 of inst : label is "2C70C00DC2AC81A549B732F5E6B07C2CB165962D22A17BD21854A93252B01B9B";
    attribute INIT_12 of inst : label is "1DCD309839722D610ACA4B24ACE4C726E2624D658B4A16FF27402DFE6E250ACD";
    attribute INIT_13 of inst : label is "8A9948DB600924E68A119EEE4B5252D5E673CCF3841B8225C3058C21E839AC21";
    attribute INIT_14 of inst : label is "C3BE440A00036A204A021991D96C9B2962444A2111CE4925E389214B2C55E333";
    attribute INIT_15 of inst : label is "0015DDD4001F84780003263800042328000577100001D560000033801C41F00D";
    attribute INIT_16 of inst : label is "00064570000712F400158EDC00115A40000E1DC8001F117800034D4800012CCC";
    attribute INIT_17 of inst : label is "CCE27367898E479E79E79E79E79E3F7C000060800003B6200001B2B0000C7210";
    attribute INIT_18 of inst : label is "349503BE8ED9311BB095D2A481908F591AA29291139E79CDE62388DC9E666639";
    attribute INIT_19 of inst : label is "17AB20AD5D0421087340208421C80400888923424B82B96EED6EA4211DC96004";
    attribute INIT_1A of inst : label is "00800B230BA02C2155165989209D201F3045092DB70B1B7FFF1626F21C0C6912";
    attribute INIT_1B of inst : label is "AA842A50040D4341692591502140000F00E808C0408C960450E191458B1105D0";
    attribute INIT_1C of inst : label is "4088188031A9015008CA00948969200901A969614882B13005135846AA692901";
    attribute INIT_1D of inst : label is "01ECC2074D9672C9D17FBB37598D52836100A0829908C200000005442304C504";
    attribute INIT_1E of inst : label is "F6CF91F17C92A8F76BA4D00B50BDB48B6B50BDB7F9CE7CF0644CA74C60ED9730";
    attribute INIT_1F of inst : label is "0EFB43E01604A0089270493489B270D9335CA1960EA0F266223C19FB36C06315";
    attribute INIT_20 of inst : label is "27B2B46895B374ECBECE5D24576C8A6A808FCEF3B1802300557FF87EBBC41111";
    attribute INIT_21 of inst : label is "C48285A68106500C99BA66E9DA246C5898D6A8BCC6356A89CC6B545E6468952B";
    attribute INIT_22 of inst : label is "B7B68EB8DBCE77FC2E0000105560A469AC0A8D0502A044062CA4015AB5885534";
    attribute INIT_23 of inst : label is "AD4AD4B52B52D6A56A65713316AA4E2662D549C4CC58893B993312CACB435AF7";
    attribute INIT_24 of inst : label is "7265B8E468B935875F606D399B2C4D71FD86F39376E3971C82000000A56A56D4";
    attribute INIT_25 of inst : label is "872E9781DE0B966F262CB65B9999B0C0038E4D2C9AC6BEC0DA726964D63FB0DE";
    attribute INIT_26 of inst : label is "47284228936498649B3DE55B4AB0E576CCEAB331C1A7C93CD3324DD22DCAAAB5";
    attribute INIT_27 of inst : label is "5024A16CDA940492825B737864A4A366D7F22096DAFF45C920D23CCB4FFED527";
    attribute INIT_28 of inst : label is "AB68447F19B942715131FC62200523225A1362A1DAA482A8295658F26652D4AB";
    attribute INIT_29 of inst : label is "5005050811111111BBB2107F1A955B41223F8D636D4851368447F1AC6DAA132A";
    attribute INIT_2A of inst : label is "2080E6290E60C2728C276AD2F6AC272CE376AD3C36A5012524B26D7F27AA9050";
    attribute INIT_2B of inst : label is "0A50BDF0336CD0286754FE96BA90847725AE302549474192D92F0E6290E60806";
    attribute INIT_2C of inst : label is "8D0A504453153316276940D421D9DBDC25FA67306C7B557F02DDDADD444B492A";
    attribute INIT_2D of inst : label is "ECCD944A6A2AE4E2C212EC45848C58999984EB94544791B2E2ACA4B02C7A6EC2";
    attribute INIT_2E of inst : label is "5AD99B391BB74234D886B22650DDFBCC0E266562971918CCCDCA892890B8F7FF";
    attribute INIT_2F of inst : label is "44921CB844222222665C50AF7AD6F7AD6CD95CBC5849C25E68912689126C9932";
    attribute INIT_30 of inst : label is "76B5FD222C512645FA59088F249917FFA58165830331353E84D401A8432E5CC2";
    attribute INIT_31 of inst : label is "766C395D13996022588002B098B29D928B6366E588224182082BDE60FF115B8B";
    attribute INIT_32 of inst : label is "47A50108C4421C6324DC91999989994230C46CB090F0A08C16920ED9C8E57970";
    attribute INIT_33 of inst : label is "0C989312624C498931FD210C8A52199ECC38521C8D90D40D20057EFEDEF90000";
    attribute INIT_34 of inst : label is "1400101989316624C551191158FB2ACACACAC809C410C10888A2213B12D8FA01";
    attribute INIT_35 of inst : label is "B2091CB102804192D30001532924C803004005AD22F991DB600B304842875455";
    attribute INIT_36 of inst : label is "B13600248C7C8BF20096F892F0D7A47091C8487A06024C805844596CB21B016C";
    attribute INIT_37 of inst : label is "E4367A449F691B2D9B72C12229607BFB4B2328CB320972232E6136B60A61BFB0";
    attribute INIT_38 of inst : label is "E80117AFAE45B6ABF6AA8610188AA099612002A22896510A06D0C368009528A9";
    attribute INIT_39 of inst : label is "454510C00000002A40000002A43882828044CBA69A20612130BB893F155F41A9";
    attribute INIT_3A of inst : label is "57770083691F110C245440BC747040ADAE8E02440242FBD59FDEACFD61E01144";
    attribute INIT_3B of inst : label is "8F8825E1E20095672A8E8E8104420573F167E21D12A09500B901C90A89520B92";
    attribute INIT_3C of inst : label is "48812353526BC018C2254B90C54923CD0318480811792063022921F01307C111";
    attribute INIT_3D of inst : label is "0A6048881822E820603436CB04454081442E9A222A06685A4044658A07201DC8";
    attribute INIT_3E of inst : label is "2AE5827604AB025416000950030C307659A00ECF1004BB1119628EC103370520";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555808055CB04E0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "5555AAAE5555AAAA5555AAAA5571F0B3092FDFE9CA31FAC73C52A8A85052A8A1";
    attribute INIT_01 of inst : label is "665BA333A5F2F41A9CD70465625328FDB6F32C93B1B620D88D0B25724134E9F0";
    attribute INIT_02 of inst : label is "D2797A0F4966F5966F5162F5966F591652F10E61C6CC85064141926CA799CCE3";
    attribute INIT_03 of inst : label is "2495C36EDB65E18BD716C9786275C5925E189D7391CD965E32E5B7A0F49E5E83";
    attribute INIT_04 of inst : label is "6F5C6716DD6294630A466CDB74F0C31267733B87647B3E6CC496DCB59A5B72CA";
    attribute INIT_05 of inst : label is "04E38E388138E38E1BEADF59A66CEB8BED6CEB8BEF5B769CA3646DEBCE799B33";
    attribute INIT_06 of inst : label is "0AB5E0AB5855AA576D1D47E2DF715D2A956CB56B206A00A0C8C32DAAA4F65BE2";
    attribute INIT_07 of inst : label is "8AF233339259934ECFBFEB6E6B3BCDC72737091E798EB0798EA31D956AF9569F";
    attribute INIT_08 of inst : label is "A4B00C010A13E023B7318F732496C391D93C739264D33D873E0B66D8D9A73C66";
    attribute INIT_09 of inst : label is "72FFFEBDD36313926E0A5418B30201CAEDBD18180E30C38E8843A4910D570463";
    attribute INIT_0A of inst : label is "5983E92BC8C7B7A95AA5FE3368C78E38C38E7905EE05F6EC2EBDC48BBDCF635E";
    attribute INIT_0B of inst : label is "C35EBCFBDAF3B6DB48E7F7B57DFAF58A6474375988EBE427599B314899920CA4";
    attribute INIT_0C of inst : label is "AF390A6C6C64F24DBFEF7AFAD2B6EF6F6FD6CC9D6B365DFDD9ECFEDB6BDC376D";
    attribute INIT_0D of inst : label is "CC27C0EE3279FDE395FE1DB9F3AC739FCEB1CE5DB59B35C9FAFB397DBE5F6F27";
    attribute INIT_0E of inst : label is "1537F041978C6039E4E04604604E84E84CC7624215F714CA8B2A0D84B690918C";
    attribute INIT_0F of inst : label is "FF80E0722A5C38E38E940A5034B2E2AA0A22888D28234D119F7E05F56BE1AB4C";
    attribute INIT_10 of inst : label is "32C72D98CB66967195FF7FE26D06DE1C772ABCBAC65E32CD2CE327F7F8FFFE7F";
    attribute INIT_11 of inst : label is "B0C4A9DF98B0076DE7236336C9E25E36D982CB30A7E162BD36DE6CE4B0C65C8C";
    attribute INIT_12 of inst : label is "4CCDC334A85031C6531312363926F79C7F7339CF36765C7E840CB8FD08D0A265";
    attribute INIT_13 of inst : label is "DFB3FEFDBFDFB6F2F35FECEC61667B258809A5BCF6AF2E664E477EFFEA228429";
    attribute INIT_14 of inst : label is "433C8C07B541CE4A1AD49991EDB6FDAFCB46633199CF7DE6CBCDF16DBED8F3BB";
    attribute INIT_15 of inst : label is "001156480014801C00017110000251300002C4A00001A6C000000F0037C01401";
    attribute INIT_16 of inst : label is "0008375000102084000C2C1400119ECC001395C00010E080001395C400107500";
    attribute INIT_17 of inst : label is "01A40006800A029A69A69A69A69885790000EF800000B2A0000045C000084530";
    attribute INIT_18 of inst : label is "96DCC880229CA539FA1E9898E02112604EACECE5999A6911A44290001A004068";
    attribute INIT_19 of inst : label is "9BC229CC33294A53334BBDA96CC973A4CCCC29C30F349D21454B0C4B4CC9D0F7";
    attribute INIT_1A of inst : label is "000038420323480D5994A9F2481001401941CED2498B9DA4931632729C59E923";
    attribute INIT_1B of inst : label is "2680A489395C2C34E84510D316E292140EC8D08003810E3424CBE285152E0190";
    attribute INIT_1C of inst : label is "9164964D739711093B10480B8D170C8C9220EBCB485CC42D2A029B929A504C92";
    attribute INIT_1D of inst : label is "022F1A5939E3DDBD09BB201D76BA8A3271A6234A10529080000005694B625BAB";
    attribute INIT_1E of inst : label is "E38E66E1899CA769BF571B757F314365957F314DD27789B1B36B3939FF2F5C2B";
    attribute INIT_1F of inst : label is "C736718C8627B7E9F9D0FCE7E9F9D0FCE2673D58CBA5E276206C4BD428E3D6FF";
    attribute INIT_20 of inst : label is "3603972E582840A4F80CD00C55080E2A2225D39E3E236446DDDDDF22360DC9C9";
    attribute INIT_21 of inst : label is "091AB5C66D4F50085420528502042EDA5D72E4FA03070E0FA038706C072C5831";
    attribute INIT_22 of inst : label is "C8C8D3CE76B5A9D09204445509422375281301E004C3900A4F0900F15691C164";
    attribute INIT_23 of inst : label is "CE7318C6339CE7398C7A3BBB9B3BD777736772EEEE6CCF51B3111337B65EF79C";
    attribute INIT_24 of inst : label is "D8464BB28DC146095E7B916CA372518279E936CA992EE9773F4444FF398C6718";
    attribute INIT_25 of inst : label is "1BCB6DE6B78CB653ED39A8768CF4C08044BB1170A308BCF722D88B85184F3D26";
    attribute INIT_26 of inst : label is "57BCB72CCE6498649A24AF495BB0657C7AB33C3E02688E453946079D32355555";
    attribute INIT_27 of inst : label is "1DCFFE7ED1C74F3FE79F902F5388F3E7F562611CFEAC4F897A9FB6537CC77FF5";
    attribute INIT_28 of inst : label is "C3EB279B513D599B798E6D4732FE7C780B3996F0CA6C87E821F418FB22715304";
    attribute INIT_29 of inst : label is "500055020505050505070F9B53D61F5F93CDABB271FB583EB279B5764E2ACC7A";
    attribute INIT_2A of inst : label is "11884308001398C7A9285B9AC7AA3099AA43C830B471D3CDEF177697FD5FD005";
    attribute INIT_2B of inst : label is "9F5C9957C631154795921B12AC312D3327300E3D6DC9FB6D249B085398C70800";
    attribute INIT_2C of inst : label is "C5CBE476799D9999D18D67610CE6F2F79E7226B2318EBB6E8A428A964F716DAB";
    attribute INIT_2D of inst : label is "89D9976B6B2BB6F32B18C4564F0F0CC4CCC6F19666721EC6B3B637F03E578BE7";
    attribute INIT_2E of inst : label is "6260CB9139397AAE56F598308471CA67A383397CC1CE1E49CE7AC9AC9CEDC679";
    attribute INIT_2F of inst : label is "AE38BEFD67236323627C7EB33DC6798EC6E176DE656FE36F52E54D2E54D6ED5A";
    attribute INIT_30 of inst : label is "DAD6E983391DB76F7072C469C6DDBD5D273DB7CE5BBBA7AF20D632C2118B9779";
    attribute INIT_31 of inst : label is "9D31CDD09B41868B7E053FDAACDADEDFCD7667073AE49726BD48533CFD450601";
    attribute INIT_32 of inst : label is "7021013A996EE6BDD30898D9C9D8CEEFD000BED5BB32F13883CE338E2331DD91";
    attribute INIT_33 of inst : label is "D84A0941082104A09414214DC8D29BBF28801BD20950517D09070686D4780090";
    attribute INIT_34 of inst : label is "36573ECB21646C8D918189C980D6BDB5B5B5B56E042041082B7C725E1B6F606A";
    attribute INIT_35 of inst : label is "DB6DCBEB6391B6DBDBA9767C55BDE839A39FE639C3919152450AA86D50875620";
    attribute INIT_36 of inst : label is "69DCDBBD8F30DF5F6CDAE7FFCD5CBDD2DB8B6D769F6FFFDBEC26EFB6DB7FBBB6";
    attribute INIT_37 of inst : label is "36FF17F6C5DFDFEC7FFF76FBAFBB6B6BFFB4DDFEDB6DE6EFFAB8A4953087CDE9";
    attribute INIT_38 of inst : label is "42BAA91441AE4D540EBBE9145BBB37ACA5E9444711D1718F9F5B77AE5E5EBC44";
    attribute INIT_39 of inst : label is "055510F0582C16050582C16050135151504849659602A10050B18BBF44002F17";
    attribute INIT_3A of inst : label is "1282E002AB02120A2C20042C202E04288525E2AA01538A04945024A010181044";
    attribute INIT_3B of inst : label is "4D5A0019410802A785010100048020820164020B101C02C414003025400C0060";
    attribute INIT_3C of inst : label is "E01103A3B2D010B0A6075F944042C2C1371628A0885186A29422C0003C14800E";
    attribute INIT_3D of inst : label is "0248AC004122C122803C28A280ECA80840359607E546C208A8C585903C221040";
    attribute INIT_3E of inst : label is "02AD4154402920159410A2560145145440248FCA0840393161640B0810520784";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA55558000055A82A0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA7F57AABB7755AAAE55FE90B35F6C924DF33621B7D756AEAE5456ACA1";
    attribute INIT_01 of inst : label is "AC5D622BE7C471B28A5AA906CB3A6058B2DBB75B394D82BC8903B1A361A7E8A0";
    attribute INIT_02 of inst : label is "D6E338C71B02713267530271B2275016C1696D6DAD588184404190658B5DA6D7";
    attribute INIT_03 of inst : label is "3621F349FDEB51E5B2FF7AD4796CBFDEB51E5B2FD5F7DAB51C5C338C71BACEB1";
    attribute INIT_04 of inst : label is "390EB20D97D84E77E1273F926E1FC679766D9D47CDF58B48C54D936F9D364FB2";
    attribute INIT_05 of inst : label is "C9C51C51F271471479E3CF19E72449996D2449996E7BAEDCCE3AC721C7B4E1C2";
    attribute INIT_06 of inst : label is "0798E079803CC3029104FB2DB2410F8B358B6E46D3484C21CABF3D300E9110A7";
    attribute INIT_07 of inst : label is "A8FE5AB7936B9FC59FBDDFBE4D55CCBE32DF0B5A2805302805412E0F3038F307";
    attribute INIT_08 of inst : label is "74D62D100597D1633ADBF75335D65B71995B2D536D6BDA9ED4FDFDCB914AFB66";
    attribute INIT_09 of inst : label is "736FECEFD371FBDBAA2648ADD68994B3E6FF940C1F3DF7E71841401307FB8279";
    attribute INIT_0A of inst : label is "61B1A72B4ADEB42858B7A6724FEB7CB7CB7EB9D6E71ED75DE7FDDEB1EDE65F5A";
    attribute INIT_0B of inst : label is "C27EA4DA7A92924905D274B6ACD9B38E4E2C36EF1C5A8F33C8F93BCB9ABF68E5";
    attribute INIT_0C of inst : label is "A913CF7FD565F764C9F319FC9324A921324272DD2193C8DC49249249389DA709";
    attribute INIT_0D of inst : label is "5A2FA2E7B2BA7959657C9955331B29E7CC6CA78890C990E9BA363148A4D26926";
    attribute INIT_0E of inst : label is "1E2420D7F6CED05686506D06D06D06D06ED7AC108423349C9A7A49E9A734D5EF";
    attribute INIT_0F of inst : label is "FF404860AE08AAAAA4112044BEDAA000A200821A044A807396434D297A514BEC";
    attribute INIT_10 of inst : label is "3F52BFFF99B5D7699D8E76A2EA2C6D4E66B0BF965CC2976BAED327E3F0FFFC3F";
    attribute INIT_11 of inst : label is "969428D698944CE6F68ABB6E485C149659B6DB34DBD043EA6C6E8ED4D2D34F4F";
    attribute INIT_12 of inst : label is "2EAAFD68992234BAD15150A297B2BBDB9151B4E6E4637A4CB146F4994263A275";
    attribute INIT_13 of inst : label is "CB3D9367D26CFA32C6768D57DD7BB97B0F0103B8BDAD3F4FBF6F94AD0C1895AD";
    attribute INIT_14 of inst : label is "426484316664C6A563083931E4B26C85CF2A359A8CAB2CFE4DC4BF6597D8FA88";
    attribute INIT_15 of inst : label is "000560380004348800087758000611200006D5C0000197800000FF8004F31098";
    attribute INIT_16 of inst : label is "00096310001CA41800033B5000003948000BEC38001018000013C7C400014640";
    attribute INIT_17 of inst : label is "98B22222D89B46CB2CB2CB2CB2C984F000001600000365400003D5F0000C5418";
    attribute INIT_18 of inst : label is "D65B6C0039AF29DDDF398F34606733A8C69858594FCB2C88B226C8888B22222C";
    attribute INIT_19 of inst : label is "7A254036A2F9CE72BAAAD7BDCAED5AEC444418A5170A7AE99D2919EF2EACB9C3";
    attribute INIT_1A of inst : label is "00000A4203618804611C0D8007C498E5C58252492454A49248A80041AD0738E0";
    attribute INIT_1B of inst : label is "43814005308E1018700798714241830408D86080008902100050C007018401B0";
    attribute INIT_1C of inst : label is "0C22900637850D05089126428A050C6850447145610008A0400A4C230E4A0850";
    attribute INIT_1D of inst : label is "4B072851B55B9894CBA6915E2E800532146E1F4550D6B180000006400B284913";
    attribute INIT_1E of inst : label is "A14E4520E8DCCABEF1F38DAB369BF5B9EB3699F432E5C207595EB1B6D3BE8BBD";
    attribute INIT_1F of inst : label is "7A1F0BD2A8158938CDB866D938CDB866D7BD6BEF7F1F42EF9B547B7DFE7CE77B";
    attribute INIT_20 of inst : label is "3D05132448992260D4102CBA1A265D22AA19138FDA8EED1DD7D7D75F4A2D7C29";
    attribute INIT_21 of inst : label is "0208A425042660120400120448110010142060F40102060F4010307A0B264898";
    attribute INIT_22 of inst : label is "ECEC98776EB5AD28FA04454465E269633C002B2800091C0206070050000061E5";
    attribute INIT_23 of inst : label is "0F83E0F83C1F07C1F07FCCA88911999151223B322A2447555D5D5DE3246C6318";
    attribute INIT_24 of inst : label is "EB7AE7D7C3F9E3FFA2A1B875F03E78F78AABA75B2B1F78FBDB2828FFC1F0781F";
    attribute INIT_25 of inst : label is "365CC874E1D762FCC936BF2EBBFCF0408E7D78FCF1FF454370EBC1E78EF15574";
    attribute INIT_26 of inst : label is "119EF56C6DCE76F697B81C313A7E55BBD33C3FC006798DCF3DC7165993AAAAB3";
    attribute INIT_27 of inst : label is "7C42FA17F51F0D0BE6858631E1432B3B62BD9C736C57BB544F0CC29436B498B3";
    attribute INIT_28 of inst : label is "6519A3F28C96CFE5B8FFCA351B5FFEFFAB95AB75BD2FFAF5F5653F5ABB3D4A14";
    attribute INIT_29 of inst : label is "05000050AAFFAAFFAAFD29F28DFB28CAD1F946992A39ECD19A3F28D324467FDF";
    attribute INIT_2A of inst : label is "318842004210C21090C7398852814B5AB19CB1DF7D47C343ED299DBD94CAC000";
    attribute INIT_2B of inst : label is "6F1E9813F2B7144FEF6E9516A467BCBAB297299E6589A649249B4A52908410C6";
    attribute INIT_2C of inst : label is "C5F96EBB5AAEAAAB9DEEEF6BCCECE9FD1D7A440E15A7EBC9D5D33A526E3D65F3";
    attribute INIT_2D of inst : label is "BCCCFBFDBDBDD339398FFFEAE53365656D61BD562B374DD6F15352529A7D47B6";
    attribute INIT_2E of inst : label is "FFFCF7DF7DDFD287F5A5DE9CED7DE87D31F5289A7A8A66EABCBF48F48DDED7FF";
    attribute INIT_2F of inst : label is "FFC0726D73AABFBFAB34B2EF7EFFF5BFF77FBA4727247123F7EF5F3E74F7EF5D";
    attribute INIT_30 of inst : label is "EB5A9789198893270AF2E65CA24C9C42AF24B2FE78888DA36FAED2D790A14BD1";
    attribute INIT_31 of inst : label is "EAB6ED2CBEC8BF812D04CBD686486648FC6AEBF333F7DFBEFD2943E910170606";
    attribute INIT_32 of inst : label is "630083B3DDEE8CEF402E9AAEFAAEE8CEF009D345B6277122C5FAFD6D3331D8D7";
    attribute INIT_33 of inst : label is "18C0180300600C018042DCBEA7397D7686A00A5841004CC511373044A8588313";
    attribute INIT_34 of inst : label is "7203315302600C01824A0202412DB0FA78FA7BB78C10400C631FB94B4B2F4808";
    attribute INIT_35 of inst : label is "CB45A6DA4E5712C998AD646A14B06C272320A69CE944453D350B9D2F9B735665";
    attribute INIT_36 of inst : label is "FD8A9299FBE4C51B265A224B479A3D985F622F28CBB492C92F23AEBAEB45ACB2";
    attribute INIT_37 of inst : label is "568B8C9BE3B265A0B6F552ECDAA9B536BEBD4D6D4B45A489B48EF4FF9AD9743C";
    attribute INIT_38 of inst : label is "EEEEEFABEBEBABBAFEAABF2443B5332C9CCD55D7D5E136CF135F25A76BCF9FDE";
    attribute INIT_39 of inst : label is "100000B0482412080482412081E3C3C3C0150D041027004280191D2FFBBEAEAE";
    attribute INIT_3A of inst : label is "5A0700028914000B245C042C545840208B8B0288144308041040208159404111";
    attribute INIT_3B of inst : label is "8D0201D1208097450F0B8F80000001C35127A21412E09764B805500A81704BA2";
    attribute INIT_3C of inst : label is "E0810383D24000F480015D144042C2413E1041F8084823C20422C1003914D10B";
    attribute INIT_3D of inst : label is "8240E08041024122A0382C9244B0E0804034102507064208E0C5C5123D001008";
    attribute INIT_3E of inst : label is "2601905C04BA025D1A2809740228A07C403C8B890404BE3171448F4102524784";
    attribute INIT_3F of inst : label is "7555AAAB5555AAAB7555BAAA5555AAAA5555AAAA5154AAAA554480804C0320B0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA5555AAAB5555AAAA554BE8A64441011595A640265656AEAC5454ACA0";
    attribute INIT_01 of inst : label is "49424A22C850A5446614F545C30CE489B24AAB070501B362D3B490C92A4B2779";
    attribute INIT_02 of inst : label is "858952AA5604A1E00A1E20A5624A5424035A6B4D609280410110D0480AD56AB1";
    attribute INIT_03 of inst : label is "34B98B604921396D7492484E5B5D24921396D74B19649213AE98150AA160542A";
    attribute INIT_04 of inst : label is "2CD8550131152B5ED4ADBB65D905042045D8DAC5B56EA5128001308E8804C024";
    attribute INIT_05 of inst : label is "49965145D265945145102886596CDB592D6CDB592C4F4922A66ECDBB09257162";
    attribute INIT_06 of inst : label is "0804008048402CA08D5430182024178C4E260980D62859A06A81A62003D0AC57";
    attribute INIT_07 of inst : label is "304D852C65B264092803348094AC3168B5E8A8609422809422A896D00B0100A0";
    attribute INIT_08 of inst : label is "41240B094B54751A75D521A68308924D39125A665A431CE48A60491625523219";
    attribute INIT_09 of inst : label is "5B801B102D884724CEAF5E836DABD52C14B29D1E19261649294C49253550994A";
    attribute INIT_0A of inst : label is "69730313ACBC92AB56BA18E4910AD0AD0AD20D41490305B3490268224035B495";
    attribute INIT_0B of inst : label is "41412AAC04AA4924B380781858306039B35821B2C6B016B602A07793322FC1E6";
    attribute INIT_0C of inst : label is "2E758FD75749E54D9B473A2303025FF7FFFFE40BF7FF0581FDFDFFFF30541505";
    attribute INIT_0D of inst : label is "B6A8FA492CB783105A83E72C0A620A582988295DFBFFB1A50BE4A371B8DC6E94";
    attribute INIT_0E of inst : label is "000480CC786A7C24027C27427427427C0C845ED6B453744F913E64D993761148";
    attribute INIT_0F of inst : label is "0009F45A8B4492492F57AD5E8B68822A008A0284303906C9804816356C61AB32";
    attribute INIT_10 of inst : label is "2498CDC62C41179C26B5A86A8EA16BD39DCA93249174CC022F38480401000040";
    attribute INIT_11 of inst : label is "A4D5AAA552A7505D798222E82E90084F396DF72F32C1700685D7BF3D98BC3979";
    attribute INIT_12 of inst : label is "08C9B6DEB56A2D2D9CDCDCA5A44675E63B33CD35894A7206AD54E40D5A7BCA47";
    attribute INIT_13 of inst : label is "FB55B725B6C492F2F5A9691105F75A41C60CE072C14AB144B144EB52083C94A5";
    attribute INIT_14 of inst : label is "417D0C54DE09CEE739DE77D56DBFEFFDAC0E67B3DBEBEDA82AEFB96DF65AB1BB";
    attribute INIT_15 of inst : label is "000885A400030EEC000606700002262000012300000060800000FF00231650B1";
    attribute INIT_16 of inst : label is "000F44300013A6640002AB840010298400183C04001F907C000386380000C38C";
    attribute INIT_17 of inst : label is "88A22222888A029A69A69A69A69BF47C4000EF800003E7600007A670000A2618";
    attribute INIT_18 of inst : label is "5FF9A4D5572BAD78499026F48D42854D6A431312079A6888A22288888A222228";
    attribute INIT_19 of inst : label is "302533C08485294A234AE42108895C9CCDDC8D049084DD9A5420529488CD290F";
    attribute INIT_1A of inst : label is "03803001B890E6E00080D07368A0D6D8E70C436DB64086DB6C804494FF261B80";
    attribute INIT_1B of inst : label is "8C5CAED48851624509200188B082100912243861C300140070A913801A211C48";
    attribute INIT_1C of inst : label is "91CA4EA104221014B0024891016260854B8908AC01C2311D2E114024B128254B";
    attribute INIT_1D of inst : label is "68847305CD3662C5EB02BD56490D588005083C08E01000000000012C60168214";
    attribute INIT_1E of inst : label is "F0CF117023C2A420B5149B7038B81B7D3038B81D908E220EC40985CE645592A6";
    attribute INIT_1F of inst : label is "55EA017CE40EB37A4E6927337A4E69273A4C71121A10E8AAA9119551027B399E";
    attribute INIT_20 of inst : label is "0743C78D1E3C78F01F009AA297AF5912AAA5ACCB5DA58B4B157FD5FF55F802A9";
    attribute INIT_21 of inst : label is "8D8010008040100952AD589122C58099007AF41F0356AD41D03D7A0E868F1A34";
    attribute INIT_22 of inst : label is "B6B6E415598C63806C0454440800001A000A800C02A2000DE980012AA1190000";
    attribute INIT_23 of inst : label is "F003FF001FE007FE007F599B9B331B3733666266E66CCC5555119ACAC9635AD6";
    attribute INIT_24 of inst : label is "2755904D3E999CB26AA067934DE6E62CAAA6493A16C11608821AB00001FF801F";
    attribute INIT_25 of inst : label is "6C0932838849C446A7EEA25B2ADA91CF0104C7A4CE72D540CF26372E639554C9";
    attribute INIT_26 of inst : label is "042C032DF31DD574D20E944C2837142163C03FFFF8A2E914551BB443A6D11102";
    attribute INIT_27 of inst : label is "101EE0F6C684347B8A3DA884143BE307702B2760EE0567D0850042A500A47BB5";
    attribute INIT_28 of inst : label is "F3A9CF63453F4C635B858D03721637366B9166BCCC76C6CF7B618C59BAE60C3A";
    attribute INIT_29 of inst : label is "00000000000055550000756342D79D4DE7B1A1FB63B95E3A9CF6343F6C626332";
    attribute INIT_2A of inst : label is "00042118C631CA529084214E73884214E218821031A10D1F3457F455FC7EC000";
    attribute INIT_2B of inst : label is "5B78D959322C582275D9A04C814A522334A51079FFA209B6DB654A5290840000";
    attribute INIT_2C of inst : label is "E5BF70775B9D99BC0909F88E60C8CCDAB25327892669010C0B34A841A4F5FFAF";
    attribute INIT_2D of inst : label is "0FBBDFEFAFEFFE33CB18CCDF9446D1D1D1C2A9176EEDBB62FBFC7EF73C00CF0E";
    attribute INIT_2E of inst : label is "CA4893999332A954E952130679894D4A8927A23693A88DBFFABBD9BD99FFAD29";
    attribute INIT_2F of inst : label is "324977F56FEEEEAABA7AAD12918D610A6CC9FFC6797D63EB2C18328102281022";
    attribute INIT_30 of inst : label is "DAD6C3CBB55DF3E626EB8CC077CF9D084EB1BED16399DDCF9ADFFD1CC972E4AB";
    attribute INIT_31 of inst : label is "662E161EA3A9299BEE6230B90CFFC7F8D0267678A31518B8C58E6A55B98FC201";
    attribute INIT_32 of inst : label is "F73420A25128E3109B089A33277776310007FFC62CBEB2A372E4ECC9884D7967";
    attribute INIT_33 of inst : label is "4598330640C819833086B5AAEF7F55A5080751B0E8069D84F20F7726E67D2120";
    attribute INIT_34 of inst : label is "D9EC9B888110220441E1E1A1E301C69C9C1E1ECBC2922826A1B63906C925BC4B";
    attribute INIT_35 of inst : label is "DB44C9338416364B1BAE53679490C4B2C2EAA5AD7A44460005A0046F99F7ED8E";
    attribute INIT_36 of inst : label is "0466DC952CFB4F5C6C4846CB8F5EB5604A222764B96DB25B25A66DB6DB44A9B6";
    attribute INIT_37 of inst : label is "3689D1B275C6C4866CAFBE0477DF7E7F24DCEDC35B44E70B0F4B0BA0A8793D05";
    attribute INIT_38 of inst : label is "BEBEEFEEFAAAAFEAEAAAAE1A4CB2B6AED8A959184619774C961C170D6A58B113";
    attribute INIT_39 of inst : label is "511114804020100804020100817757575441490410059142C091966BBABFFFFB";
    attribute INIT_3A of inst : label is "1207D00208165008205D4420555C40200BABA080040208041040208151D01000";
    attribute INIT_3B of inst : label is "A9020175200105840F2FABA8040223E5F502E81640F805D43E81E12B287D42C0";
    attribute INIT_3C of inst : label is "AA8103EBAA4002AA800116D00043C2081E1040EA004103820423C800BA84801A";
    attribute INIT_3D of inst : label is "4240FA8041024102E83C208200F3AA80402410071D560200AAD484102CA21040";
    attribute INIT_3E of inst : label is "26810075082C0416120010580208207440240EA900082C3521040E21821B0714";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA555580804D0200E0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA5557AEAA5555AAAA7559F366520821139526022E7850A8A85050A8A1";
    attribute INIT_01 of inst : label is "C9424AAACD48220E6615C4DD4B070000048449470511A62297264808924C16F3";
    attribute INIT_02 of inst : label is "8A051342281422010220142201422020005A4B016392A6106984984902D168B4";
    attribute INIT_03 of inst : label is "BB991A80492CB5616D924B2D585B6492CB5616D9DD6492CB6DB05134228144D0";
    attribute INIT_04 of inst : label is "3CCB5DB13B110BDEC425BB75DB8C108555DADED5B56EE59699513A88ED44AA28";
    attribute INIT_05 of inst : label is "5B24924916C92492451428A2496ED9936F6ED9936CCF5B76AB3567B96B2D79AF";
    attribute INIT_06 of inst : label is "70420F042182100202173252240833286C2489189EA8FAA268B1A74003CA8D64";
    attribute INIT_07 of inst : label is "18CC0CAD0806709B6A001040BA6D3B61AD802880021047021000368084020840";
    attribute INIT_08 of inst : label is "D1A40B0DE812411AF59561C2CA28B2CD7956DAD25C5210A58B924B166502B69C";
    attribute INIT_09 of inst : label is "DA0202106DCA4F6E482040802408936834B690440B2D36FB6BDCD92535519B5A";
    attribute INIT_0A of inst : label is "656241013AB4D020488000E59812C12C12C34D014B890C120B47604AC235B009";
    attribute INIT_0B of inst : label is "01C81388004EDB6D9288301050A14229E258488010B01EB48390779F323F83F5";
    attribute INIT_0C of inst : label is "2057AD77554D65CD9B47BC204C114FE7FFCFF869E7FFF4A3F9FCFE7F68701C07";
    attribute INIT_0D of inst : label is "B024824B2EB722965293C76C1A624AD269892B19F3FFB1871840A30180C0601C";
    attribute INIT_0E of inst : label is "E03E1A42706A402D0A482482402402402AA55A9084C20108042030A442835D48";
    attribute INIT_0F of inst : label is "008B41124AC0C3041480020000248AAA20A0A82431250E11A3E0E4176824BB3C";
    attribute INIT_10 of inst : label is "2D942DA668C2141834A5280249234B161DAFF36FB34581842830601008000200";
    attribute INIT_11 of inst : label is "2D10210272AC4175418AAAC43AB0AB041164922C3285E6971754A83014B00B1B";
    attribute INIT_12 of inst : label is "2AAFB24481022D648C5C4C6CAC6455062A220D65995A93048109260922800A55";
    attribute INIT_13 of inst : label is "8A77A448048900A2A5294888954AD2C19638B4F6C004E9DC89DDCA5288888020";
    attribute INIT_14 of inst : label is "4405A28241E9EE108421575F4DAFEB9D3A0462B15AAAE9243AAFA54D7456A112";
    attribute INIT_15 of inst : label is "FFE4F99FFFEBFB6FFFF3BAAFFFFBFFFFFFF87F7FFFFE9FFFFFFFFF7FD11ED1F7";
    attribute INIT_16 of inst : label is "FFFAC9EFFFF763FFFFE1BFCFFFFE1FB7FFFBD907FFFF687FFFFC1807FFEFBCF7";
    attribute INIT_17 of inst : label is "00000000000000000000000000028E72BFFFE87FFFFD689FFFFBBA8FFFF1FBE7";
    attribute INIT_18 of inst : label is "549193FFCE29E53BF9A9A6FEC118C7C95B829395170000000000000000000000";
    attribute INIT_19 of inst : label is "9031A2045B461184AAD7284612AAE124CDDC0B126AD69DE4140000002AAD7225";
    attribute INIT_1A of inst : label is "FFFDC4187C0411E08241000410D004E29505232CB3224659664585D89C400D1A";
    attribute INIT_1B of inst : label is "003C10200220000002002400000C442060010317EC5021428100042840007E06";
    attribute INIT_1C of inst : label is "221001108800A220040481205000F110041200108200024200A4200040801204";
    attribute INIT_1D of inst : label is "048A406D0DB076864902C917D9802040881000300200003FFFFFF09004812000";
    attribute INIT_1E of inst : label is "CACC115922C2AC0924549245608A124925608A12CC88208E45188D0D2865B600";
    attribute INIT_1F of inst : label is "0000ABFC8C4002489060483248906048364A133251287E6E891511514202318A";
    attribute INIT_20 of inst : label is "64800102000810019209048311204983DDFAAEDB5DF093E115557FFF5557FFFC";
    attribute INIT_21 of inst : label is "3020021810108FE40C103060818209140200219010800219010010C801000008";
    attribute INIT_22 of inst : label is "92B6CE355BDEF7D76FF54444021C000043E00010F80023F00010FE0008620008";
    attribute INIT_23 of inst : label is "0003FFFFE00007FFFF805511122222A222444C5444488891115556DAD9515A56";
    attribute INIT_24 of inst : label is "23DC9844239590F3EAB5271108A5E43CAAF2511ED2611308A6ACC00001FFFFE0";
    attribute INIT_25 of inst : label is "645A13198C29DEC6972CA2DB8ADA91CE01844464C852D56A4E22212E42955E4A";
    attribute INIT_26 of inst : label is "E72B4228832D942DB62D342A6836943583FFC00000E3E91C75173EA367444456";
    attribute INIT_27 of inst : label is "C1508284D53055421AA1000000252B1A552F04A14AA4E5CF8CF0E5EACCE75022";
    attribute INIT_28 of inst : label is "EB2F457FF5FF7A655125FFC225A4A2A6AA557AA8EE24CA9CA540295132552A55";
    attribute INIT_29 of inst : label is "00000000FFFFFFFFAAA4D77FF297597922BFF92BE92F5D72F457FF257D23D32A";
    attribute INIT_2A of inst : label is "2108421084214E7398C6318C630E739CE210C210354C15521542A595248A8000";
    attribute INIT_2B of inst : label is "0A529DF732ACDC1E6DBE4840800000AAB5AE74AB493798924927CE7398C61084";
    attribute INIT_2C of inst : label is "956F4054D1151114D1CB468436CEDECAE673A7D5AE0B017EABC828005955493A";
    attribute INIT_2D of inst : label is "8BEF954A6A2AAE2B8B1955453550D89A909555D564EDB96EABA82E973FD2FA8A";
    attribute INIT_2E of inst : label is "5B5A95FFFFF72E65DA5E56A712918E5ACB222A82B12AA1DDDE1A9DA99AA8E739";
    attribute INIT_2F of inst : label is "224935FF5E777733327F182318C6339EFFD955C5717C43E2489124C993489123";
    attribute INIT_30 of inst : label is "56B5E9533719F2E4B54F8CD167CB92AD54E1AE89D111654A10F42D086D7A74AE";
    attribute INIT_31 of inst : label is "67AD1C0492496483E8702491CCF9C5F8882AAEECE49C64E1278C72D7BFE9C201";
    attribute INIT_32 of inst : label is "7EA404E476394210922A9000000004210004248059B2B4E1B2D6ECCB88ED7B77";
    attribute INIT_33 of inst : label is "2184308610C2184308C633AA8C63556F3C3C44B1C228BC96C056EFA6E6790605";
    attribute INIT_34 of inst : label is "11010BCC4188310620808080C211860E0E0C0A098608400080A2ADACC048D850";
    attribute INIT_35 of inst : label is "D3E969B58E2424DA5B5489636922846F8673C5AD62C00A004B944225F5F30000";
    attribute INIT_36 of inst : label is "0323A9136CBA0A5648904482CB54A23290A54817134926D26D444D34D3EDF134";
    attribute INIT_37 of inst : label is "27D2D124B5448906492B248CC5925E5F012CA28193E94B1207122384653919A3";
    attribute INIT_38 of inst : label is "BBAEFAAFABEEBBFEFFBFBF18AC52B66D109B93334CD65A2E641C0A0CF6972D33";
    attribute INIT_39 of inst : label is "00000080402010080402010081D747474451090410075152A8B31D6BBEBAAABF";
    attribute INIT_3A of inst : label is "1A078442081D510820594020785944200B2B00220512080410402081E5641111";
    attribute INIT_3B of inst : label is "890201F1200905040B2BAB28844201656502C01F50B205803CA5E50F885D42C8";
    attribute INIT_3C of inst : label is "AA8103EBFA4010AA80011E100042A208361041B2084106A20423C8042C84812A";
    attribute INIT_3D of inst : label is "0240F88041024103A03C208200EBA28840241007DD164200A2D4041038201040";
    attribute INIT_3E of inst : label is "26011079483C241F1200907D0208205040240F090048283501040F0190130504";
    attribute INIT_3F of inst : label is "5557AABA5D55AAAA5555AAAAD555AAAA5545AAAA5555AAAA555580804C0220A0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "57DDAEEA5D57BAAA7555AAAA557BE9F999659259C31A67C73E53A9A95353A9A2";
    attribute INIT_01 of inst : label is "241D2023A3306CB99CDB44064331225DB6F33472703E90B84C91216E4930CDF9";
    attribute INIT_02 of inst : label is "A030340680C2688C2688C6688C26899259716E2DC448391C8E47A324BB8DC6E2";
    attribute INIT_03 of inst : label is "3415C3E12486E1CDC34921B87370D2486E1CDC3499D2486E18630340680C0D01";
    attribute INIT_04 of inst : label is "60DEA35EDDECE425319614C33639C210473311A760591A4C663EC9F110FB67DA";
    attribute INIT_05 of inst : label is "80BAEBAEA02CB2CB38E7C73DB664DB692D64DB492F7AB6CC626A4C1BD6BAD346";
    attribute INIT_06 of inst : label is "0FBDE0FBDC7DEF82BDD0E937D26B091A3D0DF74F520A4929C01E18300EC39CD2";
    attribute INIT_07 of inst : label is "883A1238B259C2C6C165D96E6398E0C70333837EFDEFB0FDEFF9081F7BF9F7BF";
    attribute INIT_08 of inst : label is "9C522E1846B32B71AB51CF0965976BB8D51C3589734A52B7168B64EDD09AFC71";
    attribute INIT_09 of inst : label is "70D92D8CDA2338D96548911CB712A0D662FC4A91BEB9EB868432F4D08AAF6675";
    attribute INIT_0A of inst : label is "79C1811868E700C18B13661345CB9CB9CB9E782E362DB2DE767CC5C58BE362C3";
    attribute INIT_0B of inst : label is "236D869A161B24DB48F014346C1830872AB416D9016DCE3B080121C0898709C4";
    attribute INIT_0C of inst : label is "81018C446660536DDB37399F23C827EFFFDFE344EFFFF215F8FC7E3F0CD2348D";
    attribute INIT_0D of inst : label is "6D664636982CCDEBAC66CC18319DF5ACC677D688F7FFB59D60382C0603018075";
    attribute INIT_0E of inst : label is "24371041D4C12B5B312B12B12312B12B0894B3E739D89262498926249892112B";
    attribute INIT_0F of inst : label is "0066235626479C79C23468912D925F57DF5F7DD028440D35AF702D097A004BE5";
    attribute INIT_10 of inst : label is "B8423D9DC12DD6718D18C656646E2E6CF3308E186E0B12DBACE3000000000000";
    attribute INIT_11 of inst : label is "DBF2E5B8D859E6866702238669685AB6DDD2CBB9FAE1E15D2866CCE6D6E2EE2E";
    attribute INIT_12 of inst : label is "088C6B712244BAD6F33322025B03699D11113AD77431DE03972FBC070EC02145";
    attribute INIT_13 of inst : label is "EB31B66DB6CDB73AD8C6300001621D838D07A7AC3061AF470F46318C80630C62";
    attribute INIT_14 of inst : label is "5006A18B6005CE21084211336DBFCFBDEB233118888BED966CC7B16DF75CB88C";
    attribute INIT_15 of inst : label is "001E491C00180204000C20080004011000074070000163400000FF001DF25490";
    attribute INIT_16 of inst : label is "000001180004201400193F6C0010198400105B0400007804001FA0040011C4C4";
    attribute INIT_17 of inst : label is "000000000000000000000000000285F18000018000000340000000F000004010";
    attribute INIT_18 of inst : label is "16DF48D5668CC4356F5E8D942631B936CE1CEDEB5D0000000000000000000000";
    attribute INIT_19 of inst : label is "D8436022763DCE7A223F9F39E88FF3E44554193BCDB85AE044010842088ED676";
    attribute INIT_1A of inst : label is "00003BE383F3EE0F7D9EFDFBEFD400459107C6DB6DC70924930F13719C010D4F";
    attribute INIT_1B of inst : label is "EFC1EFDFBDDF7F7DF9F799FBF7E39B9F1EFCF8E0038F9E3C7CFBF3C79FBF01F8";
    attribute INIT_1C of inst : label is "DDEFDEEF77BF5DDFBBFB6EDFAF7F0EEDFBEDFBEF7DDFFDBDEF5BDFF7BF7BEDFB";
    attribute INIT_1D of inst : label is "0A2F18183BEBCC3D1981A35C343FDFBB77EFBFCFFBDEF7800000076F7B7EDFBF";
    attribute INIT_1E of inst : label is "C38DC4D180C85355BABA0B6B2E19CB658B2E19CDAA6188A5B30F1839B7174D1B";
    attribute INIT_1F of inst : label is "55555403823B9B68D9C06CEB68D9C06CE3B1098DFFA6E046604848AC3805EF75";
    attribute INIT_20 of inst : label is "12B6B468D1AB56AC4ADC310C0C68CF00A09DB9141722E645D5555555FFFFFFFD";
    attribute INIT_21 of inst : label is "CFDEFDE7EF6F7018952A448912A54C0A8DD68C4ACE346AC4ACEB46246C68D1AB";
    attribute INIT_22 of inst : label is "684C58E876B5ADA8D9F000007DE3FF7FBC1FEFEF07FBDC0FEFEF01FBF79DFDF7";
    attribute INIT_23 of inst : label is "0003FFFFFFFFF8000000C8888B11D11111623222222C4640001111B1B41E210C";
    attribute INIT_24 of inst : label is "DC7367B8C9E1E70C3823DB6EB33AF9D360AD96E36D9EECF749CF00FFFE000000";
    attribute INIT_25 of inst : label is "1BCDE87661DEF47B6CBAFC3600B0E1CE0E7BB9FAF3AD7047B6DDCDDF9D6C15B2";
    attribute INIT_26 of inst : label is "38CC91AC4EBFD297739C8C19186E4439FC00000006185CC301C10459136AAAB3";
    attribute INIT_27 of inst : label is "4FC2DE17A353CF0B678580000062033172D99C502E5A37C0FC0FD8B032949CB1";
    attribute INIT_28 of inst : label is "652762DB0C1B39D998DB6C311E7618180B11C33ACD96E2C631708C591163068C";
    attribute INIT_29 of inst : label is "00000000555555550009DEDB0CF32938B16D85B92107CC12762DB0B72421CEB6";
    attribute INIT_2A of inst : label is "318C6318C6318C631CE739CE738C6318C318C21068D4F3C6CF1BB045B022C000";
    attribute INIT_2B of inst : label is "AB98DA1CEA3B8449C70E0A02842108223B5ADE306DFC3E4924918C631CE718C6";
    attribute INIT_2C of inst : label is "C58F6E33588C88896D68716319F1E3F59B5A469259B6ABED55C0880253616DC3";
    attribute INIT_2D of inst : label is "6C9DD679B9F99EB931CCCCF2670326646444711623F37CC4B1931EC8BC2B8362";
    attribute INIT_2E of inst : label is "7470C911111D59B70EB31C318C652B75A291B819488E0655513668E688CE94A5";
    attribute INIT_2F of inst : label is "A249A7F46B155511117A265AD6B5AD69447733D7263D79EBB76EDB76EDB76EDC";
    attribute INIT_30 of inst : label is "DAD6D5891D8CF3E7687AEECDC3CF9D5A87ADBEEF5888B5B36EC712C632851B59";
    attribute INIT_31 of inst : label is "DC39C531991AD689ED87D846267BD7FAECB32387BAF497A4BD6B5BADBFEFD305";
    attribute INIT_32 of inst : label is "F21813BBD9ECB18C6D88980000000318C00CB6C1231331A5ACCC1BAE7798D0C0";
    attribute INIT_33 of inst : label is "DC7B8F71EE3DC7B8F73631998C63332E64278D8E06CB0EF5A10F264A48B61210";
    attribute INIT_34 of inst : label is "EEFEE153BA774EE9DF5B5B5B1A3EA1E1E1E1E374C000410B221819035B6E2B2B";
    attribute INIT_35 of inst : label is "DBED92CE4079B6DB5AF9F67D55B3647023BFF7528580002DFFF33D6D1B60FFFF";
    attribute INIT_36 of inst : label is "7CDDF3BD9104C59B6CD832CB659939CEDB676D2ADB6DB6DB6F236DB6DBEDFDB6";
    attribute INIT_37 of inst : label is "B7DB65B6D996CD832C84B7BFC25B14946DB66F66DBEDBC9D989CDD4F98D0E67C";
    attribute INIT_38 of inst : label is "411155500110510051101127432493A485EFE44791F17185BB1B358F7F5EBE45";
    attribute INIT_39 of inst : label is "0000008040201008040201008084A0A0A0100904100280014033035440100415";
    attribute INIT_3A of inst : label is "12028402080A1008202544200108442001010208100208041040208090804111";
    attribute INIT_3B of inst : label is "090220A5200082C400000008040220303500480B005082C006803001800D0062";
    attribute INIT_3C of inst : label is "088101495A4002508001015000400A080A5040500841014A0420280080048100";
    attribute INIT_3D of inst : label is "0240528041024101401020820048508840241002C286020050CCC41001221040";
    attribute INIT_3E of inst : label is "2201102D04020200120008010208200540240509000416333104004910120000";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555808044022000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "5555AAAA5555AAAA5555AAAA555AD1E00B6D92D9A7022D06BE51A9A95353ABA3";
    attribute INIT_01 of inst : label is "400E00228710E4A290DC4007422322CC9242382A286881B4000201240085A4B1";
    attribute INIT_02 of inst : label is "8220704E0886E0086E0082E0082E01B6D9536A6D4C8030180C0681249A8D46A2";
    attribute INIT_03 of inst : label is "240489E12482A145444920A8515112482A1454449952482A28820704E0881C13";
    attribute INIT_04 of inst : label is "409080480C88C0042314301000218000451312850040080000681B4001A06D18";
    attribute INIT_05 of inst : label is "C9208208B248208221870C30002E4903652E4903646AC0104642C81218A34202";
    attribute INIT_06 of inst : label is "0000000000000002B8148B351660151A3D0D474414085021000C111008439CCA";
    attribute INIT_07 of inst : label is "9828322892CB1248016DDB2C09A1A90C04170000000000000060100000000000";
    attribute INIT_08 of inst : label is "08E22A10060320402C510D4B6DB78A201510460B515A56B4329964F1009A7045";
    attribute INIT_09 of inst : label is "50596C840852A0036408101DB342011202F0CA50A8A08A08420282404AA82646";
    attribute INIT_0A of inst : label is "5150810C28A60085020364000D8A98A98A9A68277864B25E383144C61BA10261";
    attribute INIT_0B of inst : label is "2164D29A134A920000C01434640810056AC632C9858DCC290000210900061984";
    attribute INIT_0C of inst : label is "9401084444444164C97211BF6BDA612922525B0C2912F6304E271389C4521485";
    attribute INIT_0D of inst : label is "AC0640788A24418A242240200031462400C51888948914B5351026A351A8D4D4";
    attribute INIT_0E of inst : label is "2403004354432963132932932132932908B5D3C631C800200080020008001129";
    attribute INIT_0F of inst : label is "FFC2A15226061A61AA040850AC9208222882883008640935A4312D0D3A0069AD";
    attribute INIT_10 of inst : label is "A0833CB5036DD2D31D08424064082A30513A0A20881C365BA5A62FF7F9FFFE7F";
    attribute INIT_11 of inst : label is "E3C081985060AEA72D022282298808B2CD5249A9CA40A9556872E5A256A6E828";
    attribute INIT_12 of inst : label is "08892B342850AB165212020462232CB591916B154001D802040FB00428D08144";
    attribute INIT_13 of inst : label is "693112249244939A4842100001224E02A50286201030A54405441084806A8420";
    attribute INIT_14 of inst : label is "4003808B6004842108421111249244A4A9223118899924922E4491249348988E";
    attribute INIT_15 of inst : label is "001980CC00171874000E5128000C37180007B6F0000377600000FF801DF410A0";
    attribute INIT_16 of inst : label is "000E3238001B1E6C001CC09C0001D04400000404001F087C0000000000100404";
    attribute INIT_17 of inst : label is "000000000000000000000000000280E48000FF800003F7E000076370000E6238";
    attribute INIT_18 of inst : label is "124B00400688C434056A85A40200A342C291818AD50000000000000000000000";
    attribute INIT_19 of inst : label is "D80069276371AD6A227FBE31888FF7E44444183906B8536044C00000088B1672";
    attribute INIT_1A of inst : label is "00000000000000000000000001CE420582070000010684924A8D01518C010D4F";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "012A98006BA9103101802050408000000000000003DEF7800000000000000000";
    attribute INIT_1E of inst : label is "428CAA55418073D492AC092A0D00A92D4A0D00A8A91148A209040068B634500B";
    attribute INIT_1F of inst : label is "FFFFFFFF843B19284B4025A9284B4025A1C31891652EAA0224A4A42A14048420";
    attribute INIT_20 of inst : label is "32960408102850A0CA58348A0D2A4D0000B8EA101502E205D555555555555557";
    attribute INIT_21 of inst : label is "000000000000001A50A142850A952A0A4CD0A0CA4E040A0CA4E850642D0A1420";
    attribute INIT_22 of inst : label is "24204080500000AA0A0000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "FFFC0000000000000000888889111911112223222224444000111280800A1080";
    attribute INIT_24 of inst : label is "0024060009830410482903800220410420801801701800C059F000FFFFFFFFFF";
    attribute INIT_25 of inst : label is "204484C05310822200A2D04080808FC0086021E38231905207010D1411841003";
    attribute INIT_26 of inst : label is "3DE491A45ABFD39771D45818B06A083E0000000005144AA281A91004292AAAA0";
    attribute INIT_27 of inst : label is "4F465A33B113C519628C8000006382133A9A9C606752528448448A111294C990";
    attribute INIT_28 of inst : label is "6627624148293B41C8C905311EF230300911439BD89FA64A73209CC911310204";
    attribute INIT_29 of inst : label is "00000000555555550009DE414E733138B120A4914107CC22762414922821DA9E";
    attribute INIT_2A of inst : label is "42108421084210842108421084318C631CE73DEFEC44F14CC539186C98364000";
    attribute INIT_2B of inst : label is "A9C8D34CAA2A0C0942160A09000000222C62CE1124B13C000002000000002108";
    attribute INIT_2C of inst : label is "44892F33C88C888B656933631BC3C3C4895A62166198018516C08980532124E9";
    attribute INIT_2D of inst : label is "2CCCD239F9B99291718C4462E5062C6C6C4451122321484091171240942A8922";
    attribute INIT_2E of inst : label is "4440A111111149B4469110298C6D6B449251A831888A0C4443666CE6886694A5";
    attribute INIT_2F of inst : label is "DDB6825423111111112A725AD6B5AD6B444732522E253129972E5972E5972E5C";
    attribute INIT_30 of inst : label is "8842548115889932282A66454264C80A82A49265488894996E9312C633061C48";
    attribute INIT_31 of inst : label is "44288D301903128125A048C6844A524A64A22222A25412A095295A25B989C214";
    attribute INIT_32 of inst : label is "540802A351A890842488880000000108400C924038139025A65E48A836205152";
    attribute INIT_33 of inst : label is "0000000000000000002421088842110EEC269D884E0116F0A005425C49D20200";
    attribute INIT_34 of inst : label is "1101114000000000034343434268A3535353533A840040092134391989256808";
    attribute INIT_35 of inst : label is "49E492CE463992494AF9D2255493207B229FF5630600003FBFF1152553B00110";
    attribute INIT_36 of inst : label is "F545F395318644CB2448125924CB955E4A47250AC92492492723249249E4FC92";
    attribute INIT_37 of inst : label is "93C924924C9244832585928882C939B824924722C9E49C9C889DF04E88482254";
    attribute INIT_38 of inst : label is "54405400011551550544142442A5B2A484AFC4459171208EB90914855F4A9644";
    attribute INIT_39 of inst : label is "00011080402010080402010080A0000000000904100040002033000501405040";
    attribute INIT_3A of inst : label is "1202C402080A1008202C04202820402004040000000208041040208010101111";
    attribute INIT_3B of inst : label is "090020B1200882C4058505080400208091010003001800C004003001800C0060";
    attribute INIT_3C of inst : label is "088101414240105880230A100041420800104000804100020060200400048000";
    attribute INIT_3D of inst : label is "024050804102410140142082001800804024100040060200004C441002201040";
    attribute INIT_3E of inst : label is "2201002C4416220B1200882C0208202C40240009004402131104008800120004";
    attribute INIT_3F of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555808044020000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
