-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_7M is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_7M is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_7M_0 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"2A8A2FFFA000F80002AA2FFFA000F8000B8000AA2E00800002A802FFAA00E800",
		INIT_02 => x"00AA002F82A8FFF8000A002FA2A8FFF8000A002FAA80FFF82A822FFFAA00F800",
		INIT_03 => x"00000F0C00000F000000003F0000FF00002A0F3C80000F00002A0F3CAA000F3C",
		INIT_04 => x"00000F0C00000F000000003F0000F000002A0F3C80000F00002A0F3CAA00003C",
		INIT_05 => x"00000F0C00000F000000003F0000FA00002A0F3C80000F00002A0F3CAA000A3C",
		INIT_06 => x"0000005200002000000002FB0000BE0000000B40000007800000014000000500",
		INIT_07 => x"0000000800008500000000020000200000000002000020000000001200002000",
		INIT_08 => x"00280700A0000340000000080000800000000008000080000000000800008400",
		INIT_09 => x"002A00E1000085000000010002801BD000000052A8000B00002801A0A0002900",
		INIT_0A => x"00000EBF0000FF1C00000E3F0020FFFC00000EBF0003FE1F028007E4000000C0",
		INIT_0B => x"000003EF0008FFCC0000303C000000030000203C800000020000003CC0000000",
		INIT_0C => x"00000B400000078000000000000035500000014000000500200033FF0000FBC0",
		INIT_0D => x"20823D7F0800F40000003FFF0000FFE007D43E971700D2A000003E970000D2A0",
		INIT_0E => x"002A0265A200AE00002A0206A880FC00002A026FA220F600002A026DA8886B00",
		INIT_0F => x"00000FEF0000BFF0000000000000000000000A820000C0000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"000001FF0000FD000080047F0800F440000007FF0000FF4000000B4000000780",
		INIT_13 => x"000000000000000000003FFF0000FFC00000000000000000002A0380A0000B00",
		INIT_14 => x"002507FF6000FC00002503FF6000FC00002517FF6000FC00002557FF6000FC00",
		INIT_15 => x"000000BA0000B000000000830000AB000000008000003AB000001080000003A0",
		INIT_16 => x"00001080000003A000000B800000003000001AB000000004000003AB00000000",
		INIT_17 => x"00003F0000000FC000003FC000003FC000003FE00000BFC000003FF80000FFC0",
		INIT_18 => x"00000AAA0000AA8000000AAA0000AA8000000AAA0000AA8000000AAA0000AA80",
		INIT_19 => x"00003FE000002FC0000000000000000000000AAA0000AA0000000AAA0000A800",
		INIT_1A => x"00003FD000001FC0000020BF0000FE000002003F8000F000000035FE0000FD58",
		INIT_1B => x"00003C000000FFE800083D070000FFE800023F7F0000FBD400083FE000000FD8",
		INIT_1C => x"000000FE0000FFFF0000007F0000FFFF0000007F0000FFFF0000003C0000FFFF",
		INIT_1D => x"00003CFF0000FFFF000000FF0000FFFF00003CFF0000FFFF000000FE0000FFFF",
		INIT_1E => x"0000FFFF0000FFFF00007FFF0000FFFF00007FFF0000FFFF00003C7F0000FFFF",
		INIT_1F => x"000044FE00000000000044FD000000000000447F000000000000447F00000000",
		INIT_20 => x"00000000000000C000550009054F00030000030000000000F150C00055006000",
		INIT_21 => x"0000000000026181150500004000010380000249000000000000C04054540000",
		INIT_22 => x"20005000800300005450000900000000C0030000000800140000000005156000",
		INIT_23 => x"20005000800300005400000000000000C0030000000800140000000000150000",
		INIT_24 => x"00000000000003AF00000000007E00000000FEB000000000EF40000000000000",
		INIT_25 => x"00000000000003AF00000000003E00000000FEB000000000EF00000000000000",
		INIT_26 => x"00000000000007FD0000000001E300020000DFF400000000F2D0A00000000000",
		INIT_27 => x"00000000000007FD0000003F00BF80020000DFF4000000007F80A0000000BF00",
		INIT_28 => x"33FF33FFFF00000033FF33FFFE3FFFFF0000000000000BFFFFFFFFFFFF54FFFF",
		INIT_29 => x"33FF33FCFFFF000133FC33FF0000E3FFFFFF557FFFFFFFFF0000FC0200001FFF",
		INIT_2A => x"0000FFE000003FAA02BFFFFFD000FFFF00000000BFFF000000170388F3F41EAF",
		INIT_2B => x"FFFFFFFFFFFFFFFF0000F00000000000FFFFFFFFFFFFFFFF00000000000C3501",
		INIT_2C => x"00002D5E000002E000000B5F00003C0F00003D540000F2F400003C0F00003D54",
		INIT_2D => x"000BFF40FFFF0000FF007FF800000000FFFF0000E00001FF0000000000FF2FFD",
		INIT_2E => x"00000000FFFFFFFF00000000FFFF00000000000000000000FFFF0000FFFF0000",
		INIT_2F => x"0000000000000000FFFF0000FFFF0000FFFFFFFF00000000FFFF000000000000",
		INIT_30 => x"000000000000FFFF00000000FFFFFFFF0000FFFF0000FFFF0000000000000000",
		INIT_31 => x"0000FFFF0000FFFF00000000000000000000FFFF00000000FFFFFFFF00000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"FF542C01002F400002BFFFFFF1F0FFFFC030B000BD2380000028FFFF402FFFFF",
		INIT_35 => x"FFFFFFFFC07FFFFF0000500000000000F805FFFF0FFFFFFF0AAA007FA0005400",
		INIT_36 => x"4CCF002084BFFF00C0FCFFFF02FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_37 => x"E103FFCCCB00D2D0033A34C8EB55A0800BC00315008F00030000AAAA0AA8BFFF",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_39 => x"510087F10000FF54FFFCFFFF087FFFFF31CB01FD3FFF0000FFFFFFFFE07FFFFF",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCCFFCCFFFFFFFFFFCCFFCC",
		INIT_3B => x"CBFF0000FC2F0000FF80FFFF8FFFFFFFFFFF1FFFFFCCFFCCF800FFFF7FCCFFCC",
		INIT_3C => x"000000000000001F002F00007FFF77FF8000800000000000F8009D0000000000",
		INIT_3D => x"00000000000000000000000000B4000000000000000000007000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000040100000004040000080000000008000010000000008001001000100000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7M_1 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"1D513FC05500C00009543FC00000C0003C1A03D7B5605600003E03C3FC000300",
		INIT_02 => x"0015000C417F03FC0055000C457403FC0000000C156003FCFD413FC05400C000",
		INIT_03 => x"0000078528005500000000170000F40002D5079578007D0002F507F557E056F4",
		INIT_04 => x"0000078528005500000000170000F50002D5079578007D0002F507F557E057F4",
		INIT_05 => x"0000078528005500000000070000F40002D5078578007D0002F507E557E056F4",
		INIT_06 => x"00BE002C2FC0388003FA0FFFBF00FFC000BE01A8F800A90000BE00A2F8002800",
		INIT_07 => x"03F8022CBE0038000001002CFA803880002E002C2FC03880000F002CFA803880",
		INIT_08 => x"00FF02F6FC007E0002BF022C4000380003F8022CB800380002AF022CF0003800",
		INIT_09 => x"02FF0ABAFC00F00002BF2FF2EFF02800003F002FFF80AEA000FF0BFFFC00FF80",
		INIT_0A => x"0000553F0200FFE40000550B0030FD5500005501000F55440FFB0028FE008F38",
		INIT_0B => x"00001569002C05440000183DC000FA090002183DC000FA090003003DC000F800",
		INIT_0C => x"00BE01A8F800A90003FA0202BF00BE0000BE00A0F80028003800115000006954",
		INIT_0D => x"27161FE961006AF000000FFF0000FFF001000FFE0000BFF000000FFE0000BFF0",
		INIT_0E => x"2FFF000FD000D6C02FFF005DD1006B802FFF0055D440AF802FFF004BD190FD00",
		INIT_0F => x"00BF07FFFE00FFD00000000000000000000F03EAFA00A0000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000007C0000F40003D000001F00000000BE0FFFF800FFC000BE01A8F800A900",
		INIT_13 => x"000000000000000002AA0FFF0000FFC0000000000000000002FF02FEFE00FE00",
		INIT_14 => x"0BC801570C00FD000BC801FF0C00FD000BC801FF0C0055000BC809F50C007D00",
		INIT_15 => x"0000007800000000000000780000000000000078000000000000007800000000",
		INIT_16 => x"0000007800000000000000780000000000000078000000000000007800000000",
		INIT_17 => x"02AA0FE000003FC002AA0FFA0000BFC002AA0FFE0000FFC002AA0FFF0000FFC0",
		INIT_18 => x"000006AB0000EA90000002AF0000AAD0000002BE0000ABC0000002FA0000AF80",
		INIT_19 => x"003A057E0C00BF500000000000000000000003EA0000BE00000007AA0000FA80",
		INIT_1A => x"00AA0FE002802FC002A00FF524007FC0028400BF1800FE0000AA001F8000F000",
		INIT_1B => x"001A06000000FD0000030E000580F500000B0C072800FC000013057E0000AD00",
		INIT_1C => x"0000005400005454000000540000545400000054000054540000005000005454",
		INIT_1D => x"0000505400005454000000540000545400005054000054540000005400005454",
		INIT_1E => x"0000545400005454000054540000545400005454000054540000505400005454",
		INIT_1F => x"0000005400000000000000400000000000000054000000000000005400000000",
		INIT_20 => x"000002A00200061300000090A48203030080C49000000A80821AC0C000000600",
		INIT_21 => x"06000542080384000000009020000801C0300012009085400008003000000600",
		INIT_22 => x"06000050400100000000000000000C0340000000009005000000C03000000000",
		INIT_23 => x"0600000040010000000000000000000040000000009000000000000000000000",
		INIT_24 => x"00000000000001FF00000000003F00000000FFD000000000FF00000000000000",
		INIT_25 => x"00000000000001FE0000000000BF000000006FD000000000FF80000000000000",
		INIT_26 => x"00000000000003FF00000000001502A700007FF0000000005500B6A000000000",
		INIT_27 => x"0000000000000BFF000000050054FFA700007FF8000000000540B6BF0000D400",
		INIT_28 => x"33FF33FFFFC08AFF33FF187FFF85FFFF0000FFFF0000FFFF5FFDFFFF400AFFFF",
		INIT_29 => x"33FF33C0FFFF000033FE33FF0000F1FFFFFF0000FFFF057F0000FF010000C7FF",
		INIT_2A => x"0000FFF00000BFFFBFFDFFFF5400FFFF00004000FFFD002B0007E3EFFAAAEAFF",
		INIT_2B => x"FFFFFFFFFFFFFFFF0000F00000000000FFFFFFFFFFFFFFFF00000000000C0000",
		INIT_2C => x"00003C0F00002F7E00003CAF00003D5F00003EA00000F5E800003EEF00003EA0",
		INIT_2D => x"00BFFF00FFFF0000FF0007FF00008000FFFF0000FE0000FF0000000200FFFFD0",
		INIT_2E => x"00000000FFFFFFFF00000000FFFF00000000000000000000FFFF0000FFFF0000",
		INIT_2F => x"0000000000000000FFFF0000FFFF0000FFFFFFFF00000000FFFF000000000000",
		INIT_30 => x"000000000000FFFF00000000FFFFFFFF0000FFFF0000FFFF0000000000000000",
		INIT_31 => x"0000FFFF0000FFFF00000000000000000000FFFF00000000FFFFFFFF00000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"5000FC0C0BFF000BABFFFFFFFEAAFFFF4038F402D0B8FD02AABFFFFFA015FFFF",
		INIT_35 => x"FFFFFFFFC001FFFF000000000000AAFFFF80FFFF2FFFFFFF000000100555A400",
		INIT_36 => x"2CC5F0F0401F7F80404AFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_37 => x"FC0FF5454F402D02519A84F1AAAF9F80050001C200C48A00FFFCFFFF07FFFFFF",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_39 => x"0000415402A00000FFFCFFFF0F87FFFF0E2F00503FFF0000FFFFFFFFF83FFFFF",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCCFFCCFFFFFFFFFFCCFD24",
		INIT_3B => x"EF55000A007FAAA0FFC0FFFF21FFFFFFFFFF07FFFFCCFFCCFF80FFFF07CCFFCC",
		INIT_3C => x"0000000000000FFB00140000BFFF0FFFB000400000000000FF80000000000000",
		INIT_3D => x"000000000000000C000000000040000000000800000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000100040800000000000004000100020100000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7M_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"0FFF1FFABD00E0000FFF1FFABD00E4000FFB03EBFFC083000FE301FFFF80EB00",
		INIT_02 => x"007E000EFFF0AFF4007E000EFFF0AFF4007E001EFFF0AFF40FFF1FFABD00E000",
		INIT_03 => x"0F0D00785F000000003F0003FE00F0000F3D007F5F00D0000F7D007F5E7CFF40",
		INIT_04 => x"0F0D00785F000000003F0003F500F0000F3D007F5F00D0000F7D007F557CFF40",
		INIT_05 => x"0F0D00785F000000002F0003FE00F0000F2D007F5F00D0000F6D007F5E7CFF40",
		INIT_06 => x"003F00BFFD00FEC02AF7041F7EA0D04000FF0BF3FC003F8000FF0BFBFC00BF80",
		INIT_07 => x"007F03BFFC00FF00002A00FFBF40FEC0001F00BFFD00FEC000AB00BFFF40FEC0",
		INIT_08 => x"00FF0FFBFC00BFC001FE03BFAA00FF00007F03BFF400FF0001FF03BFEA00FF00",
		INIT_09 => x"20FF0CFFF400FC0028FFFFFFFF40BE00001F00FFFF08FF3000F70D7F7C00F5C0",
		INIT_0A => x"8000005501C055548000003F00F8FFE88000002B003CEA8001FF00BEFF28FFFF",
		INIT_0B => x"200000BE00BC2FA00003055080000154000301508000015000031A3080000629",
		INIT_0C => x"00FF0BF3FC003F80007F0FBBFC00FFC0087F0BFBF480BF803E000AF80008BE00",
		INIT_0D => x"0A0407FF0000D1D02FEA01FFA000FF40278001FF0000FF40278001FF0000FF40",
		INIT_0E => x"35FC000020001F50157F000020005D6035FC0000200055B035FC000000004BF0",
		INIT_0F => x"0B50007F05E0FD0000000000000000000007005FFFC0F0000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"02EB0000BA00000003FA0008BF00200000FF047FFC00F44000FF0BF3FC003F80",
		INIT_13 => x"00000000000000000FFF01FFF800FF40000000000000000001FF0FFBFD00BFC0",
		INIT_14 => x"0FE50095240056000FE50017240050000FE50255240058000FE5101524005000",
		INIT_15 => x"002A0000A000000000020000AA000000000000002AA000000000000002A00000",
		INIT_16 => x"0000000002A000000A000000002000000AA000000000000002AA000000000000",
		INIT_17 => x"0FFF01FFF800FF400FFF01FFF800FF400FFF01FFF800FF400FFF01FFF800FF40",
		INIT_18 => x"2F80005F0000F500000B005FE000F5000000005F02F8F5002F80005F0000F500",
		INIT_19 => x"00FD003F7820F0000000000000000000000B005FE000F5000000005F02F8F500",
		INIT_1A => x"003F007EF000FD0005FE01C0BA500F400FE001D02C001F400FD000BD18007E00",
		INIT_1B => x"002F006AF800C000002F01E28030F000082C01AB0180FF00002B002FF800FE00",
		INIT_1C => x"002A00002A2A0000002A00002A2A0000002A00002A2A0000002A00002A2A0000",
		INIT_1D => x"2A2A00002A2A0000002A00002A2A00002A2A00002A2A0000002A00002A2A0000",
		INIT_1E => x"2A2A00002A2A00002A2A00002A2A00002A2A00002A2A00002A2A00002A2A0000",
		INIT_1F => x"222A0000000000002202000000000000222A000000000000222A000000000000",
		INIT_20 => x"00600000030358410150000009230100C0C0412509000000C860004005400000",
		INIT_21 => x"006000000C00100002A1090048000C0380100004090000000021C01042A00060",
		INIT_22 => x"000000000C03000000A0090000000002C030000000000000000080020A000060",
		INIT_23 => x"0000000000000000000009000000000200000000000000000000800200000060",
		INIT_24 => x"000000000000021400000000001F000000000520000000007D00000000000000",
		INIT_25 => x"0000000000000094000000000074000000000580000000000740000000000000",
		INIT_26 => x"0000000000000060000000000000BFC00000024000000000400000FF00008000",
		INIT_27 => x"00000000000001E00000000000000000000002D0000000004000000000000000",
		INIT_28 => x"33FF33FFF540E3FF33FF0785FFFF55550000FFFF0000FFFFEAAA5555AFFF5555",
		INIT_29 => x"33FF33C0FFFF000033FF33FF1FFFFCFFFFFF0000FFFF0000F05FFF00FFFF4155",
		INIT_2A => x"A800FFD20000F874FFFF5555EA80555500020002F5408BFF000051557FFF5555",
		INIT_2B => x"FFFF57D4FFFF0000F000500000000000FFFF0000FFFF003F00000000FC0C0000",
		INIT_2C => x"00003C0F00003C0F00001E0000001E2D00003C000000F03C00003F7F00003C00",
		INIT_2D => x"0BFFFF0040000000FF00007F0000FFFF00010000FFE000FF0000FFFF00FFFD00",
		INIT_2E => x"00000000FFFFFFFF00000000FFFF00000000000000000000FFFF0000FFFF0000",
		INIT_2F => x"0000000000000000FFFF0000FFFF0000FFFFFFFF00000000FFFF000000000000",
		INIT_30 => x"000000000000FFFF00000000FFFFFFFF0000FFFF0000FFFF0000000000000000",
		INIT_31 => x"0000FFFF0000FFFF00000000000000000000FFFF00000000FFFFFFFF00000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"0002FC2FFFD000BFFFFF5555FFFF5555003CD00702F0F403FFFF5555FFFF5555",
		INIT_35 => x"FFFFC0FFCA00555FFE03AAFEFFFC3FF51FF0FFFF3FFFFFFF03FF400DF5550080",
		INIT_36 => x"00E3F0F0E0073F43FFFF5555FFFF5555FFFFFFFFFFFFFFFFFFFF5555FFFF5555",
		INIT_37 => x"FF0F50022D00D025E40A30F8AAA071C210020051817FFF000000FFFF0000FFFF",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFF5555FFFF5555FFFFFFFFFFFFFFFFFFFF5555FFFF5555",
		INIT_39 => x"A00A0000BFF800000000FFFFFFFAFFFF0FFF000A1F5502AF0000FFFF0000FFFF",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFF5555FFFF5555FFFFFFFFFFCCFFCCFFFF5555FFCC52D0",
		INIT_3B => x"0000FF01000FFFFC0000FFFF3E00FFFFFFFF007FFFCCFFCC0000FFFF03CCFFCC",
		INIT_3C => x"0000000000B7BFFE00030000FFFF07544000E00000000000FFC0000000000000",
		INIT_3D => x"00000000000000BF00000000000000000000BC00000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000441010040008100000800000004100404200000000204001000400000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_7M_3 : RAMB16_S2
	generic map (
		INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => x"03D501550000000003C501550000000001FD007F5500FD0001FD001555405400",
		INIT_02 => x"0000000053C055400000000057C055400000000053C0554003C5015500000000",
		INIT_03 => x"0F0E0000AF000000003F0000FD0000000F3E0000AF0000000F3E0000AD3C0000",
		INIT_04 => x"0F0E0000AF000000003F0000F80000000F3E0000AF0000000F3E0000A83C0000",
		INIT_05 => x"0F0A0000AF000000000B0000FD0000000F0A0000AF0000000F0A0000AD3C0000",
		INIT_06 => x"0BFF00D7DDF0FD00074000000740000000F70D7F7C00F5C00BF70D7F7F80F5C0",
		INIT_07 => x"0F77007FFFE0D700001F00D7DDC0FD00000700D7DDD0FD00007F00D7DD00FD00",
		INIT_08 => x"02D1041F1E00D0400377007FF500D7000777007FD0C0D7000077007FFD00D700",
		INIT_09 => x"7D5501FD7BC004001FFF41FFFE80D70003ED0041557DFF400B40000507804000",
		INIT_0A => x"300A0000A1780000300A0000AAFC0000300A0055A87C555502BF00D7FFF4FF41",
		INIT_0B => x"0E020055AA7C5555202F000000020000002F000000000000002F005000000140",
		INIT_0C => x"00F70D7F7C00F5C03FDD0D7FFEA0D0401EB70D7F7AD0F5C03DAA555580B05500",
		INIT_0D => x"33E8007F2A00E1003FFF0015FF8054003BFE0015BD0054003BFE0015BD005400",
		INIT_0E => x"00360000F000005F003600005800005D00340000A800005B00360000F800000F",
		INIT_0F => x"0FCA00002FF00000000000000000000000010000555000000000000000000000",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"07FF0000FF4000000FFF0054FFC054003EF500007EF0000000F70D7F7C00F5C0",
		INIT_13 => x"00000000000000003FFF0005FF00500000000000000000000BD1041F1F80D040",
		INIT_14 => x"0A1500004000004002050001400000002A05000040000000AA05000040000000",
		INIT_15 => x"0030000030000000000300000300000000000000303000003000000003000000",
		INIT_16 => x"3000000003000000030000000030000030300000000C00000303000000000000",
		INIT_17 => x"3F5000051F0050003FD500057F0050003FFD0005FF0050003FFF0005FF005000",
		INIT_18 => x"FFFF0000FC000000FFFF0000FC000000FFFF0000FC000000FFFF0000FC000000",
		INIT_19 => x"3FD000051F0050000000000000000000FFFF0000FC000000FFFF0000FC000000",
		INIT_1A => x"20BF0005FE245000003F0000F000000035FE0000BF5800003FE000002F001000",
		INIT_1B => x"3AD70005FF0040003FFF0005F80050003FFE0005004050003FD000051F005000",
		INIT_1C => x"007F0000FFFF0000007F0000FFFF000000FE0000FFFF0000007C0000FFFF0000",
		INIT_1D => x"7CFF0000FFFF000000FF0000FFFF00007CFF0000FFFF0000007F0000FFFF0000",
		INIT_1E => x"7FFF0000FFFF0000FEFF0000FFFF00007FFF0000FFFF00007CFE0000FFFF0000",
		INIT_1F => x"667F00000000000066BF000000000000667F00000000000066FE000000000000",
		INIT_20 => x"000600AA00030A8F0000000000C00000C000F2A09000AA000300000000000000",
		INIT_21 => x"00002A2A020300000000000092400001C08000020000A0A88186400000000000",
		INIT_22 => x"0006A8A000000000280010000000C0030000000090000A2A0000C001000A0004",
		INIT_23 => x"0000A80000000000280010000000C003000000000000002A0000C001000A0004",
		INIT_24 => x"00000000000207E00000000000000000A00002F4000000000000000000000000",
		INIT_25 => x"00000000000201E00000000000000000A00002D4000000000000000000000000",
		INIT_26 => x"000000000000021E000000000001BD000000AD20000000005000001F00008000",
		INIT_27 => x"000000000000003E00320000000100000000AF00000000005000000023000000",
		INIT_28 => x"33FF33FF5000F8FF33FF0015FFFF55550000FFFF04FFFFFFFFFF5555FFFF5555",
		INIT_29 => x"33FF33F0FFFF000033FF33FFCFFFFE15FFFF0000FFFF0000F8015000FFFF0000",
		INIT_2A => x"FF80D50B20008780FFFF5555FFCA55550018002F0000C7FF0006555581FF5555",
		INIT_2B => x"FFFF0000FFFF0000F000000000000000FFFF0000FFFF003C000000003C002ACF",
		INIT_2C => x"0000055400001405000001550000015000001554000055500000140500001554",
		INIT_2D => x"BFF4FF0000000000FF8000070000FFFF000000001FFE00FF0000FFFF02FFD000",
		INIT_2E => x"00000000FFFFFFFF00000000FFFF00000000000000000000FFFF0000FFFF0000",
		INIT_2F => x"0000000000000000FFFF0000FFFF0000FFFFFFFF00000000FFFF000000000000",
		INIT_30 => x"000000000000FFFF00000000FFFFFFFF0000FFFF0000FFFF0000000000000000",
		INIT_31 => x"0000FFFF0000FFFF00000000000000000000FFFF00000000FFFFFFFF00000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"0007D03FFD00C3FDFFFF5555FFFF55550010000107C0D00FFFFF5555FFFF5555",
		INIT_35 => x"FFFF0035C5400000FF80FFFFF555850000530C00FFFF001500008000AA150B40",
		INIT_36 => x"0211C0FCFC010D2FFFFF5555FFFF5555FFFFFFFFFFFFFFFFFFFF5555FFFF5555",
		INIT_37 => x"FF0D031934B008429C1A08CEA8551E0B0C25C00000370000FFFAFFFF2BFFFFFF",
		INIT_38 => x"FFFFFFFFFFFFFFFFFFFF5555FFFF5555FFFFFFFFFFFFFFFFFFFF5555FFFF5555",
		INIT_39 => x"CAC70008FFFC02AFFFFFFFFFFFFFFFFF03FFFABFC00083FFFA00FFFF0800FFFF",
		INIT_3A => x"FFFFFFFFFFFFFFFFFFFF5555FFFF5555FFFFFFFFFFCCFFCCFFFF5555FFCC5400",
		INIT_3B => x"0000FF0000017FFF0003FFFFFFC0FFFFFFFF8007FFCCFFCC0000FFFF3FCCFFCC",
		INIT_3C => x"0000000300E7FFFF00010000FFFD00000000D00000000000FF40000000000000",
		INIT_3D => x"000000000000001F00000000000000000000FD00000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000002002008000000000004000000000000000004008000400000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
