-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0000BFEA0000A00000000AFF0000F8000000002F0000FFF50000017F00000000";
    attribute INIT_01 of inst : label is "0000FFFF000000170000FF400000EAAA000000BF0000FF50000017FF0000AAFF";
    attribute INIT_02 of inst : label is "7F80FF5500005000FFFF2FF8FFFF2FF807D0000007D000000140000001400000";
    attribute INIT_03 of inst : label is "F800F5558007D00F003FAABF3FC03FEA00FF00FFF000F000F40FFC0F000B5557";
    attribute INIT_04 of inst : label is "0618000006180000000000000000000002FF0000FE000000007F0002F400BFC0";
    attribute INIT_05 of inst : label is "00030003FF00FF00BF407FC00000555507F80FF53F80BFD0C000EAAA403FC03F";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "00FF0FFF0000FFFFF000FFFFFC0FFC0F01500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "C000FFFFC03FC0FF003F003FF000F000FC0F000F000FFFFA3FC0FFFF0000F000";
    attribute INIT_0D of inst : label is "001F000AFFD0FE8000BF557F000040003FC03FC0000000000FF00FF00FFCFA00";
    attribute INIT_0E of inst : label is "FC0000004000FC001F00000000800001000000000000000000000000801F0100";
    attribute INIT_0F of inst : label is "FC2F00005401FC3FFFFF00005555000ACFC0000005418FE03F00000050053F80";
    attribute INIT_10 of inst : label is "0008000A30C3A828330C80A0030C0802AA4C2A02090C2A02030C0A8200000000";
    attribute INIT_11 of inst : label is "000000003000800030CC0A02A4C3A028000A000290C3A0280000000218C3A828";
    attribute INIT_12 of inst : label is "000000AF0AA8000045FC45F80000FA002F51000000AF3F1145F80000FA0045FC";
    attribute INIT_13 of inst : label is "D7000AA80000BC0002FF02A8FC0037FF5FF802A8A000FFFC280000003F113F51";
    attribute INIT_14 of inst : label is "EEBAAEBA7B2560C22F51000000AF3F1145F80000FA0045FC00D72AA00000003E";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "00FF00AAFF00AA000000AA2A0000AA2A00000000000000000000000000000000";
    attribute INIT_18 of inst : label is "FFCFF3FFFFCFF3FFFF3F0000FF3F000000FF0000FF000000AA00FFCF00FCFFFC";
    attribute INIT_19 of inst : label is "FFFFFF00CFFC00FCAA00FF3F00AAFFFFFFFFFF00FCFF00FFFF00000000FF0000";
    attribute INIT_1A of inst : label is "AA00FFCF00A8FFCFAA00FF3F00AAFCFFFF00FF0000FF00FFFF3FFF00FCFF00FF";
    attribute INIT_1B of inst : label is "0000FFCF0000FFCF0000FCFF0000FCFFFCFF0000FCFF0000CFFFFF00CFFF00FC";
    attribute INIT_1C of inst : label is "000000C000000300CFFF0000CFFF000000FF00AAFF00AA000000FF3F0000FF3F";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF00000000FF0000FF0000FC00545500FF00";
    attribute INIT_1E of inst : label is "000000000000000000000000000000000000000000000000FF00000000FF0000";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "2F513F1100AF2AA045FC45FCFA0000283F513F1100AF280045F845FCFA000AA8";
    attribute INIT_21 of inst : label is "0BFC3FFF07FF00803FE0FFFCFFD002000E1537FFB8152A8054B0FFDC542E02A8";
    attribute INIT_22 of inst : label is "0F87000201082AAAD2F0FE002060AAA800780002010800002D00FE0020600000";
    attribute INIT_23 of inst : label is "0FFF00020108AAA0FFF0FE0020600AAA0F87000201082AAAD2F0FE002060AAA8";
    attribute INIT_24 of inst : label is "2F513F1107FC3FF045F845FC3FD00FFC2F513F1107FC00F045F845FC3FD00F00";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "FFFFFFFFC0FF000055FCFFE0FFFC0000FFFF08000400FFFFFFF000000000FFFC";
    attribute INIT_29 of inst : label is "000F0002000F0000D57FFFFFFFFF000003C3BFFEFFFF03FFFFFF00000000FFFF";
    attribute INIT_2A of inst : label is "407FFFFF0000A2AA8000FFE0003C8000FFFF08000400FFFFFFF000000000FFFC";
    attribute INIT_2B of inst : label is "FFFF17D603EF2AA800BFFFFF000000AA000300000000000FFFFF00000000FFFF";
    attribute INIT_2C of inst : label is "000FFFFFFFFF000A0000FA00FFF00000FF5FFFAFFFFFFFFFFFFCFFD0D500FFFC";
    attribute INIT_2D of inst : label is "000000AF0FFF0000F000FFFFFFFFA0003FFF07FF00573FFFF5FFFAFFFFFFFFFF";
    attribute INIT_2E of inst : label is "000FFDFF5455000AF000DFFC4554AA80FF00FFAAFFFFFCFF3FFCBFD0D500CFFC";
    attribute INIT_2F of inst : label is "000F3FF7155102AAF000FF7F5515A0003FFC07FE00573FF300FFAAFFFFFFFF3F";
    attribute INIT_30 of inst : label is "0BFF3FFF07FF0080FFE0FFFCFFD002003CF33EFB07FF2A80CF3CEFBCFFD002A8";
    attribute INIT_31 of inst : label is "00C0003E00000AA0033CBC00000000283C0C003E000028003000BC0000000AA8";
    attribute INIT_32 of inst : label is "0BF33FC107FF2AA0CFFC43FCFFD000283FF33FC107FF2800CFE043FCFFD00AA8";
    attribute INIT_33 of inst : label is "08033FC107FF2AA0C03C43FCFFD000283C033FC107FF2800C02043FCFFD00AA8";
    attribute INIT_34 of inst : label is "0202630C0000000080A0330C00000000AA82818C0000000080A0330C00000000";
    attribute INIT_35 of inst : label is "0020000F00000000A0280CC3000000002A02958C0000000080A0330C00000000";
    attribute INIT_36 of inst : label is "76C007FF000002A80038FFFCA00002A802FF37FFFC0000085FF8FFFCA0000200";
    attribute INIT_37 of inst : label is "3FFF000200002AAAFFFC80000000AAA82D5507FF00012A805578FFD0400002A8";
    attribute INIT_38 of inst : label is "0002000000002AAA800000000000AAA801FF000100002AAAFF4040000000AAA8";
    attribute INIT_39 of inst : label is "00020000000002A0800000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000300001000002A00C00400000000A80";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "000000000000000000000000000000000A000124000000180140600000009200";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0000555500005000000005550000540000000015000055000000000100000000";
    attribute INIT_01 of inst : label is "0000155000000000000050000000555500000055000050000000001500005550";
    attribute INIT_02 of inst : label is "1FFAFF00000000001FF4FFFF1FF4FFFF00000BE000000BE00000028000000280";
    attribute INIT_03 of inst : label is "FFA0F000C001000F003F55F83FC03FD500FF00FFF000F000D00FFC0F02BF0003";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000000000000000000017002AFFC0A000000002BF0000FF40";
    attribute INIT_05 of inst : label is "AAAB0003FFAAFF00FD003FC0A02B000001FF0FF03FC0F800C000D555003FC03F";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "00FF00FF00000007F000F000FC0FFC0F00000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "C000C000C03FC03FAABF003FFAAAF000FC0FF00F000F001F3FC03FC000000000";
    attribute INIT_0D of inst : label is "0005002FFD40FFE02BFD003F00000000BFC03FC0AAAA00000FFA0FF00FFC1FF0";
    attribute INIT_0E of inst : label is "FC00A8000000F400BD00A800007A00030000000000000000000000007ABD03A8";
    attribute INIT_0F of inst : label is "FC3FA8020000FC1F0005AAAA0000FFFF4FC00A800000CFDF3F002A000000FF7F";
    attribute INIT_10 of inst : label is "00060001706930C391A4330CEAC60C0CEA8640CCAB8640CC0706030C00000000";
    attribute INIT_11 of inst : label is "00000000900030001A4630CCA8690CC3000E0004B8690CC3000A0004A46980C3";
    attribute INIT_12 of inst : label is "00000155AF540000EFD044FC000055403F5102BF015507FB44FCFE805540EFD0";
    attribute INIT_13 of inst : label is "550085540000140003FF003E540031FFAFFCABC05000FFF43DFA000007FB3F51";
    attribute INIT_14 of inst : label is "0410AEBB240606E43F5102BF015507FB44FCFE805540EFD00055155200000014";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "00FF00FFFF00FF000000FF3F0000FF3F00000000000000000000000000000000";
    attribute INIT_18 of inst : label is "5545515555455155FF3F0000FF3F000000FF0000FF000000FF00FFCF00FCFFFC";
    attribute INIT_19 of inst : label is "5555FF0045540054FF00FF3F00FFFFFF55555500545500555500000000550000";
    attribute INIT_1A of inst : label is "FF00FFCF00FCFFCFFF00FF3F00FFFCFFFF00550000FF0055FF3F5500FCFF0055";
    attribute INIT_1B of inst : label is "0000FFCF0000FFCF0000FCFF0000FCFFFCFF0000FCFF00004555550045550054";
    attribute INIT_1C of inst : label is "0000001A0000A400455500004555000000FF00FFFF00FF000000FF3F0000FF3F";
    attribute INIT_1D of inst : label is "00FD0000FF000000000000FF0000FF00000000FF0000FF0000FC00FCFF00FF00";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000005500000000550000";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "3F5107FB015515FA44FCEFD05540AFFC3F5107FB01553DFA44FCEFD05540AF54";
    attribute INIT_21 of inst : label is "3FFF1FFF001500EAFFFCFFF45400AB003FFF31FFCC0003E8FFFCFF4C00332BC0";
    attribute INIT_22 of inst : label is "015F008100100ABEFF40FD141000BEA000000081001000010000FD1410004000";
    attribute INIT_23 of inst : label is "01FF008100104E15FF40FD14100054B1015F008100100ABFFF40FD141000FEA0";
    attribute INIT_24 of inst : label is "3F510FFB000502FA44FCEFF05000AF803F510FFB000502FA44FCEFF05000AF80";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "FFFFC0FFFFFFFFFFF054FFF0FFFCFFFCFFFF3F000000FFFFFF4000000000FFFC";
    attribute INIT_29 of inst : label is "00050003000F000F43FFFFFFFFFFFFFF03C0FFFF7FFD03DF7FFF00000000FFFF";
    attribute INIT_2A of inst : label is "FFFF0000FFFFF3FDF800003CFFFC4000FFFF3F000000FFFFFF4000000000FFFC";
    attribute INIT_2B of inst : label is "FFFF03CF03FFFFFF0BFF0000FFFF005F000000000000000F7FFF00000000FFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFF000F0000FFC0FFFC0000FF0FFFFF5540FFFFFFF4FF400000FFFC";
    attribute INIT_2D of inst : label is "000003FF3FFF0000FFFFFFFFFFFFF0001FFF01FF00003FFFF0FFFFFF0155FFFF";
    attribute INIT_2E of inst : label is "AAAFFCFFFCFF000FFAA8CFFCCFFCFFC0FF00FFFF5500FFFF3FF4FF400000FFFC";
    attribute INIT_2F of inst : label is "2AAF3FF33FF303FFFAAAFF3FFF3FF0001FFC01FF00003FFF00FFFFFF0055FFFF";
    attribute INIT_30 of inst : label is "3FFF1FCF001500EAFFFCF3F45400AB0028A21F0F00152BEA8A28F0F45400ABE8";
    attribute INIT_31 of inst : label is "00550014000005FA550014000000AA3C0005001400003C0A500014000000A554";
    attribute INIT_32 of inst : label is "3FFA1FEB001515F0AFFCEBF454000F7C3FFA1FEB00153DF0AFFCEBF454000F54";
    attribute INIT_33 of inst : label is "3FAA1FEB00151550AAFCEBF45400057C3FAA1FEB00153D50AAFCEBF454000554";
    attribute INIT_34 of inst : label is "AB8C070600000000330C91A400000000180C6A4600000000330C91A400000000";
    attribute INIT_35 of inst : label is "0033000D000000000CC3A46900000000C0CC6A4600000000330C91A400000000";
    attribute INIT_36 of inst : label is "3BEA01FF0000FCBEAABCFFF45000ABE003FF31FF5400002EAFFCFFF45000AB80";
    attribute INIT_37 of inst : label is "07FF000100001B55FFD04000000055E43FFF000200000070FFFC800000000D00";
    attribute INIT_38 of inst : label is "00010000000010EA400000000000AB0400020000000012D58000000000005784";
    attribute INIT_39 of inst : label is "00010000000000304000000000000D400000000000000003000000000000C000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000020000000000308000000000000C00";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000800000000001800600000000000400";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "0000BFEA0000A00000000AFF0000F8000000002F0000FFF50000017F00000000";
    attribute INIT_01 of inst : label is "0000FFFF000000170000FF400000EAAA000000BF0000FF50000017FF0000AAFF";
    attribute INIT_02 of inst : label is "7F80FF5500005000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "F800F5558007D00F003FAABF3FC03FEA00FF00FFF000F000F40FFC0F000B5557";
    attribute INIT_04 of inst : label is "0618000006180000000000000000000002FF0000FE000000007F0002F400BFC0";
    attribute INIT_05 of inst : label is "00030003FF00FF00BF407FC00000555507F80FF53F80BFD0C000EAAA403FC03F";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "00FF0FFF0000FFFFF000FFFFFC0FFC0F01500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "C000FFFFC03FC0FF003F003FF000F000FC0F000F000FFFFA3FC0FFFF0000F000";
    attribute INIT_0D of inst : label is "001F000AFFD0FE8000BF557F000040003FC03FC0000000000FF00FF00FFCFA00";
    attribute INIT_0E of inst : label is "FC0000004000FC001F00000000800001000000000000000000000000801F0100";
    attribute INIT_0F of inst : label is "FC2F00005401FC3FFFFF00005555000ACFC0000005418FE03F00000050053F80";
    attribute INIT_10 of inst : label is "0008000A30C3A828330C80A0030C0802AA4C2A02090C2A02030C0A8200000000";
    attribute INIT_11 of inst : label is "000000003000800030CC0A02A4C3A028000A000290C3A0280000000218C3A828";
    attribute INIT_12 of inst : label is "000000000AA80000BA00BA000000000000AE0000000000EEBA0000000000BA00";
    attribute INIT_13 of inst : label is "E8E00AA8FFD0FFFC02FF02A8FFFF37F5FFF802A85FFCF5FC2800000000EE3CAE";
    attribute INIT_14 of inst : label is "EEBAAEBA7EF578C200AE0000000000EEBA0000000000BA000B2B2AA007FF3FFF";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "00FF00AAFF00AA000000AA2A0000AA2A00000000000000000000000000000000";
    attribute INIT_18 of inst : label is "FFCFF3FFFFCFF3FFFF3F0000FF3F000000FF0000FF000000AA00FFCF00FCFFFC";
    attribute INIT_19 of inst : label is "FFFFFF00CFFC00FCAA00FF3F00AAFFFFFFFFFF00FCFF00FFFF00000000FF0000";
    attribute INIT_1A of inst : label is "AA00FFCF00A8FFCFAA00FF3F00AAFCFFFF00FF0000FF00FFFF3FFF00FCFF00FF";
    attribute INIT_1B of inst : label is "0000FFCF0000FFCF0000FCFF0000FCFFFCFF0000FCFF0000CFFFFF00CFFF00FC";
    attribute INIT_1C of inst : label is "000000FF0000FF00CFFF0000CFFF000000FF00AAFF00AA000000FF3F0000FF3F";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF00000000FF0000FF0000FC00545500FF00";
    attribute INIT_1E of inst : label is "000000000000000000000000000000000000000000000000FF00000000FF0000";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "00AE00EE00002AA0BA3CBA00000000283CAE00EE00002800BA00B80000000AA8";
    attribute INIT_21 of inst : label is "0BF33FFF07FF0080CFE0FFFCFFD0020001EA3787B8152A80AB40D2DC542E02A8";
    attribute INIT_22 of inst : label is "00780002010800002D00FE00206000000FFF000201082AAAFFF0FE002060AAA8";
    attribute INIT_23 of inst : label is "0EAA00020108A000AAB0FE002060000A00000002010800000000FE0020600000";
    attribute INIT_24 of inst : label is "00AE00EE07FF3FF0BA00BA00FFD00FFC00AE00EE07FF00F0BA00BA00FFD00F00";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFF000055FCFFE0FFFC0000FFFFF7FFFBD5FFFFAFF0FFC05400FFFC";
    attribute INIT_29 of inst : label is "000F0002000F0000D57FFFFFFFFF000003C3BFFEFFFF03FFFEBFFFFF0555FFFF";
    attribute INIT_2A of inst : label is "407FFFFFFFFFA2AA8000FFE0FFFC8000FFF8F7FFFBD57F550FF0FFC054005FFC";
    attribute INIT_2B of inst : label is "FFFF17D603EF2AA800BFFFFFFFFF00AA000300000000000FFC0BFFFF0555FD55";
    attribute INIT_2C of inst : label is "000F003FF03F000A0000FA00FFF00000F5F7FF53FFFF003FFFFCFFD0D500FFFC";
    attribute INIT_2D of inst : label is "000000AF0FFF0000F000FC00FC0FA0003FFF07FF00573FFFDF5FC5FFFFFFFC00";
    attribute INIT_2E of inst : label is "000F5755ABAA000AF0007554BAA8AA80F0FFF055FFFF0300C3FC43D0D5003000";
    attribute INIT_2F of inst : label is "000F155D2AAE02AAF00055D5AAEAA0003FC307C10057000CFF0F550FFFFF00C0";
    attribute INIT_30 of inst : label is "0BC23FEA07BF008083E0ABFCFED00200030C2BAE07AF2A8030C0BAE8FAD002A8";
    attribute INIT_31 of inst : label is "0B3F3FFF07FF0AA0FCFCFFFCFFD000283FF33FFF07FF2800CFE0FFFCFFD00AA8";
    attribute INIT_32 of inst : label is "000C00FF00002AA0303CFF00000000283C0C00FF000028003000FF0000000AA8";
    attribute INIT_33 of inst : label is "03FF000000002AA0FFFC0000000000283FFF000000002800FFC0000000000AA8";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "76FF07C203FF02A8FFF8F83C5FFC02A802FF37F5FFFF0008FFF8F5FC5FFC0200";
    attribute INIT_37 of inst : label is "3F5F0FFD00002AAAF5FC7FF00000AAA82FFF07EB015E2A80FFF8EBD0B54002A8";
    attribute INIT_38 of inst : label is "0FFD000000002AAA7FF000000000AAA801FF015E00002AAAFF40B5400000AAA8";
    attribute INIT_39 of inst : label is "0FFD0000000002A07FFC0000000000000005000000000AAA500000000000AAA0";
    attribute INIT_3A of inst : label is "000000000000000000000000000000000030015E000002A00C00B54000000A80";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "000000000000000000000000000000000A000124000000180140600000009200";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0000555500005000000005550000540000000015000055000000000100000000";
    attribute INIT_01 of inst : label is "0000155000000000000050000000555500000055000050000000001500005550";
    attribute INIT_02 of inst : label is "1FFAFF0000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "FFA0F000C001000F003F55F83FC03FD500FF00FFF000F000D00FFC0F02BF0003";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000000000000000000017002AFFC0A000000002BF0000FF40";
    attribute INIT_05 of inst : label is "AAAB0003FFAAFF00FD003FC0A02B000001FF0FF03FC0F800C000D555003FC03F";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "00FF00FF00000007F000F000FC0FFC0F00000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "C000C000C03FC03FAABF003FFAAAF000FC0FF00F000F001F3FC03FC000000000";
    attribute INIT_0D of inst : label is "0005002FFD40FFE02BFD003F00000000BFC03FC0AAAA00000FFA0FF00FFC1FF0";
    attribute INIT_0E of inst : label is "FC00A8000000F400BD00A800007A00030000000000000000000000007ABD03A8";
    attribute INIT_0F of inst : label is "FC3FA8020000FC1F0005AAAA0000FFFF4FC00A800000CFDF3F002A000000FF7F";
    attribute INIT_10 of inst : label is "00060001706930C391A4330CEAC60C0CEA8640CCAB8640CC0706030C00000000";
    attribute INIT_11 of inst : label is "00000000900030001A4630CCA8690CC3000E0004B8690CC3000A0004A46980C3";
    attribute INIT_12 of inst : label is "00000000075400001000BB000000000000AE000000000004BB00000000001000";
    attribute INIT_13 of inst : label is "AAFCAF545400FFF403FF003E545731FAFFFCABC0AD50FAF43D500000000400AE";
    attribute INIT_14 of inst : label is "0410AEBB2D1E2D9C00AE000000000004BB000000000010003FAA15FA00151FFF";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "00FF00FFFF00FF000000FF3F0000FF3F00000000000000000000000000000000";
    attribute INIT_18 of inst : label is "5545515555455155FF3F0000FF3F000000FF0000FF000000FF00FFCF00FCFFFC";
    attribute INIT_19 of inst : label is "5555FF0045540054FF00FF3F00FFFFFF55555500545500555500000000550000";
    attribute INIT_1A of inst : label is "FF00FFCF00FCFFCFFF00FF3F00FFFCFFFF00550000FF0055FF3F5500FCFF0055";
    attribute INIT_1B of inst : label is "0000FFCF0000FFCF0000FCFF0000FCFFFCFF0000FCFF00004555550045550054";
    attribute INIT_1C of inst : label is "0000001F0000F400455500004555000000FF00FFFF00FF000000FF3F0000FF3F";
    attribute INIT_1D of inst : label is "00FD0000FF000000000000FF0000FF00000000FF0000FF0000FC00FCFF00FF00";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000005500000000550000";
    attribute INIT_1F of inst : label is "FFFFFFFF00000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "00AE0004000015D0BB0010000000057C00AE000400003D50BB00100000000754";
    attribute INIT_21 of inst : label is "3FFA1FEB001500E0AFFCEBF454000B003EAA31FFCC000140AABCFF4C00330140";
    attribute INIT_22 of inst : label is "00000081001000010000FD1410004000015F008100100ABEFF40FD141000BEA0";
    attribute INIT_23 of inst : label is "01AB0081001041EAEA40FD141000AB4100000081001000010000FD1410004000";
    attribute INIT_24 of inst : label is "00AE0AAE00050000BB00BAA05000000000AE0AAE00050000BB00BAA050000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFF054FFF0FFFCFFFCFFFFC0FF0000FFE0FF40FFC000001FFC";
    attribute INIT_29 of inst : label is "00050003000F000F43FFFFFFFFFFFFFF03C0FFFF7FFD03DF7FFFFFFF0000FD02";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFF3FDF800FFFCFFFC4000FFFFC0FF0000BF80AF40FFC000000FFC";
    attribute INIT_2B of inst : label is "FFFF03CF03FFFFFF0BFFFFFFFFFF005F000000000000000F7EBFFFFF0000FC00";
    attribute INIT_2C of inst : label is "FFFFA03F503F000F0000FFC0FFFC0000F8F3FFE35540FFFFFFF4FF400000FFFC";
    attribute INIT_2D of inst : label is "000003FF3FFF0000FFFFFC0AFC05F0001FFF01FF00003FFFCF2FCBFF0155FFFF";
    attribute INIT_2E of inst : label is "AAAF03000300000FFAA830003000FFC0F0FFFFAA5500FFFFC3F4BF400000FFFC";
    attribute INIT_2F of inst : label is "2AAF000C000C03FFFAAA00C000C0F0001FC301FE00003FFFFF0FAAFF0055FFFF";
    attribute INIT_30 of inst : label is "3FC11F3B001500C043FCECF454000300175D1CF300152BEA75D4CF345400ABE8";
    attribute INIT_31 of inst : label is "3FAA1FFF00150550AAFCFFF45400057C3FFA1FFF00153DF0AFFCFFF454000F54";
    attribute INIT_32 of inst : label is "00AF00FF0000155AFA00FF000000A03C00AF00FF00003C5AFA00FF000000A554";
    attribute INIT_33 of inst : label is "00550000000015FA550000000000AA3C0055000000003CAA550000000000AF54";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "3BFF01EF0057FCBEFFFCFFB4AD50ABE003FF31FA5457002EFFFCFAF4AD50AB80";
    attribute INIT_37 of inst : label is "07EB015E00001BFFEBD0B5400000FFE43FFF0FFD00000070FFFC7FF000000D00";
    attribute INIT_38 of inst : label is "015E0000000010FFB54000000000FF040FFD0000000012FF7FF000000000FF84";
    attribute INIT_39 of inst : label is "015E000000000030B540000000000D4000000000000007FC0000000000003FD0";
    attribute INIT_3A of inst : label is "000000000000000000000000000000000FFD0000000000307FF0000000000C00";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000800000000001800600000000000400";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
