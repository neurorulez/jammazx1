-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0000000700000000FC3FFC3F00000000003F003FFC00FC000000D00000000000";
    attribute INIT_01 of inst : label is "06E401D007F402E03F7F02E0FFFFFFFF0000FFFF00000000AAAA00000000D007";
    attribute INIT_02 of inst : label is "000707FFF400FFF4FFE0E0001FFDFFFFFF8080001FFD3FFF00BF000007F409D8";
    attribute INIT_03 of inst : label is "FE00C7F4000000010000D000007F1FFFFF40FFFD2FFEF4002FFE000702FF0002";
    attribute INIT_04 of inst : label is "00B000000BD600000BD600005F80000000030000C003D5570FF0014000000000";
    attribute INIT_05 of inst : label is "00000000000003C000000000000000000BDE000001F800002F5800000B600000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0000000000F400E009D818C907C002C0F82FC003014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC6832558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "0000000003FF03FC2FFDFFFFFFFF000003FF0000201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "FFD08880A1FF0008F500F7FD0017AA4703FF03C107C0FFC000F408FF03C303FF";
    attribute INIT_0D of inst : label is "2FC30FC303FF03FF3C00FFFF0FF0FFFF0000F0C00000FFFF0000FFFFFFC0FFC0";
    attribute INIT_0E of inst : label is "7FFFFFFFFFFFFFFFFD00FFFFABC00BC0C1FF07FF402FFF03FFF5FC001F003C00";
    attribute INIT_0F of inst : label is "FC07FC00FE00300000020000FFFF8200FFFF0020743FFC3F68F050A803CA0A81";
    attribute INIT_10 of inst : label is "14F480FF001500F2FD3FFEBFFFC0FFFC03FD1FD0FEBF003F47FFFFE0FFFF02BF";
    attribute INIT_11 of inst : label is "00023F4003FF03FF4000FF003FFF3FFF01FF03FFFFFF003FFFFF02BEFFFF002A";
    attribute INIT_12 of inst : label is "04C0000000C40000FD7FFFFFFFFFFFE0FFFF00BFFDFDFFFFA83F083FFF000200";
    attribute INIT_13 of inst : label is "FFFF0000FFC0FAC0FF04AF00E00000BF0000FFC00000001F0000FD00FFC003C0";
    attribute INIT_14 of inst : label is "07FD007E9696F69FD5008000015F000B2CC31D96000000070000F400002F07F4";
    attribute INIT_15 of inst : label is "0000000F0000FC03020001E006BA03E080003F005F570F007F7D00F000A000A0";
    attribute INIT_16 of inst : label is "5FF400C0FC000000540003C00000001F00000000000000004000F000000201F0";
    attribute INIT_17 of inst : label is "7FF40A8077740A807FF40200FFFC02000000000000000000000000000F0000AA";
    attribute INIT_18 of inst : label is "B57C2AA0B5782AA001E00A00F5502AA0F5502AA078F002A801782AA005F8AAA8";
    attribute INIT_19 of inst : label is "0000000001400000283C03C0F0F0A0A03DE0A828F13C2A8803C02A00330CA8A0";
    attribute INIT_1A of inst : label is "C3C0ABC13023980009080C40F828F00000010003000000000000000000000000";
    attribute INIT_1B of inst : label is "009807FDC026000000B50000F5F00000000000000000000000000000BC00E000";
    attribute INIT_1C of inst : label is "015F021E0000000055E00000D82F0000260200002D60000063E090000BDA1900";
    attribute INIT_1D of inst : label is "000078FCAE00F000000107C00000003C00003F03007C03E0021C00F0C3C903C0";
    attribute INIT_1E of inst : label is "0000400000002400000000B4000000240500C0F000000003000000000034000F";
    attribute INIT_1F of inst : label is "FFFCFFDC0FFC0FC057F000000000000003C0A00000980000E6C0000000B80000";
    attribute INIT_20 of inst : label is "0000000700000000FC3FFC3F00000000003F003FFC00FC000000D00000000000";
    attribute INIT_21 of inst : label is "06E401D007F402E03F7F02E0FFFFFFFF0000FFFF00000000AAAA00000000D007";
    attribute INIT_22 of inst : label is "000707FFF400FFF4FFE0E0001FFDFFFFFF8080001FFD3FFF00BF000007F409D8";
    attribute INIT_23 of inst : label is "FE00C7F4000000010000D000007F1FFFFF40FFFD2FFEF4002FFE000702FF0002";
    attribute INIT_24 of inst : label is "00B000000BD600000BD600005F80000000030000C003D5570FF0014000000000";
    attribute INIT_25 of inst : label is "00000000000003C000000000000000000BDE000001F800002F5800000B600000";
    attribute INIT_26 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_27 of inst : label is "0000000000F400E009D818C907C002C0F82FC003014003C03C0F2D5E3C0F2D5E";
    attribute INIT_28 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC6832558";
    attribute INIT_29 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_2A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_2B of inst : label is "0000000003FF03FC2FFDFFFFFFFF000003FF0000201E3D573C3C07D00B781E2D";
    attribute INIT_2C of inst : label is "FFD08880A1FF0008F500F7FD0017AA4703FF03C107C0FFC000F408FF03C303FF";
    attribute INIT_2D of inst : label is "2FC30FC303FF03FF3C00FFFF0FF0FFFF0000F0C00000FFFF0000FFFFFFC0FFC0";
    attribute INIT_2E of inst : label is "7FFFFFFFFFFFFFFFFD00FFFFABC00BC0C1FF07FF402FFF03FFF5FC001F003C00";
    attribute INIT_2F of inst : label is "FC07FC00FE00300000020000FFFF8200FFFF0020743FFC3F68F050A803CA0A81";
    attribute INIT_30 of inst : label is "14F480FF001500F2FD3FFEBFFFC0FFFC03FD1FD0FEBF003F47FFFFE0FFFF02BF";
    attribute INIT_31 of inst : label is "00023F4003FF03FF4000FF003FFF3FFF01FF03FFFFFF003FFFFF02BEFFFF002A";
    attribute INIT_32 of inst : label is "04C0000000C40000FD7FFFFFFFFFFFE0FFFF00BFFDFDFFFFA83F083FFF000200";
    attribute INIT_33 of inst : label is "FFFF0000FFC0FAC0FF04AF00E00000BF0000FFC00000001F0000FD00FFC003C0";
    attribute INIT_34 of inst : label is "07FD007E9696F69FD5008000015F000B2CC31D96000000070000F400002F07F4";
    attribute INIT_35 of inst : label is "0000000F0000FC03020001E006BA03E080003F005F570F007F7D00F000A000A0";
    attribute INIT_36 of inst : label is "5FF400C0FC000000540003C00000001F00000000000000004000F000000201F0";
    attribute INIT_37 of inst : label is "7FF40A8077740A807FF40200FFFC02000000000000000000000000000F0000AA";
    attribute INIT_38 of inst : label is "B57C2AA0B5782AA001E00A00F5502AA0F5502AA078F002A801782AA005F8AAA8";
    attribute INIT_39 of inst : label is "0000000001400000283C03C0F0F0A0A03DE0A828F13C2A8803C02A00330CA8A0";
    attribute INIT_3A of inst : label is "C3C0ABC13023980009080C40F828F00000010003000000000000000000000000";
    attribute INIT_3B of inst : label is "009807FDC026000000B50000F5F00000000000000000000000000000BC00E000";
    attribute INIT_3C of inst : label is "015F021E0000000055E00000D82F0000260200002D60000063E090000BDA1900";
    attribute INIT_3D of inst : label is "000078FCAE00F000000107C00000003C00003F03007C03E0021C00F0C3C903C0";
    attribute INIT_3E of inst : label is "0000400000002400000000B4000000240500C0F000000003000000000034000F";
    attribute INIT_3F of inst : label is "FFFCFFDC0FFC0FC057F000000000000003C0A00000980000E6C0000000B80000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "00000000E0000000FC3FFC3F000B0000003F003FFC00FC000000000000000000";
    attribute INIT_01 of inst : label is "00402EEE00402FFE04042FFEFFFFFFFF00005555E00B0000FFFF000000000000";
    attribute INIT_02 of inst : label is "0000007F4000FF40FFFEFE000150FFFFFFF8F80001503FFF0BFF000B00403FFF";
    attribute INIT_03 of inst : label is "FF00E0000000000000004000000707FFF400FFF4FFFFC2A03FFF02A02FFF002F";
    attribute INIT_04 of inst : label is "005000803F0000000F0400A043E0280000000000EAABC003014003C000000000";
    attribute INIT_05 of inst : label is "000000000000000000000AA8C000000007810000001E0000FC0300000F000000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0000000000402AFE10412BFA00402FEAFFFFE00B0000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C943";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "0000000003FF03FE3D005555501FAAAA03FF02AA155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "FFE004E058FF02C43E00E2F0002FFFEF03FF03E081C01FC000D01DFD03C303D7";
    attribute INIT_0D of inst : label is "3F430FC303FF03FF3C007D550FF05FF50000FFC00000FFFF0000FFC3FFC0FFC0";
    attribute INIT_0E of inst : label is "1FF5FFFF7FFDFFFFFC00FFD0FFC00BC040FF03FF0015FC0FFC00FEBF0FF03F00";
    attribute INIT_0F of inst : label is "FC01FC0AFF80BC00000F0000FFFF0000FFFF0000303FFC3F00C094F400C007C5";
    attribute INIT_10 of inst : label is "2FF040FC000E0070D03FFFFF7F40FFF001FC032A5FFF803F01FFDFFEFFFDBFFF";
    attribute INIT_11 of inst : label is "002F340003F403FF0000F4003FF43FFF003F03FFFFFFE03FFFFFFFFFFFFF02FF";
    attribute INIT_12 of inst : label is "FFC0800000FF0000FC3FFFFF7FFFFFFEFFFF2BFFFC00FFFFFC3F083FFF002F00";
    attribute INIT_13 of inst : label is "FFFFAAAAFFC0FFC0FF00FF2EFE00017F0000FFC00000FFFF0000FFFFFFC08BC0";
    attribute INIT_14 of inst : label is "00000A0FF96F69694000F800000500BF04140CC30000000000000000003F0002";
    attribute INIT_15 of inst : label is "000006B700001FA4464002D000300070400007E90F82AFA8003E92FE00F00050";
    attribute INIT_16 of inst : label is "02000002F0002F5E00038F400000000700000000000000000000F0000000EB40";
    attribute INIT_17 of inst : label is "0740BBB80740232007402FE074742FE000000000000000000000000007EA4B40";
    attribute INIT_18 of inst : label is "7AB4503C7AB4F03CEABC0F007AB4F03CFAA8503C07F0AAF87AB4503C7AB47E04";
    attribute INIT_19 of inst : label is "00000000028002801FF401F81F40FAF0BC3C3ED07AB4F0B82BE8F3C071A4330C";
    attribute INIT_1A of inst : label is "01E0D3C07605E003080107007E13F00000000003000000000000000000000000";
    attribute INIT_1B of inst : label is "03C0000000F0000003D1000A147C2A80000000000000000000000000D0003C00";
    attribute INIT_1C of inst : label is "00030EAF00000000001CA800C0FC0002F00300001E04000000F040003F030000";
    attribute INIT_1D of inst : label is "6000B41E0C423C000000AD00000006B7000007EB603C01F8005D007CC3E0FFFE";
    attribute INIT_1E of inst : label is "0000000000000000000000400000000000007AD000000000000000000000A40F";
    attribute INIT_1F of inst : label is "EFFCFFFC0FFE0FEA000002A000000000B7DA0E0043C000000000808000000020";
    attribute INIT_20 of inst : label is "00000000E0000000FC3FFC3F000B0000003F003FFC00FC000000000000000000";
    attribute INIT_21 of inst : label is "00402EEE00402FFE04042FFEFFFFFFFF00005555E00B0000FFFF000000000000";
    attribute INIT_22 of inst : label is "0000007F4000FF40FFFEFE000150FFFFFFF8F80001503FFF0BFF000B00403FFF";
    attribute INIT_23 of inst : label is "FF00E0000000000000004000000707FFF400FFF4FFFFC2A03FFF02A02FFF002F";
    attribute INIT_24 of inst : label is "005000803F0000000F0400A043E0280000000000EAABC003014003C000000000";
    attribute INIT_25 of inst : label is "000000000000000000000AA8C000000007810000001E0000FC0300000F000000";
    attribute INIT_26 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_27 of inst : label is "0000000000402AFE10412BFA00402FEAFFFFE00B0000028005540AAF05541EAD";
    attribute INIT_28 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C943";
    attribute INIT_29 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_2A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_2B of inst : label is "0000000003FF03FE3D005555501FAAAA03FF02AA155507A014140BE0140501D0";
    attribute INIT_2C of inst : label is "FFE004E058FF02C43E00E2F0002FFFEF03FF03E081C01FC000D01DFD03C303D7";
    attribute INIT_2D of inst : label is "3F430FC303FF03FF3C007D550FF05FF50000FFC00000FFFF0000FFC3FFC0FFC0";
    attribute INIT_2E of inst : label is "1FF5FFFF7FFDFFFFFC00FFD0FFC00BC040FF03FF0015FC0FFC00FEBF0FF03F00";
    attribute INIT_2F of inst : label is "FC01FC0AFF80BC00000F0000FFFF0000FFFF0000303FFC3F00C094F400C007C5";
    attribute INIT_30 of inst : label is "2FF040FC000E0070D03FFFFF7F40FFF001FC032A5FFF803F01FFDFFEFFFDBFFF";
    attribute INIT_31 of inst : label is "002F340003F403FF0000F4003FF43FFF003F03FFFFFFE03FFFFFFFFFFFFF02FF";
    attribute INIT_32 of inst : label is "FFC0800000FF0000FC3FFFFF7FFFFFFEFFFF2BFFFC00FFFFFC3F083FFF002F00";
    attribute INIT_33 of inst : label is "FFFFAAAAFFC0FFC0FF00FF2EFE00017F0000FFC00000FFFF0000FFFFFFC08BC0";
    attribute INIT_34 of inst : label is "00000A0FF96F69694000F800000500BF04140CC30000000000000000003F0002";
    attribute INIT_35 of inst : label is "000006B700001FA4464002D000300070400007E90F82AFA8003E92FE00F00050";
    attribute INIT_36 of inst : label is "02000002F0002F5E00038F400000000700000000000000000000F0000000EB40";
    attribute INIT_37 of inst : label is "0740BBB80740232007402FE074742FE000000000000000000000000007EA4B40";
    attribute INIT_38 of inst : label is "7AB4503C7AB4F03CEABC0F007AB4F03CFAA8503C07F0AAF87AB4503C7AB47E04";
    attribute INIT_39 of inst : label is "00000000028002801FF401F81F40FAF0BC3C3ED07AB4F0B82BE8F3C071A4330C";
    attribute INIT_3A of inst : label is "01E0D3C07605E003080107007E13F00000000003000000000000000000000000";
    attribute INIT_3B of inst : label is "03C0000000F0000003D1000A147C2A80000000000000000000000000D0003C00";
    attribute INIT_3C of inst : label is "00030EAF00000000001CA800C0FC0002F00300001E04000000F040003F030000";
    attribute INIT_3D of inst : label is "6000B41E0C423C000000AD00000006B7000007EB603C01F8005D007CC3E0FFFE";
    attribute INIT_3E of inst : label is "0000000000000000000000400000000000007AD000000000000000000000A40F";
    attribute INIT_3F of inst : label is "EFFCFFFC0FFE0FEA000002A000000000B7DA0E0043C000000000808000000020";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "0000000700000000FC3FFC3F00000000003F003FFC00FC000000D00000000000";
    attribute INIT_01 of inst : label is "06E401D007F402E03F7F02E0FFFFFFFF0000FFFF00000000AAAA00000000D007";
    attribute INIT_02 of inst : label is "000707FFF400FFF4FFE0E0001FFDFFFFFF8080001FFD3FFF00BF000007F409D8";
    attribute INIT_03 of inst : label is "FE00C7F4000000010000D000007F1FFFFF40FFFD2FFEF4002FFE000702FF0002";
    attribute INIT_04 of inst : label is "00B000000BD600000BD600005F80000000030000C003D5570FF0014000000000";
    attribute INIT_05 of inst : label is "00000000000003C000000000000000000BDE000001F800002F5800000B600000";
    attribute INIT_06 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_07 of inst : label is "0000000000F400E009D818C907C002C000000000014003C03C0F2D5E3C0F2D5E";
    attribute INIT_08 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC0032558";
    attribute INIT_09 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_0A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_0B of inst : label is "FFF407F8000000032FFD0000EA03000003FF0000201E3D573C3C07D00B781E2D";
    attribute INIT_0C of inst : label is "FFD0F780A1FF0037A0000800000200B803FF03C107C0FFC0200008000000003F";
    attribute INIT_0D of inst : label is "003F003F03FF03FFC000FFFF000FFFFF00000F0000003D1E00000154FFC0FFC0";
    attribute INIT_0E of inst : label is "FFF800002BFF000001FF03FFFEC0FC00FE0AF800BFFF00FFFC0AFC00E000C000";
    attribute INIT_0F of inst : label is "000701FF00000000000000000000FFF800000BFF00000000BF00AE00003F002E";
    attribute INIT_10 of inst : label is "FF007F00000F000DFD00FFC07FFF007F001F1FFF003F003FFFE0F800003F0000";
    attribute INIT_11 of inst : label is "0002FF4003F003F000020000F800C00003C003C0FFFF003FFFFFFD40FFFF0005";
    attribute INIT_12 of inst : label is "FBC07E0000FB002F014003C001FFFFFF3FD0FFFF01FF03FF03C00BC0E0FF00FF";
    attribute INIT_13 of inst : label is "FFFF000014000A00000450001FFFFF400000FFC00000FFE0000002FFFFC003C0";
    attribute INIT_14 of inst : label is "07FD007E1FF40280D5008000015F000B2CC31D96000000070000F400002F07F4";
    attribute INIT_15 of inst : label is "0000000F0000FC03020001E006BA03E080003F005F570F007F7D00F000A000A0";
    attribute INIT_16 of inst : label is "5FF400C0FC000000540003C00000001F00000000000000004000F000000201F0";
    attribute INIT_17 of inst : label is "7FF40A8077740A807FF40200FFFC02000000000000000000000000000F0000AA";
    attribute INIT_18 of inst : label is "B57C2AA0B5782AA001E00A00F5502AA0F5502AA078F002A801782AA005F8AAA8";
    attribute INIT_19 of inst : label is "0000000001400000283C03C0F0F0A0A03DE0A828F13C2A8803C02A00330CA8A0";
    attribute INIT_1A of inst : label is "C3C0ABC13023980009080C40F828F00000010003000000000000000000000000";
    attribute INIT_1B of inst : label is "009807FDC026000000B50000F5F00000000000000000000000000000BC00E000";
    attribute INIT_1C of inst : label is "015F021E0000000055E00000D82F0000260200002D60000063E090000BDA1900";
    attribute INIT_1D of inst : label is "000078FCAE00F000000107C00000003C00003F03007C03E0021C00F0C3C903C0";
    attribute INIT_1E of inst : label is "0000400000002400000000B4000000240500C0F000000003000000000034000F";
    attribute INIT_1F of inst : label is "F8BCFFFC0003003F17F000000000000003C0A00000980000E6C0000000B80000";
    attribute INIT_20 of inst : label is "0000000700000000FC3FFC3F00000000003F003FFC00FC000000D00000000000";
    attribute INIT_21 of inst : label is "06E401D007F402E03F7F02E0FFFFFFFF0000FFFF00000000AAAA00000000D007";
    attribute INIT_22 of inst : label is "000707FFF400FFF4FFE0E0001FFDFFFFFF8080001FFD3FFF00BF000007F409D8";
    attribute INIT_23 of inst : label is "FE00C7F4000000010000D000007F1FFFFF40FFFD2FFEF4002FFE000702FF0002";
    attribute INIT_24 of inst : label is "00B000000BD600000BD600005F80000000030000C003D5570FF0014000000000";
    attribute INIT_25 of inst : label is "00000000000003C000000000000000000BDE000001F800002F5800000B600000";
    attribute INIT_26 of inst : label is "201E03C03C0A2D5E3C002D5E07BC007D280F2D5E281F3F570BC007D03C1F2D5E";
    attribute INIT_27 of inst : label is "0000000000F400E009D818C907C002C000000000014003C03C0F2D5E3C0F2D5E";
    attribute INIT_28 of inst : label is "1E0A0B5F0F121F400F121F570F0F1F5E1E0A0B5E0F0F1F5E1EB43C3CC0032558";
    attribute INIT_29 of inst : label is "1E2D0B783F4F3C0F3F7F3C0F0F001F570F1E1F2D00F02DE003C007D03C3C3C3C";
    attribute INIT_2A of inst : label is "3C4F0FBC3C0F02E03C3C2D7823C807D03C0A2D5E0F0F1F2D3C0F2D590F0F1F40";
    attribute INIT_2B of inst : label is "FFF407F8000000032FFD0000EA03000003FF0000201E3D573C3C07D00B781E2D";
    attribute INIT_2C of inst : label is "FFD0F780A1FF0037A0000800000200B803FF03C107C0FFC0200008000000003F";
    attribute INIT_2D of inst : label is "003F003F03FF03FFC000FFFF000FFFFF00000F0000003D1E00000154FFC0FFC0";
    attribute INIT_2E of inst : label is "FFF800002BFF000001FF03FFFEC0FC00FE0AF800BFFF00FFFC0AFC00E000C000";
    attribute INIT_2F of inst : label is "000701FF00000000000000000000FFF800000BFF00000000BF00AE00003F002E";
    attribute INIT_30 of inst : label is "FF007F00000F000DFD00FFC07FFF007F001F1FFF003F003FFFE0F800003F0000";
    attribute INIT_31 of inst : label is "0002FF4003F003F000020000F800C00003C003C0FFFF003FFFFFFD40FFFF0005";
    attribute INIT_32 of inst : label is "FBC07E0000FB002F014003C001FFFFFF3FD0FFFF01FF03FF03C00BC0E0FF00FF";
    attribute INIT_33 of inst : label is "FFFF000014000A00000450001FFFFF400000FFC00000FFE0000002FFFFC003C0";
    attribute INIT_34 of inst : label is "07FD007E1FF40280D5008000015F000B2CC31D96000000070000F400002F07F4";
    attribute INIT_35 of inst : label is "0000000F0000FC03020001E006BA03E080003F005F570F007F7D00F000A000A0";
    attribute INIT_36 of inst : label is "5FF400C0FC000000540003C00000001F00000000000000004000F000000201F0";
    attribute INIT_37 of inst : label is "7FF40A8077740A807FF40200FFFC02000000000000000000000000000F0000AA";
    attribute INIT_38 of inst : label is "B57C2AA0B5782AA001E00A00F5502AA0F5502AA078F002A801782AA005F8AAA8";
    attribute INIT_39 of inst : label is "0000000001400000283C03C0F0F0A0A03DE0A828F13C2A8803C02A00330CA8A0";
    attribute INIT_3A of inst : label is "C3C0ABC13023980009080C40F828F00000010003000000000000000000000000";
    attribute INIT_3B of inst : label is "009807FDC026000000B50000F5F00000000000000000000000000000BC00E000";
    attribute INIT_3C of inst : label is "015F021E0000000055E00000D82F0000260200002D60000063E090000BDA1900";
    attribute INIT_3D of inst : label is "000078FCAE00F000000107C00000003C00003F03007C03E0021C00F0C3C903C0";
    attribute INIT_3E of inst : label is "0000400000002400000000B4000000240500C0F000000003000000000034000F";
    attribute INIT_3F of inst : label is "F8BCFFFC0003003F17F000000000000003C0A00000980000E6C0000000B80000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "00000000E0000000FC3FFC3F000B0000003F003FFC00FC000000000000000000";
    attribute INIT_01 of inst : label is "00402EEE00402FFE04042FFEFFFFFFFF00005555E00B0000FFFF000000000000";
    attribute INIT_02 of inst : label is "0000007F4000FF40FFFEFE000150FFFFFFF8F80001503FFF0BFF000B00403FFF";
    attribute INIT_03 of inst : label is "FF00E0000000000000004000000707FFF400FFF4FFFFC2A03FFF02A02FFF002F";
    attribute INIT_04 of inst : label is "005000803F0000000F0400A043E0280000000000EAABC003014003C000000000";
    attribute INIT_05 of inst : label is "000000000000000000000AA8C000000007810000001E0000FC0300000F000000";
    attribute INIT_06 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_07 of inst : label is "0000000000402AFE10412BFA00402FEA000000000000028005540AAF05541EAD";
    attribute INIT_08 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C003";
    attribute INIT_09 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_0A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_0B of inst : label is "FF400AFF000A00013F800000FFEB000A03FF02AA155507A014140BE0140501D0";
    attribute INIT_0C of inst : label is "0000FBE0500002FBFE001D00002F001003FF03E081C01FC074001D0000000014";
    attribute INIT_0D of inst : label is "00BF003F03FF03FFC000D555000F555F00005000000050000000003DFFC0FFC0";
    attribute INIT_0E of inst : label is "FFF4FA007FFF02AF000503FFFC00FC80550CFC00FF5503FFFFFFFC00F000C000";
    attribute INIT_0F of inst : label is "0001001F20000000000000000000D75F00003D7500000000FF006B00003F003A";
    attribute INIT_10 of inst : label is "D000BF000001000FD000FFC007FFAA3F000301FFA03F003FFFFEFE00ABFF000B";
    attribute INIT_11 of inst : label is "0007C40003FB03F0002F0000FF80E00003C003C0FFFF003FFFFF0000FFFF0000";
    attribute INIT_12 of inst : label is "FFC0FF0000FF003F000003C0001F1FFFBD00FFFD000503FF03C00BC0FEFF00FF";
    attribute INIT_13 of inst : label is "FFFFAAAA0000AF000000002E81FFFE800000FFC00000000000000000FFC08BC0";
    attribute INIT_14 of inst : label is "00000A0F01402FF84000F800000500BF04140CC30000000000000000003F0002";
    attribute INIT_15 of inst : label is "000006B700001FA4464002D000300070400007E90F82AFA8003E92FE00F00050";
    attribute INIT_16 of inst : label is "02000002F0002F5E00038F400000000700000000000000000000F0000000EB40";
    attribute INIT_17 of inst : label is "0740BBB80740232007402FE074742FE000000000000000000000000007EA4B40";
    attribute INIT_18 of inst : label is "7AB4503C7AB4F03CEABC0F007AB4F03CFAA8503C07F0AAF87AB4503C7AB47E04";
    attribute INIT_19 of inst : label is "00000000028002801FF401F81F40FAF0BC3C3ED07AB4F0B82BE8F3C071A4330C";
    attribute INIT_1A of inst : label is "01E0D3C07605E003080107007E13F00000000003000000000000000000000000";
    attribute INIT_1B of inst : label is "03C0000000F0000003D1000A147C2A80000000000000000000000000D0003C00";
    attribute INIT_1C of inst : label is "00030EAF00000000001CA800C0FC0002F00300001E04000000F040003F030000";
    attribute INIT_1D of inst : label is "6000B41E0C423C000000AD00000006B7000007EB603C01F8005D007CC3E0FFFE";
    attribute INIT_1E of inst : label is "0000000000000000000000400000000000007AD000000000000000000000A40F";
    attribute INIT_1F of inst : label is "FFFCF47C000B00BFA80A02A000000000B7DA0E0043C000000000808000000020";
    attribute INIT_20 of inst : label is "00000000E0000000FC3FFC3F000B0000003F003FFC00FC000000000000000000";
    attribute INIT_21 of inst : label is "00402EEE00402FFE04042FFEFFFFFFFF00005555E00B0000FFFF000000000000";
    attribute INIT_22 of inst : label is "0000007F4000FF40FFFEFE000150FFFFFFF8F80001503FFF0BFF000B00403FFF";
    attribute INIT_23 of inst : label is "FF00E0000000000000004000000707FFF400FFF4FFFFC2A03FFF02A02FFF002F";
    attribute INIT_24 of inst : label is "005000803F0000000F0400A043E0280000000000EAABC003014003C000000000";
    attribute INIT_25 of inst : label is "000000000000000000000AA8C000000007810000001E0000FC0300000F000000";
    attribute INIT_26 of inst : label is "155501E005543EAD15552AAD00543D7D055400AD055407E8014003C005543D8F";
    attribute INIT_27 of inst : label is "0000000000402AFE10412BFA00402FEA000000000000028005540AAF05541EAD";
    attribute INIT_28 of inst : label is "01543C2F15550FB015550FB015540F0F01543C0015540FAD01403D7C1AA4C003";
    attribute INIT_29 of inst : label is "01503C0F14053CBF14053EEF15400F0015050FF0055514F0055003C014143EBC";
    attribute INIT_2A of inst : label is "14053CCF14052D1E14143C3C155403C005540AAD15540FF805543C1F15540FA8";
    attribute INIT_2B of inst : label is "FF400AFF000A00013F800000FFEB000A03FF02AA155507A014140BE0140501D0";
    attribute INIT_2C of inst : label is "0000FBE0500002FBFE001D00002F001003FF03E081C01FC074001D0000000014";
    attribute INIT_2D of inst : label is "00BF003F03FF03FFC000D555000F555F00005000000050000000003DFFC0FFC0";
    attribute INIT_2E of inst : label is "FFF4FA007FFF02AF000503FFFC00FC80550CFC00FF5503FFFFFFFC00F000C000";
    attribute INIT_2F of inst : label is "0001001F20000000000000000000D75F00003D7500000000FF006B00003F003A";
    attribute INIT_30 of inst : label is "D000BF000001000FD000FFC007FFAA3F000301FFA03F003FFFFEFE00ABFF000B";
    attribute INIT_31 of inst : label is "0007C40003FB03F0002F0000FF80E00003C003C0FFFF003FFFFF0000FFFF0000";
    attribute INIT_32 of inst : label is "FFC0FF0000FF003F000003C0001F1FFFBD00FFFD000503FF03C00BC0FEFF00FF";
    attribute INIT_33 of inst : label is "FFFFAAAA0000AF000000002E81FFFE800000FFC00000000000000000FFC08BC0";
    attribute INIT_34 of inst : label is "00000A0F01402FF84000F800000500BF04140CC30000000000000000003F0002";
    attribute INIT_35 of inst : label is "000006B700001FA4464002D000300070400007E90F82AFA8003E92FE00F00050";
    attribute INIT_36 of inst : label is "02000002F0002F5E00038F400000000700000000000000000000F0000000EB40";
    attribute INIT_37 of inst : label is "0740BBB80740232007402FE074742FE000000000000000000000000007EA4B40";
    attribute INIT_38 of inst : label is "7AB4503C7AB4F03CEABC0F007AB4F03CFAA8503C07F0AAF87AB4503C7AB47E04";
    attribute INIT_39 of inst : label is "00000000028002801FF401F81F40FAF0BC3C3ED07AB4F0B82BE8F3C071A4330C";
    attribute INIT_3A of inst : label is "01E0D3C07605E003080107007E13F00000000003000000000000000000000000";
    attribute INIT_3B of inst : label is "03C0000000F0000003D1000A147C2A80000000000000000000000000D0003C00";
    attribute INIT_3C of inst : label is "00030EAF00000000001CA800C0FC0002F00300001E04000000F040003F030000";
    attribute INIT_3D of inst : label is "6000B41E0C423C000000AD00000006B7000007EB603C01F8005D007CC3E0FFFE";
    attribute INIT_3E of inst : label is "0000000000000000000000400000000000007AD000000000000000000000A40F";
    attribute INIT_3F of inst : label is "FFFCF47C000B00BFA80A02A000000000B7DA0E0043C000000000808000000020";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
