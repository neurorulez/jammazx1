-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_8K is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(11 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_8K is

	signal rom_addr : std_logic_vector(11 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(11 downto 0) <= ADDR;
	end process;

	ROM_8K_0 : RAMB16_S4
	generic map (
		INIT_00 => x"FFFFFFFF00000000FFFFFFFF0000000000000000000000000000000000000000",
		INIT_01 => x"0000DFFC000023F7FFD00000F3200000FFFFFFFF00000000FFFFFFFF00000000",
		INIT_02 => x"FF333333FF00FF0033333333FF333333FF00FF00FF00FFCCFF00FFFFCCCCCCCC",
		INIT_03 => x"FFFF00FFCCCCCCCC00FF00FFCCFF00FF33333333333333FF333333FF00FF00FF",
		INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => x"000000000660000000000000000000000000000000000000026C800000008C62",
		INIT_06 => x"000EE0000CE222EC046222EC08888EE8046222EC06EEAA22022EE22008C622C8",
		INIT_07 => x"00AA00000EE0000000000000EE00AAEE0C2EAA2C0C2AAA2C002226C80CE222EC",
		INIT_08 => x"08C622EE0EE000000EE222200EE226C808C622640EE222EC0EE888EE00000000",
		INIT_09 => x"0CE222EC0EE08CEE0EE080EE0EE222200EE8CE62046222EC022EE2200EE000EE",
		INIT_0A => x"0CEC8CEC008CEC800CE222EC000EE000046222EC0EE8CE620CE2AECA0EE88880",
		INIT_0B => x"F1111111F00000001111111F0000000F0000000006EEA222000EE00006EC8CE6",
		INIT_0C => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_0D => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_0E => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_0F => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_10 => x"00000000000000130000000037300000000000080000037C8000000081200000",
		INIT_11 => x"0084211178000000111248000000008700000844003480004480000000084300",
		INIT_12 => x"00088033000933776EC800007003180000000EFF00408FFF000000004C880000",
		INIT_13 => x"0000000000000000000000000000000000088033004137776EC8000038039000",
		INIT_14 => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_15 => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_16 => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_17 => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_18 => x"333BBBBB00066FF0B333FFFF0000FFFFFFFF3333FFFF0000B33333B321000120",
		INIT_19 => x"333BBBBB00888BBBBB33FFFFFFC0FFFF33BBBBBB00EEC889BBB3FFFFDFF0FFFF",
		INIT_1A => x"333BBBBB00FFBBBBBB33FFFFBB10FFFF33333333000137ECBB33FFFFFF00FFFF",
		INIT_1B => x"FFFF0000FFFF0000FFFF0000FF00000000000000FFFF0000FFFF0000FFFF0000",
		INIT_1C => x"000000000000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFF0000FF000000",
		INIT_1D => x"0000FFFF0000FFFF0000FFFF000000FF0000FFFF0000FFFF0000FFFF000000FF",
		INIT_1E => x"8800000088888888000000080F0F0F00000F0F0FAB4B4300AAAAAAAA00034B4B",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"000000000000000045300100EF3004F008F313E8223333760000880000000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"FF00FF00FF00FF00FF00FFFFFF00FFFFFFFFFFFFCCCCCCCCFFFFFFFFCCCCCCCC",
		INIT_23 => x"FFFF00FFFFFF00FF00FF00FF00FF00FF33333333333333333333333333333333",
		INIT_24 => x"111119990000000099999999000000000C623111F00800001111111100000000",
		INIT_25 => x"99999999FFFFFFFF99911111FFFFFFFF9999999901113377999999997FFFFFFF",
		INIT_26 => x"99111111C800017F11111111FE80003F11111999FFEC800099999999001339CE",
		INIT_27 => x"1999999908EFFF70999911110008888F11111199F000FFE09999111100000100",
		INIT_28 => x"11111999CEFFFFEC1111111100FFFFF011199999FFFF7310999991110000088C",
		INIT_29 => x"111119994CEFFFFF991326C0FFFFF00F11111111000C60001111111100004447",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_2D => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_2E => x"F00F0F0FF00F0F0FE00F0F0EF00F0F0F55555555555555555555555445555555",
		INIT_2F => x"5555555554070745544F0F0FF00F074555555D1FF11D555554470F0FF00F0745",
		INIT_30 => x"00000000000036C8000000008C63000000000000005570740000000070747000",
		INIT_31 => x"0084211178000000111248000000008700000844003480004480000000084300",
		INIT_32 => x"0000484000EAA0E2044C0000E0E2E0000000484000EAA0E20C440000E0E2E000",
		INIT_33 => x"0000484000EAA0E2044C0000E0E2E0000000484000EAA0E2000C0000E0E2E000",
		INIT_34 => x"F1111F1FF1F33F1FF1333F1FF1D5F51F3333333333333333333333FFFF333333",
		INIT_35 => x"F1F1111FF1F3331FF1F33F1FF1F3371FF1F33F1FF1F11F1FF1333F1FF1F33F1F",
		INIT_36 => x"F1111F1FF1F33F1FF1333F1FF1D5F51FF1733F1FF1FBBB1FF113F31FF1F33F1F",
		INIT_37 => x"F1F1111FF1F3331FF1F33F1FF1F3371FF1F33F1FF1F11F1FF1333F1FF1F33F1F",
		INIT_38 => x"0000000400001337C8000000F001000000000EFF00000FFF000000004C800000",
		INIT_39 => x"00088033000133776EC8000070031000000880330001337F6EC8000030031000",
		INIT_3A => x"0000CEEF00000113FEEC000031100000000000CC00000073EE0C000031430000",
		INIT_3B => x"0000CEEF00000113FEEC0000311000000000CEEF00000113FEEC000031100000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0000",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8K_1 : RAMB16_S4
	generic map (
		INIT_00 => x"FFFFFFFF00000000FFFFFFFF0000000000000000000000000000000000000000",
		INIT_01 => x"037EE6670000000066EE730000000000FFFFFFFF00000000FFFFFFFF00000000",
		INIT_02 => x"FF00FF33FF00FF0033333333FF00FFFFFF00FF00FFCCCCCCFFCCCCCCCCCCCCCC",
		INIT_03 => x"CCCCCCFFCCCCCCCC00FF00FFCCCCCCFF33333333FFFF00FF33FF00FF00FF00FF",
		INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => x"00000000000000000111111000000000000000000000000008C73000000037C8",
		INIT_06 => x"0CC89BEC037D99900EEAAAB90136CFF00089BFD804C99BF6004FF00003788C73",
		INIT_07 => x"00FFF00007755702000CE00077203322078BAB87078BAA8706F999F706F999F6",
		INIT_08 => x"037C89990FF999980FF999800FF88C73037C88C40FF999F6037C8C7300000000",
		INIT_09 => x"07F888F70FF731FF0FF737FF0FF000000FF136C8000000FF088FF8800FF111FF",
		INIT_0A => x"0FF131FF0FF101FF0FF000FF088FF88006F999D40FF889F707F888F70FF88887",
		INIT_0B => x"F0000000F88888880000000F8888888F000000000889BFEC0CF11FC00CE737EC",
		INIT_0C => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_0D => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_0E => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_0F => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_10 => x"000004EE00000000EEC000000000000000002EC1000000003C00000000000000",
		INIT_11 => x"E1000000001248880000001E8884210000C210000000012200012C0022100000",
		INIT_12 => x"007FFFFE00008050803FE4002050800000000FFF20200A250000000025A28002",
		INIT_13 => x"00000000000000000000000000000000007FFFFE20128212803FE4004A500400",
		INIT_14 => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_15 => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_16 => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_17 => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_18 => x"00011FF1CCCCCDDC1000FFFFCCCCFFFFFFFF0000FFFFCCCC01A4A100CCCCCCCC",
		INIT_19 => x"00773113CCDDDDDDFFF0FFFFDDDCFFFF00137FFDCCCDDDDD9910FFFFDDCCFFFF",
		INIT_1A => x"00773111CCDDDDDDBFF0FFFFDDCCFFFF00EEE666CCCCCCCDFF60FFFFDDCCFFFF",
		INIT_1B => x"FFFF0000FFFF0000FFFF0000FF00000000000000FFFF0000FFFF0000FFFF0000",
		INIT_1C => x"000000000000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFF0000FF000000",
		INIT_1D => x"0000FFFF0000FFFF0000FFFF000000FF0000FFFF0000FFFF0000FFFF000000FF",
		INIT_1E => x"AA5A4800AAAAAAAA00084A5A0F0F0F00000F0F0F221000002222222200000012",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"000000000000000001EC0000136CC2000D100CD5000000002201100000000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"FF00FF00FF00FF00FF00FFFFFF00FFFFCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC",
		INIT_23 => x"FFFF00FFFFFF00FF00FF00FF00FF00FF33333333FFFFFFFF33333333FFFFFFFF",
		INIT_24 => x"00000001888800001133777F00000000F1000000F00FFFFF00000000EEEECCCC",
		INIT_25 => x"FFFFFFFF777FFFFFFFFFEEC8FFFFFFFFFFFFFFFF00000000FFFFFFFF00011133",
		INIT_26 => x"3100CCEE7FFE8000800006EE3772888180000013FFFFFFFE7FFFFFF7C0000013",
		INIT_27 => x"000888806FFF310800310008CEF3FFF7E00080007000FFF01373888008E00000",
		INIT_28 => x"00000001137FF7304CCCCC0003111000888888883100008C00000000CEEFFF30",
		INIT_29 => x"0000EFFFFFFFFFFFFFFEC01FFFFFF00F0000000000010000C444000E0000008C",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_2D => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_2E => x"F00F0F0FF00F0F0FF00F0F0F700F0F0799999999999999999999999119999999",
		INIT_2F => x"911F1F1999999999911F0F0FF00F0D19911F0F0FF00F0F199999998FF8899999",
		INIT_30 => x"0000C63100000000136C00000000000000C440C400000000C0C4C00000000000",
		INIT_31 => x"E1000000001248880000001E8884210000C210000000012200012C0022100000",
		INIT_32 => x"0000101000223032055700003032300000001010002230320557000030323000",
		INIT_33 => x"0000101000223032075500003032300000001010002230320717000030323000",
		INIT_34 => x"F8CCCF8FF8FDDD8FF8FDDD8FF8F8988FCCCCCCCCCCCCCCCCCCCCCCFFFFCCCCCC",
		INIT_35 => x"F8FDDC8FF8FDDC8FF8999F8FF8FCCE8FF8F9998FF8FDDF8FF8FDDF8FF8FDDF8F",
		INIT_36 => x"F8CCCF8FF8FDDD8FF8FDDD8FF8F8988FF8ECDF8FF8ECCF8FF88AF88FF8FCCF8F",
		INIT_37 => x"F8FDDC8FF8FDDC8FF8999F8FF8FCCE8FF8F9998FF8FDDF8FF8FDDF8FF8FDDF8F",
		INIT_38 => x"0006FFEC00000005837E00002000000000000FFF000000170000000001000000",
		INIT_39 => x"007FFFFE00000000803FE40000000000007FFFFE00000002803FE40010000000",
		INIT_3A => x"0003FFFF00000000FFFF300000000000000000FF00000000FF5F500000000000",
		INIT_3B => x"0003FFFF00000000FFFF3000000000000003FFFF00000000FFFF300000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "0000",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
