-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"c4080b0b",
    10 => x"0bb5c808",
    11 => x"0b0b0bb5",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5cc0c0b",
    16 => x"0b0bb5c8",
    17 => x"0c0b0b0b",
    18 => x"b5c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafb0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5c470bf",
    57 => x"f4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"88be0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5d40c9f",
    65 => x"0bb5d80c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"d808ff05",
    69 => x"b5d80cb5",
    70 => x"d8088025",
    71 => x"eb38b5d4",
    72 => x"08ff05b5",
    73 => x"d40cb5d4",
    74 => x"088025d7",
    75 => x"38800bb5",
    76 => x"d80c800b",
    77 => x"b5d40c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"b5d40825",
    97 => x"8f3882bc",
    98 => x"2db5d408",
    99 => x"ff05b5d4",
   100 => x"0c82fe04",
   101 => x"b5d408b5",
   102 => x"d8085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038b5",
   107 => x"d408a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34b5d808",
   111 => x"8105b5d8",
   112 => x"0cb5d808",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"b5d80cb5",
   116 => x"d4088105",
   117 => x"b5d40c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134b5d8",
   122 => x"088105b5",
   123 => x"d80cb5d8",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800bb5d8",
   127 => x"0cb5d408",
   128 => x"8105b5d4",
   129 => x"0c028c05",
   130 => x"0d0402e8",
   131 => x"050d7779",
   132 => x"5656880b",
   133 => x"fc167771",
   134 => x"2c8f0654",
   135 => x"52548053",
   136 => x"72722595",
   137 => x"387153fb",
   138 => x"e0145187",
   139 => x"71348114",
   140 => x"ff145454",
   141 => x"72f13871",
   142 => x"53f91576",
   143 => x"712c8706",
   144 => x"53517180",
   145 => x"2e8b38fb",
   146 => x"e0145171",
   147 => x"71348114",
   148 => x"54728e24",
   149 => x"95388f73",
   150 => x"3153fbe0",
   151 => x"1451a071",
   152 => x"348114ff",
   153 => x"14545472",
   154 => x"f1380298",
   155 => x"050d0402",
   156 => x"ec050d80",
   157 => x"0bb5dc0c",
   158 => x"f68c08f6",
   159 => x"90087188",
   160 => x"2c565481",
   161 => x"ff065273",
   162 => x"72258838",
   163 => x"7154820b",
   164 => x"b5dc0c72",
   165 => x"882c7381",
   166 => x"ff065455",
   167 => x"7473258b",
   168 => x"3872b5dc",
   169 => x"088407b5",
   170 => x"dc0c5573",
   171 => x"842b86a0",
   172 => x"71258371",
   173 => x"31700b0b",
   174 => x"0bb2980c",
   175 => x"81712bff",
   176 => x"05f6880c",
   177 => x"fdfc13ff",
   178 => x"122c7888",
   179 => x"29ff9405",
   180 => x"70812cb5",
   181 => x"dc085258",
   182 => x"52555152",
   183 => x"5476802e",
   184 => x"85387081",
   185 => x"075170f6",
   186 => x"940c7109",
   187 => x"8105f680",
   188 => x"0c720981",
   189 => x"05f6840c",
   190 => x"0294050d",
   191 => x"0402f405",
   192 => x"0d745372",
   193 => x"70810554",
   194 => x"80f52d52",
   195 => x"71802e89",
   196 => x"38715182",
   197 => x"f82d8683",
   198 => x"04810bb5",
   199 => x"c40c028c",
   200 => x"050d0402",
   201 => x"fc050d81",
   202 => x"808051c0",
   203 => x"115170fb",
   204 => x"38028405",
   205 => x"0d0402fc",
   206 => x"050d84bf",
   207 => x"5186a32d",
   208 => x"ff115170",
   209 => x"8025f638",
   210 => x"0284050d",
   211 => x"0402fc05",
   212 => x"0dec5183",
   213 => x"710c86a3",
   214 => x"2d82710c",
   215 => x"0284050d",
   216 => x"0402fc05",
   217 => x"0dec5192",
   218 => x"710c86a3",
   219 => x"2d82710c",
   220 => x"0284050d",
   221 => x"0402fc05",
   222 => x"0dec51a2",
   223 => x"710c86a3",
   224 => x"2d82710c",
   225 => x"0284050d",
   226 => x"0402dc05",
   227 => x"0d805984",
   228 => x"0bec0ca0",
   229 => x"0bec0c7a",
   230 => x"52b5e051",
   231 => x"a6ec2db5",
   232 => x"c408792e",
   233 => x"80eb38b5",
   234 => x"e40879ff",
   235 => x"12565956",
   236 => x"73792e8b",
   237 => x"38811874",
   238 => x"812a5558",
   239 => x"73f738f7",
   240 => x"18588159",
   241 => x"80762580",
   242 => x"c8387752",
   243 => x"7351848a",
   244 => x"2db6ac52",
   245 => x"b5e051a9",
   246 => x"a22db5c4",
   247 => x"08802e9a",
   248 => x"38b6ac57",
   249 => x"83fc5576",
   250 => x"70840558",
   251 => x"08e80cfc",
   252 => x"15557480",
   253 => x"25f13888",
   254 => x"8104b5c4",
   255 => x"08598480",
   256 => x"56b5e051",
   257 => x"a8f52dfc",
   258 => x"80168115",
   259 => x"555687c4",
   260 => x"04b5e408",
   261 => x"f80c86b6",
   262 => x"2d805186",
   263 => x"f52d7880",
   264 => x"2e8d38b2",
   265 => x"9c518fca",
   266 => x"2d8dcd2d",
   267 => x"88b504b3",
   268 => x"94518fca",
   269 => x"2d78b5c4",
   270 => x"0c02a405",
   271 => x"0d0402f0",
   272 => x"050d840b",
   273 => x"ec0c8dae",
   274 => x"2d89fd2d",
   275 => x"81f72d83",
   276 => x"528d932d",
   277 => x"815184ef",
   278 => x"2dff1252",
   279 => x"718025f1",
   280 => x"38840bec",
   281 => x"0cb0cc51",
   282 => x"85fd2d9e",
   283 => x"892db5c4",
   284 => x"08802e80",
   285 => x"f3388789",
   286 => x"51afa92d",
   287 => x"b29c518f",
   288 => x"ca2d8dcd",
   289 => x"2d8a892d",
   290 => x"8fda2db2",
   291 => x"b00b80f5",
   292 => x"2db48008",
   293 => x"70810654",
   294 => x"55537180",
   295 => x"2e853872",
   296 => x"81075373",
   297 => x"812a7081",
   298 => x"06515271",
   299 => x"802e8538",
   300 => x"72820753",
   301 => x"73822a70",
   302 => x"81065152",
   303 => x"71802e85",
   304 => x"38728407",
   305 => x"5373832a",
   306 => x"70810651",
   307 => x"5271802e",
   308 => x"85387288",
   309 => x"075372fc",
   310 => x"0c8652b5",
   311 => x"c4088338",
   312 => x"845271ec",
   313 => x"0c898504",
   314 => x"800bb5c4",
   315 => x"0c029005",
   316 => x"0d047198",
   317 => x"0c04ffb0",
   318 => x"08b5c40c",
   319 => x"04810bff",
   320 => x"b00c0480",
   321 => x"0bffb00c",
   322 => x"0402f405",
   323 => x"0d8b8b04",
   324 => x"b5c40881",
   325 => x"f02e0981",
   326 => x"06893881",
   327 => x"0bb3f80c",
   328 => x"8b8b04b5",
   329 => x"c40881e0",
   330 => x"2e098106",
   331 => x"8938810b",
   332 => x"b3fc0c8b",
   333 => x"8b04b5c4",
   334 => x"0852b3fc",
   335 => x"08802e88",
   336 => x"38b5c408",
   337 => x"81800552",
   338 => x"71842c72",
   339 => x"8f065353",
   340 => x"b3f80880",
   341 => x"2e993872",
   342 => x"8429b3b8",
   343 => x"05721381",
   344 => x"712b7009",
   345 => x"73080673",
   346 => x"0c515353",
   347 => x"8b810472",
   348 => x"8429b3b8",
   349 => x"05721383",
   350 => x"712b7208",
   351 => x"07720c53",
   352 => x"53800bb3",
   353 => x"fc0c800b",
   354 => x"b3f80cb5",
   355 => x"ec518c8c",
   356 => x"2db5c408",
   357 => x"ff24fef8",
   358 => x"38800bb5",
   359 => x"c40c028c",
   360 => x"050d0402",
   361 => x"f8050db3",
   362 => x"b8528f51",
   363 => x"80727084",
   364 => x"05540cff",
   365 => x"11517080",
   366 => x"25f23802",
   367 => x"88050d04",
   368 => x"02f0050d",
   369 => x"75518a83",
   370 => x"2d70822c",
   371 => x"fc06b3b8",
   372 => x"1172109e",
   373 => x"06710870",
   374 => x"722a7083",
   375 => x"0682742b",
   376 => x"70097406",
   377 => x"760c5451",
   378 => x"56575351",
   379 => x"5389fd2d",
   380 => x"71b5c40c",
   381 => x"0290050d",
   382 => x"0402fc05",
   383 => x"0d725180",
   384 => x"710c800b",
   385 => x"84120c02",
   386 => x"84050d04",
   387 => x"02f0050d",
   388 => x"75700884",
   389 => x"12085353",
   390 => x"53ff5471",
   391 => x"712ea838",
   392 => x"8a832d84",
   393 => x"13087084",
   394 => x"29148811",
   395 => x"70087081",
   396 => x"ff068418",
   397 => x"08811187",
   398 => x"06841a0c",
   399 => x"53515551",
   400 => x"515189fd",
   401 => x"2d715473",
   402 => x"b5c40c02",
   403 => x"90050d04",
   404 => x"02f8050d",
   405 => x"8a832de0",
   406 => x"08708b2a",
   407 => x"70810651",
   408 => x"52527080",
   409 => x"2e9d38b5",
   410 => x"ec087084",
   411 => x"29b5f405",
   412 => x"7381ff06",
   413 => x"710c5151",
   414 => x"b5ec0881",
   415 => x"118706b5",
   416 => x"ec0c5180",
   417 => x"0bb6940c",
   418 => x"89f62d89",
   419 => x"fd2d0288",
   420 => x"050d0402",
   421 => x"fc050d8a",
   422 => x"832d810b",
   423 => x"b6940c89",
   424 => x"fd2db694",
   425 => x"085170fa",
   426 => x"38028405",
   427 => x"0d0402fc",
   428 => x"050db5ec",
   429 => x"518bf92d",
   430 => x"8ba32d8c",
   431 => x"d05189f2",
   432 => x"2d028405",
   433 => x"0d04b698",
   434 => x"08b5c40c",
   435 => x"0402fc05",
   436 => x"0d8dd704",
   437 => x"8a892d80",
   438 => x"f6518bc0",
   439 => x"2db5c408",
   440 => x"f33880da",
   441 => x"518bc02d",
   442 => x"b5c408e8",
   443 => x"38b5c408",
   444 => x"b4840cb5",
   445 => x"c4085184",
   446 => x"ef2d0284",
   447 => x"050d0402",
   448 => x"ec050d76",
   449 => x"54805287",
   450 => x"0b881580",
   451 => x"f52d5653",
   452 => x"74722483",
   453 => x"38a05372",
   454 => x"5182f82d",
   455 => x"81128b15",
   456 => x"80f52d54",
   457 => x"52727225",
   458 => x"de380294",
   459 => x"050d0402",
   460 => x"f0050db6",
   461 => x"98085481",
   462 => x"f72d800b",
   463 => x"b69c0c73",
   464 => x"08802e81",
   465 => x"8038820b",
   466 => x"b5d80cb6",
   467 => x"9c088f06",
   468 => x"b5d40c73",
   469 => x"08527183",
   470 => x"2e963871",
   471 => x"83268938",
   472 => x"71812eaf",
   473 => x"388fb004",
   474 => x"71852e9f",
   475 => x"388fb004",
   476 => x"881480f5",
   477 => x"2d841508",
   478 => x"b0e45354",
   479 => x"5285fd2d",
   480 => x"71842913",
   481 => x"70085252",
   482 => x"8fb40473",
   483 => x"518dff2d",
   484 => x"8fb004b4",
   485 => x"80088815",
   486 => x"082c7081",
   487 => x"06515271",
   488 => x"802e8738",
   489 => x"b0e8518f",
   490 => x"ad04b0ec",
   491 => x"5185fd2d",
   492 => x"84140851",
   493 => x"85fd2db6",
   494 => x"9c088105",
   495 => x"b69c0c8c",
   496 => x"14548ebf",
   497 => x"04029005",
   498 => x"0d0471b6",
   499 => x"980c8eaf",
   500 => x"2db69c08",
   501 => x"ff05b6a0",
   502 => x"0c0402e8",
   503 => x"050db698",
   504 => x"08b6a408",
   505 => x"57558751",
   506 => x"8bc02db5",
   507 => x"c408812a",
   508 => x"70810651",
   509 => x"5271802e",
   510 => x"a0389080",
   511 => x"048a892d",
   512 => x"87518bc0",
   513 => x"2db5c408",
   514 => x"f438b484",
   515 => x"08813270",
   516 => x"b4840c70",
   517 => x"525284ef",
   518 => x"2d80fe51",
   519 => x"8bc02db5",
   520 => x"c408802e",
   521 => x"a638b484",
   522 => x"08802e91",
   523 => x"38800bb4",
   524 => x"840c8051",
   525 => x"84ef2d90",
   526 => x"bd048a89",
   527 => x"2d80fe51",
   528 => x"8bc02db5",
   529 => x"c408f338",
   530 => x"86e12db4",
   531 => x"84089038",
   532 => x"81fd518b",
   533 => x"c02d81fa",
   534 => x"518bc02d",
   535 => x"96900481",
   536 => x"f5518bc0",
   537 => x"2db5c408",
   538 => x"812a7081",
   539 => x"06515271",
   540 => x"802eaf38",
   541 => x"b6a00852",
   542 => x"71802e89",
   543 => x"38ff12b6",
   544 => x"a00c91a2",
   545 => x"04b69c08",
   546 => x"10b69c08",
   547 => x"05708429",
   548 => x"16515288",
   549 => x"1208802e",
   550 => x"8938ff51",
   551 => x"88120852",
   552 => x"712d81f2",
   553 => x"518bc02d",
   554 => x"b5c40881",
   555 => x"2a708106",
   556 => x"51527180",
   557 => x"2eb138b6",
   558 => x"9c08ff11",
   559 => x"b6a00856",
   560 => x"53537372",
   561 => x"25893881",
   562 => x"14b6a00c",
   563 => x"91e70472",
   564 => x"10137084",
   565 => x"29165152",
   566 => x"88120880",
   567 => x"2e8938fe",
   568 => x"51881208",
   569 => x"52712d81",
   570 => x"fd518bc0",
   571 => x"2db5c408",
   572 => x"812a7081",
   573 => x"06515271",
   574 => x"802ead38",
   575 => x"b6a00880",
   576 => x"2e893880",
   577 => x"0bb6a00c",
   578 => x"92a804b6",
   579 => x"9c0810b6",
   580 => x"9c080570",
   581 => x"84291651",
   582 => x"52881208",
   583 => x"802e8938",
   584 => x"fd518812",
   585 => x"0852712d",
   586 => x"81fa518b",
   587 => x"c02db5c4",
   588 => x"08812a70",
   589 => x"81065152",
   590 => x"71802eae",
   591 => x"38b69c08",
   592 => x"ff115452",
   593 => x"b6a00873",
   594 => x"25883872",
   595 => x"b6a00c92",
   596 => x"ea047110",
   597 => x"12708429",
   598 => x"16515288",
   599 => x"1208802e",
   600 => x"8938fc51",
   601 => x"88120852",
   602 => x"712db6a0",
   603 => x"08705354",
   604 => x"73802e8a",
   605 => x"388c15ff",
   606 => x"15555592",
   607 => x"f004820b",
   608 => x"b5d80c71",
   609 => x"8f06b5d4",
   610 => x"0c81eb51",
   611 => x"8bc02db5",
   612 => x"c408812a",
   613 => x"70810651",
   614 => x"5271802e",
   615 => x"ad387408",
   616 => x"852e0981",
   617 => x"06a43888",
   618 => x"1580f52d",
   619 => x"ff055271",
   620 => x"881681b7",
   621 => x"2d71982b",
   622 => x"52718025",
   623 => x"8838800b",
   624 => x"881681b7",
   625 => x"2d74518d",
   626 => x"ff2d81f4",
   627 => x"518bc02d",
   628 => x"b5c40881",
   629 => x"2a708106",
   630 => x"51527180",
   631 => x"2eb33874",
   632 => x"08852e09",
   633 => x"8106aa38",
   634 => x"881580f5",
   635 => x"2d810552",
   636 => x"71881681",
   637 => x"b72d7181",
   638 => x"ff068b16",
   639 => x"80f52d54",
   640 => x"52727227",
   641 => x"87387288",
   642 => x"1681b72d",
   643 => x"74518dff",
   644 => x"2d80da51",
   645 => x"8bc02db5",
   646 => x"c408812a",
   647 => x"70810651",
   648 => x"5271802e",
   649 => x"81a638b6",
   650 => x"9808b6a0",
   651 => x"08555373",
   652 => x"802e8a38",
   653 => x"8c13ff15",
   654 => x"555394af",
   655 => x"04720852",
   656 => x"71822ea6",
   657 => x"38718226",
   658 => x"89387181",
   659 => x"2ea93895",
   660 => x"cc047183",
   661 => x"2eb13871",
   662 => x"842e0981",
   663 => x"0680ed38",
   664 => x"88130851",
   665 => x"8fca2d95",
   666 => x"cc04b6a0",
   667 => x"08518813",
   668 => x"0852712d",
   669 => x"95cc0481",
   670 => x"0b881408",
   671 => x"2bb48008",
   672 => x"32b4800c",
   673 => x"95a20488",
   674 => x"1380f52d",
   675 => x"81058b14",
   676 => x"80f52d53",
   677 => x"54717424",
   678 => x"83388054",
   679 => x"73881481",
   680 => x"b72d8eaf",
   681 => x"2d95cc04",
   682 => x"7508802e",
   683 => x"a2387508",
   684 => x"518bc02d",
   685 => x"b5c40881",
   686 => x"06527180",
   687 => x"2e8b38b6",
   688 => x"a0085184",
   689 => x"16085271",
   690 => x"2d881656",
   691 => x"75da3880",
   692 => x"54800bb5",
   693 => x"d80c738f",
   694 => x"06b5d40c",
   695 => x"a05273b6",
   696 => x"a0082e09",
   697 => x"81069838",
   698 => x"b69c08ff",
   699 => x"05743270",
   700 => x"09810570",
   701 => x"72079f2a",
   702 => x"91713151",
   703 => x"51535371",
   704 => x"5182f82d",
   705 => x"8114548e",
   706 => x"7425c638",
   707 => x"b4840852",
   708 => x"71b5c40c",
   709 => x"0298050d",
   710 => x"0402f405",
   711 => x"0dd45281",
   712 => x"ff720c71",
   713 => x"085381ff",
   714 => x"720c7288",
   715 => x"2b83fe80",
   716 => x"06720870",
   717 => x"81ff0651",
   718 => x"525381ff",
   719 => x"720c7271",
   720 => x"07882b72",
   721 => x"087081ff",
   722 => x"06515253",
   723 => x"81ff720c",
   724 => x"72710788",
   725 => x"2b720870",
   726 => x"81ff0672",
   727 => x"07b5c40c",
   728 => x"5253028c",
   729 => x"050d0402",
   730 => x"f4050d74",
   731 => x"767181ff",
   732 => x"06d40c53",
   733 => x"53b6a808",
   734 => x"85387189",
   735 => x"2b527198",
   736 => x"2ad40c71",
   737 => x"902a7081",
   738 => x"ff06d40c",
   739 => x"5171882a",
   740 => x"7081ff06",
   741 => x"d40c5171",
   742 => x"81ff06d4",
   743 => x"0c72902a",
   744 => x"7081ff06",
   745 => x"d40c51d4",
   746 => x"087081ff",
   747 => x"06515182",
   748 => x"b8bf5270",
   749 => x"81ff2e09",
   750 => x"81069438",
   751 => x"81ff0bd4",
   752 => x"0cd40870",
   753 => x"81ff06ff",
   754 => x"14545151",
   755 => x"71e53870",
   756 => x"b5c40c02",
   757 => x"8c050d04",
   758 => x"02fc050d",
   759 => x"81c75181",
   760 => x"ff0bd40c",
   761 => x"ff115170",
   762 => x"8025f438",
   763 => x"0284050d",
   764 => x"0402f405",
   765 => x"0d81ff0b",
   766 => x"d40c9353",
   767 => x"805287fc",
   768 => x"80c15196",
   769 => x"e72db5c4",
   770 => x"088b3881",
   771 => x"ff0bd40c",
   772 => x"8153989e",
   773 => x"0497d82d",
   774 => x"ff135372",
   775 => x"df3872b5",
   776 => x"c40c028c",
   777 => x"050d0402",
   778 => x"ec050d81",
   779 => x"0bb6a80c",
   780 => x"8454d008",
   781 => x"708f2a70",
   782 => x"81065151",
   783 => x"5372f338",
   784 => x"72d00c97",
   785 => x"d82db0f0",
   786 => x"5185fd2d",
   787 => x"d008708f",
   788 => x"2a708106",
   789 => x"51515372",
   790 => x"f338810b",
   791 => x"d00cb153",
   792 => x"805284d4",
   793 => x"80c05196",
   794 => x"e72db5c4",
   795 => x"08812e93",
   796 => x"3872822e",
   797 => x"bd38ff13",
   798 => x"5372e538",
   799 => x"ff145473",
   800 => x"ffb03897",
   801 => x"d82d83aa",
   802 => x"52849c80",
   803 => x"c85196e7",
   804 => x"2db5c408",
   805 => x"812e0981",
   806 => x"06923896",
   807 => x"992db5c4",
   808 => x"0883ffff",
   809 => x"06537283",
   810 => x"aa2e9d38",
   811 => x"97f12d99",
   812 => x"c304b0fc",
   813 => x"5185fd2d",
   814 => x"80539b91",
   815 => x"04b19451",
   816 => x"85fd2d80",
   817 => x"549ae304",
   818 => x"81ff0bd4",
   819 => x"0cb15497",
   820 => x"d82d8fcf",
   821 => x"53805287",
   822 => x"fc80f751",
   823 => x"96e72db5",
   824 => x"c40855b5",
   825 => x"c408812e",
   826 => x"0981069b",
   827 => x"3881ff0b",
   828 => x"d40c820a",
   829 => x"52849c80",
   830 => x"e95196e7",
   831 => x"2db5c408",
   832 => x"802e8d38",
   833 => x"97d82dff",
   834 => x"135372c9",
   835 => x"389ad604",
   836 => x"81ff0bd4",
   837 => x"0cb5c408",
   838 => x"5287fc80",
   839 => x"fa5196e7",
   840 => x"2db5c408",
   841 => x"b13881ff",
   842 => x"0bd40cd4",
   843 => x"085381ff",
   844 => x"0bd40c81",
   845 => x"ff0bd40c",
   846 => x"81ff0bd4",
   847 => x"0c81ff0b",
   848 => x"d40c7286",
   849 => x"2a708106",
   850 => x"76565153",
   851 => x"729538b5",
   852 => x"c408549a",
   853 => x"e3047382",
   854 => x"2efee238",
   855 => x"ff145473",
   856 => x"feed3873",
   857 => x"b6a80c73",
   858 => x"8b388152",
   859 => x"87fc80d0",
   860 => x"5196e72d",
   861 => x"81ff0bd4",
   862 => x"0cd00870",
   863 => x"8f2a7081",
   864 => x"06515153",
   865 => x"72f33872",
   866 => x"d00c81ff",
   867 => x"0bd40c81",
   868 => x"5372b5c4",
   869 => x"0c029405",
   870 => x"0d0402e8",
   871 => x"050d7855",
   872 => x"805681ff",
   873 => x"0bd40cd0",
   874 => x"08708f2a",
   875 => x"70810651",
   876 => x"515372f3",
   877 => x"3882810b",
   878 => x"d00c81ff",
   879 => x"0bd40c77",
   880 => x"5287fc80",
   881 => x"d15196e7",
   882 => x"2d80dbc6",
   883 => x"df54b5c4",
   884 => x"08802e8a",
   885 => x"38b1b451",
   886 => x"85fd2d9c",
   887 => x"b10481ff",
   888 => x"0bd40cd4",
   889 => x"087081ff",
   890 => x"06515372",
   891 => x"81fe2e09",
   892 => x"81069d38",
   893 => x"80ff5396",
   894 => x"992db5c4",
   895 => x"08757084",
   896 => x"05570cff",
   897 => x"13537280",
   898 => x"25ed3881",
   899 => x"569c9604",
   900 => x"ff145473",
   901 => x"c93881ff",
   902 => x"0bd40c81",
   903 => x"ff0bd40c",
   904 => x"d008708f",
   905 => x"2a708106",
   906 => x"51515372",
   907 => x"f33872d0",
   908 => x"0c75b5c4",
   909 => x"0c029805",
   910 => x"0d0402e8",
   911 => x"050d7779",
   912 => x"7b585555",
   913 => x"80537276",
   914 => x"25a33874",
   915 => x"70810556",
   916 => x"80f52d74",
   917 => x"70810556",
   918 => x"80f52d52",
   919 => x"5271712e",
   920 => x"86388151",
   921 => x"9cef0481",
   922 => x"13539cc6",
   923 => x"04805170",
   924 => x"b5c40c02",
   925 => x"98050d04",
   926 => x"02ec050d",
   927 => x"76557480",
   928 => x"2ebb389a",
   929 => x"1580e02d",
   930 => x"51a9f82d",
   931 => x"b5c408b5",
   932 => x"c408bcdc",
   933 => x"0cb5c408",
   934 => x"5454bcb8",
   935 => x"08802e99",
   936 => x"38941580",
   937 => x"e02d51a9",
   938 => x"f82db5c4",
   939 => x"08902b83",
   940 => x"fff00a06",
   941 => x"70750751",
   942 => x"5372bcdc",
   943 => x"0cbcdc08",
   944 => x"5372802e",
   945 => x"9938bcb0",
   946 => x"08fe1471",
   947 => x"29bcc408",
   948 => x"05bce00c",
   949 => x"70842bbc",
   950 => x"bc0c549e",
   951 => x"8404bcc8",
   952 => x"08bcdc0c",
   953 => x"bccc08bc",
   954 => x"e00cbcb8",
   955 => x"08802e8a",
   956 => x"38bcb008",
   957 => x"842b539e",
   958 => x"8004bcd0",
   959 => x"08842b53",
   960 => x"72bcbc0c",
   961 => x"0294050d",
   962 => x"0402d805",
   963 => x"0d800bbc",
   964 => x"b80c8454",
   965 => x"98a72db5",
   966 => x"c408802e",
   967 => x"9538b6ac",
   968 => x"5280519b",
   969 => x"9a2db5c4",
   970 => x"08802e86",
   971 => x"38fe549e",
   972 => x"ba04ff14",
   973 => x"54738024",
   974 => x"db38738c",
   975 => x"38b1c451",
   976 => x"85fd2d73",
   977 => x"55a3c304",
   978 => x"8056810b",
   979 => x"bce40c88",
   980 => x"53b1d852",
   981 => x"b6e2519c",
   982 => x"ba2db5c4",
   983 => x"08762e09",
   984 => x"81068738",
   985 => x"b5c408bc",
   986 => x"e40c8853",
   987 => x"b1e452b6",
   988 => x"fe519cba",
   989 => x"2db5c408",
   990 => x"8738b5c4",
   991 => x"08bce40c",
   992 => x"bce40880",
   993 => x"2e80f638",
   994 => x"b9f20b80",
   995 => x"f52db9f3",
   996 => x"0b80f52d",
   997 => x"71982b71",
   998 => x"902b07b9",
   999 => x"f40b80f5",
  1000 => x"2d70882b",
  1001 => x"7207b9f5",
  1002 => x"0b80f52d",
  1003 => x"7107baaa",
  1004 => x"0b80f52d",
  1005 => x"baab0b80",
  1006 => x"f52d7188",
  1007 => x"2b07535f",
  1008 => x"54525a56",
  1009 => x"57557381",
  1010 => x"abaa2e09",
  1011 => x"81068d38",
  1012 => x"7551a9c8",
  1013 => x"2db5c408",
  1014 => x"569fe904",
  1015 => x"7382d4d5",
  1016 => x"2e8738b1",
  1017 => x"f051a0aa",
  1018 => x"04b6ac52",
  1019 => x"75519b9a",
  1020 => x"2db5c408",
  1021 => x"55b5c408",
  1022 => x"802e83c7",
  1023 => x"388853b1",
  1024 => x"e452b6fe",
  1025 => x"519cba2d",
  1026 => x"b5c40889",
  1027 => x"38810bbc",
  1028 => x"b80ca0b0",
  1029 => x"048853b1",
  1030 => x"d852b6e2",
  1031 => x"519cba2d",
  1032 => x"b5c40880",
  1033 => x"2e8a38b2",
  1034 => x"845185fd",
  1035 => x"2da18a04",
  1036 => x"baaa0b80",
  1037 => x"f52d5473",
  1038 => x"80d52e09",
  1039 => x"810680ca",
  1040 => x"38baab0b",
  1041 => x"80f52d54",
  1042 => x"7381aa2e",
  1043 => x"098106ba",
  1044 => x"38800bb6",
  1045 => x"ac0b80f5",
  1046 => x"2d565474",
  1047 => x"81e92e83",
  1048 => x"38815474",
  1049 => x"81eb2e8c",
  1050 => x"38805573",
  1051 => x"752e0981",
  1052 => x"0682d038",
  1053 => x"b6b70b80",
  1054 => x"f52d5574",
  1055 => x"8d38b6b8",
  1056 => x"0b80f52d",
  1057 => x"5473822e",
  1058 => x"86388055",
  1059 => x"a3c304b6",
  1060 => x"b90b80f5",
  1061 => x"2d70bcb0",
  1062 => x"0cff05bc",
  1063 => x"b40cb6ba",
  1064 => x"0b80f52d",
  1065 => x"b6bb0b80",
  1066 => x"f52d5876",
  1067 => x"05778280",
  1068 => x"290570bc",
  1069 => x"c00cb6bc",
  1070 => x"0b80f52d",
  1071 => x"70bcd40c",
  1072 => x"bcb80859",
  1073 => x"57587680",
  1074 => x"2e81a338",
  1075 => x"8853b1e4",
  1076 => x"52b6fe51",
  1077 => x"9cba2db5",
  1078 => x"c40881e7",
  1079 => x"38bcb008",
  1080 => x"70842bbc",
  1081 => x"bc0c70bc",
  1082 => x"d00cb6d1",
  1083 => x"0b80f52d",
  1084 => x"b6d00b80",
  1085 => x"f52d7182",
  1086 => x"802905b6",
  1087 => x"d20b80f5",
  1088 => x"2d708480",
  1089 => x"802912b6",
  1090 => x"d30b80f5",
  1091 => x"2d708180",
  1092 => x"0a291270",
  1093 => x"bcd80cbc",
  1094 => x"d4087129",
  1095 => x"bcc00805",
  1096 => x"70bcc40c",
  1097 => x"b6d90b80",
  1098 => x"f52db6d8",
  1099 => x"0b80f52d",
  1100 => x"71828029",
  1101 => x"05b6da0b",
  1102 => x"80f52d70",
  1103 => x"84808029",
  1104 => x"12b6db0b",
  1105 => x"80f52d70",
  1106 => x"982b81f0",
  1107 => x"0a067205",
  1108 => x"70bcc80c",
  1109 => x"fe117e29",
  1110 => x"7705bccc",
  1111 => x"0c525952",
  1112 => x"43545e51",
  1113 => x"5259525d",
  1114 => x"575957a3",
  1115 => x"bc04b6be",
  1116 => x"0b80f52d",
  1117 => x"b6bd0b80",
  1118 => x"f52d7182",
  1119 => x"80290570",
  1120 => x"bcbc0c70",
  1121 => x"a02983ff",
  1122 => x"0570892a",
  1123 => x"70bcd00c",
  1124 => x"b6c30b80",
  1125 => x"f52db6c2",
  1126 => x"0b80f52d",
  1127 => x"71828029",
  1128 => x"0570bcd8",
  1129 => x"0c7b7129",
  1130 => x"1e70bccc",
  1131 => x"0c7dbcc8",
  1132 => x"0c7305bc",
  1133 => x"c40c555e",
  1134 => x"51515555",
  1135 => x"80519cf8",
  1136 => x"2d815574",
  1137 => x"b5c40c02",
  1138 => x"a8050d04",
  1139 => x"02ec050d",
  1140 => x"7670872c",
  1141 => x"7180ff06",
  1142 => x"555654bc",
  1143 => x"b8088a38",
  1144 => x"73882c74",
  1145 => x"81ff0654",
  1146 => x"55b6ac52",
  1147 => x"bcc00815",
  1148 => x"519b9a2d",
  1149 => x"b5c40854",
  1150 => x"b5c40880",
  1151 => x"2eb338bc",
  1152 => x"b808802e",
  1153 => x"98387284",
  1154 => x"29b6ac05",
  1155 => x"70085253",
  1156 => x"a9c82db5",
  1157 => x"c408f00a",
  1158 => x"0653a4af",
  1159 => x"047210b6",
  1160 => x"ac057080",
  1161 => x"e02d5253",
  1162 => x"a9f82db5",
  1163 => x"c4085372",
  1164 => x"5473b5c4",
  1165 => x"0c029405",
  1166 => x"0d0402e0",
  1167 => x"050d7970",
  1168 => x"842cbce0",
  1169 => x"0805718f",
  1170 => x"06525553",
  1171 => x"728938b6",
  1172 => x"ac527351",
  1173 => x"9b9a2d72",
  1174 => x"a029b6ac",
  1175 => x"05548074",
  1176 => x"80f52d56",
  1177 => x"5374732e",
  1178 => x"83388153",
  1179 => x"7481e52e",
  1180 => x"81ef3881",
  1181 => x"70740654",
  1182 => x"5872802e",
  1183 => x"81e3388b",
  1184 => x"1480f52d",
  1185 => x"70832a79",
  1186 => x"06585676",
  1187 => x"9838b488",
  1188 => x"08537288",
  1189 => x"3872baac",
  1190 => x"0b81b72d",
  1191 => x"76b4880c",
  1192 => x"7353a6e3",
  1193 => x"04758f2e",
  1194 => x"09810681",
  1195 => x"b438749f",
  1196 => x"068d29ba",
  1197 => x"9f115153",
  1198 => x"811480f5",
  1199 => x"2d737081",
  1200 => x"055581b7",
  1201 => x"2d831480",
  1202 => x"f52d7370",
  1203 => x"81055581",
  1204 => x"b72d8514",
  1205 => x"80f52d73",
  1206 => x"70810555",
  1207 => x"81b72d87",
  1208 => x"1480f52d",
  1209 => x"73708105",
  1210 => x"5581b72d",
  1211 => x"891480f5",
  1212 => x"2d737081",
  1213 => x"055581b7",
  1214 => x"2d8e1480",
  1215 => x"f52d7370",
  1216 => x"81055581",
  1217 => x"b72d9014",
  1218 => x"80f52d73",
  1219 => x"70810555",
  1220 => x"81b72d92",
  1221 => x"1480f52d",
  1222 => x"73708105",
  1223 => x"5581b72d",
  1224 => x"941480f5",
  1225 => x"2d737081",
  1226 => x"055581b7",
  1227 => x"2d961480",
  1228 => x"f52d7370",
  1229 => x"81055581",
  1230 => x"b72d9814",
  1231 => x"80f52d73",
  1232 => x"70810555",
  1233 => x"81b72d9c",
  1234 => x"1480f52d",
  1235 => x"73708105",
  1236 => x"5581b72d",
  1237 => x"9e1480f5",
  1238 => x"2d7381b7",
  1239 => x"2d77b488",
  1240 => x"0c805372",
  1241 => x"b5c40c02",
  1242 => x"a0050d04",
  1243 => x"02cc050d",
  1244 => x"7e605e5a",
  1245 => x"800bbcdc",
  1246 => x"08bce008",
  1247 => x"595c5680",
  1248 => x"58bcbc08",
  1249 => x"782e81ae",
  1250 => x"38778f06",
  1251 => x"a0175754",
  1252 => x"738f38b6",
  1253 => x"ac527651",
  1254 => x"8117579b",
  1255 => x"9a2db6ac",
  1256 => x"56807680",
  1257 => x"f52d5654",
  1258 => x"74742e83",
  1259 => x"38815474",
  1260 => x"81e52e80",
  1261 => x"f6388170",
  1262 => x"7506555c",
  1263 => x"73802e80",
  1264 => x"ea388b16",
  1265 => x"80f52d98",
  1266 => x"06597880",
  1267 => x"de388b53",
  1268 => x"7c527551",
  1269 => x"9cba2db5",
  1270 => x"c40880cf",
  1271 => x"389c1608",
  1272 => x"51a9c82d",
  1273 => x"b5c40884",
  1274 => x"1b0c9a16",
  1275 => x"80e02d51",
  1276 => x"a9f82db5",
  1277 => x"c408b5c4",
  1278 => x"08881c0c",
  1279 => x"b5c40855",
  1280 => x"55bcb808",
  1281 => x"802e9838",
  1282 => x"941680e0",
  1283 => x"2d51a9f8",
  1284 => x"2db5c408",
  1285 => x"902b83ff",
  1286 => x"f00a0670",
  1287 => x"16515473",
  1288 => x"881b0c78",
  1289 => x"7a0c7b54",
  1290 => x"a8ec0481",
  1291 => x"1858bcbc",
  1292 => x"087826fe",
  1293 => x"d438bcb8",
  1294 => x"08802eae",
  1295 => x"387a51a3",
  1296 => x"cc2db5c4",
  1297 => x"08b5c408",
  1298 => x"80ffffff",
  1299 => x"f806555b",
  1300 => x"7380ffff",
  1301 => x"fff82e92",
  1302 => x"38b5c408",
  1303 => x"fe05bcb0",
  1304 => x"0829bcc4",
  1305 => x"080557a6",
  1306 => x"ff048054",
  1307 => x"73b5c40c",
  1308 => x"02b4050d",
  1309 => x"0402f405",
  1310 => x"0d747008",
  1311 => x"8105710c",
  1312 => x"7008bcb4",
  1313 => x"08065353",
  1314 => x"718e3888",
  1315 => x"130851a3",
  1316 => x"cc2db5c4",
  1317 => x"0888140c",
  1318 => x"810bb5c4",
  1319 => x"0c028c05",
  1320 => x"0d0402f0",
  1321 => x"050d7588",
  1322 => x"1108fe05",
  1323 => x"bcb00829",
  1324 => x"bcc40811",
  1325 => x"7208bcb4",
  1326 => x"08060579",
  1327 => x"55535454",
  1328 => x"9b9a2d02",
  1329 => x"90050d04",
  1330 => x"02f4050d",
  1331 => x"7470882a",
  1332 => x"83fe8006",
  1333 => x"7072982a",
  1334 => x"0772882b",
  1335 => x"87fc8080",
  1336 => x"0673982b",
  1337 => x"81f00a06",
  1338 => x"71730707",
  1339 => x"b5c40c56",
  1340 => x"51535102",
  1341 => x"8c050d04",
  1342 => x"02f8050d",
  1343 => x"028e0580",
  1344 => x"f52d7488",
  1345 => x"2b077083",
  1346 => x"ffff06b5",
  1347 => x"c40c5102",
  1348 => x"88050d04",
  1349 => x"02f4050d",
  1350 => x"74767853",
  1351 => x"54528071",
  1352 => x"25973872",
  1353 => x"70810554",
  1354 => x"80f52d72",
  1355 => x"70810554",
  1356 => x"81b72dff",
  1357 => x"115170eb",
  1358 => x"38807281",
  1359 => x"b72d028c",
  1360 => x"050d0402",
  1361 => x"e8050d77",
  1362 => x"56807056",
  1363 => x"54737624",
  1364 => x"b138bcbc",
  1365 => x"08742eaa",
  1366 => x"387351a4",
  1367 => x"ba2db5c4",
  1368 => x"08b5c408",
  1369 => x"09810570",
  1370 => x"b5c40807",
  1371 => x"9f2a7705",
  1372 => x"81175757",
  1373 => x"53537476",
  1374 => x"248838bc",
  1375 => x"bc087426",
  1376 => x"d83872b5",
  1377 => x"c40c0298",
  1378 => x"050d0402",
  1379 => x"f0050db5",
  1380 => x"c0081651",
  1381 => x"aac32db5",
  1382 => x"c408802e",
  1383 => x"9b388b53",
  1384 => x"b5c40852",
  1385 => x"baac51aa",
  1386 => x"942dbce8",
  1387 => x"08547380",
  1388 => x"2e8638ba",
  1389 => x"ac51732d",
  1390 => x"0290050d",
  1391 => x"0402dc05",
  1392 => x"0d80705a",
  1393 => x"5574b5c0",
  1394 => x"0825af38",
  1395 => x"bcbc0875",
  1396 => x"2ea83878",
  1397 => x"51a4ba2d",
  1398 => x"b5c40809",
  1399 => x"810570b5",
  1400 => x"c408079f",
  1401 => x"2a760581",
  1402 => x"1b5b5654",
  1403 => x"74b5c008",
  1404 => x"258838bc",
  1405 => x"bc087926",
  1406 => x"da388055",
  1407 => x"78bcbc08",
  1408 => x"2781cd38",
  1409 => x"7851a4ba",
  1410 => x"2db5c408",
  1411 => x"802e81a2",
  1412 => x"38b5c408",
  1413 => x"8b0580f5",
  1414 => x"2d70842a",
  1415 => x"70810677",
  1416 => x"1078842b",
  1417 => x"baac0b80",
  1418 => x"f52d5c5c",
  1419 => x"53515556",
  1420 => x"73802e80",
  1421 => x"c6387416",
  1422 => x"822badf3",
  1423 => x"0bb49412",
  1424 => x"0c547775",
  1425 => x"3110bcec",
  1426 => x"11555690",
  1427 => x"74708105",
  1428 => x"5681b72d",
  1429 => x"a07481b7",
  1430 => x"2d7681ff",
  1431 => x"06811658",
  1432 => x"5473802e",
  1433 => x"89389c53",
  1434 => x"baac52ac",
  1435 => x"f4048b53",
  1436 => x"b5c40852",
  1437 => x"bcee1651",
  1438 => x"adaa0474",
  1439 => x"16822bab",
  1440 => x"8b0bb494",
  1441 => x"120c5476",
  1442 => x"81ff0681",
  1443 => x"16585473",
  1444 => x"802e8938",
  1445 => x"9c53baac",
  1446 => x"52ada204",
  1447 => x"8b53b5c4",
  1448 => x"08527775",
  1449 => x"3110bcec",
  1450 => x"05517655",
  1451 => x"aa942dad",
  1452 => x"c5047490",
  1453 => x"29753170",
  1454 => x"10bcec05",
  1455 => x"5154b5c4",
  1456 => x"087481b7",
  1457 => x"2d811959",
  1458 => x"748b24a2",
  1459 => x"38abfc04",
  1460 => x"74902975",
  1461 => x"317010bc",
  1462 => x"ec058c77",
  1463 => x"31575154",
  1464 => x"807481b7",
  1465 => x"2d9e14ff",
  1466 => x"16565474",
  1467 => x"f33802a4",
  1468 => x"050d0402",
  1469 => x"fc050db5",
  1470 => x"c0081351",
  1471 => x"aac32db5",
  1472 => x"c408802e",
  1473 => x"8838b5c4",
  1474 => x"08519cf8",
  1475 => x"2d800bb5",
  1476 => x"c00cabbd",
  1477 => x"2d8eaf2d",
  1478 => x"0284050d",
  1479 => x"0402fc05",
  1480 => x"0d725170",
  1481 => x"fd2ead38",
  1482 => x"70fd248a",
  1483 => x"3870fc2e",
  1484 => x"80c438ae",
  1485 => x"fe0470fe",
  1486 => x"2eb13870",
  1487 => x"ff2e0981",
  1488 => x"06bc38b5",
  1489 => x"c0085170",
  1490 => x"802eb338",
  1491 => x"ff11b5c0",
  1492 => x"0caefe04",
  1493 => x"b5c008f0",
  1494 => x"0570b5c0",
  1495 => x"0c517080",
  1496 => x"259c3880",
  1497 => x"0bb5c00c",
  1498 => x"aefe04b5",
  1499 => x"c0088105",
  1500 => x"b5c00cae",
  1501 => x"fe04b5c0",
  1502 => x"089005b5",
  1503 => x"c00cabbd",
  1504 => x"2d8eaf2d",
  1505 => x"0284050d",
  1506 => x"0402fc05",
  1507 => x"0d800bb5",
  1508 => x"c00cabbd",
  1509 => x"2d8dc62d",
  1510 => x"b5c408b5",
  1511 => x"b00cb48c",
  1512 => x"518fca2d",
  1513 => x"0284050d",
  1514 => x"0471bce8",
  1515 => x"0c040000",
  1516 => x"00ffffff",
  1517 => x"ff00ffff",
  1518 => x"ffff00ff",
  1519 => x"ffffff00",
  1520 => x"20202020",
  1521 => x"3d5a5844",
  1522 => x"4f533d20",
  1523 => x"20202000",
  1524 => x"20202020",
  1525 => x"20202020",
  1526 => x"20202020",
  1527 => x"20202000",
  1528 => x"52657365",
  1529 => x"74000000",
  1530 => x"5363616e",
  1531 => x"6c696e65",
  1532 => x"73000000",
  1533 => x"53696420",
  1534 => x"38353830",
  1535 => x"00000000",
  1536 => x"436f6c6f",
  1537 => x"72204365",
  1538 => x"50436572",
  1539 => x"6f000000",
  1540 => x"4e747363",
  1541 => x"00000000",
  1542 => x"43617267",
  1543 => x"61722044",
  1544 => x"6973636f",
  1545 => x"20100000",
  1546 => x"45786974",
  1547 => x"00000000",
  1548 => x"43617267",
  1549 => x"61206465",
  1550 => x"2044534b",
  1551 => x"2046616c",
  1552 => x"6c696461",
  1553 => x"00000000",
  1554 => x"4f4b0000",
  1555 => x"496e6974",
  1556 => x"69616c69",
  1557 => x"7a696e67",
  1558 => x"20534420",
  1559 => x"63617264",
  1560 => x"0a000000",
  1561 => x"16200000",
  1562 => x"14200000",
  1563 => x"15200000",
  1564 => x"53442069",
  1565 => x"6e69742e",
  1566 => x"2e2e0a00",
  1567 => x"53442063",
  1568 => x"61726420",
  1569 => x"72657365",
  1570 => x"74206661",
  1571 => x"696c6564",
  1572 => x"210a0000",
  1573 => x"53444843",
  1574 => x"20657272",
  1575 => x"6f72210a",
  1576 => x"00000000",
  1577 => x"57726974",
  1578 => x"65206661",
  1579 => x"696c6564",
  1580 => x"0a000000",
  1581 => x"52656164",
  1582 => x"20666169",
  1583 => x"6c65640a",
  1584 => x"00000000",
  1585 => x"43617264",
  1586 => x"20696e69",
  1587 => x"74206661",
  1588 => x"696c6564",
  1589 => x"0a000000",
  1590 => x"46415431",
  1591 => x"36202020",
  1592 => x"00000000",
  1593 => x"46415433",
  1594 => x"32202020",
  1595 => x"00000000",
  1596 => x"4e6f2070",
  1597 => x"61727469",
  1598 => x"74696f6e",
  1599 => x"20736967",
  1600 => x"0a000000",
  1601 => x"42616420",
  1602 => x"70617274",
  1603 => x"0a000000",
  1604 => x"4261636b",
  1605 => x"00000000",
  1606 => x"00000002",
  1607 => x"00000002",
  1608 => x"000017c0",
  1609 => x"00000000",
  1610 => x"00000002",
  1611 => x"000017d0",
  1612 => x"00000000",
  1613 => x"00000002",
  1614 => x"000017e0",
  1615 => x"0000034d",
  1616 => x"00000001",
  1617 => x"000017e8",
  1618 => x"00000000",
  1619 => x"00000001",
  1620 => x"000017f4",
  1621 => x"00000001",
  1622 => x"00000001",
  1623 => x"00001800",
  1624 => x"00000002",
  1625 => x"00000001",
  1626 => x"00001810",
  1627 => x"00000003",
  1628 => x"00000002",
  1629 => x"00001818",
  1630 => x"00001789",
  1631 => x"00000002",
  1632 => x"00001828",
  1633 => x"000006cd",
  1634 => x"00000000",
  1635 => x"00000000",
  1636 => x"00000000",
  1637 => x"00000004",
  1638 => x"00001830",
  1639 => x"00001994",
  1640 => x"00000004",
  1641 => x"00001848",
  1642 => x"0000191c",
  1643 => x"00000000",
  1644 => x"00000000",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"00000000",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000002",
  1668 => x"00001e6c",
  1669 => x"0000158b",
  1670 => x"00000002",
  1671 => x"00001e8a",
  1672 => x"0000158b",
  1673 => x"00000002",
  1674 => x"00001ea8",
  1675 => x"0000158b",
  1676 => x"00000002",
  1677 => x"00001ec6",
  1678 => x"0000158b",
  1679 => x"00000002",
  1680 => x"00001ee4",
  1681 => x"0000158b",
  1682 => x"00000002",
  1683 => x"00001f02",
  1684 => x"0000158b",
  1685 => x"00000002",
  1686 => x"00001f20",
  1687 => x"0000158b",
  1688 => x"00000002",
  1689 => x"00001f3e",
  1690 => x"0000158b",
  1691 => x"00000002",
  1692 => x"00001f5c",
  1693 => x"0000158b",
  1694 => x"00000002",
  1695 => x"00001f7a",
  1696 => x"0000158b",
  1697 => x"00000002",
  1698 => x"00001f98",
  1699 => x"0000158b",
  1700 => x"00000002",
  1701 => x"00001fb6",
  1702 => x"0000158b",
  1703 => x"00000002",
  1704 => x"00001fd4",
  1705 => x"0000158b",
  1706 => x"00000004",
  1707 => x"00001910",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"0000171d",
  1712 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

