-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "05110414441051105504415414B26841541692F9A105505A1055044D1415695A";
    attribute INIT_01 of inst : label is "68820BC9AAA489A52658B6E10414441051104144410511041444105110414441";
    attribute INIT_02 of inst : label is "EAE2341459A76966C5D4E84EB4EA4EB4E64E54E44E57258E3ADBADB6FB2B86AA";
    attribute INIT_03 of inst : label is "6A8FABA9D224D459A75DA59B97559628A6A8FA778505146966D5D5624AA29AA3";
    attribute INIT_04 of inst : label is "49BD06926841B8524B665962492A8A6E8FAB9A0E08F59166A96E155A59BD758A";
    attribute INIT_05 of inst : label is "37DA7D87D37DB41056CB2C91414524D051499A55DA59B175BF274B6FC9D4B558";
    attribute INIT_06 of inst : label is "6D5D71E24159A7925A246B91AB46A51A446911AC46811A8768A668FA4AAE58BD";
    attribute INIT_07 of inst : label is "EC525146966F5DACAAFABBA0E28F59146966E5D72EB8A298A3E9D61493514696";
    attribute INIT_08 of inst : label is "A3EAEA149341451A59B976FE46966D5DDFA0E08F59146966C5D629AA3E9DACAA";
    attribute INIT_09 of inst : label is "1A59B57776D8F6A3D6451A59B1758A628FABA8D05155905251A59BD743D66298";
    attribute INIT_0A of inst : label is "9D56455E554E00002801545146966F5D72A45146966E5D6298A3EAEA14934145";
    attribute INIT_0B of inst : label is "59D56455E654E3939393A4E4E42B90B9393E4E4E4D59954E559954E55A956A55";
    attribute INIT_0C of inst : label is "FFCEA9F95F557D55F557D55A556955FD57F55FD57F559954E559954E55A956A5";
    attribute INIT_0D of inst : label is "F1E87EF155F557D55F557D55A556955FD57F55FE97FEA73FFCFFFFFFDFFF7FFF";
    attribute INIT_0E of inst : label is "190006403190086401FFD5D5D5D5BC6AAAEA2AD5D5D5D5FF6AAAEA2A6BF11F1E";
    attribute INIT_0F of inst : label is "AAAAAAAAAA190186405190106407190186405190106401190006403190086401";
    attribute INIT_10 of inst : label is "02002E00000F85FB308DE04405E6CDB409FB609990F3C2FF9F50707FFFF00002";
    attribute INIT_11 of inst : label is "62C49A58B125A58B1E6962C796962C41A58B105A58B1C6962C71930000000000";
    attribute INIT_12 of inst : label is "A598D75A598156966355A7981755595A859AA5989759AA5985759AA59B175E69";
    attribute INIT_13 of inst : label is "A906133802C67DFB06A04909A5968069A0069A4BA11692E4456966351A598165";
    attribute INIT_14 of inst : label is "76741595EB651CB8EDCBEE3E60AACFC6741DCD9D05CF0F12BE565953BA3AA712";
    attribute INIT_15 of inst : label is "161E2D4DA78A5361EAC4DA7AAD35B8B2FB95657ACAE69AD5B9CBEE69A2EA9AC5";
    attribute INIT_16 of inst : label is "97EC107089742009074C5C0544D16251AFC1300175DB4400000061E2E45A78B1";
    attribute INIT_17 of inst : label is "293C826939A06938F00E35CE4E6C4008040C00000000000C0408000400040A65";
    attribute INIT_18 of inst : label is "10448D88E74D30624A38F14008A24108C10929F34F34F04B2CB20B2361642A93";
    attribute INIT_19 of inst : label is "0613CE6884AF3581DBCD6E0627ADB80EF35A47B1FD2DEA018EB45D1044D11449";
    attribute INIT_1A of inst : label is "7C98817C988D7C9881B7C988D167C98817C9881A2F6D4B81E8AEF7F2F3B0D6A2";
    attribute INIT_1B of inst : label is "7C98857C98859F26225F26215F26235F26216DF2623459F26215F262167C9881";
    attribute INIT_1C of inst : label is "6205F26206DF2620459F26205F262067C98897C98897C98897C9885B7C988916";
    attribute INIT_1D of inst : label is "23547C988D7C98897C988D7C9881B7C988D167C98817C98819F26205F26215F2";
    attribute INIT_1E of inst : label is "C9889FC9885FC9885FC9885FC9885FC9881FC9881FC9881FC988187C9350E47A";
    attribute INIT_1F of inst : label is "88DFC988DFC9885FC9885FC988DFC988DFC9885FC9885FC9885FC9885FC9889F";
    attribute INIT_20 of inst : label is "D0515495AC891BC9885FC9881FC988DFC989DFC988DFC9881FC988DFC988DFC9";
    attribute INIT_21 of inst : label is "ECB5313D2A69B1769A6B5DA489D36922745A48ADF6922B7564A9A6C51A69A544";
    attribute INIT_22 of inst : label is "B6D46D551B6D46D55174D46D951B5D45D151B7D46D751B75EEB20ACBE82FBA00";
    attribute INIT_23 of inst : label is "EA2E94565669C943EEB36060A0E020FA33B2B2B1091FCBCE8A89D54A3146D951";
    attribute INIT_24 of inst : label is "809D8C510731B8DE86ACB88ABAAAAA8AFB2AAA8EE43AAAACAAF2AAACA2CAAAB8";
    attribute INIT_25 of inst : label is "E136B53E70437CE20F4E80121182751000031401288450005214C2161F44C036";
    attribute INIT_26 of inst : label is "569252A0AE7A4E4A4669D2964B9C4ACEA8383AA5923425996499CE001265BC04";
    attribute INIT_27 of inst : label is "19189E5A46421A23A01A68849DD28DD3B6B060EE7F094DFE25F7018986866E61";
    attribute INIT_28 of inst : label is "1199E7A4646191B9E6A464E19199E5A46461A382291A9E6A464A191A9E4A464A";
    attribute INIT_29 of inst : label is "9E0BE9684B5B829E0AE780BFFF5B9E4BE9674B5B829E4A279292A49516B655E7";
    attribute INIT_2A of inst : label is "441E796F552569087F4505087F450638002F6B2D95BF291209922FFFE9684B5B";
    attribute INIT_2B of inst : label is "D6FFFFCA790F434022D1069AFC2ED176BDA7D67B6BDA487D07B493DA5D05008B";
    attribute INIT_2C of inst : label is "426115091C242636D5E7F2D59FC943516F5908C5BD6C215BD6C5F805BD6FAE23";
    attribute INIT_2D of inst : label is "609271B7B04927F3B5EE77E57B2249C9967E6DEFE492662CEE619654450271C2";
    attribute INIT_2E of inst : label is "E27709DE2610659C927789DC277898419672499EDD8EDDC09782719640256682";
    attribute INIT_2F of inst : label is "B186ACB5B185AF628C54D565EE27709DE2610659C927789DC27789841967249D";
    attribute INIT_30 of inst : label is "236146A59157423688D951A96455D08DA236956BE0FB095820BE095B95B5ACB5";
    attribute INIT_31 of inst : label is "614AA59257423688D952A96495D08DA23694AA59257423688DB51A96455D08DA";
    attribute INIT_32 of inst : label is "F7FFFED25DFFFF3794EA5935748DA23694EA59357423688DB53A964D5D08DA23";
    attribute INIT_33 of inst : label is "953DD1994CD09EFD3994F765337BF6536666AA2D5195DDEF9D157EA59BA35359";
    attribute INIT_34 of inst : label is "8555445B6DD8412D5554FB94FD117F4FBB1264994D4452FED59253CE5855F1CB";
    attribute INIT_35 of inst : label is "E44D1C39383C056FB470E40566D83D8A505E4405610CFE405624FB653FAEE509";
    attribute INIT_36 of inst : label is "4930981061826490E74B71F0CD1C3019D8FE47180440E3662754E60560F10158";
    attribute INIT_37 of inst : label is "E11E17BC7F401001901402E719900003634F6040513D820178F6C4051B271EF1";
    attribute INIT_38 of inst : label is "0000FC40000000FC00038000FCC0030000FC80038000FC40030000FCB40F4783";
    attribute INIT_39 of inst : label is "210916940F4783E11E2480008000FC4000C000FC00004000FCC0008000FC8000";
    attribute INIT_3A of inst : label is "B98BA98BA98846C6C6C6C6C6C693939393939394E4E471F08765DF6623E02BAE";
    attribute INIT_3B of inst : label is "6D8AF1B606D9962DAE6AAA2A89E789A27AEF4EEC62F50BF97B4E8EA2ED4E6001";
    attribute INIT_3C of inst : label is "9AAE790925EE77D999191E909962C605846C2A42658B1A105AB09FABAB6BC61B";
    attribute INIT_3D of inst : label is "BD90939AE6424E6B5909391230DEFCDEFCDEFCDEFCDAB856599BADA190952509";
    attribute INIT_3E of inst : label is "24E6BD90939AE6424E6B590939AC6424E6BD90939AE6424E6B590939AC6424E6";
    attribute INIT_3F of inst : label is "9C6464E47D909391E6424E475909391C6424E47D909391E6424E47590939AF64";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C18303060C0C183230B0C8E2CE3AF0C4C24FB0DB43138936313090C4E2C5CD7B";
    attribute INIT_01 of inst : label is "8E30C3E1FC7C1FCF0BF0F8F303060C0C18303060C0C18303060C0C18303060C0";
    attribute INIT_02 of inst : label is "EB8F8EBBE75AD793708B8D38E38C38F38C38E38C38C34CBCF8E34D30E30F38E3";
    attribute INIT_03 of inst : label is "CF07AE2E75BE3BE758EB5E4DC22C383F3CB07A9C6BAEF9D793508B83D2FCF2C1";
    attribute INIT_04 of inst : label is "F4D8417D34006D38C34BC383D3CBF3CF07AE0CA9BE9CAF9D57D39005E4D422F3";
    attribute INIT_05 of inst : label is "00F00F30F20F00008134125C002BBE3AEF56758E35E4D022605F2E18174AE707";
    attribute INIT_06 of inst : label is "3608A2D5900618696D02F40BD02F4CBD12F4CBD22F48BD138F3CB07AD2F4E0CF";
    attribute INIT_07 of inst : label is "8EBBEF9D79360801C07AE0CA9BE9CAF9D793408B83E3FCF2C1EA75AEF8EF9D79";
    attribute INIT_08 of inst : label is "C1EB8BAEF8EBBE75E4D420859D79370810EAB8E9CAF9D793508BCF0C1EA75E0F";
    attribute INIT_09 of inst : label is "75E4D020471A863A72BE75E4D822F3CB07AE2E3AEF5EDABBE75E4DC229B2BCF2";
    attribute INIT_0A of inst : label is "A154055FD57A00002C00A5EF9D793408B835EF9D793608BCF1C1EB8BAEF8EBBE";
    attribute INIT_0B of inst : label is "5A154055FC17A3FEA95440FFAA6555803FEFFAA55150954E55F957A55A956A55";
    attribute INIT_0C of inst : label is "FFF3FF0D5095425509542555155455015405501540550954E55F957A55A956A5";
    attribute INIT_0D of inst : label is "0802000655095425509542555155455015405503D40FFC3FFCFFFFFF6FFDBFFF";
    attribute INIT_0E of inst : label is "D5C075700D5C035700FFEAEAEAEAABAA2A2AAAEAEAEAEAFF2A2A2A6A55088060";
    attribute INIT_0F of inst : label is "0000000000D5C075701D5C075700D5C035700D5C035702D5C0B5701D5C075701";
    attribute INIT_10 of inst : label is "02000188004325C7B401001995C80079107C34610F0BD0C81050736AAAAAAAA8";
    attribute INIT_11 of inst : label is "5741C5D5DC325D5D87175750C97574145D5DC125D5D851757504830000800000";
    attribute INIT_12 of inst : label is "5F4E0325F4E8217D3A045E4E0025ED7B41FB5E4E861FB5E4E061FB5E4DC61197";
    attribute INIT_13 of inst : label is "E5E3DA8FC3AFCCC303C00DA43A2F22FB492DA5F5DC617D760897D3A085F4E812";
    attribute INIT_14 of inst : label is "A0D9069ED1279D16DBDB01F290FEE220E809E83A01A86718F207CD6170F28E8B";
    attribute INIT_15 of inst : label is "01F979185E5C821F939145E4C012D0F8D1D775F8C3CF34ED3EE347F347E0FCB2";
    attribute INIT_16 of inst : label is "E410D502417400419760D30534642086CC11400D90EC763400009F979105E5E8";
    attribute INIT_17 of inst : label is "D10D00401C13810311F00BFA900140000404000000000004040000040004226C";
    attribute INIT_18 of inst : label is "5116003EBE4A30F30A28E38F34F38C38C3CD2082083493CE38E3092A12021203";
    attribute INIT_19 of inst : label is "01E9C0578217014011C05C00FAFA5D017015031ED101C4C0EB29485114451140";
    attribute INIT_1A of inst : label is "5D16085D16005D160815D1600D05D16085D16084FEB44840C7FB2A747050055C";
    attribute INIT_1B of inst : label is "5D160C5D160C57458117458217458317458205745833417458217458215D1604";
    attribute INIT_1C of inst : label is "58117458005745813417458017458015D160C5D16045D160C5D160C15D160CD0";
    attribute INIT_1D of inst : label is "F6B25D16085D160C5D16085D160415D1608D05D16045D1604574581174582174";
    attribute INIT_1E of inst : label is "D16041D16041D16041D16041D16041D16001D16001D16081D16083B21D121030";
    attribute INIT_1F of inst : label is "6041D16041D16041D16041D16041D16041D16001D16001D16041D16041D16041";
    attribute INIT_20 of inst : label is "3AEF5ED7BF2ED5D16001D16001D16041D16081D16041D16001D16041D16041D1";
    attribute INIT_21 of inst : label is "B3BC703B25F4DC517D31045D5C4317571085D5C4317571087FD7D37145F4C412";
    attribute INIT_22 of inst : label is "10C3C420710C1C420F10C1C420710C3C420710C1C430F108924DA93492D2496E";
    attribute INIT_23 of inst : label is "AAEAA1C7D3975C200F8BEAFEF2B6FAFA9ACBEBCABCA6CB4FEBC5C18C7C1C4207";
    attribute INIT_24 of inst : label is "C011D22914842BBABEBBABBAAAAAAABAAAEAAABAAFEBAAABAAAEAAABAEBAAAAB";
    attribute INIT_25 of inst : label is "C23E44E005C070090F1CE451260855203031A5E23416504B4315C2E510044847";
    attribute INIT_26 of inst : label is "1E41C2FCBDC9B1C1E1E64073FCF1C723FB0D2F1CF96F4D144911035420BADC47";
    attribute INIT_27 of inst : label is "DAD1E1C1C1E7D80AF8AFFB474228F20A6FAE327DC8078C201EF2A8CFCF23A1C7";
    attribute INIT_28 of inst : label is "ED0E1C1C1E3DAD0E1C1C1E3DAD1E1C1C1E7DB0DB8ED0E1C1C1E3DAD1E1C1C1E7";
    attribute INIT_29 of inst : label is "F4D46F86CDEADAF4D6BD88E446EAF4D46F84CDEADAF4D63DA9334CC9336C1F03";
    attribute INIT_2A of inst : label is "C2BAE38D9735CE00D3104200D30002A3B806D89B0D8C793501FB5111AF86CDEA";
    attribute INIT_2B of inst : label is "B27BBB874E4C934803B0AEB8DABBB09C1B2B78E3C1B2F2B62E9FB9B28A01200E";
    attribute INIT_2C of inst : label is "78B1B20E3FA7892EB88F71983DC5930B06CB8EEC1B2A3AC1B20CA22C1B277889";
    attribute INIT_2D of inst : label is "E9F7F2B3DA977D951A934D9CF9C7DF51F7DCACF5E977D4A4F56977EC6C83A3FA";
    attribute INIT_2E of inst : label is "21DCC7731FAA5DF577DC47711DC07EA977D5DF73BC51BC6078C1D9F7DA1E38E1";
    attribute INIT_2F of inst : label is "29AD92CF29AD9163EFCF07EBCE1DCC7731FAA5DF577DC47711DC07EA977D5DF7";
    attribute INIT_30 of inst : label is "52F8C47EF039C92DD4BF311FBC0E724B752F0ED18AB50AD0109D0AD3EF0D32CF";
    attribute INIT_31 of inst : label is "F4C87EF139C92DD4BE321FBC4E724B752FCC87EF139C92DD4BC311FBC0E724B7";
    attribute INIT_32 of inst : label is "1FBBB877C7EEEE1CF8C7EF239E4B752F8CC7EF239C92DD4BF331FBC8E724B752";
    attribute INIT_33 of inst : label is "F241717C9179730707C905F245CC1F24226AA226E2A22E6391B91B1CFA32E5DF";
    attribute INIT_34 of inst : label is "1C729E71E078C8101DC924C92279C0924C6B9EF8909E7188927BE405E1C7978D";
    attribute INIT_35 of inst : label is "F441D13D305C32430744F4324B110EC453205932401C0C43240905F248593207";
    attribute INIT_36 of inst : label is "DD702DD540D18415F44B8621C1D1705ED00C482C663CD1A04934D43241710C90";
    attribute INIT_37 of inst : label is "F66F61F181400000100400F415200003B403B003200EC00C803B00322C446F0C";
    attribute INIT_38 of inst : label is "C0007D000180007D400180007D000180007D000140007D000140007D3C3C1BC0";
    attribute INIT_39 of inst : label is "0190370C3C1BC0F66F014001C0007D400180007D4001C0007D000180007D0001";
    attribute INIT_3A of inst : label is "03322221111100156ABFC0156AA95403FEA9540A5500A3A8E9FE6DFD92B2B85C";
    attribute INIT_3B of inst : label is "821F4208C823FA72B43FB83EAFED8FABDB0E672873B831E80E4E3EB9BC47E000";
    attribute INIT_3C of inst : label is "DBA5CF277E934DAFD707237D3FFA72C3F0A72DF4FFE9CB4C3D9CB8BDACAD0820";
    attribute INIT_3D of inst : label is "427A797D09E9E5F427A7173330CCCDDDDEEEEFFFFCCCCDB5ED7F9BE070791E47";
    attribute INIT_3E of inst : label is "9E5F4A7A717D29C9E5F4A72797D29E9E5F4672797D19E9C5F4672717D19C9C5F";
    attribute INIT_3F of inst : label is "A29EDC5C8672717219E9E5C8672797219C9E5C827A717209E9C5C827A797D29C";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "246E1051B84046E10D2B8414A0CB0F840420CF2CFE10908FE1050B8034A50D07";
    attribute INIT_01 of inst : label is "F3C70E0CCF30DC7CB31DC3FE1051B84046E10D1B84246E1051B84046E10D1B84";
    attribute INIT_02 of inst : label is "0CF33041000018031810ED8AD86E82D8ED8AD86E82F8B1C3CB2CB2CB0C33CF3C";
    attribute INIT_03 of inst : label is "F32833CCC000C1000300600CA041CF33CF32833008104018032810F31ECF3CCA";
    attribute INIT_04 of inst : label is "10C60584338102833CB30CB71CF33CF32833DC808E01C4001803085600CE043C";
    attribute INIT_05 of inst : label is "384184084284289D63AE39E0850800C104000000C600C2048AF180A2BCE28867";
    attribute INIT_06 of inst : label is "30813530009D75D78B18ECE3B38ECA3B18ECA3B08ECA3B08B3CF32831ECF3FC4";
    attribute INIT_07 of inst : label is "F880040180318101C0833DC808E01C4018031810333CCF3DCA0CC02003040180";
    attribute INIT_08 of inst : label is "CA0CF3200304100600CE04C00180328111D819E01C4018032810F3DCA0CC00CC";
    attribute INIT_09 of inst : label is "0600C6044710047807100600C2043CF72833CCC10450C48000600CE058070F3D";
    attribute INIT_0A of inst : label is "55555550154080001800000401803281033004018031810F3ECA0CF320030410";
    attribute INIT_0B of inst : label is "55555555001403FFFFFF7FAAAA56A96A955AAAAAA95A55655555555555555555";
    attribute INIT_0C of inst : label is "00000001501540550154055555555501540550154055A5565555555555555555";
    attribute INIT_0D of inst : label is "5555555555015405501540555555555015405500140000400100000040010000";
    attribute INIT_0E of inst : label is "0400C10030400C10030000000000555555555500000000005555555555555555";
    attribute INIT_0F of inst : label is "00000000000403C100F0403C100F0403C100F0403C10030400C10030400C1003";
    attribute INIT_10 of inst : label is "0104001001440400044051150015444004010004005011014441041555555554";
    attribute INIT_11 of inst : label is "03281600C204600C2258033891803281600C204600C225803389400000000040";
    attribute INIT_12 of inst : label is "600C604600CE15803285600CA3450D071103600C20503600C20503600CA04018";
    attribute INIT_13 of inst : label is "F023C58F232BCD0E08F00C44B0C0F70CFCF3C610CA158432851803285600CE14";
    attribute INIT_14 of inst : label is "20B000330BCCF0B9060832C308CF5690A088982820D629D8C3240E0883C3208C";
    attribute INIT_15 of inst : label is "15C43081610DE05C43081610D2043DCB2CD075030CF0CF83FC2CB30CF30DC208";
    attribute INIT_16 of inst : label is "15441510400011441005000400001104114054005000400400001C43085610C6";
    attribute INIT_17 of inst : label is "0000144340340094180040C000000C090401000C0804040D080508000C041110";
    attribute INIT_18 of inst : label is "01000003044C34E24C34E34938A38830C30C34A30B34934A30938C1501110408";
    attribute INIT_19 of inst : label is "200CE0000003C00C00F0000000200C103C0000000000000C300000020080000C";
    attribute INIT_1A of inst : label is "0C00040C00000C000400C0000000C00040C000400C0004000020403038010000";
    attribute INIT_1B of inst : label is "0C000C0C000C03000303000203000003000200300000003000203000200C0008";
    attribute INIT_1C of inst : label is "00103000300300010003000303000300C00040C000C0C00040C000C00C000400";
    attribute INIT_1D of inst : label is "080C0C00000C00040C00000C000800C0000000C00080C0008030001030002030";
    attribute INIT_1E of inst : label is "C000C0C00040C00040C00000C00000C000C0C000C0C00040C000400000010000";
    attribute INIT_1F of inst : label is "0080C00080C00000C00000C00000C00000C000C0C000C0C00040C00040C000C0";
    attribute INIT_20 of inst : label is "C10450D070CC00C000C0C00080C00000C00000C00000C00080C00000C00000C0";
    attribute INIT_21 of inst : label is "B0C2C6207600CA3580368D610DE05843781600D60580348143D803289600DE24";
    attribute INIT_22 of inst : label is "78161605468151205878151E05448161E054581516058481BAEB1BAEB5BAEB63";
    attribute INIT_23 of inst : label is "A59A452423180DB650C431F1F5F5F50D9EE7DBDDBFB01C7FE7D11518C251A054";
    attribute INIT_24 of inst : label is "014415FF10147ABD7D7AAAA565655565AAA5956DAFA7956A59AA556A99A6556A";
    attribute INIT_25 of inst : label is "1001040514010450001104001401100000010104005000500041051011040054";
    attribute INIT_26 of inst : label is "36C359F776E72343535CDC926CD343233DCCCF249004E4005154545400050044";
    attribute INIT_27 of inst : label is "0C0CE34363430DF8CE8F08CC251CF52A00A27636DC0D047034D0D8CDF737234D";
    attribute INIT_28 of inst : label is "00CE34343430C0CE34343430C0CE34343430D8FD8C0CE34363430C0CE3436343";
    attribute INIT_29 of inst : label is "CFD4DCE42F39D9CFD473E4EEEE39CFD4DCE62F39D9CFD433D54B50D1C3019837";
    attribute INIT_2A of inst : label is "18C71C7810350C4FB301084FB301095169383CA063DC45444D0353BB9CE40F39";
    attribute INIT_2B of inst : label is "0733333BCC542635320631C78D330631C073C71E1C071F3DF1C1C807292AD4C8";
    attribute INIT_2C of inst : label is "4F25078FA0F4F105429BD1A16F4504147C1D8F11F0763C1F076F67A1F070B5EB";
    attribute INIT_2D of inst : label is "4CF34FC7D7C7355D1A9962163D934F64D3D1F1F51C7359F1F59C734941E3EA0F";
    attribute INIT_2E of inst : label is "03500D4034CB14F053D00D403500D32C73414F400E400ED4D0C34CF3743430D3";
    attribute INIT_2F of inst : label is "A433C903A433C9C3D0EC68E0F93504D4134CB1CD073504D413504D32C53C1CD4";
    attribute INIT_30 of inst : label is "004E533545B41905401194CD516D06415004243E0B084C3FE4C24C3FC3A3F903";
    attribute INIT_31 of inst : label is "4A533545B41905401094CD516D06415004A533545B41905401194CD516D06415";
    attribute INIT_32 of inst : label is "3F3330F34FCCCC3CD133545B404150046533545B41905401394CD516D0641500";
    attribute INIT_33 of inst : label is "D948D01E50D01B8D01E52379436E3794951D55D5DD551E9669866324950043CD";
    attribute INIT_34 of inst : label is "34D834D354D78435A665266524D36A5266CB24955234D3BB94925483434D8D3C";
    attribute INIT_35 of inst : label is "005401000450411450040041104500010411014113114104113523794939980D";
    attribute INIT_36 of inst : label is "0041410510001015050054010401444114410100400001111400114111415044";
    attribute INIT_37 of inst : label is "0040000507FF3FFFFFFFFC050450000405C000C4130003105C004C4101544050";
    attribute INIT_38 of inst : label is "000000C003000000C003000000C003000000C003000000C00300000040001000";
    attribute INIT_39 of inst : label is "30540040001000004000C003000000C003000000C003000000C003000000C003";
    attribute INIT_3A of inst : label is "011111111110000000001555555555540000000000003B60F350CF507588F401";
    attribute INIT_3B of inst : label is "73ED41C7CF3DDDB3D433D1747C755D1F3C702872CB02C20F4022F2C90E68F200";
    attribute INIT_3C of inst : label is "45014D053699620D8D4DB043961487197AC8710E58520DA09720DC751CF5073C";
    attribute INIT_3D of inst : label is "C0D8D0D70363535C0DCD4DA98876547654765476554765334CD50020D0D0340D";
    attribute INIT_3E of inst : label is "3735C0D8DCD70373435C0DCD8D70373735C0DCD4D70373635C0D8D8D70363535";
    attribute INIT_3F of inst : label is "3037F636C0DCD0DB0373736C0D8DCDB0363436C0D8D4DB0363436C0DCD0D7036";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "424B01092C0424B01492C052451052C0528510410B010A10B010A2C07241C078";
    attribute INIT_01 of inst : label is "C71862401C040101405310CB01892C0624B01492C0524B01492C0524B01092C0";
    attribute INIT_02 of inst : label is "41C0AEBAE309C700918D43142141140103102101100106101041041041071C71";
    attribute INIT_03 of inst : label is "C0090702B0BEBAE309E71C02463510471C0090AC2FAEB8C700918D08511C7002";
    attribute INIT_04 of inst : label is "C02450700B14F61441005100510071C00907001C01D62B8C07009141C0246371";
    attribute INIT_05 of inst : label is "727527727727400C3020413400EFBEBAEBC230AE71C02863F04537FC11407D81";
    attribute INIT_06 of inst : label is "0A18F00000F0C30CF863214C85321CC843210C853218C851071C0090511C4027";
    attribute INIT_07 of inst : label is "CAFBEB8C700A189C27907001C01D62B8C700A18D00701C700242B0BEFAEB8C70";
    attribute INIT_08 of inst : label is "0241C0BEFAEBAE31C02862B08C700A18BC21E01D62B8C700A18DC700242B0401";
    attribute INIT_09 of inst : label is "31C02C62F0BDEF0758AE31C02C6371C0090702BAEB1C02FBE31C028601D8DC70";
    attribute INIT_0A of inst : label is "00000000000080002800F8EB8C700B18D008EB8C700B18DC700241C0BEFAEBAE";
    attribute INIT_0B of inst : label is "000000000280095555551555552154955550000000008002000800200A802A00";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000008002000800200A802A0";
    attribute INIT_0D of inst : label is "FFFFFFFF00000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "5555155545555155540000000000FFEAEAEAEA0000000000EAEAEAEAFFFFFFFF";
    attribute INIT_0F of inst : label is "0000000000555415550555415550555415550555415554555515554555515554";
    attribute INIT_10 of inst : label is "0208032D00555555555555555555555555555555555555555555554000000000";
    attribute INIT_11 of inst : label is "008141C020531C02440700810C7008141C020531C02440700810400000000080";
    attribute INIT_12 of inst : label is "1C020531C020507008141C020531C078CCF01C02060F01C02060F01C02C630C7";
    attribute INIT_13 of inst : label is "C747411D0F0F584251C01000CF351E51042431C02050700914C7008141C02053";
    attribute INIT_14 of inst : label is "FDD00F9D41E7741847410310E1DC808DF00F8F7C03800800D0F3C3C0D0109D39";
    attribute INIT_15 of inst : label is "50700A141C02850700A141C028537310400701D041C510B733410051004018B3";
    attribute INIT_16 of inst : label is "5555555555555555555555555555555555555555555555555555C700A141C020";
    attribute INIT_17 of inst : label is "5015095055195215055155C00000000100010400000004010001040400000055";
    attribute INIT_18 of inst : label is "01000404100F34C38F38D30C30D38F3CE38F3CE38C30C34D38E38F0025529505";
    attribute INIT_19 of inst : label is "1000F0000003C00400F0001018500C103C0000000000000C4100000100802000";
    attribute INIT_1A of inst : label is "0C00040C00040C000400C0004000C00040C00040180000000051403038000000";
    attribute INIT_1B of inst : label is "0C00040C000403000103000103000103000100300010003000103000100C0004";
    attribute INIT_1C of inst : label is "00103000100300010003000103000100C00040C00040C00040C000400C000400";
    attribute INIT_1D of inst : label is "18200C00040C00040C00040C000400C0004000C00040C0004030001030001030";
    attribute INIT_1E of inst : label is "C00040C00080C00080C00080C00080C00040C00040C00040C000402000000000";
    attribute INIT_1F of inst : label is "0080C00080C00080C00080C000C0C000C0C00080C00080C00080C00080C00040";
    attribute INIT_20 of inst : label is "BAEB1C07842000C00080C000C0C000C0C00000C000C0C000C0C000C0C000C0C0";
    attribute INIT_21 of inst : label is "B41010DD81C02C407009101C02C60700B181C024407009103C0700B101C02442";
    attribute INIT_22 of inst : label is "818BE062B810AE042FB18AE062B810BEC62B910AE062F9108208082080820800";
    attribute INIT_23 of inst : label is "AAAABAF3F0C743E0040100000000004002C000C00C1741030B4343EF10AE042B";
    attribute INIT_24 of inst : label is "5555540055554A82828AAAAAAAAAAAAAAAAAAAA2A0A8AAAAAAAAAAAAAAAAAAAA";
    attribute INIT_25 of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_26 of inst : label is "1E00C2D43348E0D0D0E34071EC70F303702C2D1C7D3DCD555555555555555555";
    attribute INIT_27 of inst : label is "434020D0E0F34100D00D60310AF1DAF3763030336703009C0CF000C70F4FE0C7";
    attribute INIT_28 of inst : label is "74020D0E0F3434020D0D0F3434020D0C0F3430C00F4020D0F0F3434020D0D0F3";
    attribute INIT_29 of inst : label is "1C0341C1C17000DC0337310444701C0341C3C17000DC033730701E3C70B60F73";
    attribute INIT_2A of inst : label is "63986189C741C372D1145372D114500331C7701D870F1CB070F00D1101C1D170";
    attribute INIT_2B of inst : label is "D84CCCFDC336CDB1CDD8E6189CDFD8C62D8C186263D861C0261601D8FC03C737";
    attribute INIT_2C of inst : label is "DCF0BF0DB5CDCF3C7FDC10FF7043CDB18F630DC63D8C3762D8C301061D84D041";
    attribute INIT_2D of inst : label is "C0B1C25B108B1C408BD13CCC7032C70CB1C396C438B1CF96C4F8B1FC2FC34B5C";
    attribute INIT_2E of inst : label is "C0CF033C0C022C74B1CF033C0CF03008B1D2C73FDC3FDCC03C00C0B1F00F0C00";
    attribute INIT_2F of inst : label is "00E5103700E510F343B60DCDC80CF033C0C022C74B1CF033C0CF03008B1D2C73";
    attribute INIT_30 of inst : label is "D3D0D41C7532C13C74F435071D4CB04F1D3D0F73C1CD5372F513437337071037";
    attribute INIT_31 of inst : label is "D8D41C7532C13C74F635071D4CB04F1D3D4D41C7532C13C74F535071D4CB04F1";
    attribute INIT_32 of inst : label is "1CCCCC71C733331C7D41C7532F4F1D3DCD41C7532C13C74F635071D4CB04F1D3";
    attribute INIT_33 of inst : label is "7CB078772C7871078772C1DCB1C41DCBC8844400CCCCCB4130F20D1C71D3F1C7";
    attribute INIT_34 of inst : label is "1C7F1C71C072C003FFF2F472F071C02F44021C732F1C70113C71CB00F1C70308";
    attribute INIT_35 of inst : label is "5555555555555555555555555555555555555555545555555542C1DCBC0D1F03";
    attribute INIT_36 of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_37 of inst : label is "5555555554004000000001555555555555155515545554555155515555555555";
    attribute INIT_38 of inst : label is "5555551554555555155455555515545555551554555555155455555555555555";
    attribute INIT_39 of inst : label is "4555555555555555555515545555551554555555155455555515545555551554";
    attribute INIT_3A of inst : label is "06666666666005555555555555555555555555500000F00CDC0F300C30002015";
    attribute INIT_3B of inst : label is "043037101C430FF4033703B0DD43ECF7514F094001D02E403F040401D809C580";
    attribute INIT_3C of inst : label is "2CB2C7CB1FD13CC783030C3731C79863203980DCC71E608630E60F80ED00DC71";
    attribute INIT_3D of inst : label is "303C3C30C0F0E0C303C3C3000033332222111100000333E0F832DD80303C0F03";
    attribute INIT_3E of inst : label is "0E0C303C3830C0F0F0C303C3830C0F0E0C303C3C30C0F0E0C303C3830C0F0F0C";
    attribute INIT_3F of inst : label is "0C0F4C0C303C3030C0F0C0C303C3030C0F0C0C303C3030C0F0D0C303C3030C0F";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
