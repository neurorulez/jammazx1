library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_3 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"A9",X"00",X"A2",X"07",X"95",X"9B",X"CA",X"10",X"FB",X"8D",X"08",X"2C",
		X"60",X"2C",X"FF",X"01",X"10",X"01",X"40",X"48",X"98",X"48",X"8A",X"48",X"D8",X"AD",X"FF",X"01",
		X"0D",X"D0",X"01",X"D0",X"FE",X"E6",X"78",X"A5",X"78",X"29",X"03",X"D0",X"0D",X"E6",X"75",X"A5",
		X"75",X"C9",X"03",X"90",X"05",X"D0",X"FE",X"8D",X"00",X"38",X"A6",X"22",X"D0",X"1D",X"A5",X"42",
		X"25",X"43",X"10",X"17",X"8E",X"0F",X"2C",X"A2",X"04",X"CA",X"D0",X"FD",X"A2",X"07",X"8E",X"0F",
		X"2C",X"8E",X"0B",X"2C",X"AD",X"08",X"2C",X"49",X"FF",X"85",X"8D",X"20",X"42",X"77",X"A2",X"02",
		X"BD",X"00",X"24",X"0A",X"B5",X"96",X"29",X"1F",X"90",X"37",X"F0",X"10",X"C9",X"1B",X"B0",X"0A",
		X"A8",X"A5",X"78",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",X"01",X"95",X"96",X"AD",X"06",
		X"20",X"29",X"80",X"F0",X"04",X"A9",X"F0",X"85",X"8E",X"A5",X"8E",X"F0",X"08",X"C6",X"8E",X"A9",
		X"00",X"95",X"96",X"95",X"93",X"18",X"B5",X"93",X"F0",X"23",X"D6",X"93",X"D0",X"1F",X"38",X"B0",
		X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"96",X"69",X"20",X"90",X"D1",X"F0",X"01",X"18",X"A9",X"1F",
		X"B0",X"CA",X"95",X"96",X"B5",X"93",X"F0",X"01",X"38",X"A9",X"78",X"95",X"93",X"90",X"2A",X"A9",
		X"00",X"E0",X"01",X"90",X"16",X"F0",X"0C",X"A5",X"8D",X"29",X"0C",X"4A",X"4A",X"F0",X"0C",X"69",
		X"02",X"D0",X"08",X"A5",X"8D",X"29",X"10",X"F0",X"02",X"A9",X"01",X"38",X"48",X"65",X"99",X"85",
		X"99",X"68",X"38",X"65",X"8F",X"85",X"8F",X"F6",X"90",X"CA",X"30",X"03",X"4C",X"A0",X"78",X"A5",
		X"8D",X"4A",X"4A",X"4A",X"4A",X"4A",X"A8",X"A5",X"99",X"38",X"F9",X"A5",X"77",X"30",X"0A",X"85",
		X"99",X"E6",X"9A",X"C0",X"03",X"D0",X"02",X"E6",X"9A",X"A5",X"8D",X"29",X"03",X"A8",X"F0",X"1A",
		X"4A",X"69",X"00",X"49",X"FF",X"38",X"65",X"8F",X"B0",X"08",X"65",X"9A",X"30",X"0E",X"85",X"9A",
		X"A9",X"00",X"C0",X"02",X"B0",X"02",X"E6",X"8C",X"E6",X"8C",X"85",X"8F",X"A5",X"78",X"4A",X"B0",
		X"27",X"A0",X"00",X"A2",X"02",X"B5",X"90",X"F0",X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",
		X"95",X"90",X"CA",X"10",X"F0",X"98",X"D0",X"10",X"A2",X"02",X"B5",X"90",X"F0",X"07",X"18",X"69",
		X"EF",X"95",X"90",X"30",X"03",X"CA",X"10",X"F2",X"A5",X"90",X"8D",X"05",X"3C",X"A5",X"91",X"8D",
		X"06",X"3C",X"A5",X"92",X"8D",X"07",X"3C",X"A5",X"85",X"49",X"03",X"6A",X"6A",X"8D",X"00",X"3C",
		X"6A",X"8D",X"01",X"3C",X"A5",X"8E",X"F0",X"0A",X"A9",X"08",X"A0",X"AF",X"8D",X"00",X"2C",X"8C",
		X"01",X"2C",X"A9",X"00",X"0E",X"04",X"20",X"90",X"05",X"A5",X"FE",X"09",X"08",X"0A",X"85",X"FE",
		X"68",X"AA",X"68",X"A8",X"68",X"40",X"A9",X"D0",X"D0",X"02",X"A9",X"B0",X"A0",X"00",X"91",X"03",
		X"C8",X"91",X"03",X"D0",X"70",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",X"0F",X"18",X"69",X"01",
		X"08",X"0A",X"A8",X"20",X"F8",X"79",X"28",X"60",X"C0",X"4A",X"90",X"02",X"A0",X"00",X"BE",X"F9",
		X"56",X"B9",X"F8",X"56",X"4C",X"D5",X"7C",X"4A",X"29",X"0F",X"09",X"E0",X"A0",X"01",X"91",X"03",
		X"88",X"8A",X"6A",X"91",X"03",X"C8",X"D0",X"3D",X"4A",X"29",X"0F",X"09",X"C0",X"D0",X"ED",X"A0",
		X"00",X"84",X"06",X"84",X"08",X"0A",X"26",X"06",X"0A",X"26",X"06",X"85",X"05",X"8A",X"0A",X"26",
		X"08",X"0A",X"26",X"08",X"85",X"07",X"A2",X"05",X"B5",X"02",X"A0",X"00",X"91",X"03",X"B5",X"03",
		X"29",X"0F",X"09",X"A0",X"C8",X"91",X"03",X"B5",X"00",X"C8",X"91",X"03",X"B5",X"01",X"29",X"0F",
		X"05",X"01",X"C8",X"91",X"03",X"98",X"38",X"65",X"03",X"85",X"03",X"90",X"02",X"E6",X"04",X"60",
		X"A2",X"00",X"A5",X"06",X"C9",X"80",X"90",X"0A",X"8A",X"E5",X"05",X"85",X"05",X"8A",X"E5",X"06",
		X"85",X"06",X"26",X"09",X"A5",X"08",X"C9",X"80",X"90",X"0A",X"8A",X"E5",X"07",X"85",X"07",X"8A",
		X"E5",X"08",X"85",X"08",X"26",X"09",X"05",X"06",X"F0",X"08",X"C9",X"02",X"B0",X"24",X"A0",X"01",
		X"D0",X"10",X"A0",X"02",X"A2",X"09",X"A5",X"05",X"05",X"07",X"F0",X"16",X"30",X"04",X"C8",X"0A",
		X"10",X"FC",X"98",X"AA",X"A5",X"06",X"06",X"05",X"2A",X"06",X"07",X"26",X"08",X"88",X"D0",X"F6",
		X"85",X"06",X"8A",X"38",X"E9",X"0A",X"49",X"FF",X"0A",X"66",X"09",X"2A",X"66",X"09",X"2A",X"0A",
		X"85",X"09",X"A0",X"00",X"A5",X"07",X"91",X"03",X"A5",X"09",X"29",X"F4",X"05",X"08",X"C8",X"91",
		X"03",X"A5",X"05",X"C8",X"91",X"03",X"A5",X"09",X"29",X"02",X"0A",X"05",X"02",X"05",X"06",X"C8",
		X"91",X"03",X"4C",X"55",X"7A",X"20",X"1F",X"7A",X"A9",X"70",X"A2",X"00",X"A0",X"01",X"91",X"03",
		X"88",X"98",X"91",X"03",X"C8",X"C8",X"91",X"03",X"C8",X"8A",X"91",X"03",X"4C",X"55",X"7A",X"A5",
		X"78",X"29",X"0C",X"D0",X"21",X"A5",X"CD",X"F0",X"1A",X"10",X"1C",X"A6",X"CB",X"A9",X"06",X"8D",
		X"00",X"3A",X"9D",X"00",X"32",X"A9",X"0E",X"C6",X"CB",X"C6",X"CC",X"D0",X"06",X"A2",X"40",X"86",
		X"CD",X"E6",X"CB",X"8D",X"00",X"3A",X"60",X"A4",X"CC",X"D0",X"02",X"84",X"CF",X"0A",X"10",X"35",
		X"B9",X"C0",X"7B",X"10",X"0C",X"85",X"CC",X"E6",X"CE",X"E6",X"CE",X"E6",X"CE",X"A5",X"CF",X"90",
		X"0B",X"65",X"CE",X"AA",X"B5",X"23",X"65",X"CF",X"85",X"CF",X"B5",X"23",X"E6",X"CC",X"A6",X"CB",
		X"9D",X"00",X"32",X"A9",X"04",X"8D",X"00",X"3A",X"A9",X"0C",X"E8",X"E0",X"15",X"90",X"C2",X"A2",
		X"00",X"86",X"CD",X"F0",X"BE",X"A6",X"CB",X"A9",X"08",X"9D",X"00",X"32",X"8D",X"00",X"3A",X"A9",
		X"09",X"8D",X"00",X"3A",X"A9",X"08",X"8D",X"00",X"3A",X"A2",X"00",X"B9",X"C0",X"7B",X"10",X"2A",
		X"86",X"CC",X"AD",X"40",X"2C",X"8E",X"00",X"3A",X"45",X"CF",X"F0",X"16",X"A0",X"02",X"98",X"65",
		X"CE",X"AA",X"A9",X"00",X"95",X"23",X"95",X"44",X"CA",X"88",X"10",X"F8",X"E6",X"D0",X"A6",X"CB",
		X"10",X"B8",X"E6",X"CE",X"E6",X"CE",X"E6",X"CE",X"10",X"F4",X"65",X"CE",X"A8",X"AD",X"40",X"2C",
		X"8E",X"00",X"3A",X"99",X"23",X"00",X"65",X"CF",X"85",X"CF",X"E6",X"CC",X"A9",X"00",X"F0",X"DE",
		X"00",X"01",X"02",X"21",X"22",X"23",X"FF",X"A4",X"CD",X"D0",X"17",X"A9",X"08",X"C5",X"CE",X"90",
		X"11",X"66",X"CD",X"A5",X"D0",X"F0",X"0B",X"A2",X"15",X"86",X"CC",X"CA",X"86",X"CB",X"84",X"CE",
		X"84",X"D0",X"60",X"2C",X"02",X"20",X"30",X"FB",X"20",X"18",X"71",X"A9",X"B0",X"8D",X"03",X"40",
		X"A9",X"00",X"A2",X"03",X"95",X"61",X"95",X"64",X"CA",X"D0",X"F9",X"9D",X"00",X"02",X"E8",X"D0",
		X"FA",X"85",X"DD",X"85",X"D3",X"85",X"FA",X"85",X"FC",X"AD",X"01",X"28",X"29",X"02",X"85",X"FB",
		X"85",X"FD",X"A9",X"01",X"20",X"00",X"63",X"A9",X"98",X"8D",X"E9",X"02",X"8D",X"E8",X"02",X"A9",
		X"7F",X"8D",X"EC",X"02",X"A9",X"06",X"8D",X"EE",X"02",X"A9",X"FF",X"85",X"42",X"85",X"43",X"A9",
		X"30",X"8D",X"ED",X"02",X"20",X"CF",X"7F",X"AD",X"00",X"28",X"29",X"03",X"A8",X"B9",X"6B",X"7C",
		X"85",X"F8",X"85",X"69",X"85",X"6C",X"30",X"02",X"A9",X"01",X"85",X"6A",X"85",X"F9",X"85",X"6D",
		X"A9",X"03",X"2D",X"02",X"28",X"AA",X"E8",X"E8",X"C0",X"03",X"D0",X"01",X"E8",X"A5",X"8D",X"29",
		X"03",X"C9",X"03",X"D0",X"01",X"E8",X"86",X"6E",X"4C",X"44",X"78",X"00",X"20",X"50",X"FF",X"A2",
		X"D5",X"84",X"09",X"A0",X"E0",X"84",X"01",X"20",X"1F",X"7A",X"A9",X"70",X"20",X"EA",X"7A",X"4C",
		X"89",X"7C",X"A2",X"CA",X"A9",X"A4",X"20",X"D5",X"7C",X"C6",X"09",X"F0",X"02",X"10",X"F3",X"60",
		X"A9",X"F7",X"A0",X"03",X"38",X"08",X"86",X"1D",X"88",X"84",X"1C",X"18",X"65",X"1C",X"85",X"1B",
		X"28",X"AA",X"08",X"B5",X"00",X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"E5",X"79",X"A5",X"1C",X"D0",
		X"01",X"18",X"A6",X"1B",X"B5",X"00",X"20",X"E5",X"79",X"C6",X"1B",X"A6",X"1B",X"C6",X"1C",X"10",
		X"E1",X"60",X"20",X"C5",X"7C",X"A6",X"0C",X"C6",X"0C",X"BD",X"00",X"28",X"29",X"03",X"20",X"EB",
		X"79",X"A9",X"0A",X"A2",X"CB",X"A0",X"00",X"91",X"03",X"C8",X"8A",X"91",X"03",X"4C",X"55",X"7A",
		X"A2",X"FE",X"9A",X"D8",X"A2",X"00",X"8E",X"0F",X"2C",X"A9",X"11",X"9D",X"00",X"01",X"A8",X"5D",
		X"00",X"01",X"D0",X"54",X"98",X"0A",X"90",X"F3",X"8A",X"95",X"00",X"9D",X"00",X"01",X"9D",X"00",
		X"02",X"9D",X"00",X"03",X"9D",X"00",X"40",X"9D",X"00",X"41",X"9D",X"00",X"42",X"9D",X"00",X"43",
		X"9D",X"00",X"44",X"9D",X"00",X"45",X"9D",X"00",X"46",X"9D",X"00",X"47",X"CA",X"D0",X"CA",X"8D",
		X"00",X"34",X"8A",X"5D",X"00",X"01",X"D0",X"20",X"9D",X"00",X"01",X"E8",X"2C",X"07",X"20",X"10",
		X"05",X"8A",X"D0",X"EF",X"F0",X"06",X"E0",X"FB",X"90",X"E8",X"A2",X"00",X"8A",X"55",X"00",X"D0",
		X"07",X"A9",X"11",X"95",X"00",X"A8",X"55",X"00",X"D0",X"41",X"98",X"0A",X"90",X"F5",X"A0",X"00",
		X"94",X"00",X"CA",X"D0",X"E7",X"8D",X"00",X"34",X"A9",X"02",X"85",X"01",X"98",X"51",X"00",X"D0",
		X"2E",X"A9",X"11",X"91",X"00",X"AA",X"51",X"00",X"D0",X"25",X"91",X"00",X"8A",X"0A",X"90",X"F3",
		X"C8",X"D0",X"E9",X"8D",X"00",X"34",X"E6",X"01",X"A6",X"01",X"E0",X"04",X"90",X"DE",X"A9",X"40",
		X"E0",X"40",X"90",X"D6",X"E0",X"48",X"90",X"D4",X"B0",X"72",X"64",X"A0",X"00",X"F0",X"0E",X"A0",
		X"00",X"A6",X"01",X"E0",X"04",X"90",X"06",X"C8",X"E0",X"44",X"90",X"01",X"C8",X"C9",X"10",X"2A",
		X"29",X"1F",X"C9",X"02",X"2A",X"29",X"03",X"88",X"30",X"04",X"0A",X"0A",X"90",X"F9",X"4A",X"A0",
		X"07",X"8C",X"0F",X"2C",X"A2",X"20",X"90",X"02",X"A2",X"80",X"8E",X"00",X"2C",X"A2",X"A8",X"8E",
		X"01",X"2C",X"A2",X"00",X"2C",X"01",X"20",X"10",X"FB",X"2C",X"01",X"20",X"30",X"FB",X"CA",X"8D",
		X"00",X"34",X"D0",X"F0",X"88",X"10",X"ED",X"8E",X"01",X"2C",X"A0",X"08",X"2C",X"01",X"20",X"10",
		X"FB",X"2C",X"01",X"20",X"30",X"FB",X"CA",X"8D",X"00",X"34",X"D0",X"F0",X"88",X"D0",X"ED",X"AA",
		X"D0",X"BC",X"8D",X"00",X"34",X"AD",X"07",X"20",X"30",X"F8",X"10",X"FE",X"A9",X"00",X"A8",X"AA",
		X"A9",X"48",X"85",X"0A",X"A9",X"07",X"85",X"0C",X"A9",X"55",X"18",X"71",X"09",X"C8",X"D0",X"FB",
		X"E6",X"0A",X"C6",X"0C",X"10",X"F5",X"95",X"10",X"E8",X"8D",X"00",X"34",X"A5",X"0A",X"C9",X"58",
		X"90",X"E0",X"D0",X"02",X"A9",X"60",X"C9",X"80",X"90",X"D8",X"8D",X"00",X"03",X"8D",X"04",X"3C",
		X"CD",X"00",X"02",X"F0",X"02",X"E6",X"1A",X"AD",X"00",X"03",X"F0",X"02",X"E6",X"1A",X"A9",X"10",
		X"85",X"01",X"8D",X"04",X"3C",X"A2",X"24",X"AD",X"01",X"20",X"10",X"FB",X"AD",X"01",X"20",X"30",
		X"FB",X"CA",X"10",X"F3",X"2C",X"02",X"20",X"30",X"FB",X"8D",X"00",X"34",X"A9",X"00",X"85",X"03",
		X"A9",X"40",X"85",X"04",X"AD",X"07",X"20",X"29",X"80",X"D0",X"06",X"8D",X"FF",X"01",X"4C",X"00",
		X"60",X"A5",X"1A",X"F0",X"07",X"A2",X"CC",X"A9",X"57",X"20",X"18",X"7A",X"A2",X"96",X"86",X"0D",
		X"A2",X"05",X"B5",X"10",X"F0",X"21",X"86",X"0C",X"A6",X"0D",X"8A",X"38",X"E9",X"08",X"85",X"0D",
		X"A9",X"20",X"20",X"E5",X"7A",X"A6",X"0C",X"BC",X"EE",X"7F",X"20",X"F8",X"79",X"A6",X"0C",X"BC",
		X"F4",X"7F",X"20",X"F8",X"79",X"A6",X"0C",X"CA",X"10",X"D8",X"A9",X"57",X"A2",X"44",X"20",X"18",
		X"7A",X"A9",X"93",X"A2",X"A0",X"20",X"E5",X"7A",X"A2",X"03",X"86",X"0C",X"20",X"C2",X"7C",X"C6",
		X"0C",X"AD",X"01",X"28",X"48",X"29",X"01",X"20",X"CE",X"7C",X"68",X"29",X"02",X"4A",X"20",X"CE",
		X"7C",X"20",X"C5",X"7C",X"A9",X"93",X"A2",X"B0",X"20",X"E5",X"7A",X"A9",X"07",X"8D",X"0F",X"2C",
		X"8D",X"0B",X"2C",X"AD",X"08",X"2C",X"49",X"FF",X"85",X"0C",X"85",X"8D",X"0A",X"2A",X"2A",X"2A",
		X"26",X"0D",X"29",X"07",X"20",X"CE",X"7C",X"A5",X"0D",X"29",X"01",X"20",X"CE",X"7C",X"A5",X"0C",
		X"4A",X"4A",X"29",X"03",X"20",X"CE",X"7C",X"A5",X"0C",X"29",X"03",X"20",X"CE",X"7C",X"20",X"34",
		X"7C",X"A4",X"6E",X"A9",X"96",X"A2",X"94",X"C8",X"20",X"71",X"7C",X"A9",X"10",X"85",X"01",X"A5",
		X"F9",X"30",X"0A",X"A9",X"8E",X"A2",X"83",X"20",X"E5",X"7A",X"20",X"90",X"7C",X"A5",X"D4",X"F0",
		X"07",X"A2",X"CB",X"A9",X"F4",X"20",X"D5",X"7C",X"E6",X"76",X"AD",X"04",X"20",X"2D",X"05",X"24",
		X"2D",X"07",X"24",X"2D",X"06",X"24",X"10",X"0F",X"24",X"21",X"30",X"0B",X"85",X"CD",X"85",X"21",
		X"A2",X"15",X"86",X"CC",X"CA",X"86",X"CB",X"A5",X"21",X"F0",X"1C",X"A5",X"CD",X"F0",X"18",X"A9",
		X"94",X"A2",X"72",X"20",X"E5",X"7A",X"A2",X"F2",X"A9",X"57",X"20",X"18",X"7A",X"20",X"FF",X"7A",
		X"A5",X"78",X"18",X"69",X"04",X"85",X"78",X"A9",X"7F",X"AA",X"20",X"1F",X"7A",X"20",X"DA",X"79",
		X"A0",X"08",X"A9",X"00",X"99",X"FF",X"2B",X"88",X"D0",X"FA",X"20",X"A4",X"7F",X"05",X"88",X"05",
		X"87",X"05",X"86",X"F0",X"02",X"A9",X"A4",X"8D",X"01",X"2C",X"4A",X"8D",X"00",X"2C",X"8D",X"00",
		X"30",X"4C",X"3E",X"7E",X"20",X"A7",X"7F",X"A2",X"07",X"3E",X"00",X"24",X"6A",X"CA",X"10",X"F9",
		X"20",X"C4",X"7F",X"A2",X"04",X"3E",X"03",X"20",X"6A",X"CA",X"10",X"F9",X"8E",X"04",X"3C",X"A2",
		X"64",X"CA",X"10",X"FD",X"AA",X"59",X"16",X"00",X"99",X"86",X"00",X"96",X"16",X"C8",X"60",X"A5",
		X"76",X"29",X"03",X"AA",X"AD",X"0A",X"2C",X"95",X"D5",X"A0",X"00",X"A2",X"04",X"D5",X"D4",X"D0",
		X"01",X"C8",X"CA",X"D0",X"F8",X"C0",X"04",X"AD",X"08",X"2C",X"6A",X"85",X"D4",X"60",X"38",X"30",
		X"1C",X"1E",X"24",X"28",X"06",X"06",X"04",X"04",X"04",X"04",X"51",X"78",X"E0",X"7C",X"E0",X"7C");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
