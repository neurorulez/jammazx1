-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "95146D595204A0F241496A0500CCAEECF88036DF24976344BE57AAFF549448A9";
    attribute INIT_01 of inst : label is "4DA26F9D3CE9C2B0D385601A6A403311A69220E96571AFDECD93124ECD931249";
    attribute INIT_02 of inst : label is "667668A827B33B373674AE6CE9525D07F3A79D26CD7689B1A768D44411443475";
    attribute INIT_03 of inst : label is "4D747C204D35FB39D9BE7076B2E9D800D26BA7610349BDFBDF3A69E74D31504F";
    attribute INIT_04 of inst : label is "1B02546842C18041A10B061C5C6944094A474D36751782A0FB920ED65D1F0013";
    attribute INIT_05 of inst : label is "140828ED588806B437550742AEFA023377F08CEFF113B42B15A4045682D4A021";
    attribute INIT_06 of inst : label is "EF749AFB9B9B8B8C37FE7FE66B2682E24B0985245C497123E58A044B50804000";
    attribute INIT_07 of inst : label is "0C603E681AA8738D039C601CE340E7185DEBBFAA0D17CD7F9E183064DDFFFDFF";
    attribute INIT_08 of inst : label is "FBB9C49FE00F6E626C710000C0199644DA2A69939CCE499E1896BD545C0555C0";
    attribute INIT_09 of inst : label is "377369B6B69B3B4EB7B527A63A7B773F0FC27A778F4CF1E9D49DBD70BC39C5A9";
    attribute INIT_0A of inst : label is "271D3B9C65C25311272D238B4EE738D9BF36ECF9FFFEEDDF3FE754C759A6F65D";
    attribute INIT_0B of inst : label is "166240405DB07B9EE7B9CE7BDEE782AE7A9A49C4E12731C79C054F388A95AA9E";
    attribute INIT_0C of inst : label is "31163138C24B21100183AEB0082A741B69A7E86FD6D0DF2DE1D3C3A7076F4E80";
    attribute INIT_0D of inst : label is "1B0E131AB9B7F6BF0E1666308EB67AAF4B9A95286EEC777B0CFEDC02C502C78E";
    attribute INIT_0E of inst : label is "95ECE4DDCEFC3344556DD5805516363276F48CA001241765C6C0DB64C690D8C3";
    attribute INIT_0F of inst : label is "001D8B0BADDEAE037AB84EFED71B820D5ECE4B041CE57A63C3E3BBEF0C05FED7";
    attribute INIT_10 of inst : label is "13B5614A8F6827681A252CE4C6DFDA675A392E40312FED33AB392FEC621039C0";
    attribute INIT_11 of inst : label is "FF8AD600BB22E8721ED1C6D52A05CB846C6EFDFF1063036891AFD85B61948BC0";
    attribute INIT_12 of inst : label is "7664CC3B2E4CC1B2F40212900100100276FC004004009DA5BBABC5CB846C6D22";
    attribute INIT_13 of inst : label is "3338618606E8669866992629E927A69DFAEEB53248222AE558A91622EE548B11";
    attribute INIT_14 of inst : label is "2497484919CC7EAD42FC99A667A4000000000000000000000000000000000003";
    attribute INIT_15 of inst : label is "8D555555569B773DBCF6F8B90772AFD3EFF5C1FD837DBB5D29705FD81BEDDA97";
    attribute INIT_16 of inst : label is "7E3B2BBA42317EEC20817A221427468100B83E6561961858276A292797BF6A20";
    attribute INIT_17 of inst : label is "82366B9D7DF3EFFDF8E25203F7DF7D857A22E091BF6EBDBBF093849D1C1C2B57";
    attribute INIT_18 of inst : label is "4FFE67E9DFB4A08AF0ABF715E50AFA537073533033BDA2059ED1028CF9F55548";
    attribute INIT_19 of inst : label is "5D66D66CC7EB3EB3E9FB3EB3E976FEEE7B74D715FBFC7AFD3641E24F04584FFB";
    attribute INIT_1A of inst : label is "F4DEDC929BA897F985D43FBFB3E7374596AC9B5E984F9B3AD53F3E9FCF4E73FB";
    attribute INIT_1B of inst : label is "BB0C3FCC7DE476FEFDFFDFBE976BA54DAF4846CCF56EEA3ABCF4B3695F731BFD";
    attribute INIT_1C of inst : label is "379BCDE401898998BC7319BC4E27540D95F5F2A8C554532FD44D86537FDFDEEF";
    attribute INIT_1D of inst : label is "F4A7AE8CB78501DB3FC6FEDC9C9D8DC176B49C4FE7F2F4111111133178EFCE6F";
    attribute INIT_1E of inst : label is "E983B7B7CF36FE593EF6851FF19FDF42E93FAC0174D6D65020A525754937EC01";
    attribute INIT_1F of inst : label is "8BACD87718ECDAC0C5965AD2659B5219BF74199B745A3C3F6F4AEB59B91DE5BD";
    attribute INIT_20 of inst : label is "EFBF625C4ED004A291D36E6FB38DBEF0A9FCEAF36D5C1A354254D4E66C3B951A";
    attribute INIT_21 of inst : label is "105A2A2A844842AC456AA0C46AA07B9C854538F0072C27A192BF3CD650C3A0CB";
    attribute INIT_22 of inst : label is "37D8CDC3A3BDE47A99F7BC8F4EAEBE2D67FF4B13A6DDEF80A3A0040568A8AA01";
    attribute INIT_23 of inst : label is "F400000A3FDD6DDB4FA00031328AD7421D4FC81B7F44907FD80824FF6F389D8A";
    attribute INIT_24 of inst : label is "25220A0BFC11D2C09014C712D521565118A551E0AB117507B6D76D77BD7DBB69";
    attribute INIT_25 of inst : label is "5738417E585EF45F5D17B7D350411028E0BE76A5005FE142D227F6B12C5FEAA4";
    attribute INIT_26 of inst : label is "4F3FCEA947A0556DD9D34C4D4E54F5C5C5C0000F000000038D2BDEE2998C2ABA";
    attribute INIT_27 of inst : label is "CDBB64B54825D56497ACD2EF3EE3D42D33F1054398F760C2969878874950EEDD";
    attribute INIT_28 of inst : label is "94F4A53C5AE57AF1A5A155A297ADAD2AAD14BFD6BCAF5FEDFB46B54825C85E5F";
    attribute INIT_29 of inst : label is "04BE6730CBFE9652CDB8A4B0CE92C377BA4B33A4B3771C294F14A70A53C529C2";
    attribute INIT_2A of inst : label is "5B0BFDFDA114B5144836466DB4D24908A2556B05F55FCDF811704BF19FD9C4C6";
    attribute INIT_2B of inst : label is "0C7F0080A02D83FC3E666F61615CE05B8CCC336FCA7E4CB5D49FF513D6B97ED7";
    attribute INIT_2C of inst : label is "B7F9048269B6BE4C16FFF9AC434F64E94FEFE705BD8BCD6C2C29B832C2C29B03";
    attribute INIT_2D of inst : label is "70AE28BEF787B53E2D82BBEFB749580A2C02845820213AE4B8A88221BB7B5B3C";
    attribute INIT_2E of inst : label is "79779F7DEEF40F43335449AFE5911054D376FFF9BE750107FABF90051720EDFB";
    attribute INIT_2F of inst : label is "2F21E09E1ED8B90773E28A55A213BDF7DF9EE161601ABD2304EAF6BA11554DF7";
    attribute INIT_30 of inst : label is "25B89400A9C8117909139145EAA3077E1C8BF133A3B7DAB5E17D0493E0996293";
    attribute INIT_31 of inst : label is "9BBD59812F2FEFB7EFBB92E4CB309D5EBE613EBD7EFDFC60FFEFB84F84CF6EDD";
    attribute INIT_32 of inst : label is "DBD02331A2478C473769725C97968FBED4DDA9C62C029179762C029118D51335";
    attribute INIT_33 of inst : label is "2EFD0B276DEDF237F4D25AFED137DB141F899D7D3934D6D4EE2E39CC557157BC";
    attribute INIT_34 of inst : label is "5C2C515C8D689879AD811029F518B20E20083958BC95A6FB7DA6FB7FA6F9126E";
    attribute INIT_35 of inst : label is "75CB5CB17534D98124F94967D6D767DFE5482ED491504ED5234736CF45AB90BF";
    attribute INIT_36 of inst : label is "A4AB595D456DACAFBACAA7A8861AA8748535C152B3AAFAA233A62FA6EBB2D7AD";
    attribute INIT_37 of inst : label is "E335CCCD199633314CDF336CCCCED5ABA15D32AE815752CACEABEACEABE2B243";
    attribute INIT_38 of inst : label is "C2CCA58E6AA87083271449CB4517327425CDAC777364F0B99A332C6648CC5198";
    attribute INIT_39 of inst : label is "AEAEB66AD95B2C9252488BFE6DB61A3BEFDF709292FFFFFFFFC7FFFF8016EB34";
    attribute INIT_3A of inst : label is "7D915805DD248891160C0480000401AB6D6DB249492020F00000000800180902";
    attribute INIT_3B of inst : label is "D176EADE635BF3FA92FCFB742F43D0BFBEDD2BD2F4AFFA950CFE4C3FDAFD37BA";
    attribute INIT_3C of inst : label is "2AEAEB756EAD96492924F841681A015401510502A4069CB1AAAFB7DCF5EEB900";
    attribute INIT_3D of inst : label is "06490006400240009640A1A49B04609661C387092CB492000000009280008090";
    attribute INIT_3E of inst : label is "158027367CD272616AED20386BF952828259528282090090A498D3278C6F18C0";
    attribute INIT_3F of inst : label is "45690D25A4349610C2F1004050108094EE7E199FACE4167742415EF31F202424";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "77C7CDC66966E505CA6DE44F0000A27C0148C9100ADA4766C055AABB0AD8E9A9";
    attribute INIT_01 of inst : label is "763A9246C0121B81233726647C89A46642EBA43EE9D9C000972D3CB4972D3CB0";
    attribute INIT_02 of inst : label is "7610B31096BB40C89541312A86201B9048D802422543308CA5111988208A4087";
    attribute INIT_03 of inst : label is "9682C99332C8145762D495CB2505B3326D90924C9892D42000049291B6C2612D";
    attribute INIT_04 of inst : label is "20ED326CE6DD90CDB393667E350D9CA5695AB2C9C920313215E4BB2484966645";
    attribute INIT_05 of inst : label is "4F149EEC9916C4E62A69F66BCEC7B93B76026D101220367327B6B19ECB665B12";
    attribute INIT_06 of inst : label is "C964DBF333333329D3FFBFE26EA6F0D0034032B61A0068057A1D29A54C73364E";
    attribute INIT_07 of inst : label is "001818A4A2F00010000080000440002275BF2DB2BD730DF0ACCC9B326E8ECC8C";
    attribute INIT_08 of inst : label is "048809D40002626161700430022228884F44B63410D000814906610D6040C604";
    attribute INIT_09 of inst : label is "D9DE3DCBBB6ACC892C1CC419E441985C5514408EC8138902330CB186E308099D";
    attribute INIT_0A of inst : label is "080132C801D650BB176D04064CB25964C9D3B64CDDB364ED9223B02386622D66";
    attribute INIT_0B of inst : label is "D8E4CF323572D6F7BDEF7AD631AFFADBD6E8C402D31005A0A04941401299A08D";
    attribute INIT_0C of inst : label is "04CB4E6D1C998596EAD4F872653C9F333BF4D2B929A572D4BDA92B52D685AD5C";
    attribute INIT_0D of inst : label is "59203340B9498724882B684408D8D9D87005E399400C80032D2481B96899687E";
    attribute INIT_0E of inst : label is "5F71975DFCDB10B8BFCB5376496CA12069873B9665463B78D0626978D0120068";
    attribute INIT_0F of inst : label is "CC9A52663858FA4063E10D30E52332ECF719765AD083DD6DB0D834C6D1CF30E5";
    attribute INIT_10 of inst : label is "4B53818B989097B1A94480C0C7261CA42C65C0CAB9530E521D65C0D944CB529C";
    attribute INIT_11 of inst : label is "BB874C915B52E8633121E36F5D7C4B840E550200F9E655B152BBB2944A9B8EB2";
    attribute INIT_12 of inst : label is "66990CA24190CA2402E72908998898896913736236225A56CABE484B840E5253";
    attribute INIT_13 of inst : label is "4542824928F487248721D5EA92490528C3AE52C4744D1EC3D850B61ECC287B0B";
    attribute INIT_14 of inst : label is "3AA0692523C419C9D9FC5E96A428383A323232316C7D28387C7C3838333C3031";
    attribute INIT_15 of inst : label is "594504105124D2114A552300908CD59AD9580FB5960A5C01CA08BB593052E0E0";
    attribute INIT_16 of inst : label is "036020034A569205944ACAC162585A5899C9E377C19C18F496AEF0970C438755";
    attribute INIT_17 of inst : label is "556A9084A51D20BB7B4D9B2F25B25B3308701208DBB76295BA55F3AEAFA37040";
    attribute INIT_18 of inst : label is "D802CD1210A1CAD5AF5E8DAB4A55A5554505010004D912CF258967970E94005D";
    attribute INIT_19 of inst : label is "049900B088B2D9643602D96412602105088325A60826AE5249101681930C1006";
    attribute INIT_1A of inst : label is "0971222D616D6D04433E696AEC084918F917E0012DF125E3AF40E1239090F40C";
    attribute INIT_1B of inst : label is "B2805426B6934004A9570E43622448F091B2D9B72C12229607BFB4B27288A432";
    attribute INIT_1C of inst : label is "8F47A3D0600540105BE8F55AAD56D70A73F56DF5382C30502A8265C4804CCBE4";
    attribute INIT_1D of inst : label is "129A005300A24440C11F090B0B0B01A01013E78582C0080000088020F7DB3D1E";
    attribute INIT_1E of inst : label is "8EC91470618C7471DF7DAD159F2B17E020DFC1E82066E0A40524141E0A96A171";
    attribute INIT_1F of inst : label is "92CD1900006CA3F01A69A3F2CD2476262C702610F042D9A00ECF1004BB111962";
    attribute INIT_20 of inst : label is "0B65C580E04EF714D384482C0B2DCDB6DEDBCE056D79A1D74A8ECCB68C802399";
    attribute INIT_21 of inst : label is "DDA04EE55775BD540C73D210FBD374104D48A0A29468546300C2522ACBDBCE90";
    attribute INIT_22 of inst : label is "C74807D012CFEA5E5A19FD4BD19E7B3ACFFC254B4F2C20B3834D7226ABB11408";
    attribute INIT_23 of inst : label is "0694A61B3A22016C0034A5324BB3205B31A375E0489AA184599C28A553E72086";
    attribute INIT_24 of inst : label is "FEF77D9FFE36F5EBAC92C869B437044D7604D70ED259832EDB65B20102082D80";
    attribute INIT_25 of inst : label is "50010689A522238124E0D96D1A5DD23B1CE500D2BE3FE7CD54C81B5BB6FFEDDF";
    attribute INIT_26 of inst : label is "274D9265251179C0326C949160B5D5A083C000074000000596584422840321BA";
    attribute INIT_27 of inst : label is "9A2EA95A89B81F48A0E95405D20818F4AAE76B9C11DF46DB331356AA138FBD37";
    attribute INIT_28 of inst : label is "2B470A552C020C015540CA26E0AA0A245137016B014180BA668B4A89B8088281";
    attribute INIT_29 of inst : label is "E90753FE900404008115012D5004B5402012540125400242B5234A30A508D2A4";
    attribute INIT_2A of inst : label is "3966B48A5C8C74936ECDAD12422C84E49B705F26D0A92200A4D6A005A414EA7E";
    attribute INIT_2B of inst : label is "49226CCA57B268C6884914DE5A795CA2400900A21618C9291D4946D91EC990A4";
    attribute INIT_2C of inst : label is "01268A993691410CDB099088E400CAB49D20CA5A10942299C94F24559C94F245";
    attribute INIT_2D of inst : label is "026A3BD2606CD303763A52DB6064F349B9B66F73E664B40705912D6C000482D0";
    attribute INIT_2E of inst : label is "B6C92C968012616519136C09D71AA29F459B09908A82CB9BF2E959122026D836";
    attribute INIT_2F of inst : label is "40F2B65D716300908CA3B39ACC38996CB22C0CDE59C204DACA080B0252729285";
    attribute INIT_30 of inst : label is "97C9CA725025CE01ECF057382B42DEDEC07026C4C7649362CCF47B4B9E5C2E7A";
    attribute INIT_31 of inst : label is "A384C8108080D920D928541534E65E8101C4BF060608091BFFF2832E32E5C181";
    attribute INIT_32 of inst : label is "6A091C821C2B632594720382E0BD9022DB1592072EE528A4572E6D399B622351";
    attribute INIT_33 of inst : label is "59B56717A5D62EC882AA9C0C895CB1DE41362600B83600D0C4040AC032662041";
    attribute INIT_34 of inst : label is "71095882B3990212443289569461C960C2C48363AA4B494AA3494AA149409409";
    attribute INIT_35 of inst : label is "CDB3F2EFC0181FD40872965F2965BA414D83BB18D8EB2D5E9438671C6A904B95";
    attribute INIT_36 of inst : label is "C0C99F264C86499324996E4D88A4B8986B18A264C8CD0C84D4CC4CC8FE44FCCF";
    attribute INIT_37 of inst : label is "A402500820044021D0054025010554C0D4066A032D0064002B343353333648AC";
    attribute INIT_38 of inst : label is "0910A0686C23434BF420210003140642AD0160A9403CA3200A4030806900A201";
    attribute INIT_39 of inst : label is "404021980600D84100215355A08673F641B202DB703000000007C0007F94C50C";
    attribute INIT_3A of inst : label is "161AE35B0490D51AA80400000000004010026104008740000004000000080000";
    attribute INIT_3B of inst : label is "DA53334AB04EAB864431C8035634050C7220DD8D816341C89825654B6C16D240";
    attribute INIT_3C of inst : label is "0404020801002C208011216DCD735F9DF676C9AD965EFFBFBAD92C9281422331";
    attribute INIT_3D of inst : label is "5C309A5C1A5806960C00E70046E55CAC4A54A956186008000000409080008080";
    attribute INIT_3E of inst : label is "47A5019B2641AA506C201410530C0A802A0C0A802A0C00C0004A0006650CCA1A";
    attribute INIT_3F of inst : label is "00989312624C498931FD210C8A52199F4C38721C9D88D58920057EFEDEF90000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "A9D8DA3D8890BB533692660600CCAC7C286677EFFCE762873C56AA9FA2E24CA8";
    attribute INIT_01 of inst : label is "5BB2D9B36D9B53E3B327C7375423A03760B9380B5869F2F4D9D717DAD9D717DC";
    attribute INIT_02 of inst : label is "657CFBB8E532FEFD2B75FA56EFF014ED366DB3604A75D811475D8CCE38CE74D6";
    attribute INIT_03 of inst : label is "FB6EFD19BF6F561CB364357DD7FCDA3337FF7368CCDF6A5EB366FFFDFB6371CA";
    attribute INIT_04 of inst : label is "E7B1CC5272A54B3549CA9526B12E25319D62FB7F2D39111DB6F6ADBAFB9F4667";
    attribute INIT_05 of inst : label is "264E4E8A14446127168A348C6A99192A54AC49BD70CC293A852CE7148EDD11CC";
    attribute INIT_06 of inst : label is "061054FEDEDEDECEA1FF5FE652B5103900E048B807200C017845963361199323";
    attribute INIT_07 of inst : label is "026810860B30AB55055AA82AD50156A877B41D44CD9E8A7D8458B366CC0C4E4E";
    attribute INIT_08 of inst : label is "22A1497220026E666E710810020ADF1C9786DBD15A70F3CD31C23CB0120B0120";
    attribute INIT_09 of inst : label is "2A254D67299B124C1E2ED02EED02EEC2729D03FCE07D9C0FB34C35EEF7214977";
    attribute INIT_0A of inst : label is "449184957862C31BE1BC424F612552A7A50A8508502850A548A0622019204743";
    attribute INIT_0B of inst : label is "99517232622984231A42108DE75853908644F96C23E5B84692126D2424DB8CB0";
    attribute INIT_0C of inst : label is "D89EDA7B351B4F1C99B19DACCD36B2726F5C73BDACE77BDCD539FA73D4E7A9C8";
    attribute INIT_0D of inst : label is "16BA4C76A8FCF5D79E2F4EF71E6E716E589EB08EFB2A79D29BDBEA33DA33D801";
    attribute INIT_0E of inst : label is "1FD8F5954A8FE7CD62FDDD1865C6FF7E5CF5EE1D39782E4F1DA3BE4F1DE3B9AE";
    attribute INIT_0F of inst : label is "C8976DDA3F967EEE59FBCB9EBE7A1AE8FDCF5B73A9E3F658DE6F2E73699F9EBF";
    attribute INIT_10 of inst : label is "72F2CB4E17F8E4D9B9FB1E9E81F3D7CF363D7B32A079EBE7973D7A6F668E5AC8";
    attribute INIT_11 of inst : label is "F305E7417270A9402FF839B1E18BC285EA3FAD7F5C1218DCD8EADB6B6BB61FE8";
    attribute INIT_12 of inst : label is "10CE6A4D72F6A4D7AC4F89D9D9C8CCCF5F9A32723333D7E36F1F63C285EA3FF3";
    attribute INIT_13 of inst : label is "616B34936EBD35CD35C9726FDF77C3AC7BCA786F58E64629C13A704E208D1823";
    attribute INIT_14 of inst : label is "ACBD2E31C3A18D7DF3A993E4EFBEAD52AD56ADB6A9B2A9B24DB24DB1B24DB24D";
    attribute INIT_15 of inst : label is "C2FBEAFBE9378425F287C1ECE9E71FF3FFCF72C9459FB7F56B932594AEFDBEB9";
    attribute INIT_16 of inst : label is "946BBCE97397C01B1673B381C39C7070E96EFA53F15E51F8E5EED8E44BFEE875";
    attribute INIT_17 of inst : label is "D70ADA10F19C00ADD666E6D1B7FFEDEDD3B7A3DC76FE5FBF77879FBCFCF47B7D";
    attribute INIT_18 of inst : label is "9142AB1B74214A976575A4AEDA5765572037563446FDE19FBFF0CFC70E09D721";
    attribute INIT_19 of inst : label is "DFFFB7D84DDF6DB6FF776DB6DB4C94C7276DB7B756C8F0AB7A5062C609249FF4";
    attribute INIT_1A of inst : label is "6DA4ECF8BE492B610F88D8DB39AF7B1641BAB2D9B54FFE1EB17BA5B716DAE53E";
    attribute INIT_1B of inst : label is "8B9478CADB2572F2F5E8F36FFCFF6F5BFDFEA7FFC76FBAE3B080BFFBCDD3BDDB";
    attribute INIT_1C of inst : label is "28140A07C00500506100816030182E7F5555F7D7D7FC014EE4DEB2B7A5333D1E";
    attribute INIT_1D of inst : label is "10D0201245E7E0020912001617160141005A490582C0A000A00800A282082050";
    attribute INIT_1E of inst : label is "0B08871DD75511C74D35BD06110C128200049141020A40A08F800D0F488491C0";
    attribute INIT_1F of inst : label is "9BC9949D00A822A0186183A201E4564630744614F40388690B4A084039316164";
    attribute INIT_20 of inst : label is "EFFF66F72227359E5DF6ECCF3BC9E6ED9B7F7BAE81DD797273E6A0F4EA6CB994";
    attribute INIT_21 of inst : label is "C8B8646596294A580F7B73C0F3735ED871F0CA0CE6B7963D0B05A4B6E352D35E";
    attribute INIT_22 of inst : label is "04005010601F48AF9383E915D87E3A3E0EAA3572EDAF5EC4EAEC7326C9319658";
    attribute INIT_23 of inst : label is "D9E6304EAD85AEB7F6CF31A9B69BBD61CF3CD9B77CECBADBD49EACBE5835ED13";
    attribute INIT_24 of inst : label is "EDA7C91EAA3CD34C08D8A18CA3195A6596A618E39B3769996DBADDBEB5B5D6FE";
    attribute INIT_25 of inst : label is "C6B5960F858192E4DCBD67BAE2649C6E38F51718C49549E5977BB6D3E4F559B4";
    attribute INIT_26 of inst : label is "B6D5E55581195A652FB6DF758D73A0092D000019800000052A3B44E6184D160C";
    attribute INIT_27 of inst : label is "0F0BE0D2CEAE42ACBDD59729C0005E7FA17A2BD766401A9CA75124AE1AA3752E";
    attribute INIT_28 of inst : label is "E52139483723D7A1F1E1CBB8B92FAF2C5DC5E84DE87AE42F43C2C2EE2F48E6F5";
    attribute INIT_29 of inst : label is "BDE8AFDF5EF8A995A195ABCDBCAFB6BD32BC6F2BE6B9B6CA532539129C994A44";
    attribute INIT_2A of inst : label is "94DB4B24A66136587177EA59659A4632CB9522812E34A0F27A5DDEA9315B1DDB";
    attribute INIT_2B of inst : label is "6E9F86673DBC8928B776EA6B6B6D6CBBB64ED9CDE4276EADF5D7BCDCF6E2DEB9";
    attribute INIT_2C of inst : label is "DF6FB6E65D74BFEA0CF67F7E71F7735CE2CA6B9B2D16DD4D6D6DBC74D6D6DB87";
    attribute INIT_2D of inst : label is "DDB46E6EC99FB26CED1B9BFDBDD35E6ECF7BB79E66672F35EEEB93B1CBD76D7E";
    attribute INIT_2E of inst : label is "FBEFB7DBFBB23239131970A782C7CDA692CCF67F647323C5FBB7DCC77D3A6E5B";
    attribute INIT_2F of inst : label is "7A1CA3912FB1ECE9E7C6EAE2672C3DFFDB3FBB63665BC91332EFADEB9C709B86";
    attribute INIT_30 of inst : label is "692E731993674B9B3B34DC2F6C23E375A65EB366FBF6FDB37B4988F20790F32D";
    attribute INIT_31 of inst : label is "324F74923B326DBD6DBC9725E5B795F7CB6729EB91274DF3AA9ABBC83C8572F7";
    attribute INIT_32 of inst : label is "90CE9667963DBA3A335FDAE4BD0AE0B68DD95B042A47AC9B642A47BD95B33271";
    attribute INIT_33 of inst : label is "6CFD4665F97B346CE6BADFAEF0FFFE8F359B37D323A44E9CA8E8F4BFCF877D33";
    attribute INIT_34 of inst : label is "D4AC7176ECEE46278BE2CE77647969D263876A994673CDA3D3CDA3D3CDA0DFCD";
    attribute INIT_35 of inst : label is "AA146985A153423D4228C9628C96300165C8EB8674F1CBDB9F2D31CBDD2CCE3A";
    attribute INIT_36 of inst : label is "5F08AEE29B94D3740D3754D3F90D5F8BD0CBC6C55AD5AD1D5AD542D54C051AD9";
    attribute INIT_37 of inst : label is "58CF233AC6618CEA23388CE232306C4E6A76B5394B9DC5F36346B56B50BD44D4";
    attribute INIT_38 of inst : label is "36730611BF53CDF55CFFF737EADCCA9E6F32EF53CCEBAD66618CEB19F6338C66";
    attribute INIT_39 of inst : label is "727A8C12A056177DD5367EFCAE452C7FF3FFD9909FCFFFFFFFC03FFFFFAC81DA";
    attribute INIT_3A of inst : label is "94468662FB2E3E46820400000406006A81585DF754D9E0900000080C00080000";
    attribute INIT_3B of inst : label is "F64C3C46F1455AB1511C914776771DC72451DD9DC770B4E2485F6D5CB77BAFB2";
    attribute INIT_3C of inst : label is "0727A8D9532B6BBEEA9B9ED35BD672B722DC8B391939A452658DB6DBA40883B9";
    attribute INIT_3D of inst : label is "BBBEB3BBB3BF8CEFEF89B3AA434168666F9F6ED7DF754C0000000090C0008000";
    attribute INIT_3E of inst : label is "7021018B962751464E34C469420E0191110E00C4440C00C02A421455A12B4233";
    attribute INIT_3F of inst : label is "004A0941082104A09494214DC8D29BBFA8802BD291405179090706A6D6780090";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "CD9CA7F9C8D0323A24DA6206CCCCAFA42866BECB64F961F7D752AADDE6EE75A8";
    attribute INIT_01 of inst : label is "9B74DC9B24D906B9F58D73BEB61550ABE835DC374064FAF6489332DA489332DE";
    attribute INIT_02 of inst : label is "2FA7C88CAF179364BC7BC978F39002F993649B212F79C845E79CC46D3C456CFF";
    attribute INIT_03 of inst : label is "592525F5D9666309F3E2023F9F6A4B7FB3EDA92FAECFAB5EB9367DB7EFB5195E";
    attribute INIT_04 of inst : label is "4B998B3F5C7EF62CFD7BEFD6020EF514ADBD6D266E3D9D5FA61245B2C9696FFE";
    attribute INIT_05 of inst : label is "74CAE9C78DE55F2EADCF2FCE5F7155BF636D1C08D3441FAFF098CEC24C3B37D4";
    attribute INIT_06 of inst : label is "04480FE3A9A3A9B531FFDFF5BF23E9A02680ECBF3404C0028048BF33AF0DB3E1";
    attribute INIT_07 of inst : label is "0A002117C950799C03CCE01E6700F33828C470F86EE4B7DB64993060D0521012";
    attribute INIT_08 of inst : label is "0B463E60E008474042520010031886EE52D2CB9D962975C268C6B4400A0400A0";
    attribute INIT_09 of inst : label is "2EA4CAE6FD95767582A260A0060A00726E9A0B104162582C41D4720703E73DA6";
    attribute INIT_0A of inst : label is "029929C04162629305AE31434A70703D608103044C99224082C6204659202AAB";
    attribute INIT_0B of inst : label is "FE363888FB9ACF398C63B9E6B58E45CCE520C100030408020A004414008DC708";
    attribute INIT_0C of inst : label is "3A2D3337770A86CA078F8FBD14DE66F77199B3AEDF675D3F61FEC1EDA7DA07FA";
    attribute INIT_0D of inst : label is "5C7968F2FBBF6BDAF50D6FAF74BDBFF6BDCC36B7FBAEFDD5BBFFEE45B645A000";
    attribute INIT_0E of inst : label is "65BB6BDCCE77ADCFEA748B5F3CFADADBFF6BD75E3C730C6E3D10B2EE3CCF991E";
    attribute INIT_0F of inst : label is "B5FF3D936EBD4D5BF53D7FED7AD7745D5BB6BD616F5D6E377BBDBFBDFE9DED7B";
    attribute INIT_10 of inst : label is "57FFFF771778AF78B17274F7ECFDAF5A1EDAF3AEFB3ED7AD2FDAF3B5AE2F2B63";
    attribute INIT_11 of inst : label is "FDFFEBA86B69D9772EF8FBD468EAE7775EFAAB554552C9ECAB6D6BEBA7F57354";
    attribute INIT_12 of inst : label is "FAE64EE9FA656E9FB904A2EAAEABAAFBF7EAAFAAEABEFDEFF51BA6E7675EEFA6";
    attribute INIT_13 of inst : label is "70F828E26FFE218E2188EB53FBE4DEB6E0E7EAA23E2BC558BB162AC5FD8B1566";
    attribute INIT_14 of inst : label is "0E3DB73CF963A5659554BB2EE34F1A4B1F1B1E0AEFFAEC424FF9F441F3BDF3BE";
    attribute INIT_15 of inst : label is "C079E0F3C59E0AC46151A8EAFD23967524C673FBD3D57AF463DF3FBD1EABD73D";
    attribute INIT_16 of inst : label is "DE5D8EEDB9E1410B4579D5F9FBC73E7EF5F65C3A78E7EC9DAFD77DAE9BAF5875";
    attribute INIT_17 of inst : label is "D71E7E67D2241156AFA2F6D0936DB6C99F9B32BAA7485D6AC28616B0B0BE5D1D";
    attribute INIT_18 of inst : label is "4D42E74BF6DCF89EECEBA79DD9CEEC567562022EAA26AE09925704580001D701";
    attribute INIT_19 of inst : label is "6925925E475D75D68B5965968B97D79CAA2593315EECDC2961D85FC77FFFF05F";
    attribute INIT_1A of inst : label is "45C78BBF8EE9FF2532B27AFB9D3D3BFBF98C3E4CB484978D3873B0BEC45E5D97";
    attribute INIT_1B of inst : label is "09B67CBAE9BD335E7CF17568BD49BF3D265A6B6F752ECDBA9F776BEB94DEBD4B";
    attribute INIT_1C of inst : label is "0804020D011540114100804020106C77D55F5555D5F6613CD8CEB253B5757F3F";
    attribute INIT_1D of inst : label is "3090241207A5840208120915141401E1008A08140A01E0020A08802282082010";
    attribute INIT_1E of inst : label is "8F4004504104104104103C14180807E02484C1E0204A48F08F00169E00859160";
    attribute INIT_1F of inst : label is "CDBFADDD006882E0030C23E201207446207E4200564A0A288B890404BE317144";
    attribute INIT_20 of inst : label is "949322E726A319976F57267B9EFEFB5F91B73B23A0F5156BB8F57F6BEEEE9D7F";
    attribute INIT_21 of inst : label is "AEF5D777EBA7297F59C5EEF5C5FE6F9D2DAA42B8561D16198065B6946943965C";
    attribute INIT_22 of inst : label is "F12639612E9DE652B853BCCA4001FD6D47FE3317E6F14B4537F2ABEBF5D75EEA";
    attribute INIT_23 of inst : label is "F8C614F5B48336DB77C6303B3688F92DF72ECBBB2E65365E9D994E179D91C91D";
    attribute INIT_24 of inst : label is "A5A2A94BFF8B43470A2E6DDE1D1E973CC333CF679D77BD8FB6DB6B3DDB26DB6E";
    attribute INIT_25 of inst : label is "6318A8168206F2F778BDBCBAF32EAF55A188DB9CE7DFFD05C732D2D1545FF6B5";
    attribute INIT_26 of inst : label is "80D06536EA41B64C1B165A66A61181048100000580000007030910731540082C";
    attribute INIT_27 of inst : label is "73D4D76BF7CF7A3C3DC787B2010145D9DB1CE8D1A40015AD2B91B10F9A72F09E";
    attribute INIT_28 of inst : label is "BDF1AF7A1FA19FAA6E72AFDD3DF353B57EE9EE87EE33F7539CE57BD7CF73F5F6";
    attribute INIT_29 of inst : label is "CDC83CC45CAAA9952481A0C9D8832729D20CF620CF2D756BDEB5EFDAF7ED7BF6";
    attribute INIT_2A of inst : label is "EE92FDB7C77FABEAF6FB57FFBED347BE57BB39AFF73E8396336EFCF8BD4F0F99";
    attribute INIT_2B of inst : label is "45D5776B5ADFCFBCFB2EFF2B2B0424B9E775D99EC7F675E4F9E5DCD5740E0F39";
    attribute INIT_2C of inst : label is "B77975765D74BF4EF79B5DBE5767636ADB5F21CBFF57DF6767609F6676760996";
    attribute INIT_2D of inst : label is "DDA555BC8DC922EE591DC9B6D9DB6EF79775E32E5575FFA1ED71B355EBD6CB64";
    attribute INIT_2E of inst : label is "CB2CB3CDB3B3BB3E224AF66599C48924FB779B5DBDE36159F5E584D5591DB76D";
    attribute INIT_2F of inst : label is "721F46BB6FF8EAFD22D558F2320EE6924D5332622E6AEF11734BACC9CE71CF9A";
    attribute INIT_30 of inst : label is "6D76F38F9F578BD6172EAF2F57A12DABF45ED16A3AD24C91327F985742BA5761";
    attribute INIT_31 of inst : label is "BBE9DD8E7A7B249D249EA7B1E7AEB9F6EF5D7BEFD1A76455FFFD335D35DA3A77";
    attribute INIT_32 of inst : label is "F68F1731762C8AB561999CF63D697C31EC9BD9F77CFFA0C967CCFFB3FCB11B6B";
    attribute INIT_33 of inst : label is "F748DD2ECB9DD0FF6D7DE73357A64A89668B5199757F65F5C0E0F0EFC0111998";
    attribute INIT_34 of inst : label is "DC75BE7476B7D00111EA2F31AB15E5FA7BE7E9399C7CE780D4E7A0C4E78EA675";
    attribute INIT_35 of inst : label is "0431830E0D530231024CFDBECFDBC822A479E8FF7CB15FEFD62F22CDC90ECF4C";
    attribute INIT_36 of inst : label is "CE0D9E2648844915C49158498804909907990AAC5445440C54440444F02CE0C6";
    attribute INIT_37 of inst : label is "662418983138624408842218898D8470E38231C108E08CDC59151151111441C4";
    attribute INIT_38 of inst : label is "8B8869CC188E22CEA200E8899C2221C02888E0C0220080113E6278C4F9890313";
    attribute INIT_39 of inst : label is "BABAA92236469E7D55367E609A135C493A49DD009BFFC0003FC7C0000006B639";
    attribute INIT_3A of inst : label is "A0C48EF37FFE24448E040000040001A8D11B7DE554D9E0000000080000080002";
    attribute INIT_3B of inst : label is "3C1F8094C0C155BC3C6EFD144344511FBF4510D11446DEBF6C16166EDACBACBA";
    attribute INIT_3C of inst : label is "2BABAA991A236F3EAA9BEED3719C62E63398CE319FBD369B4924924E346A8985";
    attribute INIT_3D of inst : label is "3F2E673F37BFB9CFCBBF5FAA491722F323AF1E3D97754C000000009000008000";
    attribute INIT_3E of inst : label is "63008289932000A6428DC3E8AA515475B1515431B1010010A267510F6336E767";
    attribute INIT_3F of inst : label is "00C0180300600C0180C2DCBEA7397D7606A01A58C9184C4111373064AA588313";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "A7A6A1F06D3B4020006C9D6FED00A2FA2D4CA89202DE4066D652AA848AC8A9A8";
    attribute INIT_01 of inst : label is "59BAC9B12DC90615BAAF2AB77251333368F1250B00016204D9B6B25AD9B6B25A";
    attribute INIT_02 of inst : label is "456E499B85A2B626E044C9C0899054913625B9213844C967144C8CFDFCCDEBD7";
    attribute INIT_03 of inst : label is "C96D6D55DB245B311566504CE6DADAEBB64B6B6AAED92040E7FFC96ED923370B";
    attribute INIT_04 of inst : label is "8805000DCE9D3400373860C48ACC88C5214B49BC4671119226DA099CDB5B5D76";
    attribute INIT_05 of inst : label is "5C98BA298115404E0028A02940055524445708D6AA8806E26A529CA959325598";
    attribute INIT_06 of inst : label is "0B00430A6260686B100120030CC0EB102C4012B762058815641920A74A55224A";
    attribute INIT_07 of inst : label is "091014C492488041040208201041008222B5241831616182904489122B09090B";
    attribute INIT_08 of inst : label is "00B4AB50400A00010410A49A09A86D8E40B2496523408201E910C18969489694";
    attribute INIT_09 of inst : label is "688C914EA93244C94242D8402D84004260998502F0A00E14037D7A0D07B4A915";
    attribute INIT_0A of inst : label is "4A40870D98049520E011452421C30346B52A54AB162448B1212DA0AD824460C2";
    attribute INIT_0B of inst : label is "220658888002084200000008421082C109343822D8E091B0295B2052B64220A4";
    attribute INIT_0C of inst : label is "062906050C809596007C48639C760AA21054F60BDDEC17BFE477CAEF95FF23F3";
    attribute INIT_0D of inst : label is "90E1A4C12A2DE786A08C4F4C216FED7F7F72F8C90220A11A282091C521E52000";
    attribute INIT_0E of inst : label is "751FE7D5001F480A8A421656596F80844DE7A99725EA8C4C3028304D302E0618";
    attribute INIT_0F of inst : label is "A293106C08294B75A52529BCF0A2D7CA51BE7F5AC219460DD4E826F752E93CF0";
    attribute INIT_10 of inst : label is "426AD0C9DC5A84DEF968C08888B79E90B7F9E29F221BCF4856F9E2FFFE0B3AE3";
    attribute INIT_11 of inst : label is "955598E4626C9645B8BEA19D7870327A8898AE5583CDF4CBD693FE86EFC9721D";
    attribute INIT_12 of inst : label is "10D840AE63848AE6271423AEEEBEAFE84D9AAAAFBBFA137B68525C326A888B5E";
    attribute INIT_13 of inst : label is "617B2CBABC9F27EB37ED6C4BDC79C8AE0080626E5EE694B28254A594292A52CA";
    attribute INIT_14 of inst : label is "BEF129AD60021CFE95001304CFBEEEAEEB1EEA0D11511150E5515550020C020D";
    attribute INIT_15 of inst : label is "C079E0F3C3B78E617BD5C38891CED0DB6D9C4A901C11C305EF1CA901E08E18F1";
    attribute INIT_16 of inst : label is "11E670894AD36119C04902D1624D5A589F6B620A4C45C29784DFDA85EE326075";
    attribute INIT_17 of inst : label is "D70EDC62F39610BF81EFDB27FEDB6DB614D83E2B3075F183AA3F51F8B8B1E6E1";
    attribute INIT_18 of inst : label is "0168001BE67DD17C08C01818000C00EC9ED8EC9F8EED842916C214148901D701";
    attribute INIT_19 of inst : label is "DB64B64B4CDB6DB689536DB6899B4708286C96375C82C72921097504E7D65550";
    attribute INIT_1A of inst : label is "44C70A074E174050F273030045B1225DF69CBCD890CD979CB96A4094444ECD72";
    attribute INIT_1B of inst : label is "CBB260A0F0306B52C599B3689D9B275E6C4866CAEBE04775F5F5F24D8ED8315B";
    attribute INIT_1C of inst : label is "080402055141041041008040A0506AF55D57F757D77E6932CED8BB4225666230";
    attribute INIT_1D of inst : label is "109022120755D40208120817545541C1008A08140A05F20080A2280282082010";
    attribute INIT_1E of inst : label is "0B2806504104104104102894102813A8640481C4304360E28714040A208481D0";
    attribute INIT_1F of inst : label is "57A3D111002003A8104103A201A07D42207D4200D54208200F29000838352104";
    attribute INIT_20 of inst : label is "CDB6EBC4B08E579652CE7DC771C96FC2DF0DEC26016F39E24ADC9BE5C088A703";
    attribute INIT_21 of inst : label is "CCBC4445B3294A5EE8BF7E3EB76F461009CC0702947054F203CB6DA20852E598";
    attribute INIT_22 of inst : label is "C835B60204854F801110A9F0000002C802ABB00261AE629112662232D991168C";
    attribute INIT_23 of inst : label is "C6B4A6B3844058490635A5A24B1BF14939A15DB062EEBED0812BACB059B5A82C";
    attribute INIT_24 of inst : label is "B6B86D6000C62D336B16896B289780596505978AD25DA62E92412059604B0920";
    attribute INIT_25 of inst : label is "9084190442C243C520F18B009A48D2B329011CD6B575563DD76A9B5C37000CD7";
    attribute INIT_26 of inst : label is "8A5085253D51709C8136484521A41408224000000000000034501404A9223100";
    attribute INIT_27 of inst : label is "0B0AD852E9BC4ECCF1D9DE3961005D7F3572A1C1406AA329AF21A5CC580A2044";
    attribute INIT_28 of inst : label is "21414852B62B1629696CCBA4F16B6B445D278A6D8962C52B4ACA52C93C7EC4C5";
    attribute INIT_29 of inst : label is "F18DCAD798AD062041A1C329A70C26D13C3269C306D1475214A90AD4852A42B5";
    attribute INIT_2A of inst : label is "106CB45B25DEC59364A495820820042C932A482AD0A3330CA59710A8355AB17A";
    attribute INIT_2B of inst : label is "4910464294923AC3A8499863630E66B25449114A155889EDD5B2669798305CB5";
    attribute INIT_2C of inst : label is "4C965CB800506420B1098690C5148A209D3C73AB6356338E6E61BF6CE6E61BB6";
    attribute INIT_2D of inst : label is "16D8B388213A1389D09AFF6DB16D834B01A2CA03FDFC262788BD062408181043";
    attribute INIT_2E of inst : label is "DB6DB6D9022223A550926648997C9008211109869182CB1002D201933125FC7F";
    attribute INIT_2F of inst : label is "6392AA16B9B38891CE0B33DAEE4A4DB6FF7E2D9A59750ED2CBB4248A56708146";
    attribute INIT_30 of inst : label is "B6CB5AC6DC458F158DA8973C6B474FE04478F7EEE5BFDDB3ED922F42FA17A646";
    attribute INIT_31 of inst : label is "328CCBCE82826DB16DB09E27944A16C588942D8B1C385E15AA9AA70BF0B5E3C5";
    attribute INIT_32 of inst : label is "8509DEE75F3F82B8977C1BC4F18C9020A4914975695D829B45495D939493326D";
    attribute INIT_33 of inst : label is "FDF95404C11A73FDE6F3DE26C224D8A847BF77102CA930A280E0F0EFC0077173";
    attribute INIT_34 of inst : label is "61295F84B8C978441B3809230637616252C48921905BC0E2E3C0E2E3C0E0D79C";
    attribute INIT_35 of inst : label is "C711F1C7CA0C77721462134E2134A42148D2B1EB58B509BB963C42166CF0CBE6";
    attribute INIT_36 of inst : label is "40088222288845100451004588C47888C7880284D04D0404504480447E047C47";
    attribute INIT_37 of inst : label is "22200884111C2220089022408988847CE3E631F308F8845F412413413014C0CC";
    attribute INIT_38 of inst : label is "8F98A8C45C6420C06204008800222021D088183E223861111E22184478880110";
    attribute INIT_39 of inst : label is "E2E323A48E9199C3A06174169344517FE3FF16ED6DB00000000000000006A239";
    attribute INIT_3A of inst : label is "B17C934BB4D3E4FC90001000000000923246631E8185C0000008000000002000";
    attribute INIT_3B of inst : label is "5E200076C2D1532424316908C48C230C5A42312308C34399B348100249300864";
    attribute INIT_3C of inst : label is "0E2E32324748ECE1D03331658D63DA99A26689ED12F9E4D2FFCDB6DE280900C1";
    attribute INIT_3D of inst : label is "FCF1DEFCCE7877BE386ECE40C341682763AF5E1670C818000000001000000000";
    attribute INIT_3E of inst : label is "F73421AB57A1AB1000A107811C828A5511802A555580DD0841C620006310E71E";
    attribute INIT_3F of inst : label is "4598330640C819833086B5AAEF7F55A4080741B0E0069C04F20F7726E67D2120";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "E7A6A8D069726D809B65DA4FCCCCA67CD95DC51209DE422EF856AABF9AD9FBAA";
    attribute INIT_01 of inst : label is "D2769122491253B5A7846AB4E80560AB45A56CAA42434418DDB326DEDDB326D9";
    attribute INIT_02 of inst : label is "ED489112AD76A449880D53101AA010B624492240620D501440D5089C308BE6CE";
    attribute INIT_03 of inst : label is "124849758049901A005C30C8049092AF0092424BAC024083424012480242255A";
    attribute INIT_04 of inst : label is "B00D77C4E78F19DB12963C64E11D9DCD615A000282335556E5801900921255E0";
    attribute INIT_05 of inst : label is "CF3D9598E33458E6C069A86B51051142885718C6B2BB62762217BD884B76D5BB";
    attribute INIT_06 of inst : label is "00807100202028291001A00A448C4F507D4136B7EA0FB825783D69AED8CD6ADA";
    attribute INIT_07 of inst : label is "F087D01586D30423D8211EC108F60847A8A8073039684880A060C1830A0A0A08";
    attribute INIT_08 of inst : label is "A4A02AD80FE0808880908210002028AB6AB0123252C40895FD81000380D0380D";
    attribute INIT_09 of inst : label is "78CE1B4F6B3644D94343564235642153C47164236C846D908D4E30340A282B2D";
    attribute INIT_0A of inst : label is "80224020020908040820801090080404A54A152850A94285093C203C02605456";
    attribute INIT_0B of inst : label is "400C5800088621084210842108420644234002110008420040E08081C1001040";
    attribute INIT_0C of inst : label is "062906059CC09CB2000054E71E540AB6113656D568ADAAD0B4296852D0A5A104";
    attribute INIT_0D of inst : label is "32EF04DA6628AD0481ACCC0DC12A5D4AD110A4AB0E418364610091C521C53000";
    attribute INIT_0E of inst : label is "A690AD220109420802A17692CB248404C8AD09D3AD49ADCD36BAB2CD36A6DCBB";
    attribute INIT_0F of inst : label is "83B2006E55015544055D5915A00651D8694AD2DAC418A58C944A645242AA95A0";
    attribute INIT_10 of inst : label is "D66ACDDB7C57AC56BD69498998A2B400942B4E1666115A00642B4E49552912A2";
    attribute INIT_11 of inst : label is "5555988D66798CCDF8AC8D85692966309990DABE4B4E06C3B6BA92024A197511";
    attribute INIT_12 of inst : label is "8809919066891906E715610888AACAAAC192222AA2AAB07A68555D6630998A1F";
    attribute INIT_13 of inst : label is "4140430CAD98CDB45D93725B5861D8AE05516666DC663506A4D1A8351068D41A";
    attribute INIT_14 of inst : label is "EBA62B2520084D6C95A8B32CF7EE0E0C00E0000003BC03BEABBFBBBFFDF3FDF1";
    attribute INIT_15 of inst : label is "C079E0F3C100231B4C2D3132B2445C8B6DCDDA92302040994A29A923430204A2";
    attribute INIT_16 of inst : label is "214041B15A52C018C15806452AC9CB4AB749528AA22A26AAACB552ACAE000075";
    attribute INIT_17 of inst : label is "D708590898D800A95366C965B6DB6DB77054EA8A2800714002A41430B0A14007";
    attribute INIT_18 of inst : label is "12E510894D7C405110104C002000100010110105466DAC2A86D615370E01D701";
    attribute INIT_19 of inst : label is "924DA4DA889A69A7DBE269A7D248281C4049B4B6A512C6D24408DE0CD51459E0";
    attribute INIT_1A of inst : label is "E9081004124708CA72204506474226D54410A09120490412A14465214A902226";
    attribute INIT_1B of inst : label is "B2C17300D04067B4B96A827D20924852489004929248CC4921D1F0124A203393";
    attribute INIT_1C of inst : label is "08040202D04450004100804020100280282082820000028146D9B4026E2AAD56";
    attribute INIT_1D of inst : label is "0090201202F24402081208030303000100820804020048208888800082082010";
    attribute INIT_1E of inst : label is "01088410410410410410148410280028200480A0320260001284840520848000";
    attribute INIT_1F of inst : label is "32592336002000081041014201200006202C42102C0A08200109004804350104";
    attribute INIT_20 of inst : label is "0DB760DDA91ED51456944895255944A6534966E48329254ADA8E88B491B962B1";
    attribute INIT_21 of inst : label is "AAA157754AB18C50D9854A9D855AC4064CCF9E5291F8517307C24966D8868C13";
    attribute INIT_22 of inst : label is "54013880ACE54622B3BCA8C4580003D4A2AAB0164C6AB4B33640ABBAA555546E";
    attribute INIT_23 of inst : label is "46B5EFB3ED84806D8A35ADE64991B74979B053A458A9A2A52354E9ADD2A11464";
    attribute INIT_24 of inst : label is "B2B92726A9E26D7179321A2980524CCB329CB38AD64CC76EDB61B49204900DB1";
    attribute INIT_25 of inst : label is "0002160D8102628922A6CB088BCEF691234420529435529535450B4C97354453";
    attribute INIT_26 of inst : label is "742709E5713751E02000919960000C12001FFFC01FFFFFF04004000040104001";
    attribute INIT_27 of inst : label is "6AD2B662BBE8B309A6613441C00089527AA0A0825BFFEE2BE745DCC8D01B23A4";
    attribute INIT_28 of inst : label is "31D18C74945974C7534EAA6FA21A9A77537D3685362E8B4A9AA472BBE9A6889A";
    attribute INIT_29 of inst : label is "C13713B4137580700925601D478075162E0151E015121A631C318E18C74C63A6";
    attribute INIT_2A of inst : label is "946F345365D8FDB6EE458D900820362FB7681862D1AA2769A5D6232A26D4E256";
    attribute INIT_2B of inst : label is "799055731C922A8288C99C4A4A2C63B648D923C21450D929755A66AF9D7CD7A6";
    attribute INIT_2C of inst : label is "61A00D980448251999693499ED88CA32990C63BBB17633894945BB6494945BB6";
    attribute INIT_2D of inst : label is "627191C3522CCA3166565249262DF35BD9BAF3B35455644D36BD87A6146926DA";
    attribute INIT_2E of inst : label is "9A69A6988EDAA5AD9536EC009B4486DC01996934988A5BBC065A2BB2266C4892";
    attribute INIT_2F of inst : label is "6F16AAB2B90132B24599168A66D909B6DB36EDCACB42105E5A18C4BAD27080A6";
    attribute INIT_30 of inst : label is "93C95AC65194EA298CB132A9999B1A54C95333666DB6DDBB6DD02C5662B30CD0";
    attribute INIT_31 of inst : label is "26919BAECDC449264929744D146AB09810D561302C598855AA92E55955954498";
    attribute INIT_32 of inst : label is "812B566356AD8AB2CB5C7689A68EB289A043520D99552A920D19553BF5222643";
    attribute INIT_33 of inst : label is "6CDB562CCB1A336CEDB6D6E4960A92AAD912226169E805A580E0F0EFC0033731";
    attribute INIT_34 of inst : label is "71695B9B9CEB488C23182B020E2741244255B1219949C076B9C056B9C056B50D";
    attribute INIT_35 of inst : label is "105404141308CAB308E2934E2934B0014C8299094AAF596AD4A8731E6C712926";
    attribute INIT_36 of inst : label is "560AAEAABAA15750157501572A157AAAD7AA07556D56D5516D513D5101D50150";
    attribute INIT_37 of inst : label is "8AAB2AA25540AAA82AA0AA82AAAAAD41480A840552025520B55B55B55F597A95";
    attribute INIT_38 of inst : label is "AC2AE2D5797EABD7CAB97AAE206AABE832AAFA1CAABA045548AA815502AA6554";
    attribute INIT_39 of inst : label is "444D85F605C2B041B03B66DCB608F152449266C938B0000000000000002EAABA";
    attribute INIT_3A of inst : label is "A845835BA4DA244580000000001000D81F0AC106C0ED80000000002000000000";
    attribute INIT_3B of inst : label is "5F5FFF4A8462A7C485B1CE285E85A12C739A13A1285A41489A68B21A6DB08B26";
    attribute INIT_3C of inst : label is "0444D85F02E17820D8163364C731CA8CAA32A8E556720924001B6492CC438085";
    attribute INIT_3D of inst : label is "58200A580A582296081ECF6052534A6543AF0EB4106C0A000000001000000000";
    attribute INIT_3E of inst : label is "7EA4058B96200408110200060008000044AA8000000800806053B00869C0F28A";
    attribute INIT_3F of inst : label is "4584308610C2184308C633AA8C63556EBC3C64B1D228BC16C056EFA6E6790605";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "9D3C1E4BC4C9123664D237A52121AEFA7E2212D964F16787BE51AAD6F1F624A9";
    attribute INIT_01 of inst : label is "1B30DDB36D9BC2F13185E226340100226031103323207AE6C9B6D25AC9B6925C";
    attribute INIT_02 of inst : label is "076CD888E703B66F9421DF2843B022CDB66DB360E521D83CB21DC47CB846E4E6";
    attribute INIT_03 of inst : label is "DB6C6C319B6F7214B36C352DB6D8D82736DB63618CDB6F5CBB66DB6CDB7111CE";
    attribute INIT_04 of inst : label is "6218CC7230E1C335C9CB971D000F723AC5B649252F3D11193692A5B6DB1B04E6";
    attribute INIT_05 of inst : label is "A26F4ECE5EE00F846FC707C60CF00030677D0CCE6966B93B99CC6B632E2D8166";
    attribute INIT_06 of inst : label is "CF7CDCE787878F9477FEFFEEF3A729012484EC7D2024809AAA6DC7183191C3B3";
    attribute INIT_07 of inst : label is "0F783C070190FBDC07DEE03EF701F7B800F734E266CDDE5B8C9D3A74F8D8D8D8";
    attribute INIT_08 of inst : label is "63810876200F6F676F70000002C886064056DB81B64EE34F2846FDFC7F0FC7F0";
    attribute INIT_09 of inst : label is "0E2441E13D813204242433266332640E03833264264C84C990CE3060310909E7";
    attribute INIT_0A of inst : label is "6FDDBFDDFDF6F7BBF7DF77EF6FF77BFBA952A4489522548911E403643918220B";
    attribute INIT_0B of inst : label is "44F8B0000CF8318C6318C6318C630106308CFDEEFBF7BDF7BF1F6F7E3EDFEFBF";
    attribute INIT_0C of inst : label is "320C3231740A070C00031F9D041760234A9D719DEEE33BD8F7B1EF63DEC7BDC4";
    attribute INIT_0D of inst : label is "19983236336EC1B6046E6C23042C636C1CCB32B433BF3D93CD925F4187418000";
    attribute INIT_0E of inst : label is "CBD8C1DDBCEC2168DAE48CDC34D612126EC1941C32646E6C8C47BF6C8D99B066";
    attribute INIT_0F of inst : label is "819B1BD91C845C421171CDD8321392CCBD8C1B339846F67AC361376B188BD832";
    attribute INIT_10 of inst : label is "7366E30692DCE65CB964A4E4CDBB064216307ACEBB1D832136307B6C660E98E0";
    attribute INIT_11 of inst : label is "EECDF6437370C86725B879B265C4C3204CDCF9FF2E38CCDE4D64D8D97B3407C0";
    attribute INIT_12 of inst : label is "66EF4F4B7AF4F4B73D0580C44408C08E65D80002202399617117B4C3204CDB21";
    attribute INIT_13 of inst : label is "6168228A2CD82188A1A863439B658D8F71CC3822182240C819020640CE810320";
    attribute INIT_14 of inst : label is "0C39B4BAD1612D6C41559BE6C60FBFBFBC03BF180208020B1A0A0A0A4E4E4E4F";
    attribute INIT_15 of inst : label is "C079E0F3C70702106841A8C8CD6382E36D8760D9E9D9326673D20D9E0CC9933D";
    attribute INIT_16 of inst : label is "DC190ECDA5B150C740603181C3063470C3761C62E18E18B8E6C45CE6C92E5875";
    attribute INIT_17 of inst : label is "D71A1800D0B58D4DAE62F491B6DB6DECD383B3882E5B4972DB86DDB6B6BC1999";
    attribute INIT_18 of inst : label is "7FFCCF5B56D821A2E03FB207C103E0FFEFEEFEE5622DE68BB6F345CD6A81D701";
    attribute INIT_19 of inst : label is "DB6DB6DE46DB6DB7DBFB6DB7DB64BD80F76DB6B5F3ECFAAB6648E0C748208FFB";
    attribute INIT_1A of inst : label is "ED9D9C9999BA9F31A1C5F8F9BBEF7B22198932D9B065964936739DB6CEDA55B6";
    attribute INIT_1B of inst : label is "8B842DC8D9A47BFAF5E44B7DB25B6C996CD812C85B7BFC2DB34B46DB26F23DDB";
    attribute INIT_1C of inst : label is "08040208800004404100804020101020A882020802823D1C924E9237BF911C8F";
    attribute INIT_1D of inst : label is "1090001202929402081208080808008100820804020050088800088082082010";
    attribute INIT_1E of inst : label is "0148041041041041041010041008010A400480A1220240500000040000848014";
    attribute INIT_1F of inst : label is "0BCD9ED9002081681041002A01200002202D42002D4208200489000402333104";
    attribute INIT_20 of inst : label is "EDB666F612E509D768F76E46918E76DD012C79A2588C116224E3E0DECF4E999C";
    attribute INIT_21 of inst : label is "CCBA6665D32D6B5D17D963C1596277CF64A54AA8C2DF02D8807B6D9C614392DE";
    attribute INIT_22 of inst : label is "B5001141E7BEAE5399F7D5CA4800041E0556313364D3DF44F3602222C1199708";
    attribute INIT_23 of inst : label is "BC63786E32A16492E5E31B3D240CBDA58F0CC9BB6E4430739E140C361CB5E91B";
    attribute INIT_24 of inst : label is "4C45D81554FDD8CEC08DF7C6211C1230C4230CE181337CC124924965996C925C";
    attribute INIT_25 of inst : label is "F7BDF29220249AF658B92CB67020896EC979F38C60CABCC5863BF632ECAABB08";
    attribute INIT_26 of inst : label is "81DC7736D10196245BB6DE668FF7F1EDEFC0001FC0000007BF7BDEF7BDEF3FBE";
    attribute INIT_27 of inst : label is "9324D94AC40F5A6E39CDC7A758C1C459193220C3A46AB28CC6D1A0AE1870EC1D";
    attribute INIT_28 of inst : label is "8C24630817A1D7306460CB103DA3A3265881C925C93AF49324D94AC40E48F6E4";
    attribute INIT_29 of inst : label is "ADED6752DEFE891125B5A1CDDE87377DBA1C77A1C77D2418C30C618630C31861";
    attribute INIT_2A of inst : label is "7BD8C96CB735930C7992C6C924B6C5B863D32FC3270590B3133CCED1BFD9ACCB";
    attribute INIT_2B of inst : label is "8467065AD6D983783224476B6BAD68B92644992CC06E04258984BC0AF076D83D";
    attribute INIT_2C of inst : label is "B6CB30625B2D92EF05B2C9273AE6204CC6676B0B981788ED6D75B07AD6D75B47";
    attribute INIT_2D of inst : label is "9D8C6E2D8D81324C09199B6DBD9B0E8627458A4E848737A1C9613050E9965965";
    attribute INIT_2E of inst : label is "DB6DB6D93B223A32A10C7B678DC049219665B2CB246332E7F1248C411D106F5B";
    attribute INIT_2F of inst : label is "7A59439A25B8C8CD6246E0F0222E2DB6DB17BB20240DE90120472DED2C718316";
    attribute INIT_30 of inst : label is "6C76319D8A470BD33B068C2E6673636BB45CB16231B6DCB97B0981734B9A732B";
    attribute INIT_31 of inst : label is "B3EFF883737B6DB96DB687A1C3039CE5EE0739CBD3A66DC1555D31CD1CDA7AE6";
    attribute INIT_32 of inst : label is "B08C1731162DB8357199D8F439294B9CEDC9DBD7AC4D80DB270C4D919DB11361";
    attribute INIT_33 of inst : label is "6ED80566F9D9B42EC030E7B6F36EDE0B358B11DF3BBC0CFCE0E0F0EFC0111D98";
    attribute INIT_34 of inst : label is "CC14B0646294C833C4E80C01631365DB4B86485D2475C180C5C180C5C188866D";
    attribute INIT_35 of inst : label is "00100004051A42111A18C8A18C8A621AA048608C70B1CD8B172F04C3C18E8E0B";
    attribute INIT_36 of inst : label is "46088E22288045100451004508047888C78802C45C45C4005C401C4000C40040";
    attribute INIT_37 of inst : label is "E003000E001C0023800E003800000040400200010000C4007107117117105884";
    attribute INIT_38 of inst : label is "000010C0006C0007E000600008000003F80000FE0000E100160038007800E001";
    attribute INIT_39 of inst : label is "3A328C1A30440618511409350AC79C1B7ADB9DA4864800000000000000010000";
    attribute INIT_3A of inst : label is "06C06EB0CB6E02404200000000100168C1101861445020000000002000000002";
    attribute INIT_3B of inst : label is "B0C3BFC6C06150B2124C35C4344310D30D610D10C4259C6646923C2592CB649A";
    attribute INIT_3C of inst : label is "23A328C11822230C2880DCD238CE30F303CC0F181D800000002DB6D9B4428190";
    attribute INIT_3D of inst : label is "030C210321030840C301B8A22B4C699774C1D3A9861444000000801A00000A00";
    attribute INIT_3E of inst : label is "F21813522447FBF76EFDF7F9FFAAA40000A8045555A8AA8AA2015007008E2161";
    attribute INIT_3F of inst : label is "007B8F71EE3DC7B8F73631998C63332EE4279D8E0EC30EF1A10F264A48B61210";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "9514144940402912D24152850000A6B47A1132C96CD36506BE51AAC051D56AAB";
    attribute INIT_01 of inst : label is "49324C912489C221120442224001202228912139212122465C9206CA5C9206C8";
    attribute INIT_02 of inst : label is "42244888A221122794248F284910328192249120E5248834A248C478A846C4A6";
    attribute INIT_03 of inst : label is "492424310924660599282D64B248486212492121884924489922492449311144";
    attribute INIT_04 of inst : label is "22084420604081108181021C000D542B4DD4DB6D649111102237AC9649090C42";
    attribute INIT_05 of inst : label is "862D0C440AA006A42D45034204600012233404DEE5229019118429462A248122";
    attribute INIT_06 of inst : label is "0000C8E505050D1837FEFFE6A3A20A002800A4754005100BA12D4D0850914292";
    attribute INIT_07 of inst : label is "000030050290000000000000000000002A6010A22B45D4498000000018181818";
    attribute INIT_08 of inst : label is "03A10910200000000001041042480C0E46E24915AE0E418F4800000000000000";
    attribute INIT_09 of inst : label is "0400088114022008202033260332600A02833262264C44C988C63000012908B1";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000BA54A952A50A1428548E8086830212228";
    attribute INIT_0B of inst : label is "44A8D0000CD0318C6318C6318C63028630840000000000000000000000000000";
    attribute INIT_0C of inst : label is "2008200150840514000216940C32403182C52294E64529C87690ED21DA43B4C4";
    attribute INIT_0D of inst : label is "89A892531126449204E42425046433244CD99298623511114D92CD0105010000";
    attribute INIT_0E of inst : label is "FA884488946421685AA594D455521212264498142326E524946E9324949A926A";
    attribute INIT_0F of inst : label is "8189094B14845442115144C8921110C7A88449128C4EA22A43211329088AC892";
    attribute INIT_10 of inst : label is "5126410A1248A2C89124E464449912423211224F110C892132112324320A0840";
    attribute INIT_11 of inst : label is "488C900721244222249348932544D1284449FBFF2A2A744A15AC484929102500";
    attribute INIT_12 of inst : label is "226C450B22C450B2340500C44408C08A2CC8000220228B23391590D128444925";
    attribute INIT_13 of inst : label is "2028A08224482488248923490B2C848571446022482200400800020044000100";
    attribute INIT_14 of inst : label is "2491B8AB50402526015689224224000003FC00E3FC03FC0000000003FFFFFFFE";
    attribute INIT_15 of inst : label is "C079E0F3C60302112844A8888122825124C440D8A91366C739100D8A089B3791";
    attribute INIT_16 of inst : label is "1819088DC6B1084D0040328142065450813A0C22A08A08A8A24C48A3096CD875";
    attribute INIT_17 of inst : label is "D710080050B005C4AA225208924924A5168222896CDB4B66DA92D51696981991";
    attribute INIT_18 of inst : label is "EFFC444944EC2003803E060701038000000000002224A28A9251450C2841D701";
    attribute INIT_19 of inst : label is "4924924E46492493C9F92493C96DBD8C77249295F78042A92640F6C41C71CFFF";
    attribute INIT_1A of inst : label is "E49D9C8199E09C001005A0E203EF22671C8996489064B24993223C948E4A1192";
    attribute INIT_1B of inst : label is "890471C8582422FA54ACC93C92C924CB244832584928882491898249247211C9";
    attribute INIT_1C of inst : label is "0804020880000000410080402010142A02A80AA022A8311892C892323F33359B";
    attribute INIT_1D of inst : label is "10902012028284020812080A0A0A00A100820804020000000000000082082010";
    attribute INIT_1E of inst : label is "0180841041041041041014041008016200048001000240000000040000848000";
    attribute INIT_1F of inst : label is "09C48A1100200160104101620120284220044200040208200089004402131104";
    attribute INIT_20 of inst : label is "E493324416D4ACD3705326429087325481642A22D94411224647407A45089188";
    attribute INIT_21 of inst : label is "8890444482252948613322863322230954D5ACA5A268826583B924961001A8C8";
    attribute INIT_22 of inst : label is "B3908141A332AA5089E6554A080005544154201121D9CF2A2120222241111208";
    attribute INIT_23 of inst : label is "942168A21291649244A10914028D91D50D05C999244490738A1424924C94AB28";
    attribute INIT_24 of inst : label is "000542155465484A5095574223143651446514C0821175412492496D996C9248";
    attribute INIT_25 of inst : label is "000010521094BA46489125B6505091A2C859F284204AA484922BD212A4AAAA00";
    attribute INIT_26 of inst : label is "811445375021D564599249574000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "9926594A48244C64910C92270041C4492912264392200A8AC6C128244850E41C";
    attribute INIT_28 of inst : label is "846C21183223122121208920910909044904892C8962449926494A4824624444";
    attribute INIT_29 of inst : label is "8C886508C8FF843084E4E1ACDF86B3719E1A37E1A371040846042302118108C0";
    attribute INIT_2A of inst : label is "6B4AC9259514B51468B246DB649245A8A3532D41250481B10164C8D09FC90C80";
    attribute INIT_2B of inst : label is "882C044A52D103303640032929A529920448112D806448249C8DB40AD472C895";
    attribute INIT_2C of inst : label is "96CB10A6DB2CB26504B64B2D6A44404C82E32919883300652534912252534912";
    attribute INIT_2D of inst : label is "14A4A22CA10362081B12892491494A8A25468A4A8485122489A168698B125B6D";
    attribute INIT_2E of inst : label is "4924924B22222223B1146B678DC00494B264B6492C2217A3F2AD880111202449";
    attribute INIT_2F of inst : label is "2251C28C24988881224A22502242649249122940400D88020046248E34710112";
    attribute INIT_30 of inst : label is "2532109488450911290094244A61D12A8448912220924C99295B41518A8C4883";
    attribute INIT_31 of inst : label is "91091105232324912498922482228A448C45148912246541554F3146146E2245";
    attribute INIT_32 of inst : label is "B18813311224A82521C91244912B8B9C44C889D2A4C480C92204C49188911120";
    attribute INIT_33 of inst : label is "264905A2488B946640927232512A4A0A0489111D1990944460E0F0EFC0111198";
    attribute INIT_34 of inst : label is "5818D044A298C01345A00801651125434A84084D2C5480824480824480889265";
    attribute INIT_35 of inst : label is "D867F61BDF084003003080C3080C690AC44028845091449912262C8B43888A1B";
    attribute INIT_36 of inst : label is "99F330CCD33D9A67D9A67D9AB3D9833318330519A19A19DDA19DE19DFF19FD9F";
    attribute INIT_37 of inst : label is "EEEF3BBE777CEEEFBBBEEEFBBBBFFDBDAFECF7F67BFB19FF86686686686DA359";
    attribute INIT_38 of inst : label is "BC3B83DDC1FCEE1FCEF1FBBC386EEFEFFBBBFBFEEEFBE7777EEEF9DDFBBBE777";
    attribute INIT_39 of inst : label is "2223801E00C0041070001B340A429A09224914801248000000000000003FBFFB";
    attribute INIT_3A of inst : label is "02C12A90C96E004102000000000001780B011041C00060000000000000000002";
    attribute INIT_3B of inst : label is "500040C4406152A00058B544024010162D5100900404B8C40EB62C24925B65BE";
    attribute INIT_3C of inst : label is "22223803006022083809D849685A10D503540D0814800000002492483C438090";
    attribute INIT_3D of inst : label is "0208000200020000820288E0094628D23468D1A9041C00000000001800000000";
    attribute INIT_3E of inst : label is "540803428500000000000000005D5400005D5455555D55D5E020700210040040";
    attribute INIT_3F of inst : label is "0000000000000000002421088842110EEC269D884E011674A005425C49D20200";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
