-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "54292AA049326940A502940A502940A502940A502940A5007E532429B203E993";
    attribute INIT_01 of inst : label is "089B026254A2AE108B0803128C0B4C8AA71389C4E271383A674CE99D33A674ED";
    attribute INIT_02 of inst : label is "9679A95BD064EC6F8A80FDC8D732815B0B003001118C89225DEF666711EA3010";
    attribute INIT_03 of inst : label is "C726EC03933C9BE4CF26F933C9BE4DF26F933C9BE4CF2E7D5A959733CD4F679A";
    attribute INIT_04 of inst : label is "307C140726EC7266C726EC7266C4018CE338CE327266C726EC7266C726EC7266";
    attribute INIT_05 of inst : label is "A84D9B28D908FD08D9095909590AC4E31ADFB06185CCBF0DFF1E79F3F43E51E1";
    attribute INIT_06 of inst : label is "28FD0B3610A5D0C5942C842C9A52FCD29F431F431F50FBC54D97F85580BFC05E";
    attribute INIT_07 of inst : label is "7C99E44F27F917CE45B182A55781849450898165DAEF25976BBC965D8EF21976";
    attribute INIT_08 of inst : label is "9C89E723F85F3C8DE46F227917C99E4FF277917C9FE45F267937C8DE4FF22F93";
    attribute INIT_09 of inst : label is "79C8BE722F9C89E722F9C8DE723F9C8BE72379C8BE72279C8FE722F9C89E722F";
    attribute INIT_0A of inst : label is "5F5CF2F787FE89E4DF227933E0BE44B32FC72FDC9BE7A2F9C8DE723F9C89E723";
    attribute INIT_0B of inst : label is "4ABBD048B1F4D34DFFFE2C78A02810F5EDEAD8395B572B617AE7D5F7AFE0F57D";
    attribute INIT_0C of inst : label is "5440810AC5E993D7BC99F56C7F84C04AC8002118F5E800273014334B533652B5";
    attribute INIT_0D of inst : label is "D1432CB22A4FBD3B6C0897DB2C8213EF46D40256FC96FD6FD026D9B4CB0CB402";
    attribute INIT_0E of inst : label is "FFDC89A2605175DE7A768292026392B46D26F937CC9FDBC8307B2FD13E7FA344";
    attribute INIT_0F of inst : label is "9EB800D10BC64C9B3F385005A22A16EAFCDCF38F5F5B1B1D57EAFCAABA6E757D";
    attribute INIT_10 of inst : label is "0A4215CCCDF3F1109D6E4B5C3AF3D87D150FEBEA22BE7E4EBCEB680AD71CF9D7";
    attribute INIT_11 of inst : label is "728805804425E0169E2BCD722674A3F4947EC90C73A649EF46F4BEAAE9B7FD7F";
    attribute INIT_12 of inst : label is "79E79E79E797B55AF3791FE8F7319758A0324CA2E18843108C5E03190C7FC607";
    attribute INIT_13 of inst : label is "95F69257CA5589C635BFB87FFC30286210C42317C80C67031FF1B4BCEED5E79E";
    attribute INIT_14 of inst : label is "33C9BF47F22CE6A6AFDD237CF813C1BE44F2651C9D152791B258DA7E2761BFF9";
    attribute INIT_15 of inst : label is "5F117FF59D513E6D7D61C5AE77CF7CF7CF7CF7CB5559BC8FDE6BDCBBF4CF26F9";
    attribute INIT_16 of inst : label is "FB30FB3D27FFFFF80E79C1CBFDB9D65DB9D064B07FD6DDA9D06C35CE7E59A6FF";
    attribute INIT_17 of inst : label is "7A4FCF586C44B8B11DE7BCCE7301625EB5C0AD2782AD00B001D8E08920FF1050";
    attribute INIT_18 of inst : label is "1E3B069F0F1F834F878EC1A7C3C7E8D7E1E3B46BF0F1FA35F878EF31A300C005";
    attribute INIT_19 of inst : label is "EF4DACFDAB7D5AC6F56FB5DEDAA07D7FB7FE351CDDDFFECFFF768D7E3C7E8D7E";
    attribute INIT_1A of inst : label is "55792901F55555557CC06D5B56B5AD28CBEDB72B13FADBC93FED6F5FB54A5BAC";
    attribute INIT_1B of inst : label is "7F27F23F2655555555559F61556CB4E4836F55555555CEA3D5555B3D3901D555";
    attribute INIT_1C of inst : label is "27F2BF2BF2BF27F27F27F27F27F27F27F27F27F27F27F27F27F27F27F23F27F2";
    attribute INIT_1D of inst : label is "55555555555555555555555555555555555555555555555555555BF2BF27F27F";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "B28EB1C33A8E4BA3855555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "97B0E5C8D5AC33ECA2248525CEE5B22E75A1447395EAF578E78E3472AD9518ED";
    attribute INIT_21 of inst : label is "B3B78620A16A8033711AE039D464649E5AAEAA80002A8000000007E65500752C";
    attribute INIT_22 of inst : label is "2031D8CB10000740407004074000700007400070080740807008074080731D8C";
    attribute INIT_23 of inst : label is "37373B337360A888882023AC20596CBA855555552AAAAAB55282020022000002";
    attribute INIT_24 of inst : label is "EB74D2189A52EA5D8539C8E79E38E38E79E78F31A4269010484D068030D77737";
    attribute INIT_25 of inst : label is "0F7873C39614A4A4E464E492A4924924000000002109AEAAE8CB10897E9A6F49";
    attribute INIT_26 of inst : label is "C6AD5CC0B65A403913E1FE45F86FC73E3DE1EF0E7873E19F1CF8E7C7BE3DF1EF";
    attribute INIT_27 of inst : label is "1010C4556AE17F0BD6919680000002439545AB85FC2F5A461A108421010E555E";
    attribute INIT_28 of inst : label is "BF85E98684210842439555EB85FC2F4C34000000021C8A2F5C2FE17A61A10842";
    attribute INIT_29 of inst : label is "00012988A2E5C2FE17A65A108421094E45562E17F0BD32D00000000872A8B170";
    attribute INIT_2A of inst : label is "7937C9DE4DF87FC3FE99F0DFA6FC37E1FF4EF87FD3FE1BF0DCB85FC2F4CB4000";
    attribute INIT_2B of inst : label is "25B6DEDB727A5202520240000001F6DEDBFCCFD341C99E4FF267937C99E4DF26";
    attribute INIT_2C of inst : label is "0568AEA3337ECC151846FD182460568AE815D3472EAC4E31ADF8000000124949";
    attribute INIT_2D of inst : label is "BF31DCD80A5BA62CF8DDFF7360296E98B36377E980A58CEDF44551806FD98A46";
    attribute INIT_2E of inst : label is "9F8CE338CF702FB9B014B74C59B1BBFEE6C052DD3167C6EFFB9B014B74C59B1B";
    attribute INIT_2F of inst : label is "82FC67417E33A0BF19B6372AB8311CB5706298A0571AB8705C55C382E0A05D34";
    attribute INIT_30 of inst : label is "817F8026116AE8E5ED1968E5A3968E5A39618E6B40F0E2EE40B417E19D05F8CE";
    attribute INIT_31 of inst : label is "0230DBD49E0A1B9584468A2034D02B7332C6D4694400A0140200504A24333A85";
    attribute INIT_32 of inst : label is "A850C32AFE23DDCBCA15FC7E2B5F94554A32C60B12C4B12C4BA8B9EC217A5210";
    attribute INIT_33 of inst : label is "3E5C101F4C9821C1A6887441220E6B4087FFFEA7D4547535A9CD455677DEBDA8";
    attribute INIT_34 of inst : label is "4E633A27319D1398CE89CC6744E633BDF2ABAB1E5ABAB163A0CE3575E371575E";
    attribute INIT_35 of inst : label is "EFE8FEC807901FA8925D4B50905CEB3A572624262451A27319D1398CE89CC674";
    attribute INIT_36 of inst : label is "04FECAFF457EFECFE8817901FAA925D4B72DF98BF5124BA16D6B416FE8AFF657";
    attribute INIT_37 of inst : label is "6D2F2B55D19974BB79C9E21881BF0390E95CEAAB4AFCA2A788BF5524BA16D6B4";
    attribute INIT_38 of inst : label is "7878380052BF8BD33C74C6366CD9B90D8D890C00001970BF4B853B92C46D392C";
    attribute INIT_39 of inst : label is "07777757F75F5F777444444444444444455110CCCCCCCCCCCC00000000006478";
    attribute INIT_3A of inst : label is "55555555555551589C635BF3340C9BD2ECC90224F4BBCD2A7C90A7FFFFF80000";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555554555555555555555450555554515";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "03F0E81E96662CCBB32ECCBB32ECCBB32ECCBB32ECCBB32CC0634C91864F9187";
    attribute INIT_01 of inst : label is "2CF32666DAC6F65DBD6B7727FCDA22E66A3D1A8F46A3D124CC989332624CC99D";
    attribute INIT_02 of inst : label is "077D905D1A619C801782771508C6AA333A6672448A9198560779CEDEFB8E7279";
    attribute INIT_03 of inst : label is "FC5C0FBA2E51708B845CA2E51708B945CA2E51708B8454A6843808BBEC8477D9";
    attribute INIT_04 of inst : label is "11BB2E7C5C8FC5C8FC5C0FC5C0FD9FC0701C0700C5C8FC5C0FC5C0FC5C8FC5C8";
    attribute INIT_05 of inst : label is "7920D2428022A422802380238032824814D0B2ED8FF89D40E820820C089B74F3";
    attribute INIT_06 of inst : label is "C292201249896221230911094C00A7B62D088D888D846D0BC19FFA33239BD3C8";
    attribute INIT_07 of inst : label is "5956CA96513285B9A9462760F5535386D43F5B082710DC69BCD13082710DC69B";
    attribute INIT_08 of inst : label is "3156CC54AE6A7956CA06553289940CAB650B289942CAB650B289944CA9651328";
    attribute INIT_09 of inst : label is "33152CC5533154CC5533154CC54B3152CC55B3154CC5433154CC5533152CC55B";
    attribute INIT_0A of inst : label is "F8A945422A1342CE167033A5946CE846EB7AEB3140CCD4B3152CC55B3152CC54";
    attribute INIT_0B of inst : label is "C7ADFAC5A3192D93924869F252BDAF8A81150B268134D425C5026A04D42C9A04";
    attribute INIT_0C of inst : label is "1F651226C915026C53448B10B8D289C3ACF644999B019298C4BC48D839A4B18F";
    attribute INIT_0D of inst : label is "49B0042491C6E2812C9D8F11092471B8A046D63027B23622459212BCDA24224E";
    attribute INIT_0E of inst : label is "8F7140960492FD6DC54249B12410318E1C634B1B3D8931B259D7623319C4540C";
    attribute INIT_0F of inst : label is "2059921A6C2C31E18849327834F23EBE792C40966662222557BE792AEF901661";
    attribute INIT_10 of inst : label is "676766C48525A50067A61279E48428877990AC3B4F14B4192105E4A49E696B24";
    attribute INIT_11 of inst : label is "40459911236304521E47E0E062058890F11B58AEFFEAD872986958ABBE4DFDFF";
    attribute INIT_12 of inst : label is "2692692692644BBA2D2281B608C49FCC64E03866039147321CC7073FACFFDB9C";
    attribute INIT_13 of inst : label is "0101B0041625049029A299397AB8F0E451CC87311C1CFC6B3FF6D1D1E83E9269";
    attribute INIT_14 of inst : label is "813529A04508CB41E700495133E1960CF067C1B3529A62685622049E465C8E84";
    attribute INIT_15 of inst : label is "C82C420C73ECCCF3259B9FFCC924D34924D34922BB049140719E33708E845526";
    attribute INIT_16 of inst : label is "7002700A43FFFF0D1CB79393FAF3691AF36991C8FF691AE36991491899C4C328";
    attribute INIT_17 of inst : label is "4AE88060A59AC11666EC5D08620B413A72CB9CB30ECC85A1B3A3111D91FF5922";
    attribute INIT_18 of inst : label is "52A0792229503C9114A91E488A548720452A0390229501C8114A9079E449E42F";
    attribute INIT_19 of inst : label is "F891B20CB468A28BE68D457D155F208AFB07CBD2B12DFF92FF58F244A548F244";
    attribute INIT_1A of inst : label is "551A00E02D555555399C0B5004200802A24F47FC280036A0600F8E073F14A201";
    attribute INIT_1B of inst : label is "197597197515555555551939555DDF8FC05B55555554CDC0D5555767E3D13555";
    attribute INIT_1C of inst : label is "7597197197197597597597197597597597197597197597597597197597197597";
    attribute INIT_1D of inst : label is "5555555555555555555555555555555555555555555555555555559719759759";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "130169AC0C010BC0555555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "4B4154905394046125024A469A65121578900680590D86C01241300B0899981F";
    attribute INIT_21 of inst : label is "18F3040043A5002A6800D20DB0005457404F3300003300000000785500007858";
    attribute INIT_22 of inst : label is "02418CE1A40407004070000740407400070000700C074080740C0700807618CE";
    attribute INIT_23 of inst : label is "888C4400444075F5F4A021A6BA61AB34D0CCCCCCCCCCCCC66600000202000002";
    attribute INIT_24 of inst : label is "1FFFB5BDF6C13026FAC1A1869A698618618699E73E3EF0F9F29B3DA95D48C888";
    attribute INIT_25 of inst : label is "D8A6C536288404848444C49C12492492B6DB6DB6F6B7754702A673E049603006";
    attribute INIT_26 of inst : label is "52E7CE7BFEBF7976819D4DA967026C93609B34D9A6CD1468B3459A2C51628B14";
    attribute INIT_27 of inst : label is "3DEF1A3CFDCF1478B9C7ADCE5394F5BC6CF3F73C51E2E71EB729CA72DEF1A380";
    attribute INIT_28 of inst : label is "8A3C5CBDCA729CB7BC68E3B73C51E2E56E5394E5ADE3671DB9E28F172B7394E5";
    attribute INIT_29 of inst : label is "4E5BDE3671CB9E28F172B7394E53D6B1A3CF5CF1478B95B9CA729EB78D9E7AE7";
    attribute INIT_2A of inst : label is "B6C5960DB067933C99E4CF267933C99E0CF067833C19E0CF0173C51E2E56E539";
    attribute INIT_2B of inst : label is "B69242493B0B7B037B0B6124248212424823C0FEDBB62CB16D836C1B62DB06D8";
    attribute INIT_2C of inst : label is "2DF3E77644E1532FDD69C2A65F62DF3E7CB91AA0F12824814D149242493B6DED";
    attribute INIT_2D of inst : label is "22BB1025576C357A43B11440955DB0D5E90EC4555576DD352886F9D29C226DF6";
    attribute INIT_2E of inst : label is "F7B80E0B83E4FA204AAED86AF4876228812ABB61ABD31D88A204AAED86AF4C76";
    attribute INIT_2F of inst : label is "10A5C10852E0842970604E797DA799F2FB4F93C16679FDE6D9CFEF36CDBB6AA7";
    attribute INIT_30 of inst : label is "8C5B9A68C3955F8B592B896E25B896E25B8238ADA57EFFFC8F70851F04214B82";
    attribute INIT_31 of inst : label is "F673F03C084FB10F9EE35E75BFB57FCBBE74B2DE0C89913626C4C8DC691FC0B1";
    attribute INIT_32 of inst : label is "34EBAE8D70539999F67B350C7ECFECEEC0A99CDC771DC771DCB9C09B87235BF9";
    attribute INIT_33 of inst : label is "CED9DDAAE9753BD377DC908A9578AD851C2225001988902E373988ABA985910D";
    attribute INIT_34 of inst : label is "B8AE085C57042E2B821715C10B8AE0636797F26CF97F264E256CF3FECD673FEC";
    attribute INIT_35 of inst : label is "DA15215129D4839D6EF4ADB92AE02C0DFC4F4F4D4DAB85C57042E2B821715C10";
    attribute INIT_36 of inst : label is "892117928BCDA11251139D4839F6EF4ADBB63C5873ADDE9DB05E29B215790ABC";
    attribute INIT_37 of inst : label is "16D1C6AAABFF3B0DDF136631CA9FDADAB6F0C7FFB67F677BD5873EDDE9DB05E2";
    attribute INIT_38 of inst : label is "AAAA58003E5B56157259BD143850EBFB7FDBDBB6DB7AE7887ED2BEBD4143EE81";
    attribute INIT_39 of inst : label is "07FDD7DDD7F577DD501010010100505001141400222222220000000000014398";
    attribute INIT_3A of inst : label is "555555555555525049029A05EF2A0C01317BCA83004C7BF587BF587FFFF80000";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "55E6CAAE2745BB74EDD3B74EDD3B74EDD3B74EDD3B74EDD07C490CE4A6729C86";
    attribute INIT_01 of inst : label is "9BAA054093A4A8716ADBC21508549AF131D0E8763B1D0E5322644CA995322651";
    attribute INIT_02 of inst : label is "C451384B0321E8628501B7F40EF4381A14DDA7BB710D56358A50A8A522F26893";
    attribute INIT_03 of inst : label is "A7D0AA23EA1F40FA87D0BEA5F42EA87D4BE85F52FA17503A84A80EA289E24513";
    attribute INIT_04 of inst : label is "001D0A67D0AA7D0AA7D0AA7D0AA1181C0701C070FD02A7D02A7D02A7D0AA7D0A";
    attribute INIT_05 of inst : label is "1899D48A800AA40A800AA40B8004655050AA20AD26FA0AE1A30EBF76ED9A7051";
    attribute INIT_06 of inst : label is "4AA4085862A960AA475205401195924A8183A902A91500C2B525529529AAB4D1";
    attribute INIT_07 of inst : label is "D756BA25D1AE8D5EA077A2D868181960843B48B6D84920DB6526CA4906DB0924";
    attribute INIT_08 of inst : label is "BF52AFD4B26C5744BA25D52E8D756BAA5D12E89756BAB5D1AE8D746BA25D52E8";
    attribute INIT_09 of inst : label is "2BF52AFD42BF50AFD4ABF52AFD42BF52AFD42BF50AFD4ABF52AFD4ABF50AFD4A";
    attribute INIT_0A of inst : label is "8FA9754BEA1D50BAA5D52F897D6BA27453EC53BD42AFD02BF50AFD42BF52AFD4";
    attribute INIT_0B of inst : label is "B54BA8B541F69A4D64B2527F9DC669FA15F5293E8527D0A6750BE817D024FA84";
    attribute INIT_0C of inst : label is "A593B93085D40BAE1D40EB11EF9874B4B2332650EB84CCCEF42AE6561BA92D6A";
    attribute INIT_0D of inst : label is "70256C00EEB77E81EB156C4B093BADDFA87085ADDA5692692766B6EA14119DA5";
    attribute INIT_0E of inst : label is "7BBF40E5A76CEA3EF543CEAD3AA7AD68B45A9AD7B16EEDDA70B458EADDB7540B";
    attribute INIT_0F of inst : label is "CAF418E786E03873A289931DCF183C96D9DE116333377777FD16D9803EDA2D9E";
    attribute INIT_10 of inst : label is "939381C2007A401572EC1F8E325971DE8E3BC6F4F1AF482C964FD131E39E9592";
    attribute INIT_11 of inst : label is "87BB70EEDC5ADB8EF4D00F095892AA485549160EB9D8965B50755C00FB6FAA6A";
    attribute INIT_12 of inst : label is "0A28820A288C1350A0BEA55C4FF4848D309964558D695AC26B101ADE0B6A9D30";
    attribute INIT_13 of inst : label is "54492D513588CAA0A156212D6E889B5856B09AC5516B7D42DAA757752ABA2882";
    attribute INIT_14 of inst : label is "81F42FA97D00EB536C110B05AEE9774BBB5D903D50025BAA05BAC8E041587130";
    attribute INIT_15 of inst : label is "D13913CDCB3BBEC354ED694B145104104145145635425F50DB6B3D52EA97543E";
    attribute INIT_16 of inst : label is "D480D000419249BD0B69F15D53BBDEEBBBDCEE70AADEEBABDCEE715A9DB119CA";
    attribute INIT_17 of inst : label is "80F805508F72A13DC1EA3DA94B0286DBACF6EB631BAB01436DBBF12E29AA6180";
    attribute INIT_18 of inst : label is "499D1CA924CC8E549267472A49332B91249995C8924CEAE4492665A0E188E00A";
    attribute INIT_19 of inst : label is "04D839B73C1DE1DD3383C3A7022A82A895C56D4A5BF754FBAA6CB912933AB912";
    attribute INIT_1A of inst : label is "553D18D8D1555555344A2456B5AD63581983C0D436C6D8C8478280D80A96C06D";
    attribute INIT_1B of inst : label is "4AC0AC4AC0E5555555541325554FBBA331B455555554C3B1155557EEE8CD6555";
    attribute INIT_1C of inst : label is "C4AC4AC0AC4AC4AC4AC0AC4AC4AC4AC4AC4AC0AC4AC4AC4AC4AC4AC0AC4AC0AC";
    attribute INIT_1D of inst : label is "555555555555555555555555555555555555555555555555555556AC4AC4AC4A";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "EB9254AB435218A4855555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "3000BAA988850297E1FC693F490CEE76141536B49D6EB71922527493A75D3924";
    attribute INIT_21 of inst : label is "5CE8860021CE002C28205040A084588BA162BC00003C000000000066550014D5";
    attribute INIT_22 of inst : label is "20132C758C0C07C0807C0C078080780C0780807C08078080780C0780C07B32C7";
    attribute INIT_23 of inst : label is "6226AAAEAEE00A00AA104A2A1201040A283C3C3C0F0F0F078182020022000002";
    attribute INIT_24 of inst : label is "136491D6DB512224DA469D34514534D34D34511A224A8929CCE9DC8C52462226";
    attribute INIT_25 of inst : label is "743BA1DD0EBC98181C9818196DB6DB6CEDB6DB6CE73841160AA699C8D9223046";
    attribute INIT_26 of inst : label is "46B2DB69346948EAE15E0AB15783AA1D50EE87743BA1DF0EE07703B81DC0EE87";
    attribute INIT_27 of inst : label is "8E73DC3019BAB7D4A9699EE319CE3BCF74C066EADF52A5A63B8CE718E73FD301";
    attribute INIT_28 of inst : label is "5BEA569EE718CE7BCF74D066EADF52B47738C673CE7F86833756FA95A3B8C673";
    attribute INIT_29 of inst : label is "E31CEFB86023756FA95A3B9CE319E73FC3411BAB7D4AD1DCE718CF79EE9A08DD";
    attribute INIT_2A of inst : label is "2AED576ABA57D2BE95F4AFB57D2BE95F4AFA57DABE95F4AFA46EADF52B47719C";
    attribute INIT_2B of inst : label is "B72490925B437B037B43704909210490920A97924D576ABA55D2AED574ABB55D";
    attribute INIT_2C of inst : label is "89FDADBC1FAB9E7B152F5F3CFC489FDAD33F7680584655050AB52490925B6DED";
    attribute INIT_2D of inst : label is "EEAC7676FC36EC50CA6771D993F8DBB14329DDDB6FC370595EC3B156F57BC7C4";
    attribute INIT_2E of inst : label is "6E366D9B675850ECC9FC6DD8A1D4EEE3B3B7E1B76286533B8ECC9FC6DD8A194E";
    attribute INIT_2F of inst : label is "E8EDB3F476D9FA3B6CD2775BAF765D575EEC3B0BC7EB2F375FD979B86E99CF3D";
    attribute INIT_30 of inst : label is "245A4A5C42D13B4E90B285AB16A85AB16A97B4EECDEDDB6B0E1F4746CFD1DB67";
    attribute INIT_31 of inst : label is "D5ACADEB5E673209B981134CA491B35376E4C6ECA0E43C8390720E46E479B891";
    attribute INIT_32 of inst : label is "99BA492778FA556B7866306255DAE0FCB2A9A51485A1485A14EEFDF35B568ED3";
    attribute INIT_33 of inst : label is "EA4D88B3CDEC98C3C515DF63D334EECDDAEEE621CCCCC7331CA4CCCFFCEFA9C5";
    attribute INIT_34 of inst : label is "74ED9FBA76CFDD3B67EE9DB3F74ED95275BAFF6EABAFF6EC8D8FD65F6F7F65F6";
    attribute INIT_35 of inst : label is "F2B9AF9C3C0498B3E5A78FE3F8F45916A83C2C3C3C89FBA76CFDD3B67EE9DB3F";
    attribute INIT_36 of inst : label is "1FAFDD17EE8F2FDAFDC2C0498B1E7A7CFF1B811B167CB4F1F85420DAB9D17CE8";
    attribute INIT_37 of inst : label is "450595A272EF6903BE9B04290FB58A0A9AA02515F2D707EC19B163CF4F9F8542";
    attribute INIT_38 of inst : label is "33DC480049D7975BAF39CE3A64C9DD1D39999CC9249CDD581450510504511104";
    attribute INIT_39 of inst : label is "F82A000A0028280A82221221222AFFAAFBBFEA00040000400000000000004223";
    attribute INIT_3A of inst : label is "555555555555508CAA0A1543B63C8C1120ED8F2304486DB486DB48000007FFFF";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "D56606AA316F9FBF5AB5FBF5AB5FBF5AB5FBF5AB5FBF5AB457781AFD2D788C0A";
    attribute INIT_01 of inst : label is "BBDF2AE7C3BE2A7DEAD5EF33BC8EC0F9F1B8FC6C3E1B0F576AFD5D8BF1762FD0";
    attribute INIT_02 of inst : label is "8EEAC8E3030284FA8621F4C4029610113E9B37366F7BBEEB8948CD63713038A9";
    attribute INIT_03 of inst : label is "FB1437F5884C426293141880C4072831498A4C426213949C808802F75662EEAC";
    attribute INIT_04 of inst : label is "18450E7B14BFB14B7B14BFB14B715F8C2318C230B14BFB14B7B14BFB1437B143";
    attribute INIT_05 of inst : label is "01C194888008A4088008A408800108A62AA5DE47DD5CB84120138A142B74E581";
    attribute INIT_06 of inst : label is "88A40A5A6AA140880440044031951042A1822002201100C3F0F7F9CC1D63ECB5";
    attribute INIT_07 of inst : label is "046023111888C0562814A0B85D1B5BE0C0124D369A49A4934DB4DA4D349A6DA6";
    attribute INIT_08 of inst : label is "EC403B108370C46223911888C046023011808C046223111C88C447223111888E";
    attribute INIT_09 of inst : label is "8EC403B100EC423B108EC423B108EC403B108EC423B100EC423B100EC423B108";
    attribute INIT_0A of inst : label is "C6283141DA4C5033919C8CE04F03381678AE78AE523B948AC403B100EC423B10";
    attribute INIT_0B of inst : label is "F6E23CF5E0F4DA6D6D927B4BBCEF616296C42958852B14A7B909C85B90A57214";
    attribute INIT_0C of inst : label is "A0B05AB44AE405CC0C406314C35A7774160B56997304DED2943466CE1B291CED";
    attribute INIT_0D of inst : label is "34292900EFF15CA0CFF8E8CA403BFC572830EBBC48140040064436C60E109DBB";
    attribute INIT_0E of inst : label is "70AC407387E82712B901CFBD376B3DEF2F7899C4BBE6D8547876F9E7C5731027";
    attribute INIT_0F of inst : label is "CA2D5AE386761E3B0181A34DC7181465B19A71D93939393F7565B1FF985E3B8E";
    attribute INIT_10 of inst : label is "B0B0AD87C3925155B49A19A692793CCC8E19C66471824E249E4335B669A49493";
    attribute INIT_11 of inst : label is "93BE6CEF9AF9D34DEA5E1AA9FB88A00314003E528C39EEDE485453FE6173FEBF";
    attribute INIT_12 of inst : label is "8820820A28A892D8E49C806422952A0F2891247F9CFDF9FBE796B9EB57BFC96A";
    attribute INIT_13 of inst : label is "94699C51B782114C5549BDC6C53BCF3F6E7AF9F45AE7A95DEFF26D6502B928A2";
    attribute INIT_14 of inst : label is "84C5062031022A605AA102010C806403211B002E5043F9CA178BE8017F4C6FA4";
    attribute INIT_15 of inst : label is "B0BD198BE83BC282C7F0F2BF94514514510410442D504E40CB692E5262939098";
    attribute INIT_16 of inst : label is "9010901E2224930287A6C0740B8AEEA38AEBEBFAC1EEA39AEBEB7E52A57319E2";
    attribute INIT_17 of inst : label is "D852C334EEA669BA95A5344A5243DD959FA4E7CEB577A1EEC94A75AAADFF2DB0";
    attribute INIT_18 of inst : label is "9E394E8D4F1EA746A78F53A353C721D1A9E3D0E8D4F1E8746A78E7978781471F";
    attribute INIT_19 of inst : label is "A97C0C99DD04686511A0D0A34757DF7F58E32E5CECB3FE59FF2E9D5B3C7A9D5A";
    attribute INIT_1A of inst : label is "55480008F555555560223D58800000041FE0D225125B4C6A02A4A568927BE8B4";
    attribute INIT_1B of inst : label is "0000000000D555555555D10555741008917D5555555500915555590402257555";
    attribute INIT_1C of inst : label is "0000400000400000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "55555555555555555555555555555555555555555555555555555C0040000000";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "4314C0E050940885055555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "2820114420AA1915234044061CA4421C1132B4251848241140D410A302190944";
    attribute INIT_21 of inst : label is "BA6400000180803838287050E0A0700309824000004000000000000000001010";
    attribute INIT_22 of inst : label is "00131C6B800403004030040300403004030040300403004030000300003331C6";
    attribute INIT_23 of inst : label is "FFFBF73337200AAA000A0208082906082003FC03F00FF0180000000000000000";
    attribute INIT_24 of inst : label is "9376DBDFDB5582A0924ADD308A4926D32C229B9AF5D1D74DFCFD4FCC795BFBBF";
    attribute INIT_25 of inst : label is "3819C0CE02882C246068603169A69A68E9A69A68E7324D26C826D1E88322B454";
    attribute INIT_26 of inst : label is "F80CB479346B58CCC04E033113818E4C7267033819C0CE067833C19E0CF06783";
    attribute INIT_27 of inst : label is "CC625C20C923131C9DEDCCF73CC731897083248C4C7277B733DC731CC625C20E";
    attribute INIT_28 of inst : label is "898E5ECCF73DC73399F083248C4C72F667B9EE399C4F841924626397B33DCF31";
    attribute INIT_29 of inst : label is "E7B9CCB849824626397B33DCF73CCE65C20C123131CBD99EE7B9E6732E106091";
    attribute INIT_2A of inst : label is "8CC066033013809C046223111809C04E023111888C04E0270048C4C72F66799E";
    attribute INIT_2B of inst : label is "B7B6D2DB7B4B7B037B4B716D2DA316D2DA3029DB6A6623311988CC0660331198";
    attribute INIT_2C of inst : label is "8BAF1B6C13B88FB2DEAF791F6A38BAF1B62F66C030108A62AA55B6D2DB7B6DED";
    attribute INIT_2D of inst : label is "C87EF6649C15CDB9CCE7539D92785726E733D91B49C1704FE47B2CEAF791F6A7";
    attribute INIT_2E of inst : label is "DC6E7BD6E63D39CEC93C2B937399EC87B3B4F0AE6DCE67BA9CEED382B937399C";
    attribute INIT_2F of inst : label is "C85F73662FBDB217DCB879175A9AE44EB535CD7DF9A75A9AA6BAD4D7355DE79E";
    attribute INIT_30 of inst : label is "5CF419ACDCFBF6C58D998CC7331CCC63319B6C66C5CD9AD79F5642DDCD98BEF6";
    attribute INIT_31 of inst : label is "AFBE387F3662D78D3DE3D2CAF6D9575779F88A58B0FC3DC7F0F71FE17AB34B73";
    attribute INIT_32 of inst : label is "8CB4CB57897D2BF6D56B62A3E4B5AABFF209A7AC8BB2E8B32CEC4B7E72D6FF99";
    attribute INIT_33 of inst : label is "53E6EAB9E5DCDB72DBCAF649936C66E5B7555328844464E98DCC444C467368DD";
    attribute INIT_34 of inst : label is "6C7B9B363DED9B1EE6CD8F7B66C7B9B9917599B227599B3675F34EB3349AEB33";
    attribute INIT_35 of inst : label is "3FC8FC8FE5A3E85CF8F132DD90BC771FDDE7E7F7E7B9B363DED9B1EE6CD8F7B6";
    attribute INIT_36 of inst : label is "E5F88BBC45D3F88F88FE5A3E85CF8F132DD958F50B9F1E265AEE6E5FC8BBE45D";
    attribute INIT_37 of inst : label is "510713B7F98ADBEB758819CE336B5C479DF61FA4D9AD55F58F50B9F1E265AEE6";
    attribute INIT_38 of inst : label is "119848AAA465E19BCB1AC7F7EFDFF91919B9BCCD34DD918B0450045551005050";
    attribute INIT_39 of inst : label is "539113B113C143B1176747747677222224488AEECCCAACCCEEA38798782A85DD";
    attribute INIT_3A of inst : label is "555555555555502114C554BBB27EAD1586EC9FAA4541EF34DEF249CD5535715C";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "80583C034014AD5AB56A4489122D5AB56A4489122D5AB56A964D1896AC4876C1";
    attribute INIT_01 of inst : label is "2EC0BC57AAED485932716AB402C248E8944A05028944A0A8D50AA1546A8D5097";
    attribute INIT_02 of inst : label is "0410101CEBB0228AD7EBB5843CC724AAB2324664CE601290824001884084222F";
    attribute INIT_03 of inst : label is "9E14C99B487A53D29E90F4A7A43D29E9074A3A41D28E9470A3288CA080830001";
    attribute INIT_04 of inst : label is "9D59AC5E1449E1449E1441E1441D172A4A02A0A0E14C9E14C9E14C1E14C1E14C";
    attribute INIT_05 of inst : label is "454AC352ACB21AB22CB288B288B62B0F47148374099AE942ACA49224591A774A";
    attribute INIT_06 of inst : label is "D288B0384940EB688B44594446A4D32523ACA22CA22510AB914D551953CA89E4";
    attribute INIT_07 of inst : label is "3851C28E14F0A73D20EE370A8492922AE60105820A2006400C821024B0494082";
    attribute INIT_08 of inst : label is "38418E1047805853C29E14F0A7853C29E14F0A7851C28E1470A3851C28E1470A";
    attribute INIT_09 of inst : label is "E38418E10E38438E10638418E10638438E10E38418E10E38438E10E38418E106";
    attribute INIT_0A of inst : label is "AD29E90F083A51D29E94F4A7851D68C50B390B38538E10E78438E10E38418E10";
    attribute INIT_0B of inst : label is "102C04102B9925B6082008B2539CE5C21B843170863E14C4E90F0A6E10C5C298";
    attribute INIT_0C of inst : label is "89255326ABA43F0C7843D38A8812891124AA64C5C31A909CC6A8CC92BD86852A";
    attribute INIT_0D of inst : label is "46B814109916708729C420950D26459C29CAE084032A1AA085BA082812A82248";
    attribute INIT_0E of inst : label is "4B3A538084A6A96CE10E09042D180429564B225B242C01965D110808591694C1";
    attribute INIT_0F of inst : label is "AA23970B37BA1BB58C4972EE165DCB97018C3103B33333B2801709D5305E2410";
    attribute INIT_10 of inst : label is "2C2C2AC94736EBEA3AF11B2CB6D534F02CDE478165E6DA2DB5420E2CCB2DBDB6";
    attribute INIT_11 of inst : label is "4065D91977084EF3616025B50B494823690D42D8A520020B9D791D54C169A8EA";
    attribute INIT_12 of inst : label is "F3CF3CF1C7146B2E22B0838F1CC4BA1259C07044B739AE7339DD8E63C9AAAD59";
    attribute INIT_13 of inst : label is "48340520C0AC561E8E2AB1B171E1C5CE6B9CCE6796398E726AAB59993C20CF3C";
    attribute INIT_14 of inst : label is "83A41C20E9478C0030B60D15F4C7AE3D30E986B851EB4B0830A33400688A80D0";
    attribute INIT_15 of inst : label is "E42E0B2E632ED8FB85B83941E79E79E79E79E79AB283584341B4BA51C28E1474";
    attribute INIT_16 of inst : label is "510B51010192488351EF2B1952A34BCAA34DBCDAAA4BCAB34DBC5F9CD9146A2D";
    attribute INIT_17 of inst : label is "4C8040CCC0C9998322E8DD91C4E84922C6C9319BE441F4249223BD1091AA892B";
    attribute INIT_18 of inst : label is "4E11AF6CA708D7B653846BDB29C2B5ED94E15AF6CA70AD7B653844C214F517AA";
    attribute INIT_19 of inst : label is "564E19B31D8C6CC531B1D9A7657D7DDE69A9270A71B754DBAA6D5ED89C2B5ED9";
    attribute INIT_1A of inst : label is "5508000041555555000090500000004004B1D95436C6DEF272B2B2D8CA927C6D";
    attribute INIT_1B of inst : label is "0000004000055555555511015544180000025555555400009555510600010555";
    attribute INIT_1C of inst : label is "0000000400000000000000000000000000000000000000000000000000400000";
    attribute INIT_1D of inst : label is "5555555555555555555555555555555555555555555555555555540000000000";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "08252C0494655649555555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "08434C351A713D604C9A023987090D4B48840009400502C2502567283840B25B";
    attribute INIT_21 of inst : label is "4019FFFFFC658047014A029C15268D5068497F80007FFFFF80007FFFFFFFC841";
    attribute INIT_22 of inst : label is "0340200404080040800408004080040800408004080040800408004080040200";
    attribute INIT_23 of inst : label is "C888440444400AAAAAC10D34234808A0C00003FFFFF000000002202121020223";
    attribute INIT_24 of inst : label is "C59B6F636DA0F41E40223412092012092090400E40B30AC18732092BC048CCCC";
    attribute INIT_25 of inst : label is "3471A38D18E818105818106012D92D9292D92D9294A30C32D298657220140E81";
    attribute INIT_26 of inst : label is "0042E13658AD6974A38D1D29E3471838C1C68E3471A38D1C68E3471A38D1C68E";
    attribute INIT_27 of inst : label is "294FB10045C28E104426394A56B4A53E4201170A38411098E7295AD294F90005";
    attribute INIT_28 of inst : label is "47082229CA56B4A73E4401170A384111CA52B5A529F63008B851C2088A7295AD";
    attribute INIT_29 of inst : label is "5A529F61009B851C2088A7295AD29CB90004DC28E10445394AD694E7C8C026E1";
    attribute INIT_2A of inst : label is "7483841D20E307183843C20E1071838C1C21E1070838C1C60B70A3841114E72B";
    attribute INIT_2B of inst : label is "00000C000030000000300E00C01CE00C01C0066DB3A43C21E90F487A43D20E90";
    attribute INIT_2C of inst : label is "78863001C20198B0562C0B316017886300AC50030362B0F4714A000C00000000";
    attribute INIT_2D of inst : label is "AA0785535B9F218A105446114D667C86284111081599C70A2CEB0562C0B31601";
    attribute INIT_2E of inst : label is "4A25491A450F4B0882B73E431420A88CA29ADCF92C5082AAB2AA6B73E4B1420A";
    attribute INIT_2F of inst : label is "05B12A00D891006C48885BBC01B8EED80371DC512B6C01B8ADE00DC771112CB3";
    attribute INIT_30 of inst : label is "D69A2F8F7CC2424C43E01F017C05F017C04B64C6F5A34521C9800DA4880B6254";
    attribute INIT_31 of inst : label is "20E781A14C7508A213200498DB6C45A5DB3C2A900BC9596B6D6CAC954E60315A";
    attribute INIT_32 of inst : label is "9CB261C75E72043C0146BE70D5E002B414A6184020982608821374C0CFA1C929";
    attribute INIT_33 of inst : label is "48EE8CB32DCB9693D0C6C06E0EE4C6D5D20007C2CCCCCC4918A4CCEECCE7D1E5";
    attribute INIT_34 of inst : label is "64C9503264881932540C9922064C91003BC01BA76C01BA744596D80374B78037";
    attribute INIT_35 of inst : label is "7019819B66399C60C41492FD9EBC4B1204C3D3C3C30603264881932440C992A0";
    attribute INIT_36 of inst : label is "65819880CC47019819B66399C60C614D2ED9C7B38C18829A5E82B65819880CC4";
    attribute INIT_37 of inst : label is "0050000482EF81C4DC9B884253C0AF6398130814C30015A87338C18C2925E82B";
    attribute INIT_38 of inst : label is "01326D960018740663A0218D1A3426F6F65652B25B22E145B450015554000555";
    attribute INIT_39 of inst : label is "F94141414104014144446666646D7FD7FDDFF7888CC888CC894355555434C732";
    attribute INIT_3A of inst : label is "55555555555556C561E8E288DA3703A0F2368DC0E83C3680436804000007DBF6";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "3C5321E299DC64C993264C99326DDBB76EDDBB76E4C99324F86B28B594586D93";
    attribute INIT_01 of inst : label is "664E20C40A70694A1A352A3828A135E6582C160B0D86C3542A8550AA554AA954";
    attribute INIT_02 of inst : label is "10820154CB6488A597B3FC8684A6A33E3176EEEDD803314848021088660E2665";
    attribute INIT_03 of inst : label is "0A1A90890D487A43521A90F487A43421A90F487A43521E10F5A814A4900B4920";
    attribute INIT_04 of inst : label is "11092D4A1A90A1A90A1A90A1A90D522A8AA288A221A98A1A98A1A98A1A98A1A9";
    attribute INIT_05 of inst : label is "D137C03A013A133A133A813A8120100F802083DC1B33E447A324D3AF4D9AFF23";
    attribute INIT_06 of inst : label is "7A81380559E013A13D009D4084F4BB6F80CE84CE8075030B8B5D5763F71E9B8E";
    attribute INIT_07 of inst : label is "404A0240120094343D252504E2969712D4C4925B6D965B65965964964B65B249";
    attribute INIT_08 of inst : label is "286A0A1A00000048024012809004802401200940480240128090048024012809";
    attribute INIT_09 of inst : label is "0286A0A1A8286A0A1A028680A1A0286A0A1A0286A0A1A028680A1A028680A1A0";
    attribute INIT_0A of inst : label is "A43C21E10D0878024012009004802425452145286A0A1A028680A1A0286A0A1A";
    attribute INIT_0B of inst : label is "0D14810B129B2CB3D34CC5D2D6BDED43D087A590F4B21A95A1A10F021E164342";
    attribute INIT_0C of inst : label is "5C6CD6AF8886810B486842C6A0961B8B8D9AD5F142D2B0B4A4814CA13F804210";
    attribute INIT_0D of inst : label is "A0B45C02BB8A50F0B8F3158700AEE29434228C43337E13E135BE13A9312106DC";
    attribute INIT_0E of inst : label is "C9286A4C75A62884A1A12BE3AC84621280856429261586935918870E290A1E18";
    attribute INIT_0F of inst : label is "9A11D29A6404D42782252A4934D0A068455C42B22222222000684D55241052B2";
    attribute INIT_10 of inst : label is "656575D69C36C400A5045269B6D32882699004134D06DCEDB4C044249A6DB5B6";
    attribute INIT_11 of inst : label is "64EDD83B76C42EC0746FC5A6C663E84C7D09B19CF7AD815840F439549040A9AA";
    attribute INIT_12 of inst : label is "8208208208260299A1D0F004A4A4F908E382A0984315862B18BAE62678AABD9A";
    attribute INIT_13 of inst : label is "0C2722309C40201F0042E9A9689580C5618AC62EBB989ADE2AAF4149E5E00820";
    attribute INIT_14 of inst : label is "F486A43521E25C0485E30F0900900480240120A86A0AC50F4C53A65E670A0E98";
    attribute INIT_15 of inst : label is "8BAF0C58752EE5C62AB53421800000000000000329C2E87A6DB9286843C21E90";
    attribute INIT_16 of inst : label is "D023D0280249250599800215FAD36BAAD76ABA5CFF6BAAC76ABA58B489084D34";
    attribute INIT_17 of inst : label is "2ACD9D26F99A4DE66DC638000A8A2B7242DB90BB6CD0C515B712991595AAD963";
    attribute INIT_18 of inst : label is "8006291A4001148D20018A469000452348006291A4001148D20008E644F9262A";
    attribute INIT_19 of inst : label is "F892912A56A83483A0D56975AA8A20A19605490011A754D3AA685234000C5234";
    attribute INIT_1A of inst : label is "5508020201555555000090500020080004156A6A24A490984D55549755B48549";
    attribute INIT_1B of inst : label is "00040000002555555554B1015544180000905555555410001555510600012555";
    attribute INIT_1C of inst : label is "0000000000000000400400000400000400000400000400000400000400000400";
    attribute INIT_1D of inst : label is "5555555555555555555555555555555555555555555555555555500000000040";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "0000000000004000155555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "0000000000003C00000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000FFFFFC000001010202040406000000007F80007FFFFF80007FFFFFFF8000";
    attribute INIT_22 of inst : label is "2000000004080040800408004080040800408004080040800408004080000000";
    attribute INIT_23 of inst : label is "CCCC888CC8880000000308204100300200000000000000000020002200022002";
    attribute INIT_24 of inst : label is "ADDB6D216DF03E076D963090080092012012086F0D94365596B3C93947CCC88C";
    attribute INIT_25 of inst : label is "1E10F48784D804044004044592DB649392DB64929DAEBEE9FA13757A5CCE85D2";
    attribute INIT_26 of inst : label is "BBED0BB2DDAD2940F407A03D01E10F487843C21E90F086843D21E10F48784352";
    attribute INIT_27 of inst : label is "6BDA9249C503C21E061729CA56B5AF6A4927340F0878185CE7295AD6B5A9249B";
    attribute INIT_28 of inst : label is "E10F0129CA56B5AD6A4927140F0878094A52B5AD7B524939A07843C04E5295AD";
    attribute INIT_29 of inst : label is "5AD7B526939A07843C04A7295AD6B5A9349C503C21E025394AD6B5AD4924E681";
    attribute INIT_2A of inst : label is "80B405802D01600B405802C01600B405802D01680B405802D140F0878094E52B";
    attribute INIT_2B of inst : label is "000000000000000000000000000000000000046DB605A02C01680B405A02D016";
    attribute INIT_2C of inst : label is "2E96C4DCC10514A5A0AA02294792E96C4F288927040100F80200000000000000";
    attribute INIT_2D of inst : label is "B7439D9B130F1607045DBE766C4C3C581C1176E49110F300089A5A0AA0229479";
    attribute INIT_2E of inst : label is "466098260B4F071912261E240E08B95CE4D89878B03822EDF3B36261E2C0E08B";
    attribute INIT_2F of inst : label is "3333049999824CCCC10D4A30E4AC88E1C95996652230E4ACC887256659D529A2";
    attribute INIT_30 of inst : label is "B49BA9A94C84260823483A51E947A51E947220949567CE69AB89B9A432666609";
    attribute INIT_31 of inst : label is "38438700C46DD11353264E3ADB6CCDF5D83A2F12CAC9596B6D6DAD9148E662D2";
    attribute INIT_32 of inst : label is "1ABC51955554A2312D5FBCFDEB8A5AA20E84CC4128DA368DA3996440C639A935";
    attribute INIT_33 of inst : label is "ECCBEABA29C19393F84089A4266094B5700004610CCCCCC91084C88888E51D75";
    attribute INIT_34 of inst : label is "A09864D04C326826093413049A098204230E5AE470E5AE5F95C461CB5F221CB5";
    attribute INIT_35 of inst : label is "58110112E39BBF2CDE0C92B58CA0A53902C3C3C3C3634D04C1268260934130C9";
    attribute INIT_36 of inst : label is "6181104088258110112E39BBF2CDE0C92A589F37E59BC1925481261811040882";
    attribute INIT_37 of inst : label is "114058C84BDC277ABC139AD6B214CF57500ADAEACC52D51DFB7E59BC19A54812";
    attribute INIT_38 of inst : label is "0000132B0040682643642183060C1252525252925B7281E14815104445111444";
    attribute INIT_39 of inst : label is "55151515155155151646444464675DDFD55777CCCCC88CCCCC072D32D2612000";
    attribute INIT_3A of inst : label is "555555555555500201F00408DAB7A1703A36ADE95C0E36CB236DB27FFFFD4952";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "543422A1A067B264C993264C993B76EDDBB76EDDBB76EDDA3E7986ECC373DCC1";
    attribute INIT_01 of inst : label is "D9938372E1930471E1C1C7869E5EC0F9B3D9ECF673399CF3FE7FCFF9BF37E6DC";
    attribute INIT_02 of inst : label is "C6798C17A1301E6FC3ACB441663A06838ECD839B31099E278739CCF7B3381CD1";
    attribute INIT_03 of inst : label is "E1058E2082C406203101882C41620A105880C406203105082CCA4633CC666798";
    attribute INIT_04 of inst : label is "16648461058E1058E1058E1058E0198C6318C6301058E1058E1058E1058E1058";
    attribute INIT_05 of inst : label is "9CC196C836C836C836C8A4CCA4DFEFF07FDFB5FD83BEA985A7D24D9325A4754C";
    attribute INIT_06 of inst : label is "48B6C88874222C82441266121D9196D88C320DB20D986CE1F1F2ABC53D215E95";
    attribute INIT_07 of inst : label is "CC1460A305182C420B39D9BA1CDCDDE8431248B6D86DB29A6124824D16DB0DB6";
    attribute INIT_08 of inst : label is "8414210580006C1660A3051828C1660A3059828C1660B3059828C1660A305182";
    attribute INIT_09 of inst : label is "0841621050841421050841621050841621058841421058841421050841421058";
    attribute INIT_0A of inst : label is "920B105080C41660B305982CC1460B39F88DF884162105084162105084162105";
    attribute INIT_0B of inst : label is "73E658F1ECF6D26C6DB77A0908425A20B04161082C2105871050808101042020";
    attribute INIT_0C of inst : label is "B1D91C38F0404082C40420A0925C76F63B33875E20B4E6E63B3C731E932DBCE5";
    attribute INIT_0D of inst : label is "1A012C496671080C4F1DE2CB1259BC42031807BC5EC636636B6636159EC49DB3";
    attribute INIT_0E of inst : label is "64841637873CBF321050CE3C38213DE62879B3CC8DE6FC4276F27993C4F1010F";
    attribute INIT_0F of inst : label is "EC6E1CE386641C3B06D1C38DC718A8F4A1F251CB3B3B3B3AAAF4A1AAB65A3C59";
    attribute INIT_10 of inst : label is "9999970684B6D555BECA9B8E36DDB8CB8E19665C7196DC0DB766B8BAE38DB1B6";
    attribute INIT_11 of inst : label is "D39B34E6CC7BD9A48B7A0F6D78C630D8C61B1E08253AFEDFCC1C06AAD9775655";
    attribute INIT_12 of inst : label is "8E38E38E38ECB0C8AC082CC14639AC01809C2727ADE9DBD3E7489BD64F557C36";
    attribute INIT_13 of inst : label is "944CFC5137BFDFE0FFBF85C684800B7A76F4F9D2426F5913D55F2426228138E3";
    attribute INIT_14 of inst : label is "08404202105A24034A3D030ED82CC1660B305A0406207880C79CC86161413120";
    attribute INIT_15 of inst : label is "943110F988B1324E50C3C79E18618618618618660C4604169242041420310188";
    attribute INIT_16 of inst : label is "D6DCD6DB1B2492856E16CC43510D84190980C1652A84190980C164426471D8C3";
    attribute INIT_17 of inst : label is "D813873CCE6679B99F27E4DAD6B7D6CD9D366F6C1B8F5BEB6CDCCAC74155F5DC";
    attribute INIT_18 of inst : label is "5BBDCCEB2DDEE67596EE733ACB77399D65BBDCCEB2DDEE67596EF7337B1EB2DF";
    attribute INIT_19 of inst : label is "56DB0DB10ECCF6CD33D9EDA7BAA02A0194436CDECDB6AADB556F99D7B77B99D6";
    attribute INIT_1A of inst : label is "55084202D95555550000B650040008408D99EE3716F6D8C81FDEDCD87A06D76C";
    attribute INIT_1B of inst : label is "0004004004655555555411015544180001A45555555410011555510600014555";
    attribute INIT_1C of inst : label is "0400000400000400000400000000400000000400000000400000000400400400";
    attribute INIT_1D of inst : label is "5555555555555555555555555555555555555555555555555555500000040000";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFBFFFE55555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFF000003FFFFFEFEFDFDFBFBF9FFFFFFFF807FFF8000007FFF800000007FFF";
    attribute INIT_22 of inst : label is "017FFFFFFBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFFFFFF";
    attribute INIT_23 of inst : label is "333373733338155554BBEBBE78E3AE3BE1FFFFFFFFFFFFE00000000101200021";
    attribute INIT_24 of inst : label is "1A24908C921512B29B69C4124024004904820B923068C1A1E8CC2EC639537773";
    attribute INIT_25 of inst : label is "05882C414748040C400008186D2492496D249249621045040824818883B22046";
    attribute INIT_26 of inst : label is "054E954DA210C6180CC04603301880840420B105882840620A105082C41620A1";
    attribute INIT_27 of inst : label is "8630CC303060B105B8C8C6B1884218C332C0C182C416E3231AC621086B0CC305";
    attribute INIT_28 of inst : label is "5882DCC631884218C330C0E182C416E6358C4210C61996070C1620B731AC6210";
    attribute INIT_29 of inst : label is "210C61996070C1620B7318C62108630CC303060B105B98C63108431866581830";
    attribute INIT_2A of inst : label is "986CC3461B30D1868C3661B30D986CC3461A30D1868C3661B6182C416E6318C4";
    attribute INIT_2B of inst : label is "48492124848484FC848480921240092124000B924CC3661A30D986CC3661B30D";
    attribute INIT_2C of inst : label is "C0D90B1716C88B3A1C2D9116787C0D90B1AF76C1F9FEFF07FDE0492124849212";
    attribute INIT_2D of inst : label is "C8B8E6645C39E831E2E643999170E7A0C78B991365E39C584443A1C2D9116787";
    attribute INIT_2E of inst : label is "D92E4B92E4F0F1EEECB873D863C5CEA73B22E1CF418F17321CCC8B873D063C5C";
    attribute INIT_2F of inst : label is "C8D972E46CB972365CF87363173F0D862E7E1F81C363173F0D98B9F87E11CE3D";
    attribute INIT_30 of inst : label is "A5E4084C42F9F8C79CB7C58E163858E163930C42C598309E0C2E46CDCB91B2E5";
    attribute INIT_31 of inst : label is "C79C7CFF1762070C1CC39860E491BA0A24C4C2EC30B6168290520A6474399A97";
    attribute INIT_32 of inst : label is "88B2EBA39E3319C2B066CC50759560B9F20933BEC721C8721C66197F3A564EC1";
    attribute INIT_33 of inst : label is "FB0F88B3CDDE5CEB473CEE4BD98C42C5960016A3C4446C338DEC444C46D72985";
    attribute INIT_34 of inst : label is "4C4B972625CB9312E5C98972E4C4B9FBB6315BF6C315BF7D0586C62B7E3662B7";
    attribute INIT_35 of inst : label is "7488C8882E109431E1E326C9B6B4791C5924242424DC72625EB9312F5C98972E";
    attribute INIT_36 of inst : label is "0DC88F244797488C8882E109431E3E366C9B64D2863C3C64DDFCA0DC88F24479";
    attribute INIT_37 of inst : label is "EBEB8733F5AA5D2F6188C4210B2B05C099E60534F0AB05C2452863C7C6CDDFCA";
    attribute INIT_38 of inst : label is "000001CC002F93D98918CE7EFDFBFD8D8D8D8C6DA48C305B16BFEABEBFEBEBEB";
    attribute INIT_39 of inst : label is "5050505050454050522222220205FD7FD77F5F44444004444540504504140000";
    attribute INIT_3A of inst : label is "55555555555553FDFE0FFBF72028881515C80A230565C9269C936DCD55356D5B";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "FC1227E010228912244891224480000000000000000000007E7802AC01534C03";
    attribute INIT_01 of inst : label is "48B90720C0862450A9414503940A40C89148A45229148A12A2544A89512A254C";
    attribute INIT_02 of inst : label is "863888568100B42F82A534C1263200111A44A28911088A228F7BC6C631291541";
    attribute INIT_03 of inst : label is "43048401824C126093049804C026093009804C026013049821880631C4426388";
    attribute INIT_04 of inst : label is "1264044304843048430484304846118C6318C630304843048430484304843048";
    attribute INIT_05 of inst : label is "92438018005812580058805880400000000137998A2640C72753499325A47215";
    attribute INIT_06 of inst : label is "1880580850E025800C002C0014B0824B8496049604B024C1D092AA4D24615230";
    attribute INIT_07 of inst : label is "4C106093041820C6093189E874D4D5A040000092492490492092412090002000";
    attribute INIT_08 of inst : label is "8C10630400006C106093049820C126083041820C106093041820C10609304982";
    attribute INIT_09 of inst : label is "98C12630418C12630418C10630498C10630418C12630498C10630418C1263049";
    attribute INIT_0A of inst : label is "96013001800C126083041820C1260831A885A88C12630498C10630418C106304";
    attribute INIT_0B of inst : label is "D7A6F850A4D249016DB629488421026080C10118202304053049820304046080";
    attribute INIT_0C of inst : label is "9149142844C029820C006080925452D2292285086080A6A6313C400A170035AF";
    attribute INIT_0D of inst : label is "1801380022D11800454CA2CE0008B446001002B45A5C12C1212C129C8A4C9496";
    attribute INIT_0E of inst : label is "6C8C023285349D3230088A142A3115AE3829B14C9CA6F44252D629B944C30025";
    attribute INIT_0F of inst : label is "8D2810D152640C1F06110205A28A0A61A8D051A9999999980061A0AA94CA34DB";
    attribute INIT_10 of inst : label is "41415506849255559C5A894512519A4B4549725A28924C049472A1A251449092";
    attribute INIT_11 of inst : label is "528914A2442B08AD8B6A0D242A42E0485C090A0208486A94440406AA53365515";
    attribute INIT_12 of inst : label is "082082082084B0D9A41800C1063190A8A1B06C62A5A94B52AD48094405157492";
    attribute INIT_13 of inst : label is "9C05D470168000000001854E8C80896A52D4AB52C0251301455D2C2C27812082";
    attribute INIT_14 of inst : label is "24C12609300A600A1A9F060CD820C1060830400C000029800299806141217000";
    attribute INIT_15 of inst : label is "342301F309A0360CC086829414514514514514520DC20C0008090C0260830418";
    attribute INIT_16 of inst : label is "8015801902249385243644C6001800301800834400003018008344C764D14887";
    attribute INIT_17 of inst : label is "580B873C995679655D07A0D6B5955A54B512AD2428854AAD2558C8850155D555";
    attribute INIT_18 of inst : label is "193504890C9A8244864D41224326A0912193104890C988244864C63142382257";
    attribute INIT_19 of inst : label is "06490C911A4652641948A48298002AAB04D2249ECC92AA4955260913326A0912";
    attribute INIT_1A of inst : label is "550802020155555500008050042100000008A623127248581FCC4C4830125324";
    attribute INIT_1B of inst : label is "40000000002555555554B1015544180004925555555410049555510600012555";
    attribute INIT_1C of inst : label is "0400000000000400400000400400400400400000400400400400400000000000";
    attribute INIT_1D of inst : label is "5555555555555555555555555555555555555555555555555555500000040040";
    attribute INIT_1E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_1F of inst : label is "0000000000000000055555555555555555555555555555555555555555555555";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "3333337773240AAAAA4000008204004000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "084000180070960209090092080010412492020000A002810081680220573333";
    attribute INIT_25 of inst : label is "001804C0264C0C0444080000000000000000000000400410180051184A8600C2";
    attribute INIT_26 of inst : label is "110C35008508001800C026003001824C106003009804C006083041824C126093";
    attribute INIT_27 of inst : label is "4210C00020601300B185009084210843000081804C02C61402421084290C0004";
    attribute INIT_28 of inst : label is "0980580090842108430000A1804C02C004842108421800050C02601600242108";
    attribute INIT_29 of inst : label is "108421800050C026016002421084210C00020601300B00121084210860001030";
    attribute INIT_2A of inst : label is "1820C126083049820C126093049820C126083041820C1260821804C02C004842";
    attribute INIT_2B of inst : label is "000000000000000000000000000000000000090004C106093041820C10608304";
    attribute INIT_2C of inst : label is "40901A13324889900C24911320240901A1E55201A20000000000000000000000";
    attribute INIT_2D of inst : label is "AA1054404898A46180C55151012262918603154104898CC8444900C249113202";
    attribute INIT_2E of inst : label is "DB0C4310C5A0A0A880913148C3018AA2A20244C5230C062A8A880913148C3018";
    attribute INIT_2F of inst : label is "A04862502431281218E041A6151C068C2A380E014146151C0530A8E038114415";
    attribute INIT_30 of inst : label is "A6240C84646022C75DB50D843610D84361112C4644B063B408250249894090C4";
    attribute INIT_31 of inst : label is "02B4747D3764130110020A208002885C01840280109212424849090440400A98";
    attribute INIT_32 of inst : label is "8890C3A68E610886A0C4CC50A1354191D60016A84210842108AA0B7C28C20A11";
    attribute INIT_33 of inst : label is "B007089104D8500A022C655B002C4644860012E3C44464418DEC444446526084";
    attribute INIT_34 of inst : label is "6C4312B621895B10C4AD886256C431EB9A6149D346149D3904828C293A14C293";
    attribute INIT_35 of inst : label is "2488C888461114208141324C93946918F120202020512B621895B10C4AD88625";
    attribute INIT_36 of inst : label is "24C88E244712488C888461114208341724C964E2841028264C38B24C88E24471";
    attribute INIT_37 of inst : label is "441606804188D42A2588C842116A21C289C6082041AA0C864E28410682E4C38B";
    attribute INIT_38 of inst : label is "000001F0002C13C019000862C58B1000000000249250300B0140451110444111";
    attribute INIT_39 of inst : label is "500550055015100552222222222557FF7555FF00000440000185999998580000";
    attribute INIT_3A of inst : label is "55555555555550000000003200218030948008610C058002580121D55555715C";
    attribute INIT_3B of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
