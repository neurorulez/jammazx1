-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "C52891615CA2B20280220142410082818250B27FFFFE00A0C1FEA7A3D3F3EDB5";
    attribute INIT_01 of inst : label is "DBA998E455D27FF936B9E826B56D0834B02845CAA43E3F5B40531AB5428B026A";
    attribute INIT_02 of inst : label is "2B1F640A80DDBCBB590C4223C60050C34002133F6199B676C00F5B2E7B44B008";
    attribute INIT_03 of inst : label is "5B21D17B84731534B27721F3DC381225E8FBA01B4D36DA1F9A13C1F66B9F9CDC";
    attribute INIT_04 of inst : label is "CF44EDD1897111BAA9AF43EC2D23E2AE6FBBE4C90D74C00000000924000374AD";
    attribute INIT_05 of inst : label is "479AB02DC35800002AF731C70D385214CD4F3EAABB1404440017EAEFA2AA4E33";
    attribute INIT_06 of inst : label is "030006692D2EFB8C54C9C530293355B6C000200024006000349A577CF97840E9";
    attribute INIT_07 of inst : label is "9883B4AB0C297959DBB12134BDC99F227C81F217C81F237000260000C0009800";
    attribute INIT_08 of inst : label is "B48000916FB718C1412082495FFECF3ECB6E4D97E4B477A65297EF4FE196A2F8";
    attribute INIT_09 of inst : label is "63E8B5B42D16891B03FA1320601B2475F782F7D09084C592339B9A5DC757FEDE";
    attribute INIT_0A of inst : label is "B20003DAA2757316018600040001F0040080036401F0FE4592838CD92C69A541";
    attribute INIT_0B of inst : label is "6C4D9E7532EF532E00403093108B820B1845F5F890508B5A982888D146CA7F51";
    attribute INIT_0C of inst : label is "BB0000819020072926D4D2A84A896B572514509570074424969DEDEDE8C90236";
    attribute INIT_0D of inst : label is "C33FFCD34D34D073CF3FFFCF3CFFFC6318C3FFF9A55CB7924407759E537D8C2D";
    attribute INIT_0E of inst : label is "D284D1117117A67A45A6D04814538C7BB84D1348052000026A300B288E0840E2";
    attribute INIT_0F of inst : label is "40031AD1A0894448201547BF84D19E12AA5FAA10B5D725068812C9C25ECDF1B4";
    attribute INIT_10 of inst : label is "318C3FFC0000000000008002A802A6448C89481D94919A1A1A81B4D29A644A15";
    attribute INIT_11 of inst : label is "A2457326150079545A296DF7283452DB922FFFCD34D34D073CF3FFFCF3CFFFC6";
    attribute INIT_12 of inst : label is "FEDF9FFC540401E105E482F3E0CAEB48A90D4A7E7C5929A4115425962D4140E1";
    attribute INIT_13 of inst : label is "47686EAA83972321A226324E808E18710988D5524CA13161108324EB39B6B3FB";
    attribute INIT_14 of inst : label is "1E1F9F7F7F7F10EEF625DDDB34CB134CB2909D425E86EAAE39723131D275025D";
    attribute INIT_15 of inst : label is "4034927F0348418BF05ABA7F7DA28DF7E050CC08B4CC46239180812488FE79BE";
    attribute INIT_16 of inst : label is "24A041111F148D0220980C80D3052D984526E90624AA35705B2E29481103CC50";
    attribute INIT_17 of inst : label is "84209392E2A28124915667BA4F8FE53A8B2BFCC7E95826B626B728FA5387F887";
    attribute INIT_18 of inst : label is "806AA290805691E667979FACC64CF7F09DCB9B964D553B8411C21874954404A2";
    attribute INIT_19 of inst : label is "9DF435233A8A8EB968BFC7438F74265E3A76F01C2C1580B0300204929F7CB148";
    attribute INIT_1A of inst : label is "A59227C79B0004464C99C81D110836A87BB84D10355541A6C45117450AAA3D98";
    attribute INIT_1B of inst : label is "13285988C220046E884A16120071C1A4E94C92F14524C4095622D54DA228262D";
    attribute INIT_1C of inst : label is "431B40088C14C93D0D5267510EDC40F0E09118B23CE941292033164C668C6486";
    attribute INIT_1D of inst : label is "7F699AC9D9266FB472D09688CF6635722722A3F28520817FA17F723CF3095949";
    attribute INIT_1E of inst : label is "47BBEEEECDDDDD767B8DDDDCFBBBBEE776FBB111F76226BB5AA4A4F7989FFD8B";
    attribute INIT_1F of inst : label is "AD56DE24B9644FAA3DD36FB586224ED95276CA098893B6549DB28260C300240B";
    attribute INIT_20 of inst : label is "EEB3FC6F1EEEB3FC675CFE37DD675CFE37DD6F1EEEB3FC6F1EEEB32766B6B1A5";
    attribute INIT_21 of inst : label is "70020B2088D915585C96CFC4B28E7DEA6CD55D77679BBAEAABAEE6D9DD756F1E";
    attribute INIT_22 of inst : label is "8F39E5DEDEDEDEDEDECF4F4F4F4F4F77B7B7A3D1E8F40804D6C409B732E65B00";
    attribute INIT_23 of inst : label is "64E94BA3335B49725F29720000000000000000000000019E7D6479E7D647E5B7";
    attribute INIT_24 of inst : label is "0000000000031E531C9242C9991737D8965B789CA176DB606DCCB9A5D02E4B52";
    attribute INIT_25 of inst : label is "52E4000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "C3E9D3A6B93A69D55A8548880A6648825CA401DF4FCDC4C99D51A966B292E4BE";
    attribute INIT_27 of inst : label is "4EC00351AAA4569302A4C4A915C620060B0373A60E9B471D55815CE01D45CE5E";
    attribute INIT_28 of inst : label is "BB3E0B35D626900D34D493064003581E01054604ED533B5022001A0A4C4BF329";
    attribute INIT_29 of inst : label is "D39366E4C669A4715A6870854B9E66F6574951781AF69C730F1103A5F18BB257";
    attribute INIT_2A of inst : label is "D34A1210AA4A2AD3B649FBD9A779E5E4CD3923A6294C1C3124AFCA694D33AECD";
    attribute INIT_2B of inst : label is "6FDFFFFFFD5B42BA94CB74CEC22777DDA8E1511EF9E79ECA674B9B267CB9FAE7";
    attribute INIT_2C of inst : label is "5D362F9ADD2E3BF686E259E648D6C7BF5971A7FCF5D33B0C545444C9A6CBB63B";
    attribute INIT_2D of inst : label is "D9D9C990AE16006405445B999CEC199CD9371999CF9BE199DB62BA9F5A9BBF0A";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC00C55F001EA400EAA807554E0C01041D1919999";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "E80183E5BCF9736592B0486D6C964993D004007FFFF8592DCAFBCD6603E38D93";
    attribute INIT_01 of inst : label is "86C08117676DA8AA49802B229222EB12A6E7EE3FE16A92E52C9FBC4729633010";
    attribute INIT_02 of inst : label is "F0D03C030045438A80E512D7EF9A671F8D3C25610D99D66726CD2B6C6ED00191";
    attribute INIT_03 of inst : label is "D27DF84B1EA4D23FE4D533C4D183387F1580AA81F69960BF4369DD03CC14AD20";
    attribute INIT_04 of inst : label is "FF2DFD8CAE35DC9FF3D21A093111F790A023019B440500000092400000001511";
    attribute INIT_05 of inst : label is "B40CF01EC5A8000006EF25C82B41712496C1EEEEFAFAEEBFFEFD01054518C417";
    attribute INIT_06 of inst : label is "3F000562369EDC0CCE9A03B0080AF6DB4000A001A800A000F10D0F7C49A1C170";
    attribute INIT_07 of inst : label is "AED85198ED93312EFBD600983D813E01F803E03F80FE02F000160003C001D800";
    attribute INIT_08 of inst : label is "42124996104D39CA64B64800300010202B808925E99B188DC485957FE5BDF7F9";
    attribute INIT_09 of inst : label is "87B19292B9DEE5377A62F139642E7607C9B61B1780E8CF3B00031BFFE02804A6";
    attribute INIT_0A of inst : label is "00492600287F75A9C1F80081DFFE09F9FF0E0381FE00008016E85F8C91D201D5";
    attribute INIT_0B of inst : label is "33302015D9815D99911FEA0EBD6671407EB33E66C91B64032BB3A21A1520A005";
    attribute INIT_0C of inst : label is "01000024C2FED0F28020046DBFC4806556468A67841387FF486BAFEFE27FC8A0";
    attribute INIT_0D of inst : label is "6AFFFCD34D34D073CF3FFFCF3CCF3C630800F3C219E124F92D104D727C890B49";
    attribute INIT_0E of inst : label is "055C16A9EA9F1AACC80A0EB138E529484221A4332EC615E71E865C23712919DF";
    attribute INIT_0F of inst : label is "1EDB39442ED5EBC75C8B9484221A3E47BBE61B6806A55610D3345CD1241F7680";
    attribute INIT_10 of inst : label is "000000000000000000008008C020521AB4B8C172592C975757AC000400B1A772";
    attribute INIT_11 of inst : label is "308BC972CB24D06FB6C248255F6D849018800000000000000000000000000000";
    attribute INIT_12 of inst : label is "9868CE03965FB46C302F0817AF9BAA1115BD7E42F5F36F15A236DF4801D58BE8";
    attribute INIT_13 of inst : label is "B49A8914B240446A2D6D5F0937AA8B335C1536B0C468824BBAD7729AE29B4112";
    attribute INIT_14 of inst : label is "5757B5ADADADA602D1480434411AC015503448EE11A8914924044B6AF848AE10";
    attribute INIT_15 of inst : label is "BF02CCE66E7FBFD4DB03C788A02A05D7F558B5A3DA97AAD5EA991EBED1691297";
    attribute INIT_16 of inst : label is "F7D531ECC04354BDC30B4476FAEF91E8F3902BA221D63A9A809078C25EC822CA";
    attribute INIT_17 of inst : label is "A372725EE69ACB85C385970607B7FDAA42C2045730C0DADA49C42423C81A1651";
    attribute INIT_18 of inst : label is "48EE9ADAD898EA808164ACDB54021004415662ACF135C037DA77367E526E1190";
    attribute INIT_19 of inst : label is "43DBB24A833110F785405C0EA8091146F8A7F59D40A01402C96105C5E40472C5";
    attribute INIT_1A of inst : label is "6E00482FD4CD977BC18A8B622293DB7D484221A83D25E1F823AEAA3AE67CA04C";
    attribute INIT_1B of inst : label is "887F652D4184D6D01A235926007E006DA1EA7F93F7BEB6B6B3F91AC755427273";
    attribute INIT_1C of inst : label is "1B02196922134A71EA8F49826758DF4491C652CB4AD20C6A66A8006140C09154";
    attribute INIT_1D of inst : label is "9DB36C92524DB6DAA16B27EF1501C208408C441DD88809F77688DCA343D29212";
    attribute INIT_1E of inst : label is "9AC5BEAFB820A009D43D7DF54541415A29450EBE8A1D780EF7F7491083258C05";
    attribute INIT_1F of inst : label is "1BF53D41BA9884444E221362A09B972CD5B924162CE55B656ACB0589649A5A8C";
    attribute INIT_20 of inst : label is "BDCE338F7FDFDEB5A73DEF5A96A73DCF5A94A73DEF5A96A73DCF5A38900C4278";
    attribute INIT_21 of inst : label is "25966210E6533733034D9273A45427DCB4000000000000000104445155554E77";
    attribute INIT_22 of inst : label is "3472CB101010101010282828282828141414160B058099F05CB6B44908193659";
    attribute INIT_23 of inst : label is "1A12DC454C04C40D32540C000000000000000000000000BA358F0BA358F55B6D";
    attribute INIT_24 of inst : label is "000000000001ACB7341452D58E3D67F64DB6D329C6020033124206513981A628";
    attribute INIT_25 of inst : label is "A818000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "A2157A55E3C002C0005B757DDF0D9485D900935855D5B834A222DB980D881A64";
    attribute INIT_27 of inst : label is "C309978A15BAB98266F01B6EABA4B16F10019A55902184CC006A00AF32100901";
    attribute INIT_28 of inst : label is "40415AD009806EBB001940458997957570F771B2B0F02C36644CB9AB8A02827A";
    attribute INIT_29 of inst : label is "30C03BB01F981906E002352892E1CD3380AEBEFCC7F9EEFA1F72C26203600F80";
    attribute INIT_2A of inst : label is "304688C9B96EF12142DA0E93094A1D2A00C06A18DC01134ECBAAE002004C0077";
    attribute INIT_2B of inst : label is "BF1FFFFFF84D264F660CC70C5669FA7E998563982282281C8090044001000480";
    attribute INIT_2C of inst : label is "F2D27565965455215CBCD2E0540A4EFEB25E0381F35C31589989889EA8B6CB2C";
    attribute INIT_2D of inst : label is "999989D1E4222C440AE852AE528C9A52A1CCD5A528144D5A00064F66F7601F1C";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC00014D1C1C042A85E9542F4F5D0305191B1D9D9";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "081800E13C9372458080804949200081D11600BFFFF811D543F94D7719E99B81";
    attribute INIT_01 of inst : label is "134094866646A4AA59080A0014414A102245280EBAD508A408FDBC7708600830";
    attribute INIT_02 of inst : label is "A5D2FC0C0049D793A8D01206A41275CA49B635D96D112454C669206849420111";
    attribute INIT_03 of inst : label is "C58848A8920A950668DB27D4D5063878092A0FA0010410BF92615D2CC50AB58C";
    attribute INIT_04 of inst : label is "A00DF0542D15A48553F65A2D30FFFD8228A22A1241445200000000000000442C";
    attribute INIT_05 of inst : label is "2F54301A8A880000587421E49F24FE4845CD7BEBEBBEFAEFFFFEFFBEC1008615";
    attribute INIT_06 of inst : label is "6280084CB228324E5DB9276809F1C5B6C000640028006001265594187824C0F9";
    attribute INIT_07 of inst : label is "9445C1BAEF31121D9FB5C5BF0C3258CB630D8C463198C4680065000DA0023400";
    attribute INIT_08 of inst : label is "A98000945B350840010482001FF2D3B2EFAAA5B7EF8E2A0D8E85A47FC5BCB2F9";
    attribute INIT_09 of inst : label is "2B90A49481C0E11CB862A01E438D4611CA340B15086286A34A4231B2200854C6";
    attribute INIT_0A of inst : label is "000003F57F882919C7E60085DFFF0085FF8E3C85FFF00084A5280DCE205BA054";
    attribute INIT_0B of inst : label is "3B43EF7FDA1FFDA1FE0854855FE820B76FF43E676E1248400B82C2005402A015";
    attribute INIT_0C of inst : label is "FF00003884308010A06400A92AA10801708002850FE32F7E10801014547F42A0";
    attribute INIT_0D of inst : label is "C280000000000000000000000000000000000003A1559AB847E04504C3E5DA66";
    attribute INIT_0E of inst : label is "24069049E49FBC96DC9E10F92CB4A529720547400F07951483001E4201BE11FD";
    attribute INIT_0F of inst : label is "02425064A125FC0DE19AD29520501E43AFE62A4E80E170D0021458D0440D5185";
    attribute INIT_10 of inst : label is "000000000000000000000A0B0FE0900486AC821490090C4C4D68140080392914";
    attribute INIT_11 of inst : label is "00E1036281006F85163B37D80A2C766F78A00000000000000000000000000000";
    attribute INIT_12 of inst : label is "FFF68CA4D4842068D42E7A172AAF3F1C252D4B62E515FB9538549511A05410E8";
    attribute INIT_13 of inst : label is "35162A26AA90F0D82839172A052A8A32D04054208668084150A442820F24B74B";
    attribute INIT_14 of inst : label is "4C4D6C848484B444336884F6685A149511240923E960A26AA90F01C8B95163E9";
    attribute INIT_15 of inst : label is "904404F6786BAA8ABD42A80A80222DD5D755A52282A74AADD239153486FFEDAC";
    attribute INIT_16 of inst : label is "86837F868E840408BC4EA404114AA12C558482E8E184EAD486A030837871C824";
    attribute INIT_17 of inst : label is "E37C719EA2AAB211C9A51E5407BFFD229288DAD6118CFEFE6F55A977026B7C50";
    attribute INIT_18 of inst : label is "4862AA9488CEBA53A1B6F66FD20452E409DBB3B7D9552AA451EB7F09506F9D45";
    attribute INIT_19 of inst : label is "0A6D2629119998DAE56DD2C92427421FA1E4BDF540A09612F17D7D0432CC3482";
    attribute INIT_1A of inst : label is "6F5A6E16169C937D850A6A3337FB6EA929320543F9455F9006B0497B06F690B5";
    attribute INIT_1B of inst : label is "817861087504F47852021863E07FF84925A852065534A430174A90842802487A";
    attribute INIT_1C of inst : label is "1C8C006833B3787DCE0A404E6FD69F478D0210C20F73096A2695E3457291D392";
    attribute INIT_1D of inst : label is "D6F9B7FB7F66DB7E93B3F6A7D23DE337667777577755DE00088AF69929529C1C";
    attribute INIT_1E of inst : label is "CFDD54057FFF55FFEABAA8AB7FFEAFFBD57FA016FF402BF79D57FDDEFBF56BAE";
    attribute INIT_1F of inst : label is "5EAF0741BE1CFB466B3219F320DBFDFE9FEFB6BF3CFFEFF7FF6FAFCD74DAFEA7";
    attribute INIT_20 of inst : label is "A4231A4025210A520A33A4A33A4827218A720A33E6B3BE692F639A51CFF8E20C";
    attribute INIT_21 of inst : label is "75169B9A44D14334DFBBFF0F7F9BDA77DCC00000000000000104445155554231";
    attribute INIT_22 of inst : label is "B073EE0D040D040D040682020682068341034080D02211068EA45B3736FCEF51";
    attribute INIT_23 of inst : label is "7DD2DE676FFC837EEF7B7FDDDDDDDDDDDDDDDDDDDDDDDCAA6D688AA6D68C0EFB";
    attribute INIT_24 of inst : label is "EEEEEEEEEEED3EE526D752595FAC77FE52EFBB41E3E08214CDCDBF6DAA6FDD76";
    attribute INIT_25 of inst : label is "F6FEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE";
    attribute INIT_26 of inst : label is "3A250AB482C292CA8551621DDF14A4AC1AA001510D958CFBB8335BDFFD06FDDE";
    attribute INIT_27 of inst : label is "870807E840B1190A0234022C42B4B20FD030CAB5D0A50D4CA84B42AA34142941";
    attribute INIT_28 of inst : label is "F7C6A83436A1950A141050F44807C2157DD069DEB160AC52838031E3CE9BEA72";
    attribute INIT_29 of inst : label is "21D0FBB40790ED01F21A355DA23145E3104E5D7CEBFAFEB81F34FA4198A87710";
    attribute INIT_2A of inst : label is "216680008A0A942360924C8A092B5CAC42E04A5C3C41D04690F8E200524FA1F7";
    attribute INIT_2B of inst : label is "3F4AAAAAAF9E87F7F9E72182172CAE2B9DC061861861A692232A8CA23288CE23";
    attribute INIT_2C of inst : label is "FFF45DB7FFFB6EFFDBFF1B8659DECBFEFFFF2035F4C60858DDDCCCDB2CFF7377";
    attribute INIT_2D of inst : label is "919189911F56446413E91BBB4A68534A5967C934A5966C935F4BF7F7BFF39F16";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC00455F1C1C0400C0140600AEDA01021B9B99191";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "808D80151E11385414A00001000920D8C010013FFFFC11D7C8FE64D6D8F8F2A1";
    attribute INIT_01 of inst : label is "D102D2B7FFC6255324C809A106C3131045548418D150323508F519632046A029";
    attribute INIT_02 of inst : label is "3110CC000098D431A802AAE37700D9B380669339718BF72F339ED89EECE95DDD";
    attribute INIT_03 of inst : label is "114C223338A696831043CDC6D152AFCA4B3380A4934D3410BD3A110CF58B31AA";
    attribute INIT_04 of inst : label is "9F042C431EC3CE919990D5E5E977F48298842100131800000000000000020436";
    attribute INIT_05 of inst : label is "4585301B80C80000206459828B147001044405400145150554114055611A0519";
    attribute INIT_06 of inst : label is "220000641E08B1484CF8A3201880CC9240006000600128003204045C197440E0";
    attribute INIT_07 of inst : label is "55497413915316F76B34028B4D005C057011C007009C0060008C001080001000";
    attribute INIT_08 of inst : label is "5BC924B3EFE4358804106A20150E4E1E476EAEBBEC82ABA0D905390BF312AAF4";
    attribute INIT_09 of inst : label is "D3C8918203CE2528C8C67958640A9321E40A2633C1634D4994A7CC10220850AE";
    attribute INIT_0A of inst : label is "0124935FFF55772C0000000000000000000000000000000133208D88B1498911";
    attribute INIT_0B of inst : label is "280596BF502FF5036C0910A331C0803378E06C45A4006C128338809044022011";
    attribute INIT_0C of inst : label is "D7FFFF90801180B0A04400A02A3582506704120DFB022CEC5809A129A8590A20";
    attribute INIT_0D of inst : label is "5C400000000000000000000000000000000000398367FFB044C28A769DF7D1FF";
    attribute INIT_0E of inst : label is "0014234B74B7EC72A54FE359ACF3DE73DC077312461F9A3A2A548C96C4D4B7FF";
    attribute INIT_0F of inst : label is "014F49EAC70584E62524E73FC0535F2A1EC4280A2550674480000041640FD6D5";
    attribute INIT_10 of inst : label is "000000000000000000000208004210071EB8601488094EDA9A88140080202154";
    attribute INIT_11 of inst : label is "A04862000192540056DFFEA800ADBFFDB0080000000000000000000000000000";
    attribute INIT_12 of inst : label is "2C97882482046020616C20B62A1E3E0924096BC6C5436B1D925015D88911C0A0";
    attribute INIT_13 of inst : label is "21C88385B8C52522EE265603AC00003988905CD966B012C723B22314EFB7DF6F";
    attribute INIT_14 of inst : label is "9EDAA8FCF8FCB04423608DA7614454010B580C2ADC8A38438C525132B01C2ADC";
    attribute INIT_15 of inst : label is "805006523A0C51932616CDDD5D75D8AA8ACD1F50C2BD5FA7535DF1A69A5B6D2A";
    attribute INIT_16 of inst : label is "B0E1362A03012C625854681A0738001D5706A06AC286C71652032CE122204D20";
    attribute INIT_17 of inst : label is "0130EA2DC7B2FD10A9A0CC13379C2882C6E8CFC01499FCFE6C512C701A6D1404";
    attribute INIT_18 of inst : label is "60A5B2F69E6714E6E0B2B265A78467F80CD9B9B35965AA88938A238562A748F5";
    attribute INIT_19 of inst : label is "0C25625358888CC8F064E67BCF7C02DA93FFB8F600180100703E788A7FFA5362";
    attribute INIT_1A of inst : label is "23F6BC169FAAEAACE2C5C91116190CEE73FC0573D975BEC030130F4129073DF0";
    attribute INIT_1B of inst : label is "0169E629B414BCCE8C1279A61F800724492808C6318714F3131013E40401A11F";
    attribute INIT_1C of inst : label is "1828126399E7B22ADE238D426E96E55B18AA53CA67317B565631FE83A71265A7";
    attribute INIT_1D of inst : label is "E25ADE4F89EB792F7DBDB6D5CEB97112233223F60A0228A0A880773878480A1A";
    attribute INIT_1E of inst : label is "D64F54056800000140280201D555555EABD50ABFAA157ED58E47BD6311BA3136";
    attribute INIT_1F of inst : label is "062222688214494ABD56AEB5DE4658BA72C591DB99962ECCB16676E4D2476DD6";
    attribute INIT_20 of inst : label is "290A4290A0280202840521485214812040120024290A4290A028021066DC2265";
    attribute INIT_21 of inst : label is "9850499677A23B365E9A596612A64A265A400000000000000104445155554024";
    attribute INIT_22 of inst : label is "9A2527AD642D642D6456B212369236AB590B4C86D3217F2DA714899292F66985";
    attribute INIT_23 of inst : label is "348046AB2B6CE17A69197BF4A1F4A1F4A1F4A1F4A1F4A134696D134696D4A698";
    attribute INIT_24 of inst : label is "053AF9053AFA5276B872AF4E9919E0996069898C61618E0264A4BD64A12F4D92";
    attribute INIT_25 of inst : label is "32F5053AF9053AF9053AF9053AFBAF9053AF9053AF9053AF9051053AF9053AF9";
    attribute INIT_26 of inst : label is "10852640308280800A456ACCC296244DB38A49CE2AEAC469925508D6DCC2F4D2";
    attribute INIT_27 of inst : label is "628D22A292B574C04A9152AD5C803A45414A6640608014A800091402B2014014";
    attribute INIT_28 of inst : label is "BB14AAA15B0AD929814045215D22925F7C866A6C29590A56DEA91B95BEBF3030";
    attribute INIT_29 of inst : label is "38856221561C2654C0A8B008964441E2855B557E6AFAB282006730F3DFC2BA85";
    attribute INIT_2A of inst : label is "18EB0124CCB3191336E81743043340CD42150242981482461050C20050134AC4";
    attribute INIT_2B of inst : label is "80D555555579B494B97E31EC5B4F34CD75B1B99F3CF3CF0B333CCCF333CCCB33";
    attribute INIT_2C of inst : label is "69F4BADF496EBB95B76789EABD5695BDEBB3281888C7B16C555446530E7DB2DB";
    attribute INIT_2D of inst : label is "898989C04164ACC422E9099B9CC6EBDECE73DFB9CCE739EBFB7094B98CB9AFC6";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC05A82102A2A46B3FFF59FFEFDFAEAFB81A18989";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "289D020482510B4C528940B524924D5BC06410BFFFF855A908F96C444DEDBB8A";
    attribute INIT_01 of inst : label is "921CF38627441CFE6DC4111082A2419506640000D40442A12ADD834A256CB13B";
    attribute INIT_02 of inst : label is "311C33FFFF79E4F3C9008CDE9DAFE52ED7F5ED63CD5464419D43A64317F18931";
    attribute INIT_03 of inst : label is "000EE00D3830A3D904001CFD1F762CCAC709D83CB2CB2C4098AF71C3156BB58D";
    attribute INIT_04 of inst : label is "1A402996EFBDCB855B95B96C065410B20C89205241004000000000000001289E";
    attribute INIT_05 of inst : label is "9C40703C0D38000044E9056A7853CE6CFE80D45110411004444105110DAF898A";
    attribute INIT_06 of inst : label is "1FC00FE08092DD2683C290FDF8431FFFC000FC07FC03F803F041096C01B34148";
    attribute INIT_07 of inst : label is "254A5F7B437770110852D600143328CCA30E8C3A3068C7BC007F800FF001FE00";
    attribute INIT_08 of inst : label is "405FED628255296A49B6EC28A556C616C426D5340CA1A2FAF41C31A00A01CF02";
    attribute INIT_09 of inst : label is "24132495A5D22A79D84C4C9E078543120A200A626E620AA98C60400229AA5A04";
    attribute INIT_0A of inst : label is "117FB402AAA8882000000000000000000000000000000000E561159940922070";
    attribute INIT_0B of inst : label is "2742685F2A11F2A192192102176800143BB42DCE4A2D50409F0142049444A225";
    attribute INIT_0C of inst : label is "4D00002896D380D2C9881C56AC020813E0810A898CE27CEDA0889010145B8CA2";
    attribute INIT_0D of inst : label is "08C0000000000000000000000000000000000002227268B31B2018720C1B439A";
    attribute INIT_0E of inst : label is "1C4A026B06B01656AF6D824DAEB0842F88466443631E7C200506C6DA412A354A";
    attribute INIT_0F of inst : label is "0B48C36387168CBC66ECC2F88462E0BC3FCC95AC81D3E0B02170488084922208";
    attribute INIT_10 of inst : label is "000000000000000000002203F000580C17192366C92828080812181D03A4A520";
    attribute INIT_11 of inst : label is "08A0492302BFABFEA874D2577D50E9A452A00000000000000000000000000000";
    attribute INIT_12 of inst : label is "936899A682D8E040942CDA166E3E7E5416D22DCACDC77B38A82B562120701B40";
    attribute INIT_13 of inst : label is "A192231710D0504844D91663172A0808004168A9A3C108B223300030E6924CB6";
    attribute INIT_14 of inst : label is "08080C8480809947366083B76050E0774F0080A5212031630D0506C8B318A520";
    attribute INIT_15 of inst : label is "9286DC343A0FEE3C8944E228AA2A00280A1C350CDB353A9D4AB13487147FFF08";
    attribute INIT_16 of inst : label is "30CD38A4ACA52D4AA57CBCA3764CA80D933277532A17368654A9D4224AD5A145";
    attribute INIT_17 of inst : label is "881D65BC8F1448119AA194D1B850098444D00900C2BAFCFC6C11447800FB4547";
    attribute INIT_18 of inst : label is "518F14671EED305EE5F7376F82045FD0899BB3371E38AAACA22DF6016682501A";
    attribute INIT_19 of inst : label is "8C654AC1119999D8D66D82E105F822C467D1B1960EEB5F2A4F2180026DA2C623";
    attribute INIT_1A of inst : label is "0712FE9A2EAAA23DB36171333A5D2CCC2FE846672A28F9421A322CA3376617C0";
    attribute INIT_1B of inst : label is "1121AC71491798BB80546BAE000000493AAC008601863896274A2224800303BA";
    attribute INIT_1C of inst : label is "9CAC1BC3226F481EF20309E040EC214C940AE35C4E73F180D6111E052E3AEDC2";
    attribute INIT_1D of inst : label is "C65D96CB19765B2E19B1BCC78B65E37EEE7EEFC6228820820A08E6182D668C3C";
    attribute INIT_1E of inst : label is "CC4F015038000001C0380001C000000E01C0554380AA81B3BD4724C635B46346";
    attribute INIT_1F of inst : label is "1E2626E1868FFF0EEB3C99836C94D9BCE6CDA71B2D366F79B36BC6C964946FC6";
    attribute INIT_20 of inst : label is "8C2308C2308C2308D2B08C2308C2308C2308D6918461184611846151CDB8FA5F";
    attribute INIT_21 of inst : label is "B9585F9654863BA6F23CDB6E320BFA6769C000000000000001044451555552B0";
    attribute INIT_22 of inst : label is "F867EE2129606820283034141034B0880A18452201435734C4389B367790F397";
    attribute INIT_23 of inst : label is "F1D20EEEE6DC33C8F39BC9555400000001555555540000A10EC06A11E4020F39";
    attribute INIT_24 of inst : label is "FA9501503FA97FE4828E0838F10B40124AF39DA0BB488282CD9DE40FA1791EB6";
    attribute INIT_25 of inst : label is "B791503FABFA9501503FABFA9503FABFA9501503FABFA9501503FA9501503FAB";
    attribute INIT_26 of inst : label is "2A367CF422540E9AA50266790658B675E32AFE25B08C0DE37A7745CDBC6791E7";
    attribute INIT_27 of inst : label is "A24DB0CA5133334A6CF50A4CCEB4B92190849CF5B5029999AA7A52B2A6352951";
    attribute INIT_28 of inst : label is "4449F11524A905B0851954540DB0D365B2C6A892A588A962F12D87DDD2B68A72";
    attribute INIT_29 of inst : label is "A854A6551A545942CA92B468BCC98D2654A2A681540D28A020A64A10252A4654";
    attribute INIT_2A of inst : label is "A8BC104911E45528FC2140E011BB86ED4C07DB805951535ADBAA4C0E81CC294C";
    attribute INIT_2B of inst : label is "800AAAAAA8809DB494D461B8500CA82A51142B8186186185B296CA5BA96E85B2";
    attribute INIT_2C of inst : label is "196C1996D96208B1D2E699471CCD8300DB7343D009C6E140CCCCCCD30CDB42B4";
    attribute INIT_2D of inst : label is "898999882378C96440001B134A4293085867883085866883001DB4939C93C026";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFE000001800006000000000008000000189E98D8D";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "603D9294A25549D5539359B5B6DB6DDAC274023FFFFAD5FB5BFE82666BEB9FAB";
    attribute INIT_01 of inst : label is "80031CDAEF6406AAD903014D328A797927552084551579436AFB860B6D7DB04F";
    attribute INIT_02 of inst : label is "9203300FC045588AB21A58CC00F034487891343C2E66199866532952910E3375";
    attribute INIT_03 of inst : label is "584D430A50C4A2A422007484011AED48654CA80208208270FEA9D033235CBD1A";
    attribute INIT_04 of inst : label is "3A6E1D5C2D199BDAA0CD1F08551010C4DB364D5B5B6DC000000004100821491C";
    attribute INIT_05 of inst : label is "040010080008000000200100080040000C00105414514005050151414DB8952E";
    attribute INIT_06 of inst : label is "160002C00000100001800021C8000C9240007C073C033803200000080020C040";
    attribute INIT_07 of inst : label is "0DCA511E59538A1518300000040018002004801200480120002C00058000B000";
    attribute INIT_08 of inst : label is "6632D9A28213BDE924926E03BE92D372DE92A92409C0E488C5A615481E88D907";
    attribute INIT_09 of inst : label is "B433B6D73BDD6C7B014042BE87977E5A08A85A021AE50BBF294841FFE5A9B406";
    attribute INIT_0A of inst : label is "26CB66A280A02B360000000000000000000000000000000096B21C8844DBA498";
    attribute INIT_0B of inst : label is "E14BAEF50A5F50A4DE49138132A9164F3954A4436E6D51490211CE49D49EA075";
    attribute INIT_0C of inst : label is "0100003982729252E03D0276A65A292042924E9087E62424269ABAB234C80E84";
    attribute INIT_0D of inst : label is "4A40000000000000000000000000000000000003A42024900FE4CB214A402909";
    attribute INIT_0E of inst : label is "024E526B86A841018108A20168A0000800986749272F9030C7224E5649FE7728";
    attribute INIT_0F of inst : label is "48484148A414808404248082098220ED1A441DAE920042D2496183469C18136C";
    attribute INIT_10 of inst : label is "000000000000000000003C0BFFC0504D941819364B2ED08085116D23A060A532";
    attribute INIT_11 of inst : label is "13E4900C1365D51542404828AA84809074A40000000000000000000000000000";
    attribute INIT_12 of inst : label is "08208892B24CA4B3D4B46A52309A2A1C96DA264246132908B93B5323A49889A3";
    attribute INIT_13 of inst : label is "AD9A5B151652F2E9447D321917AD14F0A14930820A6269366631059640482000";
    attribute INIT_14 of inst : label is "80851A82868698DAD45314140782700D294138A691A5B15B652F23E990C8A690";
    attribute INIT_15 of inst : label is "4926DC0EB92504904D484575DD57D7FF5FDA94424A142A150E575092107DB6D0";
    attribute INIT_16 of inst : label is "92453E96949496247CC8651A9128A40903182A06EC96E2221EA4E11B69F280B2";
    attribute INIT_17 of inst : label is "843DE9AD07147C2984949C48587818B45858F78008CADDDD4C3645B00F88E504";
    attribute INIT_18 of inst : label is "4CA5144612EC340209A6A64D601D9001315AB2B55A28B924A3AEF2F1C3079A57";
    attribute INIT_19 of inst : label is "30412A706111115098492090C1000D6E07D806E38342684D7CBD7A312404520B";
    attribute INIT_1A of inst : label is "72364A5F24000AA81834312222110AEC08209868FA28C7846002280021240400";
    attribute INIT_1B of inst : label is "267125217D6DB1CA209849260000006DA2E1892F2C9290B2362A420C124A8612";
    attribute INIT_1C of inst : label is "DF90C9D933AB7B3BD64948C074D5002F9C3242484B52739C4E06F2D971B02D20";
    attribute INIT_1D of inst : label is "94110482504412090525245520D54224444444B557DFD5D7F5DFB4040B465050";
    attribute INIT_1E of inst : label is "8A7355555AAAAAAAD55AAAAAD5555556AAD55001AAA0012AD6AF4894A5254A54";
    attribute INIT_1F of inst : label is "2B5434DC064A92A44A2891425CD0102E808135D23C040BE0204F748D74D54854";
    attribute INIT_20 of inst : label is "AD2B4AD2B4AD2B4AC234AD2B4AD2B4AD2B4AC234AD2B4AD2B4AD2B8C89224A4A";
    attribute INIT_21 of inst : label is "A27C52D345B222A28124922920A0974496800000000000000104445155554234";
    attribute INIT_22 of inst : label is "15025639B1B9B1F8F0BCF8D85C58DCDE3C3E7A3D9E8E7D3DAA909224A4089205";
    attribute INIT_23 of inst : label is "494AE44444931A04921204AAAAAAAAAAABFFFFFFFFFFFEABAD500ABAD501892D";
    attribute INIT_24 of inst : label is "AAAAAAAA80012465455AD26BC9C920285892D15D42CD9652892902C9294092A4";
    attribute INIT_25 of inst : label is "240AAA8000000000002AAAAAAAA8000000000002AAAAAAAAAAA8000000002AAA";
    attribute INIT_26 of inst : label is "BB1428564BCE018995D3665FD60C97FCA1AD97412E8388922922588922340924";
    attribute INIT_27 of inst : label is "1E0DB2EB49B3303B6EF58A6CCB96BB65D278C856D381D088993B5AD2A2D5AD59";
    attribute INIT_28 of inst : label is "77FA0ACDBCADE5BC759956F78DB2DB777C872CDAE0C6B832DD8D95C7D6C00B69";
    attribute INIT_29 of inst : label is "4756EA959EA3FD62D2DAE62A9450CDE216262D83ED097CF330267B0F662B7616";
    attribute INIT_2A of inst : label is "C2A6276D557554AD310028D4734A6528932C68645A59D9CE49F9D613C0276DD5";
    attribute INIT_2B of inst : label is "D07FFFFFFF47FD2D288C4D29C1AB595659946B8CF3CF3CC8EDE3B58EDE397CE5";
    attribute INIT_2C of inst : label is "D04951049041802530B512D4D2892A40925AE0240974A700C88888DAE8D2D5AD";
    attribute INIT_2D of inst : label is "8D8D8D838A80F18482ED93AA0851A20853448220853448224D0D2D22D523A074";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFDF8EE3F62A2B580DB6C06DB69D3A3A3B8DAD8F8F";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "208C089223004C01C849269092492449AD10487FFFFF23A9E5FF46E2C9F9C9B8";
    attribute INIT_01 of inst : label is "8136B53223626DA9009E74F8C87104D9D264BE17814078A591D5166394249129";
    attribute INIT_02 of inst : label is "E904CC0000C9E493C8109D2F62B348D159A3036711998666E28F588E79529711";
    attribute INIT_03 of inst : label is "2164443821160980004397D3C4344CA9D278800C61871DA00139404CE1CAB5C8";
    attribute INIT_04 of inst : label is "35955EE4151699D5D1C509AC1C3210DB04C131C0208240000000048009038248";
    attribute INIT_05 of inst : label is "F3FFEFE7FFF7FFFFFF9FFCFFE7FF3FFFFBFF8055405400055001540170C8459C";
    attribute INIT_06 of inst : label is "EDFFFDBFFFFFEFFFFF7FFFDE37FFFB6DBFFF83F883FC87FC9FFFFFF7FF9F3FBF";
    attribute INIT_07 of inst : label is "98E130888419A16667CFFFFFFBFFE7FF9FFA7FE9FFA7FE9FFFDBFFFB7FFF6FFF";
    attribute INIT_08 of inst : label is "21ED2608492D8C64924922248FFACA1AC6E225B60CC13B84480DC9140F2F9C03";
    attribute INIT_09 of inst : label is "506C58D8C0E472910CC539787040932823073629C1F0E04194A73D003387F017";
    attribute INIT_0A of inst : label is "49B498AAAA2A2394000000000000000000000000000000019224C4882A005242";
    attribute INIT_0B of inst : label is "A0A4101505215052012CB88B9114CD00B88A6440012408A4084C212445222911";
    attribute INIT_0C of inst : label is "930000848DA8410823254112191154810949214B78122424114020202A49620D";
    attribute INIT_0D of inst : label is "650000000000000000000000000000000000003852CCB3906012208DA364B42C";
    attribute INIT_0E of inst : label is "412129C49C480CB3660F08DFEEBDEF799826D0A6CA96598FB09D940124090260";
    attribute INIT_0F of inst : label is "23677CC050C2A615328AF799826981F9CA44448148810909249A6EAC54429954";
    attribute INIT_10 of inst : label is "0000000000000000000010000FC302204D48E6CD26844E5E5A849460A8221088";
    attribute INIT_11 of inst : label is "C81203BA48DA04104709648A200E12C994500000000000000000000000000000";
    attribute INIT_12 of inst : label is "65B7884809B210460A640532314A2A02424099464669290204890C9452427656";
    attribute INIT_13 of inst : label is "034106C04129898413009204C01249871CA48A5DF200948DDD6EF2491B64B649";
    attribute INIT_14 of inst : label is "5E5A8C2C2C2C32663766CC96704D1105983046105C106C06129898049026105E";
    attribute INIT_15 of inst : label is "A4D924442CB940C720A59A2A0828022808E34C03A14C964B2533325D4B7FFF8E";
    attribute INIT_16 of inst : label is "4BB0B040474A4691024924421B9050188910201A3042261860530EE00408CE49";
    attribute INIT_17 of inst : label is "9850E60CF041038C86CA442720741E4125283CC3B449BCBC2CD9127019887048";
    attribute INIT_18 of inst : label is "2A50412D4A6612F221B6366D963673304D9B3B3798826C860858360F190A81B2";
    attribute INIT_19 of inst : label is "6B64032BD8888CDAC564964B2F241A4433E6879374A41483C96301E096CD29F6";
    attribute INIT_1A of inst : label is "AB802D328600022CE1C2C4111A9D4FBB79B826D82882410D2A9983A99457BC90";
    attribute INIT_1B of inst : label is "092CB294C8DEDB5E18252CB20000010060226402835D4A598B0529F4410072DD";
    attribute INIT_1C of inst : label is "186336068887CC50C32EA641A5D4C0D0C3EB29652E71A0013FBD1020B3806196";
    attribute INIT_1D of inst : label is "E65D96CB99765B2CB8B8B985964D7192332222B682A000A800A097B7790923B3";
    attribute INIT_1E of inst : label is "C63B550008000000400802AAD5555556AAD55001AAA005B39F476E6310BA3102";
    attribute INIT_1F of inst : label is "8EA686008B045B02391B8DB106025CB812E5800B8A972E54B96202E0C2002E02";
    attribute INIT_20 of inst : label is "AD2B4AD2B4AD2B4AC234AD2B4AD2B4AD2B4AC234AD2B4AD2B4AD2B2865B42306";
    attribute INIT_21 of inst : label is "BD3F0B00000980086496DB84B396DA66D8400000000000000104445155554234";
    attribute INIT_22 of inst : label is "B2216F860606060707430323A3A32331D1D18CC663301B920F4A099213265B53";
    attribute INIT_23 of inst : label is "24A1562222D8E1925B5993FFFFFFFEAAABFFFEAAAAAAAB752D4F1752D4F045B9";
    attribute INIT_24 of inst : label is "55555555555617FEBA1610D8CB3D22B80C5B9B28717041986484C9658C324B13";
    attribute INIT_25 of inst : label is "B327FFFFFFFFFFFFFFD555555555555555555557FFFFFFFFFFFFFFFFFFFFD555";
    attribute INIT_26 of inst : label is "04C28509002220844A28F100222240460C5368CB18CF464914112EC5B5C324B6";
    attribute INIT_27 of inst : label is "662E4584A47891C4912A611E20887C8B097A250808888A084480A520090A50A4";
    attribute INIT_28 of inst : label is "08A6046246523347DA642988EE45A68BF298BA01223D488B0612238183197405";
    attribute INIT_29 of inst : label is "5929220A623C809845213D80C116242229978E01D90E6824301984F890948229";
    attribute INIT_2A of inst : label is "1C20092444D10A1970C8D343872B84AD443C008708A424A124AC52A044101244";
    attribute INIT_2B of inst : label is "118AAAAAA8160DB5B24661E4424FADEB78B3B9779E79E783B20EE83B28ECA3BA";
    attribute INIT_2C of inst : label is "596C5D96D9665DBD96F659421C458B42DB7BA0748987910C444446C30EDB69B6";
    attribute INIT_2D of inst : label is "8B8B8B85F0FF01F500505B139ECE1B9EC87619B9EC87619B96F9B5BB9DBB9036";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC08EE3F02A2B42ADB6D56DB69D3A3A3B89A98D8D";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "00100080200040010000160000000081843000FFFFFEA30091FE0391C8F8C091";
    attribute INIT_01 of inst : label is "0100943222620101009A70A810C30859E045B53414107800519106244028000A";
    attribute INIT_02 of inst : label is "8102000000C89491281094A7E69309D34987024710888222E2855884314A5733";
    attribute INIT_03 of inst : label is "5124023830920182203237D3C410080B40388004C30D35AF0238002021CA1088";
    attribute INIT_04 of inst : label is "25419554150699D080470AA41C6600C280A2A8C010454000000000004003410C";
    attribute INIT_05 of inst : label is "080000000010000000400200100080000800550000555550000155542828020E";
    attribute INIT_06 of inst : label is "0400008000000000010000400000012480004000400040004000000000400000";
    attribute INIT_07 of inst : label is "1043304888119126700000000000100040010004001000400008000100002000";
    attribute INIT_08 of inst : label is "21A49280D9200000000006801FFA4A2A48E2A49204C02B8248800B180C2A1203";
    attribute INIT_09 of inst : label is "404AD4C4A0944A4400C434502000C4A021022621A140406252952DA20307F516";
    attribute INIT_0A of inst : label is "00924A02002A8354000000000000000000000000000000019200AC8820404040";
    attribute INIT_0B of inst : label is "2A94101544A1504A00AA55855012A080A809644000800A8008089000C4962030";
    attribute INIT_0C of inst : label is "B300008280000000680D04200211100101200128780A24351529A9A9A9484600";
    attribute INIT_0D of inst : label is "56000000000000000000000000000000000000384A0D9790560A4105D124B865";
    attribute INIT_0E of inst : label is "04843106906804372F25804FA799CE79B8161090181C5D0A2A5030028400A020";
    attribute INIT_0F of inst : label is "034528C06182AC15628A679B816141C10A44080100810100005848C0440A115C";
    attribute INIT_10 of inst : label is "000000000000000000000000000A02008D08D01402044E1E1A801C25A0A00010";
    attribute INIT_11 of inst : label is "8000232205495015060B2DA2AA0C165B90400000000000000000000000000000";
    attribute INIT_12 of inst : label is "6C9388001004006008750432238A2A00000803464431290000100190404040E0";
    attribute INIT_13 of inst : label is "05400A800221010002B01208800A283508801875D26050B0010AA082096C96C9";
    attribute INIT_14 of inst : label is "1E1A8A2A2A2A104622228C822046301208102C02CC00A80A22101580904402CC";
    attribute INIT_15 of inst : label is "1210000222A150A72084182AA02AA2800A538E02010C0603011110510B5B6D8E";
    attribute INIT_16 of inst : label is "2A28A020272926488140A022055048188110200200A20444404ABAD00204CD24";
    attribute INIT_17 of inst : label is "00C0C2084000010CA60C4406B860102014383D8C9649F4F46455017019806040";
    attribute INIT_18 of inst : label is "2C0000210A6610F220931324860573302C89191388000A8000422404411880B0";
    attribute INIT_19 of inst : label is "0B2C222318888CCA452486430F2C03423092470B44A014038943008096DC01D0";
    attribute INIT_1A of inst : label is "0980240682000224D1A0C0111ACD64027998161800000000AAB103AB14533C90";
    attribute INIT_1B of inst : label is "0520A31080178816081428A20000010060810040045188511A0421D40000224F";
    attribute INIT_1C of inst : label is "30020008888680C08028C45023484050028A21442421D08C15311054D218C486";
    attribute INIT_1D of inst : label is "72CCB259CB32C96431919804865D319233222212028000AA80AA333278083232";
    attribute INIT_1E of inst : label is "453900001AAA0000C01AAAAA55555002AA400000AAAAAC910A062673919B3906";
    attribute INIT_1F of inst : label is "040303007004490239180C910A00C998064C80198832664193220660C2006406";
    attribute INIT_20 of inst : label is "8C2308C2308C2308C2308C2308C2308C2308C2308C2308C2308C232064902604";
    attribute INIT_21 of inst : label is "15140941001000006C9649049686483248400000000000000104445155554230";
    attribute INIT_22 of inst : label is "A0112B8404040404044202020202022101010C86432031000B88099213665973";
    attribute INIT_23 of inst : label is "24801222224AD1B25949B3FFFFFFFFFFFEAAAAAAAAAAAB5F148415F14840C590";
    attribute INIT_24 of inst : label is "00000000000212BB9E04521142121D280C590A28312820106484D96488364B93";
    attribute INIT_25 of inst : label is "9366AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8000000000000000000000000";
    attribute INIT_26 of inst : label is "02820404100602800A81A00882860084004925DB0CC0C6491011024495A364B2";
    attribute INIT_27 of inst : label is "D6B80C0280D011A200A94034008570180102240401800808000094A000094894";
    attribute INIT_28 of inst : label is "08260A21424A102F59502504680C1059A2D48200A9752A5A8200630100997221";
    attribute INIT_29 of inst : label is "75252209463A805054A0A50080044022A51508018902420A308502E9919282A5";
    attribute INIT_2A of inst : label is "B426040000400818D0401F4107214485423C00460A9410000000C682C0500A55";
    attribute INIT_2B of inst : label is "90AAAAAAA8368C90924224E4A06707C1A463D1528A28A286AA8AA82AA8AAA2AA";
    attribute INIT_2C of inst : label is "0B2448B24B36599486524B02484489404929E074009392844444464926492912";
    attribute INIT_2D of inst : label is "99999991FCFFFE04010049B1DEC509DEC932589DEC932589B268909908998012";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFDF501417C1C0DC1249209249E0C0C0C19BBB9999";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
