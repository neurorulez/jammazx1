-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu2 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu2 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9B7746700BA8BA2E433700BA984567BA984BA2E00B389AB372D439CA8DE2D0F2";
    attribute INIT_01 of inst : label is "4570B3A98B370415637000BA9BA6756700BA982E7456788BA1D6A9BA6745600A";
    attribute INIT_02 of inst : label is "433C433CD543CADEBE8C372D043378874529BA2E7452284B374522918BEB3A2E";
    attribute INIT_03 of inst : label is "2EA2A411402D1CB50EE0140CE3450CCCCCE47BF003D9410CCDCB089AFCD5C7E1";
    attribute INIT_04 of inst : label is "CDD15C0442CCE705426AF2CB7141DB7112EA6EA2CDD5D4C00001100FB50E2680";
    attribute INIT_05 of inst : label is "CEA6A44559158DC0003400002E8888A1C01162CCDD159C00003C0000003AEA62";
    attribute INIT_06 of inst : label is "CCDE01148881AEA240105498CDD0558DC2E626E445919D4002A2899C00013558";
    attribute INIT_07 of inst : label is "455800000002444548899C0002F6A6899D04445499EEAE00115D19C0002E602C";
    attribute INIT_08 of inst : label is "159C000342E00119ECCCCECE81159C0000382EA6A4DC11499C011499C0002BA4";
    attribute INIT_09 of inst : label is "F6628899C46000131AA0115C02A62A45591D000000CDD58CCCE9C0000000CDC1";
    attribute INIT_0A of inst : label is "4444444444773FB73C022EA62E88888888888888888899D159D002E4559C0002";
    attribute INIT_0B of inst : label is "72D87250FA5072D872D852D8721CB610FA503E943E94026D54C048C044444444";
    attribute INIT_0C of inst : label is "929190939298DC8D0A36943E9432D8721CB618732D8721CB610FA503E9433E94";
    attribute INIT_0D of inst : label is "4FC6D5B692DEC8D8D8C608DB04219D163466340C227A7235B58C619392919093";
    attribute INIT_0E of inst : label is "48B1179FEF10F473CA5460A0869671C453E2B540247613DC8171C2C212794721";
    attribute INIT_0F of inst : label is "A2341F72E69C994226963521EE4ECE972D629FB0D2C45E7FBF3578BD72F14E9B";
    attribute INIT_10 of inst : label is "E199A7814E090B09158995BD696A788ADEB7B9A8DCAE90E82DAB4B9E8D4AE94E";
    attribute INIT_11 of inst : label is "61A07D061A07D061A07D061A07D058481F418481F418481F418481F416D2E6B9";
    attribute INIT_12 of inst : label is "62C28B05A7B2F71462C28B05081BEC1BD4258681F418681F418681F418681F41";
    attribute INIT_13 of inst : label is "A788A216285C952562237145C50849E4108D72C22F0518B08BC159EC64BDE464";
    attribute INIT_14 of inst : label is "5B85C7E2F8849E676490D95169651AA37A8D6C5096DA1B9C7DF790F50B963635";
    attribute INIT_15 of inst : label is "253A725237141B8EC8569662DEDAE5ADB4975DE427D09F4A26358D464BDE4608";
    attribute INIT_16 of inst : label is "72F41A5467FBA702665467A74264363439A6639A643A6250505CE7998E79906E";
    attribute INIT_17 of inst : label is "7F924BFC9C7DF798F70B9B6B968F96C509E59A5889DE7D641DE7D6623718218E";
    attribute INIT_18 of inst : label is "8C80C0509192519649351557B934BF894ADA98D08D78218714A24A08909094F2";
    attribute INIT_19 of inst : label is "BA85E033A08660ACDE3083A097378C20CE49434E8879B4E60AC0E8633A084ECC";
    attribute INIT_1A of inst : label is "727521869CE910AD12DDB747B965290EA61A4929091909298D48D4252F1CB06B";
    attribute INIT_1B of inst : label is "9D4BFB952FE9B9D4BF99418484E9927618621CE9109F798F29769AD4061A73A6";
    attribute INIT_1C of inst : label is "614234815355551975582E8BC2D2749D5D55EEEE792FEA5615E7649EED52FC9B";
    attribute INIT_1D of inst : label is "7674C234BFCB9B550D90BA55758421936FF9FDD6174A7A51E70872670534BA55";
    attribute INIT_1E of inst : label is "F1F13232F2F233F3734B736B7378507030F0F1F131310888888B48B0888888BD";
    attribute INIT_1F of inst : label is "1727C1C5C5F0F0F0704951797179517131F2F232F233F3F370487068707030F1";
    attribute INIT_20 of inst : label is "7C4C4C4C7C7C8CBC8C8C8C8C8C8CCCCCCCFCCCCC3C3C0C3C0C0C7C4C7C4F0707";
    attribute INIT_21 of inst : label is "02FC3C0C0C3C0C0C4C4C4C4C7C4C8CBC8C8CBC8CFCCCCCCCCCFC0C0C3C0C3C0C";
    attribute INIT_22 of inst : label is "EEE792FE25595E7E69EED52FE9B944BF99616464E91297498D4859473A452340";
    attribute INIT_23 of inst : label is "BAAAAAAA5D0824E4A5DBF67F45C6D29C9479C21C99D14D2958588D237155D55E";
    attribute INIT_24 of inst : label is "6C6CACFC2C6CFC6F0B0B1B2BC2C2C6F0B1B1BC2C6CEC2C6C6C2C2AAAAAAAA98A";
    attribute INIT_25 of inst : label is "22414A196A56A462594B5942D652D650B51B5265FD4D9D30B52FF2E514327C3C";
    attribute INIT_26 of inst : label is "7BF6424E5A55208E24B04F08FA501A7DFDC13D09392919093994DF87F098548D";
    attribute INIT_27 of inst : label is "3929348261523489052A5FD6DFF9D30B52FF2E5943A422A5392957114627B4BF";
    attribute INIT_28 of inst : label is "9293482615234810522537D914BFCB9750F908902E40890825AA310939291909";
    attribute INIT_29 of inst : label is "69447517968D23718955030198C9D475186A42080FA516F16539392974BB509F";
    attribute INIT_2A of inst : label is "09C4A58548D204158945F64D2FF2E5D43E63B09B5A348D550301D553549D1E7E";
    attribute INIT_2B of inst : label is "D4A42A61C55A57237815D34BFE9585D6108815354A637235AF25393929193482";
    attribute INIT_2C of inst : label is "C2C9C452C8DC41C152F9C6E246164550D619F9A79F5879A4242715615C8D2054";
    attribute INIT_2D of inst : label is "2E80B89BBE90F6EF2C20909185911CBC542D35867E69E7E692FE427CB2C45D5F";
    attribute INIT_2E of inst : label is "C86F571EE7D2FE258D8D497BA25C5CE90E64E4A361AAEBEBF2672C6F9C61E69C";
    attribute INIT_2F of inst : label is "4E7843746598484F70E798390B908D25C5750F93A5A6E61B4F9612FE24E957DF";
    attribute INIT_30 of inst : label is "27DE4A55C822D390B925C5750F93A5B5BD1827D64A5D64D27DE4A55C822D1C52";
    attribute INIT_31 of inst : label is "D264A5D264D27D2E4A55C822D08E7925C53E4E92352827D186427D264A5D264D";
    attribute INIT_32 of inst : label is "AD85B5BD19DD827D264A5D264D27D2E4A55C822D390B925C5750F93A5B58E427";
    attribute INIT_33 of inst : label is "061207D061207D05A2893B89A5818C282049B5B5DA73E692FFE253B8897E5394";
    attribute INIT_34 of inst : label is "94890537B7813FCAA1045703D44442C1224258681F418681F4161207D061207D";
    attribute INIT_35 of inst : label is "0000000030400000000000000000004C4800461045458D0E98948DC5458D0E98";
    attribute INIT_36 of inst : label is "8AA61817149E670D051A96D23A6D649D189F723568E9A59A8DABCB3A6A8D3040";
    attribute INIT_37 of inst : label is "9CE590C97928D7EC1A9C0538349E635E4A1817149E6707EC3618948D5A28D692";
    attribute INIT_38 of inst : label is "9415256E48DC9755256E48DC9715256249714A97BA25C53893A9622B59252DE6";
    attribute INIT_39 of inst : label is "9B69759349F792957208B51432497158D8D4457254948B151CEF9054E2725AE4";
    attribute INIT_3A of inst : label is "D28A0E98705C52799C34186A568AD28D1A9A98EA692D189F4235B7826909F4B8";
    attribute INIT_3B of inst : label is "418481F418481F4169E0630A0B1E6AF6DAE4B5243A8B97928D6DE69E4AD2868A";
    attribute INIT_3C of inst : label is "65277042651EFC6D2F97D0961207D061207D061207D061207D058481F418481F";
    attribute INIT_3D of inst : label is "73835B48E92742227DC2BA6963A346F2CE900000000019D95171A59676545469";
    attribute INIT_3E of inst : label is "89C95B923725D5C95B923725C5C958925C5497B925C53893A9E2225E4A352790";
    attribute INIT_3F of inst : label is "B89B697699349F4B92957208B4E7E450C925C563635115C952522C5473BE4153";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1440111221110040111122111111111115500408811266622622166277773726";
    attribute INIT_01 of inst : label is "111211111000111111122211100001112211114001111CC11511110000111221";
    attribute INIT_02 of inst : label is "21162116622166626633226222111CC011110040011115500011111110000440";
    attribute INIT_03 of inst : label is "04440000221AC9889448A984499884444448999CDC8888844441222267733226";
    attribute INIT_04 of inst : label is "000444800044598888889DEDD211DCC000444000CCC0044888A001D8888488A2";
    attribute INIT_05 of inst : label is "4444000000444448889C888884444445C444440000444488889C8888889C4444";
    attribute INIT_06 of inst : label is "0000C4444449C4440000000000044444484440CCCCC000488844000044444C44";
    attribute INIT_07 of inst : label is "44448888888844445C444488885C440000444445C44440000000444888844440";
    attribute INIT_08 of inst : label is "44448889C8444444444445C444444488889C844400CC000000444444488885C4";
    attribute INIT_09 of inst : label is "5C44000004444444C444444488440CCCCC00488888000444445C488888880004";
    attribute INIT_0A of inst : label is "CCCCCCCCCCCCC888840084444000000000000000000000044448004444448888";
    attribute INIT_0B of inst : label is "4400337722225511000031110040333722225111000001155559999DCCCCCCCC";
    attribute INIT_0C of inst : label is "71717178707CB8CB812C00733326221151000000400337322261111400011111";
    attribute INIT_0D of inst : label is "4665E36DD9B344BCB47ECCB600C3AF1F2C5D2E881BDFE32E6EC7E07272727271";
    attribute INIT_0E of inst : label is "DC63104838086AF90975D8E0F9F5F020138A78C8C8EEF3B675C7ABCBE7C700B0";
    attribute INIT_0F of inst : label is "C12D08D91E7E5FE1BFF92DA33541C29C9B727003B18C4120E9BAECE21B8886F6";
    attribute INIT_10 of inst : label is "30EF4C4482AD9EB67A0EFAAB9BD4C4C5B36CDF74B275E8FC9B76EDF34B475ECF";
    attribute INIT_11 of inst : label is "9B122FA1B132FA1B132FA1B122FA26F44BE86F40BE86F4CBE86F48BE89B37DDF";
    attribute INIT_12 of inst : label is "2982AE02FAC3AE782982AE02300E180E201E6F40BE86F44BE86F44BE86F40BE8";
    attribute INIT_13 of inst : label is "4C7C723310B68DA7B9D20CD71C0F9F1E0C4BB982BB020A60AEC0BE707C6F1C28";
    attribute INIT_14 of inst : label is "CC571E4B9AF9F1CDBE73B5D79F5C0A12E44BB80079B30DF5E381FAAF3DF92D2E";
    attribute INIT_15 of inst : label is "3F13CA7D20CF0C42BA793DF181B37DF79DFDE73C1F7379D79D2E4B67C6F1C2E8";
    attribute INIT_16 of inst : label is "D5BD0B7DCDAAFDA3FE79CDBDE3BCED2D8F9FF0F9BE13FA7434B43E7F83E6F675";
    attribute INIT_17 of inst : label is "95E007FE65E381FAAF3DF6CDF785FB80077DE4D7C57FC7FF97BC7BF1AF30370D";
    attribute INIT_18 of inst : label is "3FB7332070707878E012A79E4EC0754F84BC7CB8CB8673FB088FCA23F2A07646";
    attribute INIT_19 of inst : label is "294BBD111B4B4F1477B721BDCD1DEDC856DCE13AF4ABA474F148461111B4AF07";
    attribute INIT_1A of inst : label is "CBAFA7CFFAFFBAFB470010CA4EC207673C73C62727171707CB8CB81D3848603D";
    attribute INIT_1B of inst : label is "EC0776FA1D6F4EC0776FB7CEFEFF3BAE7CDBFAFFB379CFAE279CFFBEDF3FEBFC";
    attribute INIT_1C of inst : label is "12EB2E48B30DD784175875EE2991ACEB8A2AB193A01DD3D7F88D7D7B11A1D7F4";
    attribute INIT_1D of inst : label is "9F824E207FC6FEA766F9D731D75C2175D55F001C71CCD7DC8D0B4E4D411C5723";
    attribute INIT_1E of inst : label is "191111111911313939091D2D011236327A3A323A121A0888888B88BC888888B6";
    attribute INIT_1F of inst : label is "0F0FC363C3F830103830141438182C3058303830383830381101152509395119";
    attribute INIT_20 of inst : label is "46464E444644444646464C4E4C4644444C4E4E4E8E8C8E8C848E8C84868F8F8F";
    attribute INIT_21 of inst : label is "003C0E0404060C0C0C0E0C04060E0C0E040E0C06040C040406044646444C4E44";
    attribute INIT_22 of inst : label is "193A01DDBD4788DBE7B11A1D7F4E00777FB72E1EFCF37DEFDBEDCB2EBF3CB6C0";
    attribute INIT_23 of inst : label is "11111111A73C9C5C5D755FC0171C7337F72342D39340471C84B6CBD20CD8A2AB";
    attribute INIT_24 of inst : label is "1614161E56565C9D05850587414161D05050741014175C565696911011111011";
    attribute INIT_25 of inst : label is "9210DCBE33E3FC37E0C3E1D0B870B8343C05737EA217E093881FF1BE5D97F616";
    attribute INIT_26 of inst : label is "D55FC5C1C1CD11EDBCE4260A555400459E02402717171717070C7E2AE2E4B6CB";
    attribute INIT_27 of inst : label is "07471E4B92DB2E48433BEA217EEE093881FF1BE5D97C313E17174C9343BF9C59";
    attribute INIT_28 of inst : label is "7071C4B92DB2E48733BE517E707546F9765F0C62BBE3EF842947482717171717";
    attribute INIT_29 of inst : label is "E7004D79F74B92FAEF93BE4CF84F5C4D7CBFE10AA555555AAE4417175F75717C";
    attribute INIT_2A of inst : label is "171C1E4B6CB921CEEF985F9C1D51BE5D97E873A6DD2C4B93366C5DF9743408DB";
    attribute INIT_2B of inst : label is "C81EB3C7CB07D5B2C48BA30754F34B5D70A48B31C1F2C32DC466441717171E4B";
    attribute INIT_2C of inst : label is "8F4FA89BB4830721D388C353EB01F8741C734F1E3575DF5C281F2C1B56CB922C";
    attribute INIT_2D of inst : label is "D291D4F938F8AE646410A07AC07C72A61F2A071CD3C78D7D734281D0418C4070";
    attribute INIT_2E of inst : label is "6665E5893941D53E4B4B88EF4A71384F81BC2B12C9434447F97C101882BC3C7C";
    attribute INIT_2F of inst : label is "E22BCED65DFE7BC2DA1CF28F0CFCCBA7139765F13E4D1A8C25FA81D53C4FA96D";
    attribute INIT_30 of inst : label is "7C73C1CD44B0B8F0CFA7139765F13E6FD7089D7BC5D77D77C73C1CD44B0BAC18";
    attribute INIT_31 of inst : label is "71BC5D797D77C793C1CD44B0B861CFA71317C4FB2D04E97089C9D71BC5D797D7";
    attribute INIT_32 of inst : label is "6B9E6FD70A7289D71BC5D797D77C793C1CD44B0B8F0CFA7139765F13E6FF5C9D";
    attribute INIT_33 of inst : label is "A1B102FA1B132FA29CEF1D4F4F482A76D9EF6CD3A8097E81C753C193EFB5E174";
    attribute INIT_34 of inst : label is "9E48432D6DD0A064C04248C8A6F090803B81E6C44BE06C40BE09B132FA1B112F";
    attribute INIT_35 of inst : label is "00000000000000000000EF4A400E00C8C0088C0424CB4B44FA9F4833CB4B44FA";
    attribute INIT_36 of inst : label is "433C785C79F1CD3B820CF9B313FBDEF9CEFAF32FA24F6D744BC11993F8CB0000";
    attribute INIT_37 of inst : label is "FA3CF84F9F349EA98FFA4108EDF1F2E7CC745C79F1CD42A8ED0EF2CB943CBBB1";
    attribute INIT_38 of inst : label is "9D0CA37984BE9C8EA37984BE9C8CA379A9C0FA8DF6A71304F093171EF7BEBB1F";
    attribute INIT_39 of inst : label is "F5DF5DF5DF1CF073512C2E9D9BE9C4E4B4BA06DA369EC63B7657473253FA3BDA";
    attribute INIT_3A of inst : label is "BF4F24F1C171E7C734EE043FE50DBFCB0FFCBCF3FB19CDFAC32E6FE9CB275C54";
    attribute INIT_3B of inst : label is "E86C40BE86C4CBE893D20A9DB577F2ADBB7CD3001C3DF9FFCBBB1FF7FDB3A50D";
    attribute INIT_3C of inst : label is "5D3AE2A37E7556B41F640079BD12FA1BD22FA1BD22FA1BD12FA26C4CBE86C40B";
    attribute INIT_3D of inst : label is "008EE6DC4F0E731BEBA093DB5112C84664FAA2AAA8A82EB5D7B07D7BAD75E01F";
    attribute INIT_3E of inst : label is "4FE8DE612FA72368DE612FA723E8DE6A70328DF6A71304F0939B10E7DD277C74";
    attribute INIT_3F of inst : label is "54F5DF5C5F5DF1E4F073512C2C3C6A766FA71392D2E81B68DA7B18EDD95D1CC9";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "111111111111111111111111111111111111111CC22222222202220222220202";
    attribute INIT_01 of inst : label is "1111111111111111111111111111111111111111111110011111111111111111";
    attribute INIT_02 of inst : label is "2222222222222202202222202222200111111111111111111111111111111111";
    attribute INIT_03 of inst : label is "04444444400888808888888888888888888888888808888888A2222222222222";
    attribute INIT_04 of inst : label is "4444444028888808888888800CCC000110444444000444444441108808888880";
    attribute INIT_05 of inst : label is "4444444444444444445844444444444584444444444444444458444444584444";
    attribute INIT_06 of inst : label is "4445844444458444444444444444444444444400000444444444444444445844";
    attribute INIT_07 of inst : label is "4444444444444444584444444458444444444445844444444444444444444444";
    attribute INIT_08 of inst : label is "4444444584444444444445844444444444584444440044444444444444444584";
    attribute INIT_09 of inst : label is "5844444444444445844444444444400000444444444444444458444444444444";
    attribute INIT_0A of inst : label is "88888888888888888A2044444444444444444444444444444446204444444444";
    attribute INIT_0B of inst : label is "B11322A00222A0022002033333B3222A2222A222222222E26888888888888888";
    attribute INIT_0C of inst : label is "D0D0D0DCD0D81E81920531802208022080220233333222222222222222201133";
    attribute INIT_0D of inst : label is "24E2A43144C5201416A7641C8AE9883C043404B0AAC7E804314A70D0D0D0D0D0";
    attribute INIT_0E of inst : label is "04EE026AB2A6891DACD34CCCF45172108928AB06E65BC927734D7F7FD2490471";
    attribute INIT_0F of inst : label is "E804101E04C78D6AADF2048800E2A3344C18DEEB63B809AACADA2ACB8B2AE8D3";
    attribute INIT_10 of inst : label is "50CD004C818E8C88DB5CDB4C0C000400C53040501632D2FE4C53040501E32DEF";
    attribute INIT_11 of inst : label is "001C080401C08C4010083401008F400402010040231004C20D004C23D0C10140";
    attribute INIT_12 of inst : label is "30132C88F3CA04D130132C88B82CB22C883400742010074231004420D004423D";
    attribute INIT_13 of inst : label is "006008804D77008404206ECD36FF45142281102332884C04CCA23CF3376806B1";
    attribute INIT_14 of inst : label is "000D36DFB4F4515A249B634D4514290060813220D0C50CD34428D731CCD2060C";
    attribute INIT_15 of inst : label is "3DA3E84006ED8CA3B0D00180A0C5004D34D34D3474D0D3513404813356806B22";
    attribute INIT_16 of inst : label is "40A0ACD35A48267734D35A263736DA0CCF034CF135A3D849B57B3C0D33C4D632";
    attribute INIT_17 of inst : label is "00DA8503834428D731CCD3140128D3220D00400700D34D344D34D34804DFB231";
    attribute INIT_18 of inst : label is "E62EA600D0D0D0D000784C3265B8508D6010D812810937F712E92EBA4B80D367";
    attribute INIT_19 of inst : label is "5116147554145551C54945061471525154614744115011C5551555475541511E";
    attribute INIT_1A of inst : label is "1B8E6F8242FE42E3FDEDCCAA65960D3334D2480D0D0D4D0D81681034B26AC881";
    attribute INIT_1B of inst : label is "58851AF1282F658851AF2F8180FEC38EF80E02FE42FBFF2C2FBFFE39BE090BFB";
    attribute INIT_1C of inst : label is "754B05015266D9098C9232C4120B8CA3296A999952146FDA029ADF799A1282F6";
    attribute INIT_1D of inst : label is "3762A7F85038F40D28D0CB9A4D36A0D3403FAA34D345AEEE9AA9629A0A34CB49";
    attribute INIT_1E of inst : label is "40486458404840444C5C50546C606454506C444860547FF3FFFEFFEBFFFFFFE8";
    attribute INIT_1F of inst : label is "01C3808070E05C786C4054585C6064545C5C50484C54484C54686C6074505C64";
    attribute INIT_20 of inst : label is "1F10151D1B191F1C1F1113141A181C151B181A10191B1F1D161C1E1C1D1C4181";
    attribute INIT_21 of inst : label is "003B18131A1B16191815111F1C11191A151F1D1D1F1211171E1C1F1F1D18191E";
    attribute INIT_22 of inst : label is "99952142BDB429A9E799A1282F65F851AF2FC1D0FFC2FBEFE39BF0E0BFF2B8C0";
    attribute INIT_23 of inst : label is "FCCCCCCD0D4C343434D00BEA8D34D16ABBA6AA58A6828D3D1D52C1006E5296A9";
    attribute INIT_24 of inst : label is "0E0F0F050F0E010E82838303F0C0E0F830383D0F0E0E0B0B0E0E0CCECCCCCDCC";
    attribute INIT_25 of inst : label is "006240707FC77D77CF1D0F0F83C783C3D188C735CC8DD8A9FE140E3C34A37F0E";
    attribute INIT_26 of inst : label is "700BC343436634C6BCC98C8C0001555555A0EE0D0D0D0D0D0D34D82CC4CD52C1";
    attribute INIT_27 of inst : label is "0D0D34D3354B040189735CC8D88D8A9FE140E3C34A343AFC0D0D344D23BC3543";
    attribute INIT_28 of inst : label is "D0D34D3354B040199735E8DDD85028F0D28D0E877BC8EF0A3233EE0D0D0D0D0D";
    attribute INIT_29 of inst : label is "E709F38005010048EF387C3EF2AF31F38637C28C0000000000EE0D0D3708C0DC";
    attribute INIT_2A of inst : label is "0D3434D52C100664CD7A3776140A3C34A348A9C314040138783F33C4C36829A9";
    attribute INIT_2B of inst : label is "9035334D974D04B0C057928500DBD73CFA901726C3606A07D670EE0D0D0D34D3";
    attribute INIT_2C of inst : label is "93CF5D4B001B8F13C9222323D792E0F33CF68B2E68F3C71EA0365C7442C3405C";
    attribute INIT_2D of inst : label is "28F8C8DF30D333D67228C0F5E4B8F2C13CB0CF3DA2CB9A1C72A703F8E3B80AB5";
    attribute INIT_2E of inst : label is "3B3FA71997E14234818330001849B68D22263C207633C2C40E363992277D2496";
    attribute INIT_2F of inst : label is "8FAF2C991CD6FF28911CDD4F7CD241049B0D28D2340187E228D72142348D3F33";
    attribute INIT_30 of inst : label is "34F343EECD3004F7CD049B0D28D234304DAC3CF343CF34F34F343EECD3005F4D";
    attribute INIT_31 of inst : label is "FB343CF134F34F0343EECD3005514F049B2348D1048A70DAC3C3CF7343CF134F";
    attribute INIT_32 of inst : label is "0134304DACF9C3CFF343CF034F34F1343EECD3004F7CD049B0D28D234307343C";
    attribute INIT_33 of inst : label is "C4012083401108F4D0CD0C8D00445632234D30489F8A376141236AF4CD3340D2";
    attribute INIT_34 of inst : label is "10018B43307BC9C9C06A52B522D30E0213034004C201004C2310012080401208";
    attribute INIT_35 of inst : label is "00410010000000010000F0A0AF0000300000380666978328F21001BB978328F2";
    attribute INIT_36 of inst : label is "3334D334D4515AB60ADFF0C523748EF05EF31A077A8D303881D59CA37C410004";
    attribute INIT_37 of inst : label is "F336F2AF00530130DDF104BED892604014DF34D4515A0932DADEFE8123381380";
    attribute INIT_38 of inst : label is "126CC000203212EDC000203212AFC004212AFD0000849B0898C0100D23BC748D";
    attribute INIT_39 of inst : label is "D3CD3CD3CD3CD0FBB34C0034A34126C81831E9CC021013B7221BDBBE236C0002";
    attribute INIT_3A of inst : label is "C16F68D36CD351456AD82377C8CCC1815DFD7DF378005DF33A043043440F3CC8";
    attribute INIT_3B of inst : label is "31004C20D004823D0012048C88D37530C1014815AD4CD00181348DF004C518CC";
    attribute INIT_3C of inst : label is "25B05F3334D0037A158EE0D001F080401F08C4013083401308F40078201007C2";
    attribute INIT_3D of inst : label is "4BED83148D1003ABCC61E34C0220416728DC7FF0CFABCC134D71249304D35049";
    attribute INIT_3E of inst : label is "8DB000080C84BB3000080C84AB7001084ABF0000849B0898C018010014C02490";
    attribute INIT_3F of inst : label is "C8D3CD3C0D3CD3C4D0FBB34C013670D28D049B20E047A73008404EDC886F6EF8";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000010001000001010";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000004400000000000000000";
    attribute INIT_02 of inst : label is "0000000000000010010000010000044000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000004000000000000000000000000004000000000000000000000";
    attribute INIT_04 of inst : label is "0000001100000040000000044000444000000000000000000000000040000000";
    attribute INIT_05 of inst : label is "0000000000000000000800000000000080000000000000000008000000080000";
    attribute INIT_06 of inst : label is "0000800000008000000000000000000000000000000000000000000000000800";
    attribute INIT_07 of inst : label is "0000000000000000080000000008000000000000800000000000000000000000";
    attribute INIT_08 of inst : label is "0000000080000000000000800000000000080000000000000000000000000080";
    attribute INIT_09 of inst : label is "0800000000000000800000000000000000000000000000000008000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "455444455444455445147096644566445664456641665000C800000000000000";
    attribute INIT_0C of inst : label is "30343030303CF04F1D3FA6776667766677667260966641666416664166661944";
    attribute INIT_0D of inst : label is "0703073C00F004FCF09004FF41470B0F3E0F3C1F72D1C13F3C39043030303030";
    attribute INIT_0E of inst : label is "C03B014C3D4072C05071C1C3D071F00001C0C1C141DC3774D1C7030741C72038";
    attribute INIT_0F of inst : label is "413C00DF2CF7C7472C7F3C070043100C0F00344570EC0530FC02F07501D40873";
    attribute INIT_10 of inst : label is "0CC70C340D0C0C0C30CC70C7C700C030F03C0308F03340F40F03C030CF03340F";
    attribute INIT_11 of inst : label is "C30E0F0030E0FC030E0F3030E0FF30C383C00C383F00C343CC0C343FCCF00C03";
    attribute INIT_12 of inst : label is "0DE00743CF013C3E0DE00743500F2D0F500F0C383C00C383F00C383CC0C383FC";
    attribute INIT_13 of inst : label is "0C1200700C301C0300001CC71D3D071C044FCDF0DE4383783790F3C02CCF2D8E";
    attribute INIT_14 of inst : label is "C0071CBF2CD071DE1C7571C7071C83D3CF4FFD003CF0CC70CB20701C0C7F3F3F";
    attribute INIT_15 of inst : label is "1C21C03001CD0CD02C3C30482CF00C071C71C71C0C7031CC0F3FCF02CCF2D841";
    attribute INIT_16 of inst : label is "D33E6071DE331D431C71DE1D031D5F3C0B31C0B31C21C0373C302CC702CC7033";
    attribute INIT_17 of inst : label is "EA460103F0CB207C1F0C73C030087FD0030C30C23071C71C071C71C13C703702";
    attribute INIT_18 of inst : label is "CCC888B0303C3032C0E0071F441018C704F03CF04FC33FD38D40D45035303014";
    attribute INIT_19 of inst : label is "003C00E0003C000380000F0000E00003C0000E0003C00380003C000E0003C038";
    attribute INIT_1A of inst : label is "C17F131C30F4F44F2021201F441003031C31C30303030303CF04FC0C1D407410";
    attribute INIT_1B of inst : label is "40018D7C0697440018D7D31F0FF4FD7D31C030F4F135C707135C78FC4C70C3D3";
    attribute INIT_1C of inst : label is "F0C13C00313FFFCFC7F033770DC17F5FFCC0D1D1080631FC3FDE1C7D13C06974";
    attribute INIT_1D of inst : label is "1D009C30100C7FC3087CCDFFC71D8031EA87031C71CDE1D7DE6158DE031ECDFF";
    attribute INIT_1E of inst : label is "242424282C2C242424282C2C2C2020242C2C202028280CC0CCCCCCCCCCCCCCC3";
    attribute INIT_1F of inst : label is "8103604070E4282C2C2424242428282C2C242828282428282020202424282820";
    attribute INIT_20 of inst : label is "040A0A0B07040405050A0A0B0B08050906070B08050506070B050506060D01C1";
    attribute INIT_21 of inst : label is "0034050906060B0805090A06070805050A06070404090A0A0704080506070704";
    attribute INIT_22 of inst : label is "1D1080631FC7FDE1C7D13C0697443018D7D32F1FF43135C78FC4CB1C3D0C13C0";
    attribute INIT_23 of inst : label is "02222220C7800C0C0C7AA1C0C71C737875F798563780C7B7FC304F001CFFCC0D";
    attribute INIT_24 of inst : label is "0B0908080A09080E4282820390B080E0202C3A0A0809090A080A022122222112";
    attribute INIT_25 of inst : label is "0018C03331F31F31F3F3F3C0FCFCFCF03C0C7E1C310740270004071F0C21FB09";
    attribute INIT_26 of inst : label is "EEA1C0C0C0FF8CF31F7737400000000000071C0303038303031C7F07F83C304F";
    attribute INIT_27 of inst : label is "03031EE0F0C13C0063E1C31073340270004071F0C21F771F03031C07031D1CD1";
    attribute INIT_28 of inst : label is "3031EE0F0C13C0073E1C207420103C7C3087FFF031C3C7DD0D881C0303038303";
    attribute INIT_29 of inst : label is "C7330C3C308FD3C1C7C7E30870871F0C3071F74000000000031C03031DCC703C";
    attribute INIT_2A of inst : label is "031C0FC304F001CF87081D08040F1F0C21C0C733C33F4FC7E30B1F4070780DE1";
    attribute INIT_2B of inst : label is "4C0F31C3C3F0FC13C003C101A87FC31C76000313C0F3C13CF1471C0303431EE0";
    attribute INIT_2C of inst : label is "E0470C01C0070300C1D80331F3C1DC301C77871F7871C71D8C0F0FCBF04F000C";
    attribute INIT_2D of inst : label is "3600CC70DC701C314074303CF07430700C1C071DE1C7DE1C7058C0D000EC03F0";
    attribute INIT_2E of inst : label is "8840BC8D1040631FCFCF01C000353087432D02D3C1884C4C0F1C063D843C1C74";
    attribute INIT_2F of inst : label is "F9F0D5DF2C7090DDDF2C70CBFC704FC353C3087E1F0D10840870C0631F87C480";
    attribute INIT_30 of inst : label is "1C71C0FF6E0DFCBFC7C353C3087E1F3C07700C71C0C71C71C71C0FF6E0DFCF01";
    attribute INIT_31 of inst : label is "731C0C731C71C731C0FF6E0DFCF2C7C353E1F87D3C0DCC7700C0C731C0C731C7";
    attribute INIT_32 of inst : label is "4F0F3C07707500C731C0C731C71C731C0FF6E0DFCBFC7C353C3087E1F3C00C0C";
    attribute INIT_33 of inst : label is "C030E0F3030E0FF31CC7CCC70C38403030C73C03C3021CC06931C20CC7F0F030";
    attribute INIT_34 of inst : label is "0C00636F3C32404C44F18D70C00000C000C0F0C3C3C00C3C3F0C30F0F0030E0F";
    attribute INIT_35 of inst : label is "00410010000800810020F505000033333323EC4F18C3CF08700C0073C3CF0870";
    attribute INIT_36 of inst : label is "031C301C7071DE57000C7CF0E1C71C72CC71C13C34871C0B4F1C5021CB4F0004";
    attribute INIT_37 of inst : label is "702C7087C3002CCC0C7000255C71E3F0C0301C7071DE00CD5C0C704FD888FC78";
    attribute INIT_38 of inst : label is "0DCD070004F00D4D070004F00D4D070000D4CB1C000353CCB40300C1C71C071C";
    attribute INIT_39 of inst : label is "71C71C71C71C703FDB837F0C21F0D4FCFCF0C0C0700C03037037C63031C07000";
    attribute INIT_3A of inst : label is "F00F0870C071C1C7795C0431F620F0CFCC71FFF1C782CC71C13F3C00DF031DCC";
    attribute INIT_3B of inst : label is "F00C383CC0C383FCC30E100C0C31C71CF00C036021CC7C308FC71C70C0F00620";
    attribute INIT_3C of inst : label is "1C13C2071C36A90804F1C03C30E0F0030E0FC030E0F3030E0FF30C383C00C383";
    attribute INIT_3D of inst : label is "0255F3C3875CB771C704E1C704D3D7140872444A21AA7CF1C7301C7E3C71C007";
    attribute INIT_3E of inst : label is "C701C0013C035341C0013C035341C00035341C000353CCB40304C5F0C00B1C70";
    attribute INIT_3F of inst : label is "CC71C71CC71C71CC703FDB837F2D4C3087C353F3F3C30301C0300C0DC0DF18C0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
