library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sinistar_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sinistar_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"7E",X"2E",X"45",X"B6",X"CB",X"00",X"81",X"04",
		X"24",X"1D",X"CE",X"C0",X"10",X"DC",X"28",X"9E",X"2A",X"10",X"9E",X"2C",X"36",X"36",X"DC",X"22",
		X"9E",X"24",X"10",X"9E",X"26",X"36",X"36",X"DC",X"1E",X"9E",X"20",X"36",X"16",X"0F",X"1E",X"B6",
		X"BF",X"FF",X"34",X"02",X"8A",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"B6",X"C8",X"0C",X"86",
		X"39",X"B7",X"CB",X"FF",X"96",X"80",X"85",X"08",X"10",X"27",X"00",X"99",X"DC",X"4C",X"90",X"4F",
		X"C3",X"00",X"80",X"97",X"19",X"9B",X"4F",X"97",X"4F",X"DC",X"49",X"90",X"4E",X"C3",X"00",X"80",
		X"97",X"18",X"9B",X"4E",X"97",X"4E",X"96",X"4A",X"2A",X"04",X"86",X"F0",X"20",X"02",X"86",X"0F",
		X"97",X"1A",X"8E",X"9F",X"60",X"10",X"8E",X"00",X"00",X"4F",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",
		X"EE",X"84",X"A6",X"03",X"43",X"A4",X"C4",X"A7",X"C4",X"DC",X"18",X"AB",X"84",X"81",X"74",X"25",
		X"15",X"31",X"A4",X"26",X"06",X"31",X"21",X"96",X"2E",X"1F",X"89",X"96",X"18",X"2A",X"04",X"86",
		X"73",X"20",X"1F",X"4F",X"20",X"1C",X"5D",X"2A",X"06",X"EB",X"01",X"25",X"15",X"20",X"04",X"EB",
		X"01",X"24",X"0F",X"31",X"A4",X"26",X"0B",X"31",X"21",X"D7",X"1B",X"96",X"30",X"C6",X"74",X"3D",
		X"D6",X"1B",X"ED",X"84",X"EE",X"84",X"E6",X"C4",X"27",X"04",X"6F",X"03",X"20",X"08",X"96",X"1A",
		X"A7",X"03",X"A4",X"02",X"A7",X"C4",X"30",X"04",X"8C",X"9F",X"88",X"26",X"A3",X"86",X"05",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"0C",X"32",X"8E",X"9F",X"F6",X"E6",X"81",X"27",X"12",X"6A",X"1E",
		X"E6",X"1F",X"27",X"0C",X"96",X"5A",X"26",X"08",X"A7",X"1F",X"A7",X"1E",X"AD",X"99",X"41",X"92",
		X"8C",X"9F",X"FC",X"25",X"E5",X"96",X"5A",X"27",X"02",X"0A",X"5A",X"B6",X"C8",X"0C",X"97",X"18",
		X"98",X"59",X"27",X"09",X"D6",X"18",X"D7",X"59",X"8E",X"E1",X"97",X"8D",X"29",X"96",X"8A",X"27",
		X"16",X"96",X"96",X"26",X"12",X"0C",X"5C",X"26",X"0E",X"0C",X"5B",X"26",X"0A",X"CC",X"F1",X"F0",
		X"DD",X"5B",X"C6",X"06",X"BD",X"4A",X"8E",X"12",X"12",X"12",X"35",X"02",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"3B",X"30",X"04",X"58",X"48",X"24",X"FA",X"34",X"17",X"5D",X"2A",X"02",X"30",X"02",
		X"AD",X"94",X"35",X"17",X"26",X"ED",X"39",X"8E",X"9F",X"FA",X"20",X"12",X"8E",X"9F",X"FA",X"20",
		X"1B",X"8E",X"9F",X"F8",X"20",X"08",X"8E",X"9F",X"F8",X"20",X"11",X"8E",X"9F",X"F6",X"A6",X"84",
		X"26",X"13",X"86",X"09",X"A7",X"84",X"A7",X"01",X"39",X"8E",X"9F",X"F6",X"A6",X"84",X"27",X"05",
		X"86",X"02",X"A7",X"84",X"39",X"6F",X"84",X"6F",X"01",X"39",X"4B",X"01",X"4A",X"FB",X"4A",X"F5",
		X"86",X"78",X"97",X"5A",X"39",X"39",X"3F",X"E1",X"95",X"E1",X"95",X"E1",X"90",X"E1",X"90",X"E1",
		X"61",X"E1",X"66",X"E1",X"6B",X"E1",X"79",X"E1",X"95",X"E1",X"95",X"E1",X"57",X"E1",X"5C",X"E1",
		X"95",X"F0",X"03",X"E1",X"95",X"E1",X"95",X"FC",X"A0",X"16",X"10",X"83",X"4F",X"E2",X"26",X"01",
		X"39",X"BD",X"5D",X"A6",X"7E",X"5D",X"C1",X"CC",X"38",X"7A",X"ED",X"25",X"E7",X"27",X"6F",X"A8",
		X"10",X"6E",X"B8",X"1A",X"AE",X"9F",X"50",X"35",X"86",X"0A",X"A7",X"88",X"1D",X"DC",X"78",X"ED",
		X"88",X"11",X"86",X"FF",X"A7",X"88",X"13",X"7D",X"A0",X"13",X"39",X"01",X"02",X"E1",X"EF",X"11",
		X"11",X"BE",X"A0",X"14",X"8C",X"4F",X"B2",X"27",X"06",X"AE",X"9F",X"98",X"78",X"AE",X"0A",X"39",
		X"7E",X"8E",X"D8",X"7E",X"8F",X"18",X"7E",X"8F",X"67",X"7E",X"8E",X"D0",X"7E",X"8F",X"10",X"7E",
		X"8F",X"5F",X"7E",X"8F",X"AF",X"7E",X"8F",X"A2",X"E2",X"25",X"7E",X"8F",X"AA",X"7E",X"8F",X"9D",
		X"E2",X"8F",X"7E",X"E2",X"F9",X"D0",X"EA",X"D0",X"00",X"D0",X"1A",X"D0",X"34",X"D0",X"4E",X"D0",
		X"68",X"D0",X"82",X"D0",X"9C",X"D0",X"B6",X"D0",X"D0",X"D1",X"04",X"D1",X"1E",X"D1",X"38",X"D1",
		X"52",X"D1",X"6C",X"D1",X"86",X"D1",X"A0",X"D1",X"BA",X"D1",X"D4",X"D1",X"EE",X"D1",X"FC",X"D2",
		X"16",X"D2",X"30",X"D2",X"4A",X"D2",X"68",X"D2",X"82",X"D2",X"9C",X"D2",X"B6",X"D2",X"D0",X"D2",
		X"EA",X"D3",X"04",X"D3",X"1E",X"D3",X"38",X"D3",X"52",X"D3",X"70",X"D3",X"8A",X"D3",X"A4",X"D4",
		X"DC",X"D4",X"76",X"D3",X"BE",X"D4",X"1C",X"D3",X"DE",X"D3",X"F0",X"D4",X"06",X"D4",X"48",X"D4",
		X"BC",X"D3",X"D4",X"D4",X"5C",X"D4",X"A2",X"D4",X"32",X"D4",X"90",X"D4",X"52",X"D4",X"C6",X"D4",
		X"F6",X"D5",X"04",X"D5",X"12",X"D5",X"20",X"D5",X"2E",X"D5",X"3C",X"D5",X"4A",X"D5",X"58",X"D5",
		X"66",X"D5",X"74",X"D5",X"82",X"D5",X"88",X"D5",X"96",X"D5",X"A4",X"D5",X"B2",X"D5",X"C0",X"D5",
		X"CE",X"D5",X"DC",X"D5",X"EA",X"D5",X"F8",X"D6",X"06",X"D6",X"14",X"D6",X"22",X"D6",X"30",X"D6",
		X"42",X"D4",X"F6",X"D6",X"50",X"D6",X"5E",X"D6",X"6C",X"D5",X"3C",X"D6",X"7A",X"D6",X"88",X"D6",
		X"96",X"D6",X"A4",X"D6",X"B6",X"D6",X"C4",X"D6",X"D2",X"D6",X"E0",X"D6",X"EE",X"D6",X"F8",X"D7",
		X"02",X"D7",X"10",X"D7",X"16",X"D7",X"24",X"D7",X"32",X"D7",X"38",X"D7",X"3E",X"D7",X"44",X"D7",
		X"6A",X"D7",X"3E",X"D7",X"3E",X"D7",X"3E",X"D7",X"3E",X"34",X"76",X"CE",X"E3",X"3B",X"8E",X"D0",
		X"00",X"86",X"39",X"B7",X"CB",X"FF",X"A6",X"C0",X"27",X"1D",X"34",X"02",X"44",X"44",X"44",X"44",
		X"C6",X"0F",X"E4",X"E0",X"ED",X"81",X"3D",X"31",X"8B",X"34",X"20",X"A6",X"C0",X"8D",X"0A",X"AC",
		X"E4",X"25",X"F8",X"32",X"62",X"20",X"DA",X"35",X"F6",X"8D",X"00",X"8D",X"00",X"5F",X"48",X"24",
		X"02",X"C6",X"10",X"48",X"24",X"02",X"CA",X"01",X"E7",X"80",X"39",X"46",X"00",X"82",X"FF",X"FF",
		X"80",X"00",X"46",X"C6",X"E7",X"F1",X"D9",X"CF",X"EE",X"46",X"60",X"C3",X"C9",X"C9",X"FF",X"76",
		X"46",X"1C",X"16",X"93",X"FF",X"FF",X"90",X"46",X"69",X"CF",X"CD",X"C9",X"F9",X"70",X"46",X"7E",
		X"EB",X"C9",X"C9",X"D9",X"70",X"46",X"03",X"C1",X"F1",X"FD",X"8F",X"01",X"46",X"78",X"EF",X"C5",
		X"C5",X"EF",X"78",X"46",X"06",X"8F",X"C9",X"69",X"3F",X"1E",X"46",X"7E",X"E3",X"C1",X"C1",X"E3",
		X"7E",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"FC",X"39",X"1F",X"13",X"FE",X"70",X"46",
		X"89",X"FF",X"CD",X"89",X"DF",X"F0",X"46",X"3C",X"7E",X"E3",X"C1",X"C3",X"66",X"46",X"C9",X"FF",
		X"81",X"C1",X"FB",X"7E",X"46",X"89",X"FF",X"FD",X"C9",X"C9",X"E3",X"46",X"89",X"FF",X"FD",X"89",
		X"09",X"03",X"46",X"3C",X"7E",X"E3",X"C1",X"D3",X"76",X"46",X"E9",X"FF",X"88",X"18",X"F9",X"FF",
		X"43",X"80",X"F9",X"FF",X"46",X"70",X"C1",X"C1",X"FF",X"7F",X"05",X"46",X"E5",X"FF",X"8C",X"1A",
		X"F3",X"C1",X"46",X"89",X"FF",X"F0",X"80",X"80",X"C0",X"47",X"FF",X"87",X"0C",X"18",X"0D",X"C7",
		X"FF",X"46",X"FF",X"87",X"0C",X"38",X"FF",X"81",X"46",X"7E",X"E3",X"C1",X"C1",X"F3",X"7E",X"46",
		X"91",X"FF",X"F9",X"91",X"16",X"1C",X"46",X"3E",X"63",X"41",X"71",X"E2",X"3E",X"46",X"F1",X"FF",
		X"8D",X"11",X"FA",X"CE",X"46",X"6E",X"C7",X"CF",X"D9",X"7B",X"70",X"46",X"82",X"C3",X"FB",X"7F",
		X"03",X"01",X"46",X"FF",X"F9",X"C0",X"C0",X"C1",X"7F",X"46",X"07",X"7C",X"C0",X"E0",X"7C",X"07",
		X"47",X"FF",X"70",X"38",X"1C",X"38",X"71",X"FF",X"46",X"C1",X"E7",X"38",X"3C",X"E7",X"81",X"46",
		X"01",X"CF",X"98",X"F8",X"7F",X"0F",X"46",X"C0",X"E3",X"F1",X"99",X"CF",X"C7",X"36",X"08",X"21",
		X"86",X"10",X"40",X"16",X"F0",X"00",X"44",X"C7",X"DF",X"00",X"00",X"45",X"00",X"08",X"FF",X"81",
		X"81",X"45",X"81",X"81",X"FF",X"08",X"00",X"45",X"03",X"01",X"DD",X"CF",X"06",X"45",X"07",X"03",
		X"00",X"07",X"03",X"42",X"07",X"03",X"16",X"AA",X"A8",X"46",X"C0",X"60",X"38",X"1C",X"06",X"03",
		X"46",X"14",X"14",X"14",X"14",X"14",X"14",X"44",X"00",X"C3",X"C3",X"00",X"46",X"76",X"DB",X"C9",
		X"DE",X"70",X"D0",X"42",X"20",X"E0",X"45",X"04",X"06",X"FF",X"06",X"04",X"46",X"10",X"38",X"7C",
		X"10",X"10",X"10",X"33",X"FA",X"2F",X"80",X"33",X"93",X"E8",X"00",X"33",X"EA",X"AB",X"80",X"33",
		X"AA",X"AF",X"80",X"33",X"38",X"8F",X"80",X"33",X"BA",X"AE",X"80",X"33",X"FA",X"AE",X"80",X"33",
		X"0B",X"A1",X"80",X"33",X"FA",X"AF",X"80",X"33",X"38",X"AF",X"80",X"13",X"00",X"33",X"F8",X"AF",
		X"80",X"33",X"FA",X"AD",X"80",X"33",X"FA",X"28",X"80",X"33",X"FA",X"27",X"00",X"33",X"FA",X"A8",
		X"80",X"33",X"F8",X"A0",X"80",X"33",X"FA",X"2E",X"80",X"33",X"F8",X"8F",X"80",X"33",X"8B",X"E8",
		X"80",X"33",X"C2",X"0F",X"80",X"33",X"F8",X"8D",X"80",X"33",X"FA",X"08",X"00",X"35",X"F8",X"2F",
		X"82",X"F8",X"33",X"F8",X"2F",X"80",X"33",X"F8",X"A3",X"80",X"33",X"39",X"2B",X"80",X"33",X"F8",
		X"AD",X"80",X"33",X"0B",X"E0",X"80",X"33",X"FA",X"0F",X"80",X"33",X"3B",X"03",X"80",X"35",X"FA",
		X"0F",X"A0",X"F8",X"33",X"D8",X"8D",X"80",X"33",X"3B",X"83",X"80",X"33",X"CA",X"A9",X"80",X"33",
		X"21",X"CA",X"80",X"23",X"55",X"50",X"23",X"22",X"20",X"33",X"0A",X"A3",X"80",X"31",X"B8",X"33",
		X"21",X"48",X"80",X"33",X"89",X"42",X"00",X"31",X"18",X"11",X"C0",X"11",X"80",X"3B",X"FA",X"2F",
		X"80",X"FA",X"2F",X"80",X"FA",X"2F",X"80",X"35",X"20",X"8F",X"9C",X"20",X"00",X"13",X"18",X"13",
		X"1E",X"13",X"0B",X"16",X"0A",X"1E",X"0F",X"1D",X"1E",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",
		X"0B",X"1E",X"8F",X"0B",X"16",X"16",X"0A",X"1D",X"23",X"1D",X"1E",X"0F",X"17",X"1D",X"0A",X"11",
		X"99",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"1C",X"19",X"17",X"0A",X"0F",
		X"1C",X"1C",X"19",X"1C",X"8A",X"0B",X"16",X"16",X"0A",X"1C",X"19",X"17",X"1D",X"0A",X"19",X"95",
		X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",X"19",X"16",X"16",X"19",X"21",X"9D",
		X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"0F",X"0A",X"1E",X"19",
		X"0A",X"0F",X"22",X"13",X"9E",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"1D",
		X"0A",X"0E",X"0F",X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",X"99",X"18",X"19",X"0A",X"0D",X"17",
		X"19",X"9D",X"0D",X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",
		X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"17",X"1F",X"1D",X"1E",X"0A",
		X"0C",X"0F",X"0A",X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",
		X"1E",X"19",X"1A",X"0A",X"1C",X"0B",X"13",X"1D",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"1E",
		X"0F",X"1D",X"9E",X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",X"0F",X"0A",X"1A",X"1C",X"19",X"1E",
		X"0F",X"0D",X"1E",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"0D",X"19",X"16",X"19",X"1C",
		X"0A",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"9E",X"12",X"19",X"1C",X"13",X"24",X"19",X"18",
		X"1E",X"0B",X"16",X"0A",X"0C",X"0B",X"1C",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",
		X"0F",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"1E",X"0F",
		X"1D",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",
		X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",X"11",X"12",X"0A",X"1D",
		X"0D",X"19",X"1C",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",X"10",X"1E",X"0A",X"0D",
		X"19",X"13",X"98",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",X"13",X"98",X"1D",X"16",
		X"0B",X"17",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8B",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8C",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8D",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"0E",X"13",X"1C",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"16",X"0F",X"10",X"1E",X"27",X"1C",
		X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8B",X"16",X"0F",X"10",
		X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8C",
		X"16",X"0F",X"10",X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",
		X"12",X"0A",X"8D",X"16",X"0F",X"10",X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0E",X"13",
		X"1C",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"10",X"13",X"1C",X"8F",X"0C",X"19",X"17",X"8C",X"1D",
		X"19",X"1F",X"18",X"0E",X"0A",X"16",X"13",X"18",X"8F",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",
		X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"16",X"0F",X"10",X"1E",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",
		X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1C",X"13",X"11",X"12",X"1E",
		X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1A",X"0B",X"13",X"0E",X"0A",
		X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"9D",X"10",X"1C",X"0F",X"0F",X"0A",X"1D",X"12",X"13",X"1A",
		X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"13",X"18",X"0A",X"17",
		X"13",X"18",X"1F",X"1E",X"0F",X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1D",X"12",X"13",X"1A",
		X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",
		X"0F",X"0E",X"13",X"1E",X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",
		X"0B",X"11",X"0F",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"9E",X"11",X"0B",X"17",X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",
		X"18",X"1E",X"9D",X"10",X"13",X"1C",X"1D",X"1E",X"0A",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"1D",
		X"12",X"13",X"1A",X"0A",X"0B",X"9E",X"0B",X"0E",X"0E",X"13",X"1E",X"13",X"19",X"18",X"0B",X"16",
		X"0A",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"1D",X"12",X"13",X"1A",X"0A",X"1A",X"19",X"13",X"18",
		X"1E",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"9C",X"1D",X"12",X"13",X"1A",X"1D",X"0A",X"1A",X"0F",
		X"1C",X"0A",X"11",X"0B",X"17",X"8F",X"0E",X"13",X"10",X"10",X"13",X"0D",X"1F",X"16",X"1E",X"23",
		X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",X"0D",X"19",X"18",X"1E",X"13",X"18",X"1F",X"19",
		X"1F",X"1D",X"0A",X"10",X"13",X"1C",X"8F",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",
		X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0B",X"1E",X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",X"0F",
		X"8E",X"1A",X"1C",X"13",X"0D",X"13",X"18",X"11",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"13",
		X"19",X"98",X"0A",X"0A",X"0A",X"0A",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",
		X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1C",X"13",
		X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",
		X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",
		X"0A",X"10",X"19",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"1F",
		X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",
		X"1C",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",
		X"0A",X"0A",X"17",X"13",X"18",X"13",X"17",X"1F",X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",
		X"10",X"19",X"1C",X"0A",X"0B",X"18",X"23",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"1C",X"0F",
		X"1D",X"1E",X"19",X"1C",X"0F",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",
		X"1E",X"1E",X"13",X"18",X"11",X"9D",X"0D",X"16",X"0F",X"0B",X"1C",X"0A",X"0C",X"19",X"19",X"15",
		X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"12",X"13",X"11",
		X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",
		X"1D",X"0F",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"0D",X"23",X"0D",X"16",X"8F",X"1D",X"0F",X"1E",
		X"0A",X"0B",X"1E",X"1E",X"1C",X"0B",X"0D",X"1E",X"0A",X"17",X"19",X"0E",X"0F",X"0A",X"17",X"0F",
		X"1D",X"1D",X"0B",X"11",X"8F",X"1F",X"1D",X"0F",X"0A",X"2C",X"17",X"19",X"20",X"0F",X"2C",X"0A",
		X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"10",
		X"13",X"1C",X"0F",X"27",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",X"2C",X"0A",X"0C",X"1F",
		X"1E",X"1E",X"19",X"18",X"1D",X"0A",X"1E",X"19",X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",X"0A",
		X"1E",X"12",X"0F",X"0A",X"20",X"0B",X"16",X"1F",X"8F",X"23",X"0F",X"9D",X"0B",X"0E",X"14",X"1F",
		X"1D",X"1E",X"17",X"0F",X"18",X"9E",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"0A",X"10",X"0B",X"13",
		X"16",X"1F",X"1C",X"8F",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",X"1E",
		X"13",X"18",X"11",X"1D",X"0A",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"8E",X"0C",X"23",X"0A",
		X"19",X"1A",X"0F",X"18",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",
		X"19",X"1C",X"0A",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"9A",X"0B",
		X"18",X"0E",X"0A",X"1E",X"1F",X"1C",X"18",X"13",X"18",X"11",X"0A",X"11",X"0B",X"17",X"0F",X"0A",
		X"19",X"18",X"0A",X"0B",X"18",X"0E",X"0A",X"19",X"10",X"90",X"0A",X"0D",X"16",X"0F",X"0B",X"1C",
		X"0F",X"8E",X"0A",X"0A",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"E5",X"4D",X"E5",
		X"63",X"E5",X"71",X"E5",X"7B",X"E5",X"85",X"E5",X"90",X"E5",X"A0",X"E5",X"B5",X"E5",X"C9",X"E5",
		X"CB",X"E5",X"D2",X"E5",X"E0",X"E5",X"F7",X"E6",X"13",X"E6",X"2B",X"E6",X"39",X"E6",X"57",X"E6",
		X"62",X"E6",X"69",X"E6",X"70",X"E6",X"7A",X"E6",X"8A",X"E6",X"93",X"E6",X"9E",X"E6",X"A9",X"E6",
		X"B9",X"E6",X"C9",X"E6",X"D9",X"E6",X"E9",X"E6",X"F9",X"E7",X"0A",X"E7",X"1D",X"E7",X"30",X"E7",
		X"43",X"E7",X"57",X"E7",X"5B",X"E7",X"5F",X"E7",X"69",X"E7",X"7B",X"E7",X"8A",X"E7",X"9B",X"E7",
		X"AB",X"E7",X"B7",X"E7",X"C1",X"E7",X"D6",X"E7",X"E8",X"E7",X"FC",X"E8",X"13",X"E8",X"23",X"E8",
		X"36",X"E8",X"58",X"E8",X"66",X"E8",X"78",X"E8",X"87",X"E8",X"A1",X"E8",X"B2",X"E8",X"C5",X"E8",
		X"DA",X"E8",X"EE",X"E9",X"0B",X"E9",X"2E",X"E9",X"4E",X"E9",X"66",X"E9",X"7D",X"E9",X"93",X"E9",
		X"9D",X"E9",X"B5",X"E9",X"CA",X"E9",X"F9",X"E9",X"FC",X"EA",X"06",X"EA",X"0C",X"EA",X"14",X"EA",
		X"2D",X"EA",X"4F",X"EA",X"6A",X"EA",X"72",X"EC",X"5D",X"EC",X"62",X"EC",X"67",X"EC",X"6D",X"EC",
		X"70",X"EC",X"77",X"EC",X"79",X"EC",X"7B",X"EC",X"83",X"EC",X"89",X"EC",X"91",X"EC",X"97",X"EC",
		X"9B",X"EC",X"A0",X"EC",X"A8",X"EC",X"B1",X"EC",X"BD",X"EC",X"C4",X"EC",X"CC",X"EC",X"D3",X"EC",
		X"DC",X"EC",X"E1",X"EC",X"E8",X"EC",X"F0",X"EC",X"FB",X"ED",X"00",X"ED",X"08",X"ED",X"0F",X"ED",
		X"1F",X"ED",X"23",X"ED",X"2C",X"ED",X"30",X"ED",X"39",X"ED",X"42",X"ED",X"45",X"ED",X"4E",X"ED",
		X"52",X"ED",X"55",X"ED",X"5D",X"ED",X"63",X"ED",X"65",X"ED",X"6D",X"ED",X"6F",X"ED",X"7A",X"ED",
		X"7F",X"ED",X"82",X"ED",X"87",X"ED",X"8B",X"ED",X"92",X"ED",X"94",X"ED",X"96",X"ED",X"98",X"ED",
		X"9A",X"ED",X"9C",X"ED",X"9E",X"ED",X"A0",X"ED",X"A2",X"ED",X"A4",X"ED",X"AC",X"ED",X"B1",X"ED",
		X"B3",X"ED",X"B5",X"ED",X"B7",X"ED",X"B9",X"ED",X"BB",X"ED",X"C1",X"ED",X"C4",X"ED",X"C9",X"ED",
		X"CE",X"ED",X"DB",X"ED",X"E5",X"ED",X"EB",X"ED",X"EE",X"ED",X"F8",X"ED",X"FD",X"EE",X"06",X"EE",
		X"12",X"EE",X"16",X"EE",X"1C",X"EE",X"25",X"EE",X"29",X"EE",X"2E",X"EE",X"31",X"EE",X"36",X"EE",
		X"3E",X"EE",X"43",X"EE",X"4D",X"EE",X"54",X"EE",X"59",X"EE",X"5D",X"EE",X"64",X"EE",X"6B",X"EE",
		X"70",X"EE",X"74",X"EE",X"79",X"EE",X"81",X"EE",X"86",X"EE",X"8C",X"EE",X"91",X"EE",X"99",X"EE",
		X"9C",X"EE",X"9F",X"EE",X"A3",X"EE",X"AA",X"EE",X"AE",X"EE",X"B4",X"EE",X"B9",X"EE",X"C0",X"EE",
		X"C4",X"EE",X"C9",X"EE",X"CF",X"EE",X"D5",X"EE",X"DC",X"EE",X"E1",X"EE",X"E6",X"EE",X"EB",X"EE",
		X"EF",X"EE",X"F6",X"EE",X"FE",X"EF",X"03",X"EF",X"09",X"EF",X"0F",X"EF",X"13",X"EF",X"16",X"EF",
		X"1B",X"EF",X"1D",X"EF",X"26",X"EF",X"2F",X"EF",X"37",X"EF",X"3D",X"EF",X"41",X"EF",X"4A",X"EF",
		X"51",X"EF",X"57",X"EF",X"5D",X"EF",X"5F",X"EF",X"66",X"EF",X"6A",X"EF",X"6E",X"EF",X"72",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"0B",X"17",
		X"0F",X"8A",X"19",X"20",X"0F",X"1C",X"8A",X"0C",X"19",X"18",X"1F",X"1D",X"8A",X"0B",X"1E",X"8A",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"8A",X"01",X"8A",X"02",X"8A",X"0D",X"1C",X"0F",X"0E",X"13",
		X"1E",X"1D",X"8A",X"0F",X"17",X"1A",X"1E",X"23",X"8A",X"0D",X"1C",X"23",X"1D",X"1E",X"0B",X"16",
		X"8A",X"1D",X"0B",X"20",X"0F",X"0E",X"8A",X"10",X"19",X"1C",X"8A",X"21",X"0B",X"1C",X"1A",X"8A",
		X"0F",X"18",X"11",X"13",X"18",X"0F",X"1D",X"8A",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",
		X"8A",X"13",X"18",X"1E",X"0F",X"1C",X"0D",X"0F",X"1A",X"1E",X"0F",X"0E",X"8A",X"0B",X"1E",X"1E",
		X"0B",X"0D",X"15",X"8A",X"0E",X"0B",X"17",X"0B",X"11",X"0F",X"0E",X"8A",X"1E",X"0B",X"1C",X"11",
		X"0F",X"1E",X"8A",X"0F",X"18",X"1E",X"0F",X"1C",X"13",X"18",X"11",X"8A",X"20",X"19",X"13",X"0E",
		X"8A",X"21",X"19",X"1C",X"15",X"0F",X"1C",X"8A",X"21",X"0B",X"1C",X"1C",X"13",X"19",X"1C",X"8A",
		X"1A",X"16",X"0B",X"18",X"0F",X"1E",X"19",X"13",X"0E",X"1D",X"8A",X"24",X"19",X"18",X"0F",X"8A",
		X"1A",X"1C",X"0F",X"1A",X"0B",X"1C",X"0F",X"8A",X"0C",X"0B",X"1E",X"1E",X"16",X"0F",X"8A",X"0D",
		X"19",X"18",X"11",X"1C",X"0B",X"1E",X"1F",X"16",X"0B",X"1E",X"13",X"19",X"18",X"1D",X"8A",X"23",
		X"19",X"1F",X"8A",X"0E",X"0F",X"10",X"0F",X"0B",X"1E",X"0F",X"0E",X"8A",X"1E",X"12",X"0F",X"8A",
		X"1D",X"13",X"18",X"13",X"1D",X"1E",X"0B",X"1C",X"8A",X"0D",X"19",X"17",X"1A",X"1F",X"1E",X"0F",
		X"1C",X"8A",X"13",X"1D",X"8A",X"0F",X"18",X"11",X"0B",X"11",X"13",X"18",X"11",X"8A",X"18",X"19",
		X"21",X"8A",X"13",X"18",X"8A",X"1D",X"0D",X"0B",X"18",X"18",X"0F",X"1C",X"8A",X"1C",X"0B",X"18",
		X"11",X"0F",X"8A",X"21",X"8A",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"8A",X"0F",X"8A",X"16",
		X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"8A",X"17",X"13",X"18",X"0F",X"8A",X"1E",
		X"19",X"8A",X"17",X"0B",X"15",X"0F",X"8A",X"1D",X"0B",X"17",X"8A",X"0E",X"13",X"0D",X"15",X"0F",
		X"1C",X"8A",X"18",X"8A",X"19",X"8A",X"0B",X"8A",X"12",X"8A",X"10",X"8A",X"16",X"8A",X"1D",X"8A",
		X"1E",X"8A",X"13",X"8A",X"1C",X"13",X"0D",X"12",X"0B",X"1C",X"0E",X"8A",X"21",X"13",X"1E",X"1E",
		X"8A",X"1C",X"8A",X"0C",X"8A",X"14",X"8A",X"17",X"8A",X"0D",X"8A",X"1D",X"21",X"0B",X"1C",X"17",
		X"8A",X"19",X"10",X"8A",X"1D",X"13",X"18",X"13",X"8A",X"1D",X"1E",X"0B",X"1C",X"8A",X"1D",X"13",
		X"18",X"13",X"17",X"17",X"19",X"1C",X"1E",X"0B",X"16",X"1D",X"8A",X"1D",X"1F",X"1C",X"20",X"13",
		X"20",X"19",X"1C",X"1D",X"8A",X"1E",X"19",X"0E",X"0B",X"23",X"8A",X"1E",X"17",X"8A",X"0D",X"19",
		X"1A",X"23",X"1C",X"13",X"11",X"12",X"1E",X"8A",X"01",X"09",X"08",X"02",X"8A",X"21",X"13",X"16",
		X"16",X"13",X"0B",X"17",X"1D",X"8A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",
		X"1D",X"8A",X"13",X"18",X"0D",X"8A",X"0C",X"16",X"0B",X"1D",X"1E",X"8A",X"0D",X"1C",X"23",X"1D",
		X"1E",X"0B",X"16",X"1D",X"8A",X"19",X"10",X"10",X"8A",X"1A",X"13",X"0D",X"15",X"8A",X"1F",X"1A",
		X"8A",X"10",X"13",X"16",X"16",X"8A",X"0C",X"19",X"17",X"0C",X"0C",X"0B",X"23",X"8A",X"21",X"13",
		X"1E",X"12",X"8A",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",X"1D",X"8A",X"10",X"13",X"1C",
		X"13",X"18",X"11",X"8A",X"0E",X"19",X"0F",X"1D",X"8A",X"18",X"19",X"1E",X"8A",X"0B",X"10",X"10",
		X"0F",X"0D",X"1E",X"8A",X"17",X"13",X"11",X"12",X"1E",X"23",X"8A",X"19",X"18",X"16",X"23",X"8A",
		X"0D",X"0B",X"18",X"8A",X"1E",X"12",X"13",X"1D",X"8A",X"18",X"0F",X"17",X"0F",X"1D",X"13",X"1D",
		X"8A",X"19",X"18",X"0D",X"0F",X"8A",X"0C",X"1F",X"13",X"16",X"1E",X"8A",X"17",X"1F",X"1D",X"1E",
		X"8A",X"0E",X"0F",X"1D",X"1E",X"1C",X"19",X"23",X"8A",X"13",X"1E",X"8A",X"19",X"1C",X"8A",X"12",
		X"0B",X"0E",X"8A",X"0C",X"0F",X"1E",X"1E",X"0F",X"1C",X"8A",X"1C",X"1F",X"18",X"8A",X"1A",X"1C",
		X"0F",X"1D",X"1D",X"8A",X"10",X"13",X"1C",X"0F",X"8A",X"0C",X"1F",X"1E",X"1E",X"19",X"18",X"8A",
		X"1D",X"0F",X"0F",X"8A",X"12",X"13",X"11",X"12",X"8A",X"1D",X"0D",X"19",X"1C",X"0F",X"8A",X"1D",
		X"1E",X"0B",X"1C",X"1E",X"8A",X"13",X"18",X"1D",X"0F",X"1C",X"1E",X"8A",X"0D",X"19",X"13",X"18",
		X"8A",X"1A",X"16",X"0B",X"23",X"8A",X"12",X"0B",X"20",X"0F",X"8A",X"12",X"0B",X"1D",X"8A",X"1A",
		X"13",X"0F",X"0D",X"0F",X"1D",X"8A",X"1D",X"17",X"0B",X"1D",X"12",X"0F",X"0E",X"8A",X"23",X"19",
		X"1F",X"1C",X"8A",X"1C",X"0B",X"18",X"15",X"1D",X"8A",X"0B",X"17",X"19",X"18",X"11",X"8A",X"1E",
		X"19",X"1A",X"8A",X"03",X"00",X"8A",X"11",X"13",X"20",X"0F",X"8A",X"03",X"8A",X"13",X"18",X"13",
		X"1E",X"13",X"0B",X"16",X"1D",X"8A",X"19",X"1A",X"0F",X"1C",X"0B",X"1E",X"19",X"1C",X"8A",X"17",
		X"0F",X"1D",X"1D",X"0B",X"11",X"0F",X"8A",X"0F",X"18",X"1E",X"1C",X"23",X"8A",X"1F",X"1D",X"0F",
		X"8A",X"14",X"19",X"23",X"1D",X"1E",X"13",X"0D",X"15",X"8A",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",
		X"8A",X"1E",X"0B",X"0C",X"16",X"0F",X"8A",X"1C",X"0F",X"1D",X"0F",X"1E",X"8A",X"05",X"8A",X"1A",
		X"19",X"13",X"18",X"1E",X"1D",X"8A",X"01",X"05",X"00",X"8A",X"02",X"00",X"00",X"8A",X"05",X"00",
		X"00",X"8A",X"01",X"05",X"00",X"00",X"00",X"8A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"A6",X"EF",X"B2",
		X"EF",X"BA",X"EF",X"C2",X"EF",X"C6",X"EF",X"D6",X"EF",X"DE",X"EF",X"E2",X"EF",X"E6",X"8E",X"A0",
		X"8E",X"B0",X"8E",X"C4",X"8E",X"C8",X"68",X"55",X"99",X"04",X"42",X"43",X"33",X"05",X"39",X"34",
		X"33",X"86",X"4C",X"2F",X"99",X"08",X"00",X"00",X"99",X"87",X"4C",X"1D",X"99",X"09",X"00",X"00",
		X"99",X"87",X"4C",X"4A",X"22",X"8A",X"4C",X"4A",X"22",X"0A",X"42",X"2B",X"22",X"0D",X"39",X"2B",
		X"99",X"0B",X"34",X"1C",X"99",X"8C",X"4C",X"4B",X"33",X"0E",X"2F",X"1F",X"33",X"8F",X"85",X"57",
		X"88",X"90",X"85",X"3F",X"99",X"A5",X"85",X"43",X"99",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"0B",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"7E",X"2E",X"45",X"B6",X"CB",X"00",X"81",X"04",
		X"24",X"1D",X"CE",X"C0",X"10",X"DC",X"28",X"9E",X"2A",X"10",X"9E",X"2C",X"36",X"36",X"DC",X"22",
		X"9E",X"24",X"10",X"9E",X"26",X"36",X"36",X"DC",X"1E",X"9E",X"20",X"36",X"16",X"0F",X"1E",X"B6",
		X"BF",X"FF",X"34",X"02",X"8A",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"B6",X"C8",X"0C",X"86",
		X"39",X"B7",X"CB",X"FF",X"96",X"80",X"85",X"08",X"10",X"27",X"00",X"99",X"DC",X"4C",X"90",X"4F",
		X"C3",X"00",X"80",X"97",X"19",X"9B",X"4F",X"97",X"4F",X"DC",X"49",X"90",X"4E",X"C3",X"00",X"80",
		X"97",X"18",X"9B",X"4E",X"97",X"4E",X"96",X"4A",X"2A",X"04",X"86",X"F0",X"20",X"02",X"86",X"0F",
		X"97",X"1A",X"8E",X"9F",X"60",X"10",X"8E",X"00",X"00",X"4F",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",
		X"EE",X"84",X"A6",X"03",X"43",X"A4",X"C4",X"A7",X"C4",X"DC",X"18",X"AB",X"84",X"81",X"74",X"25",
		X"15",X"31",X"A4",X"26",X"06",X"31",X"21",X"96",X"2E",X"1F",X"89",X"96",X"18",X"2A",X"04",X"86",
		X"73",X"20",X"1F",X"4F",X"20",X"1C",X"5D",X"2A",X"06",X"EB",X"01",X"25",X"15",X"20",X"04",X"EB",
		X"01",X"24",X"0F",X"31",X"A4",X"26",X"0B",X"31",X"21",X"D7",X"1B",X"96",X"30",X"C6",X"74",X"3D",
		X"D6",X"1B",X"ED",X"84",X"EE",X"84",X"E6",X"C4",X"27",X"04",X"6F",X"03",X"20",X"08",X"96",X"1A",
		X"A7",X"03",X"A4",X"02",X"A7",X"C4",X"30",X"04",X"8C",X"9F",X"88",X"26",X"A3",X"86",X"05",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"0C",X"32",X"8E",X"9F",X"F6",X"E6",X"81",X"27",X"12",X"6A",X"1E",
		X"E6",X"1F",X"27",X"0C",X"96",X"5A",X"26",X"08",X"A7",X"1F",X"A7",X"1E",X"AD",X"99",X"41",X"92",
		X"8C",X"9F",X"FC",X"25",X"E5",X"96",X"5A",X"27",X"02",X"0A",X"5A",X"B6",X"C8",X"0C",X"97",X"18",
		X"98",X"59",X"27",X"09",X"D6",X"18",X"D7",X"59",X"8E",X"E1",X"97",X"8D",X"29",X"96",X"8A",X"27",
		X"16",X"96",X"96",X"26",X"12",X"0C",X"5C",X"26",X"0E",X"0C",X"5B",X"26",X"0A",X"CC",X"F1",X"F0",
		X"DD",X"5B",X"C6",X"06",X"BD",X"4A",X"8E",X"12",X"12",X"12",X"35",X"02",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"3B",X"30",X"04",X"58",X"48",X"24",X"FA",X"34",X"17",X"5D",X"2A",X"02",X"30",X"02",
		X"AD",X"94",X"35",X"17",X"26",X"ED",X"39",X"8E",X"9F",X"FA",X"20",X"12",X"8E",X"9F",X"FA",X"20",
		X"1B",X"8E",X"9F",X"F8",X"20",X"08",X"8E",X"9F",X"F8",X"20",X"11",X"8E",X"9F",X"F6",X"A6",X"84",
		X"26",X"13",X"86",X"09",X"A7",X"84",X"A7",X"01",X"39",X"8E",X"9F",X"F6",X"A6",X"84",X"27",X"05",
		X"86",X"02",X"A7",X"84",X"39",X"6F",X"84",X"6F",X"01",X"39",X"4B",X"01",X"4A",X"FB",X"4A",X"F5",
		X"86",X"78",X"97",X"5A",X"39",X"39",X"3F",X"E1",X"95",X"E1",X"95",X"E1",X"90",X"E1",X"90",X"E1",
		X"61",X"E1",X"66",X"E1",X"6B",X"E1",X"79",X"E1",X"95",X"E1",X"95",X"E1",X"57",X"E1",X"5C",X"E1",
		X"95",X"F0",X"03",X"E1",X"95",X"E1",X"95",X"FC",X"A0",X"16",X"10",X"83",X"4F",X"E2",X"26",X"01",
		X"39",X"BD",X"5D",X"A6",X"7E",X"5D",X"C1",X"CC",X"38",X"7A",X"ED",X"25",X"E7",X"27",X"6F",X"A8",
		X"10",X"6E",X"B8",X"1A",X"AE",X"9F",X"50",X"35",X"86",X"0A",X"A7",X"88",X"1D",X"DC",X"78",X"ED",
		X"88",X"11",X"86",X"FF",X"A7",X"88",X"13",X"7D",X"A0",X"13",X"39",X"01",X"02",X"E1",X"EF",X"11",
		X"11",X"BE",X"A0",X"14",X"8C",X"4F",X"B2",X"27",X"06",X"AE",X"9F",X"98",X"78",X"AE",X"0A",X"39",
		X"7E",X"8E",X"D8",X"7E",X"8F",X"18",X"7E",X"8F",X"67",X"7E",X"8E",X"D0",X"7E",X"8F",X"10",X"7E",
		X"8F",X"5F",X"7E",X"8F",X"AF",X"7E",X"8F",X"A2",X"E2",X"25",X"7E",X"8F",X"AA",X"7E",X"8F",X"9D",
		X"E2",X"8F",X"7E",X"E2",X"F9",X"D0",X"EA",X"D0",X"00",X"D0",X"1A",X"D0",X"34",X"D0",X"4E",X"D0",
		X"68",X"D0",X"82",X"D0",X"9C",X"D0",X"B6",X"D0",X"D0",X"D1",X"04",X"D1",X"1E",X"D1",X"38",X"D1",
		X"52",X"D1",X"6C",X"D1",X"86",X"D1",X"A0",X"D1",X"BA",X"D1",X"D4",X"D1",X"EE",X"D1",X"FC",X"D2",
		X"16",X"D2",X"30",X"D2",X"4A",X"D2",X"68",X"D2",X"82",X"D2",X"9C",X"D2",X"B6",X"D2",X"D0",X"D2",
		X"EA",X"D3",X"04",X"D3",X"1E",X"D3",X"38",X"D3",X"52",X"D3",X"70",X"D3",X"8A",X"D3",X"A4",X"D4",
		X"DC",X"D4",X"76",X"D3",X"BE",X"D4",X"1C",X"D3",X"DE",X"D3",X"F0",X"D4",X"06",X"D4",X"48",X"D4",
		X"BC",X"D3",X"D4",X"D4",X"5C",X"D4",X"A2",X"D4",X"32",X"D4",X"90",X"D4",X"52",X"D4",X"C6",X"D4",
		X"F6",X"D5",X"04",X"D5",X"12",X"D5",X"20",X"D5",X"2E",X"D5",X"3C",X"D5",X"4A",X"D5",X"58",X"D5",
		X"66",X"D5",X"74",X"D5",X"82",X"D5",X"88",X"D5",X"96",X"D5",X"A4",X"D5",X"B2",X"D5",X"C0",X"D5",
		X"CE",X"D5",X"DC",X"D5",X"EA",X"D5",X"F8",X"D6",X"06",X"D6",X"14",X"D6",X"22",X"D6",X"30",X"D6",
		X"42",X"D4",X"F6",X"D6",X"50",X"D6",X"5E",X"D6",X"6C",X"D5",X"3C",X"D6",X"7A",X"D6",X"88",X"D6",
		X"96",X"D6",X"A4",X"D6",X"B6",X"D6",X"C4",X"D6",X"D2",X"D6",X"E0",X"D6",X"EE",X"D6",X"F8",X"D7",
		X"02",X"D7",X"10",X"D7",X"16",X"D7",X"24",X"D7",X"32",X"D7",X"38",X"D7",X"3E",X"D7",X"44",X"D7",
		X"6A",X"D7",X"3E",X"D7",X"3E",X"D7",X"3E",X"D7",X"3E",X"34",X"76",X"CE",X"E3",X"3B",X"8E",X"D0",
		X"00",X"86",X"39",X"B7",X"CB",X"FF",X"A6",X"C0",X"27",X"1D",X"34",X"02",X"44",X"44",X"44",X"44",
		X"C6",X"0F",X"E4",X"E0",X"ED",X"81",X"3D",X"31",X"8B",X"34",X"20",X"A6",X"C0",X"8D",X"0A",X"AC",
		X"E4",X"25",X"F8",X"32",X"62",X"20",X"DA",X"35",X"F6",X"8D",X"00",X"8D",X"00",X"5F",X"48",X"24",
		X"02",X"C6",X"10",X"48",X"24",X"02",X"CA",X"01",X"E7",X"80",X"39",X"46",X"00",X"82",X"FF",X"FF",
		X"80",X"00",X"46",X"C6",X"E7",X"F1",X"D9",X"CF",X"EE",X"46",X"60",X"C3",X"C9",X"C9",X"FF",X"76",
		X"46",X"1C",X"16",X"93",X"FF",X"FF",X"90",X"46",X"69",X"CF",X"CD",X"C9",X"F9",X"70",X"46",X"7E",
		X"EB",X"C9",X"C9",X"D9",X"70",X"46",X"03",X"C1",X"F1",X"FD",X"8F",X"01",X"46",X"78",X"EF",X"C5",
		X"C5",X"EF",X"78",X"46",X"06",X"8F",X"C9",X"69",X"3F",X"1E",X"46",X"7E",X"E3",X"C1",X"C1",X"E3",
		X"7E",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"FC",X"39",X"1F",X"13",X"FE",X"70",X"46",
		X"89",X"FF",X"CD",X"89",X"DF",X"F0",X"46",X"3C",X"7E",X"E3",X"C1",X"C3",X"66",X"46",X"C9",X"FF",
		X"81",X"C1",X"FB",X"7E",X"46",X"89",X"FF",X"FD",X"C9",X"C9",X"E3",X"46",X"89",X"FF",X"FD",X"89",
		X"09",X"03",X"46",X"3C",X"7E",X"E3",X"C1",X"D3",X"76",X"46",X"E9",X"FF",X"88",X"18",X"F9",X"FF",
		X"43",X"80",X"F9",X"FF",X"46",X"70",X"C1",X"C1",X"FF",X"7F",X"05",X"46",X"E5",X"FF",X"8C",X"1A",
		X"F3",X"C1",X"46",X"89",X"FF",X"F0",X"80",X"80",X"C0",X"47",X"FF",X"87",X"0C",X"18",X"0D",X"C7",
		X"FF",X"46",X"FF",X"87",X"0C",X"38",X"FF",X"81",X"46",X"7E",X"E3",X"C1",X"C1",X"F3",X"7E",X"46",
		X"91",X"FF",X"F9",X"91",X"16",X"1C",X"46",X"3E",X"63",X"41",X"71",X"E2",X"3E",X"46",X"F1",X"FF",
		X"8D",X"11",X"FA",X"CE",X"46",X"6E",X"C7",X"CF",X"D9",X"7B",X"70",X"46",X"82",X"C3",X"FB",X"7F",
		X"03",X"01",X"46",X"FF",X"F9",X"C0",X"C0",X"C1",X"7F",X"46",X"07",X"7C",X"C0",X"E0",X"7C",X"07",
		X"47",X"FF",X"70",X"38",X"1C",X"38",X"71",X"FF",X"46",X"C1",X"E7",X"38",X"3C",X"E7",X"81",X"46",
		X"01",X"CF",X"98",X"F8",X"7F",X"0F",X"46",X"C0",X"E3",X"F1",X"99",X"CF",X"C7",X"36",X"08",X"21",
		X"86",X"10",X"40",X"16",X"F0",X"00",X"44",X"C7",X"DF",X"00",X"00",X"45",X"00",X"08",X"FF",X"81",
		X"81",X"45",X"81",X"81",X"FF",X"08",X"00",X"45",X"03",X"01",X"DD",X"CF",X"06",X"45",X"07",X"03",
		X"00",X"07",X"03",X"42",X"07",X"03",X"16",X"AA",X"A8",X"46",X"C0",X"60",X"38",X"1C",X"06",X"03",
		X"46",X"14",X"14",X"14",X"14",X"14",X"14",X"44",X"00",X"C3",X"C3",X"00",X"46",X"76",X"DB",X"C9",
		X"DE",X"70",X"D0",X"42",X"20",X"E0",X"45",X"04",X"06",X"FF",X"06",X"04",X"46",X"10",X"38",X"7C",
		X"10",X"10",X"10",X"33",X"FA",X"2F",X"80",X"33",X"93",X"E8",X"00",X"33",X"EA",X"AB",X"80",X"33",
		X"AA",X"AF",X"80",X"33",X"38",X"8F",X"80",X"33",X"BA",X"AE",X"80",X"33",X"FA",X"AE",X"80",X"33",
		X"0B",X"A1",X"80",X"33",X"FA",X"AF",X"80",X"33",X"38",X"AF",X"80",X"13",X"00",X"33",X"F8",X"AF",
		X"80",X"33",X"FA",X"AD",X"80",X"33",X"FA",X"28",X"80",X"33",X"FA",X"27",X"00",X"33",X"FA",X"A8",
		X"80",X"33",X"F8",X"A0",X"80",X"33",X"FA",X"2E",X"80",X"33",X"F8",X"8F",X"80",X"33",X"8B",X"E8",
		X"80",X"33",X"C2",X"0F",X"80",X"33",X"F8",X"8D",X"80",X"33",X"FA",X"08",X"00",X"35",X"F8",X"2F",
		X"82",X"F8",X"33",X"F8",X"2F",X"80",X"33",X"F8",X"A3",X"80",X"33",X"39",X"2B",X"80",X"33",X"F8",
		X"AD",X"80",X"33",X"0B",X"E0",X"80",X"33",X"FA",X"0F",X"80",X"33",X"3B",X"03",X"80",X"35",X"FA",
		X"0F",X"A0",X"F8",X"33",X"D8",X"8D",X"80",X"33",X"3B",X"83",X"80",X"33",X"CA",X"A9",X"80",X"33",
		X"21",X"CA",X"80",X"23",X"55",X"50",X"23",X"22",X"20",X"33",X"0A",X"A3",X"80",X"31",X"B8",X"33",
		X"21",X"48",X"80",X"33",X"89",X"42",X"00",X"31",X"18",X"11",X"C0",X"11",X"80",X"3B",X"FA",X"2F",
		X"80",X"FA",X"2F",X"80",X"FA",X"2F",X"80",X"35",X"20",X"8F",X"9C",X"20",X"00",X"13",X"18",X"13",
		X"1E",X"13",X"0B",X"16",X"0A",X"1E",X"0F",X"1D",X"1E",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",
		X"0B",X"1E",X"8F",X"0B",X"16",X"16",X"0A",X"1D",X"23",X"1D",X"1E",X"0F",X"17",X"1D",X"0A",X"11",
		X"99",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"1C",X"19",X"17",X"0A",X"0F",
		X"1C",X"1C",X"19",X"1C",X"8A",X"0B",X"16",X"16",X"0A",X"1C",X"19",X"17",X"1D",X"0A",X"19",X"95",
		X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",X"19",X"16",X"16",X"19",X"21",X"9D",
		X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"0F",X"0A",X"1E",X"19",
		X"0A",X"0F",X"22",X"13",X"9E",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"1D",
		X"0A",X"0E",X"0F",X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",X"99",X"18",X"19",X"0A",X"0D",X"17",
		X"19",X"9D",X"0D",X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",
		X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"17",X"1F",X"1D",X"1E",X"0A",
		X"0C",X"0F",X"0A",X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",
		X"1E",X"19",X"1A",X"0A",X"1C",X"0B",X"13",X"1D",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"1E",
		X"0F",X"1D",X"9E",X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",X"0F",X"0A",X"1A",X"1C",X"19",X"1E",
		X"0F",X"0D",X"1E",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"0D",X"19",X"16",X"19",X"1C",
		X"0A",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"9E",X"12",X"19",X"1C",X"13",X"24",X"19",X"18",
		X"1E",X"0B",X"16",X"0A",X"0C",X"0B",X"1C",X"1D",X"0A",X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",
		X"0F",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"1E",X"0F",
		X"1D",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",
		X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",X"11",X"12",X"0A",X"1D",
		X"0D",X"19",X"1C",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",X"10",X"1E",X"0A",X"0D",
		X"19",X"13",X"98",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",X"13",X"98",X"1D",X"16",
		X"0B",X"17",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",X"0A",X"1A",X"16",X"0B",
		X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8B",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8C",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8D",X"1F",X"1A",X"27",X"0E",X"19",X"21",X"18",
		X"0A",X"0E",X"13",X"1C",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"16",X"0F",X"10",X"1E",X"27",X"1C",
		X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8B",X"16",X"0F",X"10",
		X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"12",X"0A",X"8C",
		X"16",X"0F",X"10",X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"21",X"13",X"1E",X"0D",
		X"12",X"0A",X"8D",X"16",X"0F",X"10",X"1E",X"27",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0E",X"13",
		X"1C",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"10",X"13",X"1C",X"8F",X"0C",X"19",X"17",X"8C",X"1D",
		X"19",X"1F",X"18",X"0E",X"0A",X"16",X"13",X"18",X"8F",X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",
		X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"16",X"0F",X"10",X"1E",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",
		X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1C",X"13",X"11",X"12",X"1E",
		X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",X"9D",X"1A",X"0B",X"13",X"0E",X"0A",
		X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"9D",X"10",X"1C",X"0F",X"0F",X"0A",X"1D",X"12",X"13",X"1A",
		X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"13",X"18",X"0A",X"17",
		X"13",X"18",X"1F",X"1E",X"0F",X"9D",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1D",X"12",X"13",X"1A",
		X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",
		X"0F",X"0E",X"13",X"1E",X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",
		X"0B",X"11",X"0F",X"0A",X"1E",X"13",X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"9E",X"11",X"0B",X"17",X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",
		X"18",X"1E",X"9D",X"10",X"13",X"1C",X"1D",X"1E",X"0A",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"1D",
		X"12",X"13",X"1A",X"0A",X"0B",X"9E",X"0B",X"0E",X"0E",X"13",X"1E",X"13",X"19",X"18",X"0B",X"16",
		X"0A",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"1D",X"12",X"13",X"1A",X"0A",X"1A",X"19",X"13",X"18",
		X"1E",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"9C",X"1D",X"12",X"13",X"1A",X"1D",X"0A",X"1A",X"0F",
		X"1C",X"0A",X"11",X"0B",X"17",X"8F",X"0E",X"13",X"10",X"10",X"13",X"0D",X"1F",X"16",X"1E",X"23",
		X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",X"0D",X"19",X"18",X"1E",X"13",X"18",X"1F",X"19",
		X"1F",X"1D",X"0A",X"10",X"13",X"1C",X"8F",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",
		X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0B",X"1E",X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",X"0F",
		X"8E",X"1A",X"1C",X"13",X"0D",X"13",X"18",X"11",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"13",
		X"19",X"98",X"0A",X"0A",X"0A",X"0A",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",
		X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",
		X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1C",X"13",
		X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",
		X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",
		X"0A",X"10",X"19",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"1F",
		X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",
		X"1C",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",
		X"0A",X"0A",X"17",X"13",X"18",X"13",X"17",X"1F",X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",
		X"10",X"19",X"1C",X"0A",X"0B",X"18",X"23",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"1C",X"0F",
		X"1D",X"1E",X"19",X"1C",X"0F",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",
		X"1E",X"1E",X"13",X"18",X"11",X"9D",X"0D",X"16",X"0F",X"0B",X"1C",X"0A",X"0C",X"19",X"19",X"15",
		X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",X"9D",X"12",X"13",X"11",
		X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",
		X"1D",X"0F",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"0D",X"23",X"0D",X"16",X"8F",X"1D",X"0F",X"1E",
		X"0A",X"0B",X"1E",X"1E",X"1C",X"0B",X"0D",X"1E",X"0A",X"17",X"19",X"0E",X"0F",X"0A",X"17",X"0F",
		X"1D",X"1D",X"0B",X"11",X"8F",X"1F",X"1D",X"0F",X"0A",X"2C",X"17",X"19",X"20",X"0F",X"2C",X"0A",
		X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"8A",X"1F",X"1D",X"0F",X"0A",X"2C",X"10",
		X"13",X"1C",X"0F",X"27",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",X"2C",X"0A",X"0C",X"1F",
		X"1E",X"1E",X"19",X"18",X"1D",X"0A",X"1E",X"19",X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",X"0A",
		X"1E",X"12",X"0F",X"0A",X"20",X"0B",X"16",X"1F",X"8F",X"23",X"0F",X"9D",X"0B",X"0E",X"14",X"1F",
		X"1D",X"1E",X"17",X"0F",X"18",X"9E",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"0A",X"10",X"0B",X"13",
		X"16",X"1F",X"1C",X"8F",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",X"0F",X"1E",X"1E",
		X"13",X"18",X"11",X"1D",X"0A",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"8E",X"0C",X"23",X"0A",
		X"19",X"1A",X"0F",X"18",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",
		X"19",X"1C",X"0A",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"9A",X"0B",
		X"18",X"0E",X"0A",X"1E",X"1F",X"1C",X"18",X"13",X"18",X"11",X"0A",X"11",X"0B",X"17",X"0F",X"0A",
		X"19",X"18",X"0A",X"0B",X"18",X"0E",X"0A",X"19",X"10",X"90",X"0A",X"0D",X"16",X"0F",X"0B",X"1C",
		X"0F",X"8E",X"0A",X"0A",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"E5",X"4D",X"E5",
		X"63",X"E5",X"71",X"E5",X"7B",X"E5",X"85",X"E5",X"90",X"E5",X"A0",X"E5",X"B5",X"E5",X"C9",X"E5",
		X"CB",X"E5",X"D2",X"E5",X"E0",X"E5",X"F7",X"E6",X"13",X"E6",X"2B",X"E6",X"39",X"E6",X"57",X"E6",
		X"62",X"E6",X"69",X"E6",X"70",X"E6",X"7A",X"E6",X"8A",X"E6",X"93",X"E6",X"9E",X"E6",X"A9",X"E6",
		X"B9",X"E6",X"C9",X"E6",X"D9",X"E6",X"E9",X"E6",X"F9",X"E7",X"0A",X"E7",X"1D",X"E7",X"30",X"E7",
		X"43",X"E7",X"57",X"E7",X"5B",X"E7",X"5F",X"E7",X"69",X"E7",X"7B",X"E7",X"8A",X"E7",X"9B",X"E7",
		X"AB",X"E7",X"B7",X"E7",X"C1",X"E7",X"D6",X"E7",X"E8",X"E7",X"FC",X"E8",X"13",X"E8",X"23",X"E8",
		X"36",X"E8",X"58",X"E8",X"66",X"E8",X"78",X"E8",X"87",X"E8",X"A1",X"E8",X"B2",X"E8",X"C5",X"E8",
		X"DA",X"E8",X"EE",X"E9",X"0B",X"E9",X"2E",X"E9",X"4E",X"E9",X"66",X"E9",X"7D",X"E9",X"93",X"E9",
		X"9D",X"E9",X"B5",X"E9",X"CA",X"E9",X"F9",X"E9",X"FC",X"EA",X"06",X"EA",X"0C",X"EA",X"14",X"EA",
		X"2D",X"EA",X"4F",X"EA",X"6A",X"EA",X"72",X"EC",X"5D",X"EC",X"62",X"EC",X"67",X"EC",X"6D",X"EC",
		X"70",X"EC",X"77",X"EC",X"79",X"EC",X"7B",X"EC",X"83",X"EC",X"89",X"EC",X"91",X"EC",X"97",X"EC",
		X"9B",X"EC",X"A0",X"EC",X"A8",X"EC",X"B1",X"EC",X"BD",X"EC",X"C4",X"EC",X"CC",X"EC",X"D3",X"EC",
		X"DC",X"EC",X"E1",X"EC",X"E8",X"EC",X"F0",X"EC",X"FB",X"ED",X"00",X"ED",X"08",X"ED",X"0F",X"ED",
		X"1F",X"ED",X"23",X"ED",X"2C",X"ED",X"30",X"ED",X"39",X"ED",X"42",X"ED",X"45",X"ED",X"4E",X"ED",
		X"52",X"ED",X"55",X"ED",X"5D",X"ED",X"63",X"ED",X"65",X"ED",X"6D",X"ED",X"6F",X"ED",X"7A",X"ED",
		X"7F",X"ED",X"82",X"ED",X"87",X"ED",X"8B",X"ED",X"92",X"ED",X"94",X"ED",X"96",X"ED",X"98",X"ED",
		X"9A",X"ED",X"9C",X"ED",X"9E",X"ED",X"A0",X"ED",X"A2",X"ED",X"A4",X"ED",X"AC",X"ED",X"B1",X"ED",
		X"B3",X"ED",X"B5",X"ED",X"B7",X"ED",X"B9",X"ED",X"BB",X"ED",X"C1",X"ED",X"C4",X"ED",X"C9",X"ED",
		X"CE",X"ED",X"DB",X"ED",X"E5",X"ED",X"EB",X"ED",X"EE",X"ED",X"F8",X"ED",X"FD",X"EE",X"06",X"EE",
		X"12",X"EE",X"16",X"EE",X"1C",X"EE",X"25",X"EE",X"29",X"EE",X"2E",X"EE",X"31",X"EE",X"36",X"EE",
		X"3E",X"EE",X"43",X"EE",X"4D",X"EE",X"54",X"EE",X"59",X"EE",X"5D",X"EE",X"64",X"EE",X"6B",X"EE",
		X"70",X"EE",X"74",X"EE",X"79",X"EE",X"81",X"EE",X"86",X"EE",X"8C",X"EE",X"91",X"EE",X"99",X"EE",
		X"9C",X"EE",X"9F",X"EE",X"A3",X"EE",X"AA",X"EE",X"AE",X"EE",X"B4",X"EE",X"B9",X"EE",X"C0",X"EE",
		X"C4",X"EE",X"C9",X"EE",X"CF",X"EE",X"D5",X"EE",X"DC",X"EE",X"E1",X"EE",X"E6",X"EE",X"EB",X"EE",
		X"EF",X"EE",X"F6",X"EE",X"FE",X"EF",X"03",X"EF",X"09",X"EF",X"0F",X"EF",X"13",X"EF",X"16",X"EF",
		X"1B",X"EF",X"1D",X"EF",X"26",X"EF",X"2F",X"EF",X"37",X"EF",X"3D",X"EF",X"41",X"EF",X"4A",X"EF",
		X"51",X"EF",X"57",X"EF",X"5D",X"EF",X"5F",X"EF",X"66",X"EF",X"6A",X"EF",X"6E",X"EF",X"72",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"11",X"0B",X"17",
		X"0F",X"8A",X"19",X"20",X"0F",X"1C",X"8A",X"0C",X"19",X"18",X"1F",X"1D",X"8A",X"0B",X"1E",X"8A",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"8A",X"01",X"8A",X"02",X"8A",X"0D",X"1C",X"0F",X"0E",X"13",
		X"1E",X"1D",X"8A",X"0F",X"17",X"1A",X"1E",X"23",X"8A",X"0D",X"1C",X"23",X"1D",X"1E",X"0B",X"16",
		X"8A",X"1D",X"0B",X"20",X"0F",X"0E",X"8A",X"10",X"19",X"1C",X"8A",X"21",X"0B",X"1C",X"1A",X"8A",
		X"0F",X"18",X"11",X"13",X"18",X"0F",X"1D",X"8A",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",
		X"8A",X"13",X"18",X"1E",X"0F",X"1C",X"0D",X"0F",X"1A",X"1E",X"0F",X"0E",X"8A",X"0B",X"1E",X"1E",
		X"0B",X"0D",X"15",X"8A",X"0E",X"0B",X"17",X"0B",X"11",X"0F",X"0E",X"8A",X"1E",X"0B",X"1C",X"11",
		X"0F",X"1E",X"8A",X"0F",X"18",X"1E",X"0F",X"1C",X"13",X"18",X"11",X"8A",X"20",X"19",X"13",X"0E",
		X"8A",X"21",X"19",X"1C",X"15",X"0F",X"1C",X"8A",X"21",X"0B",X"1C",X"1C",X"13",X"19",X"1C",X"8A",
		X"1A",X"16",X"0B",X"18",X"0F",X"1E",X"19",X"13",X"0E",X"1D",X"8A",X"24",X"19",X"18",X"0F",X"8A",
		X"1A",X"1C",X"0F",X"1A",X"0B",X"1C",X"0F",X"8A",X"0C",X"0B",X"1E",X"1E",X"16",X"0F",X"8A",X"0D",
		X"19",X"18",X"11",X"1C",X"0B",X"1E",X"1F",X"16",X"0B",X"1E",X"13",X"19",X"18",X"1D",X"8A",X"23",
		X"19",X"1F",X"8A",X"0E",X"0F",X"10",X"0F",X"0B",X"1E",X"0F",X"0E",X"8A",X"1E",X"12",X"0F",X"8A",
		X"1D",X"13",X"18",X"13",X"1D",X"1E",X"0B",X"1C",X"8A",X"0D",X"19",X"17",X"1A",X"1F",X"1E",X"0F",
		X"1C",X"8A",X"13",X"1D",X"8A",X"0F",X"18",X"11",X"0B",X"11",X"13",X"18",X"11",X"8A",X"18",X"19",
		X"21",X"8A",X"13",X"18",X"8A",X"1D",X"0D",X"0B",X"18",X"18",X"0F",X"1C",X"8A",X"1C",X"0B",X"18",
		X"11",X"0F",X"8A",X"21",X"8A",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"8A",X"0F",X"8A",X"16",
		X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"8A",X"17",X"13",X"18",X"0F",X"8A",X"1E",
		X"19",X"8A",X"17",X"0B",X"15",X"0F",X"8A",X"1D",X"0B",X"17",X"8A",X"0E",X"13",X"0D",X"15",X"0F",
		X"1C",X"8A",X"18",X"8A",X"19",X"8A",X"0B",X"8A",X"12",X"8A",X"10",X"8A",X"16",X"8A",X"1D",X"8A",
		X"1E",X"8A",X"13",X"8A",X"1C",X"13",X"0D",X"12",X"0B",X"1C",X"0E",X"8A",X"21",X"13",X"1E",X"1E",
		X"8A",X"1C",X"8A",X"0C",X"8A",X"14",X"8A",X"17",X"8A",X"0D",X"8A",X"1D",X"21",X"0B",X"1C",X"17",
		X"8A",X"19",X"10",X"8A",X"1D",X"13",X"18",X"13",X"8A",X"1D",X"1E",X"0B",X"1C",X"8A",X"1D",X"13",
		X"18",X"13",X"17",X"17",X"19",X"1C",X"1E",X"0B",X"16",X"1D",X"8A",X"1D",X"1F",X"1C",X"20",X"13",
		X"20",X"19",X"1C",X"1D",X"8A",X"1E",X"19",X"0E",X"0B",X"23",X"8A",X"1E",X"17",X"8A",X"0D",X"19",
		X"1A",X"23",X"1C",X"13",X"11",X"12",X"1E",X"8A",X"01",X"09",X"08",X"02",X"8A",X"21",X"13",X"16",
		X"16",X"13",X"0B",X"17",X"1D",X"8A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",
		X"1D",X"8A",X"13",X"18",X"0D",X"8A",X"0C",X"16",X"0B",X"1D",X"1E",X"8A",X"0D",X"1C",X"23",X"1D",
		X"1E",X"0B",X"16",X"1D",X"8A",X"19",X"10",X"10",X"8A",X"1A",X"13",X"0D",X"15",X"8A",X"1F",X"1A",
		X"8A",X"10",X"13",X"16",X"16",X"8A",X"0C",X"19",X"17",X"0C",X"0C",X"0B",X"23",X"8A",X"21",X"13",
		X"1E",X"12",X"8A",X"1D",X"13",X"18",X"13",X"0C",X"19",X"17",X"0C",X"1D",X"8A",X"10",X"13",X"1C",
		X"13",X"18",X"11",X"8A",X"0E",X"19",X"0F",X"1D",X"8A",X"18",X"19",X"1E",X"8A",X"0B",X"10",X"10",
		X"0F",X"0D",X"1E",X"8A",X"17",X"13",X"11",X"12",X"1E",X"23",X"8A",X"19",X"18",X"16",X"23",X"8A",
		X"0D",X"0B",X"18",X"8A",X"1E",X"12",X"13",X"1D",X"8A",X"18",X"0F",X"17",X"0F",X"1D",X"13",X"1D",
		X"8A",X"19",X"18",X"0D",X"0F",X"8A",X"0C",X"1F",X"13",X"16",X"1E",X"8A",X"17",X"1F",X"1D",X"1E",
		X"8A",X"0E",X"0F",X"1D",X"1E",X"1C",X"19",X"23",X"8A",X"13",X"1E",X"8A",X"19",X"1C",X"8A",X"12",
		X"0B",X"0E",X"8A",X"0C",X"0F",X"1E",X"1E",X"0F",X"1C",X"8A",X"1C",X"1F",X"18",X"8A",X"1A",X"1C",
		X"0F",X"1D",X"1D",X"8A",X"10",X"13",X"1C",X"0F",X"8A",X"0C",X"1F",X"1E",X"1E",X"19",X"18",X"8A",
		X"1D",X"0F",X"0F",X"8A",X"12",X"13",X"11",X"12",X"8A",X"1D",X"0D",X"19",X"1C",X"0F",X"8A",X"1D",
		X"1E",X"0B",X"1C",X"1E",X"8A",X"13",X"18",X"1D",X"0F",X"1C",X"1E",X"8A",X"0D",X"19",X"13",X"18",
		X"8A",X"1A",X"16",X"0B",X"23",X"8A",X"12",X"0B",X"20",X"0F",X"8A",X"12",X"0B",X"1D",X"8A",X"1A",
		X"13",X"0F",X"0D",X"0F",X"1D",X"8A",X"1D",X"17",X"0B",X"1D",X"12",X"0F",X"0E",X"8A",X"23",X"19",
		X"1F",X"1C",X"8A",X"1C",X"0B",X"18",X"15",X"1D",X"8A",X"0B",X"17",X"19",X"18",X"11",X"8A",X"1E",
		X"19",X"1A",X"8A",X"03",X"00",X"8A",X"11",X"13",X"20",X"0F",X"8A",X"03",X"8A",X"13",X"18",X"13",
		X"1E",X"13",X"0B",X"16",X"1D",X"8A",X"19",X"1A",X"0F",X"1C",X"0B",X"1E",X"19",X"1C",X"8A",X"17",
		X"0F",X"1D",X"1D",X"0B",X"11",X"0F",X"8A",X"0F",X"18",X"1E",X"1C",X"23",X"8A",X"1F",X"1D",X"0F",
		X"8A",X"14",X"19",X"23",X"1D",X"1E",X"13",X"0D",X"15",X"8A",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",
		X"8A",X"1E",X"0B",X"0C",X"16",X"0F",X"8A",X"1C",X"0F",X"1D",X"0F",X"1E",X"8A",X"05",X"8A",X"1A",
		X"19",X"13",X"18",X"1E",X"1D",X"8A",X"01",X"05",X"00",X"8A",X"02",X"00",X"00",X"8A",X"05",X"00",
		X"00",X"8A",X"01",X"05",X"00",X"00",X"00",X"8A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"A6",X"EF",X"B2",
		X"EF",X"BA",X"EF",X"C2",X"EF",X"C6",X"EF",X"D6",X"EF",X"DE",X"EF",X"E2",X"EF",X"E6",X"8E",X"A0",
		X"8E",X"B0",X"8E",X"C4",X"8E",X"C8",X"68",X"55",X"99",X"04",X"42",X"43",X"33",X"05",X"39",X"34",
		X"33",X"86",X"4C",X"2F",X"99",X"08",X"00",X"00",X"99",X"87",X"4C",X"1D",X"99",X"09",X"00",X"00",
		X"99",X"87",X"4C",X"4A",X"22",X"8A",X"4C",X"4A",X"22",X"0A",X"42",X"2B",X"22",X"0D",X"39",X"2B",
		X"99",X"0B",X"34",X"1C",X"99",X"8C",X"4C",X"4B",X"33",X"0E",X"2F",X"1F",X"33",X"8F",X"85",X"57",
		X"88",X"90",X"85",X"3F",X"99",X"A5",X"85",X"43",X"99",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"0B",X"E0",X"00",X"E0",X"00",X"E0",X"00",
		X"7E",X"F0",X"1F",X"7E",X"F3",X"71",X"7E",X"F4",X"A1",X"7E",X"F9",X"97",X"7E",X"FF",X"57",X"00",
		X"F9",X"07",X"28",X"2F",X"00",X"A4",X"15",X"C7",X"FF",X"38",X"17",X"CC",X"81",X"81",X"2F",X"1A",
		X"FF",X"10",X"CE",X"BF",X"00",X"7F",X"C8",X"0D",X"7F",X"C8",X"0C",X"86",X"3C",X"B7",X"C8",X"0D",
		X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",X"B7",X"C8",X"0F",X"86",X"C0",X"B7",
		X"C8",X"0E",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"8E",X"F0",X"0F",X"10",X"8E",X"C0",
		X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"1F",X"25",X"F7",X"86",X"02",X"10",X"8E",X"F0",X"65",
		X"8E",X"00",X"00",X"20",X"3A",X"10",X"8E",X"F0",X"6C",X"7E",X"F2",X"BD",X"86",X"34",X"B7",X"C8",
		X"0D",X"B7",X"C8",X"0F",X"7F",X"C8",X"0E",X"86",X"BF",X"1F",X"8B",X"10",X"CE",X"BF",X"00",X"7E",
		X"FF",X"C0",X"86",X"00",X"8E",X"55",X"37",X"C6",X"99",X"BD",X"E2",X"03",X"86",X"01",X"8E",X"42",
		X"4B",X"C6",X"99",X"BD",X"E2",X"03",X"10",X"8E",X"49",X"F9",X"86",X"07",X"7E",X"F1",X"FD",X"1A",
		X"3F",X"7F",X"BF",X"FF",X"7F",X"C9",X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",X"8E",X"00",X"00",
		X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",
		X"56",X"20",X"02",X"44",X"56",X"ED",X"81",X"1E",X"10",X"5D",X"26",X"16",X"C6",X"39",X"F7",X"CB",
		X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"0A",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"03",X"7E",X"F1",
		X"EA",X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",X"03",X"8E",X"D0",X"00",X"8C",X"E0",X"00",X"26",
		X"BF",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",
		X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"10",X"A3",X"81",X"26",X"4A",
		X"1E",X"10",X"5D",X"26",X"16",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",X"C1",X"FF",X"26",X"0A",
		X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"03",X"7E",X"F1",X"EA",X"5F",X"1E",X"10",X"8C",X"C0",X"00",
		X"26",X"03",X"8E",X"D0",X"00",X"8C",X"E0",X"00",X"26",X"BC",X"1F",X"03",X"1F",X"B8",X"81",X"FF",
		X"26",X"05",X"1F",X"30",X"7E",X"F0",X"AD",X"4A",X"1F",X"8B",X"81",X"80",X"10",X"27",X"00",X"9A",
		X"4D",X"1F",X"30",X"10",X"26",X"FF",X"56",X"7E",X"F1",X"EA",X"30",X"1E",X"A8",X"84",X"E8",X"01",
		X"4D",X"26",X"07",X"5D",X"26",X"04",X"30",X"02",X"20",X"A6",X"CE",X"00",X"42",X"8C",X"D8",X"00",
		X"24",X"30",X"33",X"5F",X"8C",X"D0",X"00",X"24",X"29",X"CE",X"00",X"30",X"1E",X"10",X"5F",X"1E",
		X"10",X"8C",X"00",X"00",X"27",X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",X"10",X"11",X"83",X"00",
		X"30",X"23",X"EE",X"CE",X"00",X"10",X"20",X"E9",X"33",X"41",X"47",X"25",X"05",X"57",X"25",X"02",
		X"20",X"F6",X"1F",X"30",X"10",X"CE",X"F1",X"AA",X"20",X"67",X"86",X"BF",X"1F",X"8B",X"1F",X"A8",
		X"43",X"10",X"8E",X"F1",X"B7",X"20",X"33",X"BD",X"32",X"45",X"85",X"C0",X"26",X"0A",X"86",X"00",
		X"8E",X"55",X"37",X"C6",X"22",X"BD",X"E2",X"03",X"86",X"02",X"8E",X"42",X"52",X"C6",X"22",X"BD",
		X"E2",X"03",X"1F",X"30",X"1F",X"98",X"C6",X"22",X"BD",X"E2",X"06",X"1F",X"A8",X"85",X"40",X"26",
		X"03",X"7E",X"F9",X"29",X"10",X"8E",X"49",X"F9",X"20",X"11",X"C6",X"01",X"F7",X"BF",X"FF",X"F7",
		X"C9",X"00",X"10",X"CE",X"BF",X"00",X"BD",X"E2",X"22",X"6E",X"A4",X"86",X"20",X"8E",X"58",X"00",
		X"30",X"1F",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",X"EE",X"6E",
		X"A4",X"1F",X"03",X"86",X"02",X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"F2",X"20",X"7E",X"F2",X"9B",
		X"86",X"02",X"10",X"8E",X"F2",X"28",X"20",X"D5",X"10",X"8E",X"F2",X"2E",X"20",X"5D",X"86",X"01",
		X"10",X"8E",X"F2",X"36",X"20",X"C7",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",X"8E",
		X"F2",X"44",X"20",X"57",X"86",X"02",X"10",X"8E",X"F2",X"4C",X"20",X"B1",X"10",X"8E",X"F2",X"52",
		X"20",X"39",X"86",X"01",X"10",X"8E",X"F2",X"5A",X"20",X"A3",X"1F",X"30",X"1F",X"98",X"10",X"8E",
		X"F2",X"64",X"20",X"37",X"86",X"02",X"10",X"8E",X"F2",X"6C",X"20",X"91",X"10",X"8E",X"F2",X"72",
		X"20",X"19",X"86",X"05",X"10",X"8E",X"F2",X"7A",X"20",X"83",X"1F",X"B8",X"4A",X"1F",X"8B",X"26",
		X"96",X"10",X"8E",X"F2",X"87",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",X"B7",X"C8",X"0D",
		X"4C",X"B7",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",X"46",X"46",X"46",
		X"84",X"C0",X"B7",X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0F",
		X"86",X"34",X"C5",X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",X"1A",X"3F",X"8E",
		X"F3",X"4F",X"8C",X"F3",X"6F",X"26",X"02",X"6E",X"A4",X"A6",X"01",X"27",X"18",X"A6",X"84",X"5F",
		X"1F",X"03",X"86",X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",X"1E",X"03",X"26",
		X"F3",X"E1",X"01",X"26",X"04",X"30",X"02",X"20",X"D9",X"A6",X"84",X"44",X"44",X"44",X"44",X"81",
		X"0D",X"25",X"02",X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",X"CE",X"F3",X"03",
		X"7E",X"F2",X"11",X"86",X"BF",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"BF",X"00",
		X"BD",X"32",X"45",X"1F",X"A8",X"43",X"F7",X"BF",X"06",X"85",X"C0",X"26",X"0A",X"86",X"00",X"8E",
		X"55",X"37",X"C6",X"22",X"BD",X"E2",X"03",X"86",X"03",X"8E",X"42",X"52",X"C6",X"22",X"BD",X"E2",
		X"03",X"B6",X"BF",X"06",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"C6",X"22",X"BD",X"E2",X"06",X"1F",
		X"A9",X"C5",X"40",X"26",X"03",X"7E",X"F9",X"2E",X"10",X"8E",X"49",X"F9",X"7E",X"F1",X"FB",X"00",
		X"C6",X"10",X"62",X"20",X"20",X"30",X"33",X"40",X"EF",X"50",X"FC",X"60",X"1A",X"70",X"59",X"80",
		X"2A",X"90",X"00",X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",X"00",X"E0",X"F8",X"F0",X"57",X"00",
		X"00",X"86",X"04",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",
		X"FF",X"B7",X"BF",X"09",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"BD",X"F4",X"90",X"B6",
		X"C8",X"0C",X"46",X"10",X"25",X"06",X"10",X"BD",X"32",X"45",X"1A",X"BF",X"10",X"8E",X"F3",X"A3",
		X"7E",X"F2",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"10",
		X"8E",X"F3",X"B6",X"7E",X"F2",X"BD",X"86",X"BF",X"1F",X"8B",X"BD",X"32",X"45",X"86",X"00",X"BD",
		X"E2",X"12",X"C6",X"03",X"8E",X"70",X"00",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",
		X"02",X"26",X"16",X"30",X"1F",X"8C",X"00",X"00",X"26",X"ED",X"5A",X"26",X"E7",X"10",X"8E",X"F3",
		X"E9",X"8E",X"00",X"00",X"86",X"FF",X"7E",X"F0",X"9F",X"86",X"BF",X"1F",X"8B",X"BD",X"32",X"45",
		X"86",X"01",X"BD",X"E2",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",
		X"F4",X"8E",X"9C",X"00",X"6F",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",X"01",X"26",X"F4",
		X"CC",X"A5",X"5A",X"FD",X"BF",X"0B",X"B7",X"BF",X"09",X"8D",X"68",X"BD",X"F9",X"67",X"BD",X"FE",
		X"F0",X"86",X"02",X"24",X"24",X"C6",X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",X"10",X"CE",
		X"F4",X"37",X"86",X"03",X"7E",X"F2",X"11",X"10",X"CE",X"BF",X"00",X"8D",X"46",X"86",X"BF",X"1F",
		X"8B",X"86",X"03",X"C1",X"1F",X"22",X"02",X"86",X"04",X"BD",X"32",X"45",X"BD",X"E2",X"12",X"BD",
		X"F9",X"67",X"7F",X"BF",X"08",X"BD",X"FE",X"6C",X"BD",X"FE",X"76",X"BD",X"F9",X"8A",X"24",X"F8",
		X"86",X"3F",X"B7",X"C8",X"0E",X"4F",X"BD",X"F9",X"97",X"4F",X"B7",X"C8",X"0E",X"BD",X"F9",X"67",
		X"BD",X"F7",X"B8",X"BD",X"F9",X"67",X"BD",X"F7",X"1C",X"BD",X"F9",X"8A",X"24",X"03",X"BD",X"F9",
		X"67",X"20",X"75",X"7F",X"C8",X"0E",X"86",X"34",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"39",
		X"8E",X"F0",X"0F",X"10",X"8E",X"C0",X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"1F",X"25",X"F7",
		X"39",X"86",X"3C",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",
		X"3F",X"1F",X"8A",X"86",X"8F",X"BE",X"C5",X"01",X"30",X"89",X"12",X"34",X"10",X"8E",X"F4",X"C3",
		X"7E",X"F0",X"9F",X"10",X"8E",X"F4",X"CA",X"7E",X"F2",X"BD",X"86",X"BF",X"1F",X"8B",X"10",X"CE",
		X"BF",X"00",X"BD",X"FE",X"F0",X"24",X"16",X"86",X"04",X"8C",X"CD",X"00",X"23",X"02",X"86",X"03",
		X"BD",X"32",X"45",X"BD",X"E2",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"F9",X"8D",X"31",X"10",
		X"8E",X"F4",X"A1",X"86",X"04",X"7E",X"F1",X"FD",X"8D",X"78",X"BD",X"F9",X"67",X"BD",X"32",X"45",
		X"86",X"07",X"B7",X"C0",X"00",X"BD",X"F9",X"67",X"86",X"38",X"B7",X"C0",X"00",X"BD",X"F9",X"67",
		X"86",X"C0",X"B7",X"C0",X"00",X"BD",X"F9",X"67",X"8D",X"06",X"BD",X"F9",X"67",X"7E",X"F9",X"A7",
		X"8E",X"C0",X"00",X"10",X"8E",X"F5",X"62",X"EC",X"A1",X"ED",X"81",X"86",X"39",X"B7",X"CB",X"FF",
		X"8C",X"C0",X"10",X"25",X"F2",X"CC",X"00",X"00",X"8E",X"00",X"00",X"BF",X"BF",X"06",X"30",X"89",
		X"0F",X"00",X"ED",X"83",X"34",X"02",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"02",X"BC",X"BF",X"06",
		X"26",X"F0",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",
		X"DA",X"39",X"05",X"05",X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",
		X"85",X"85",X"BD",X"32",X"45",X"4F",X"BD",X"F7",X"AD",X"7F",X"BF",X"FF",X"7F",X"C9",X"00",X"86",
		X"FF",X"B7",X"C0",X"01",X"86",X"C0",X"B7",X"C0",X"02",X"86",X"38",X"B7",X"C0",X"03",X"86",X"07",
		X"B7",X"C0",X"04",X"10",X"8E",X"F6",X"A4",X"CC",X"01",X"01",X"AE",X"A4",X"C6",X"39",X"F7",X"CB",
		X"FF",X"C6",X"01",X"ED",X"81",X"AC",X"22",X"26",X"FA",X"31",X"24",X"10",X"8C",X"F6",X"CC",X"26",
		X"E9",X"86",X"11",X"10",X"8E",X"F6",X"84",X"AE",X"A4",X"BF",X"BF",X"06",X"A7",X"84",X"7C",X"BF",
		X"06",X"C6",X"39",X"F7",X"CB",X"FF",X"BE",X"BF",X"06",X"AC",X"22",X"26",X"EF",X"31",X"24",X"10",
		X"8C",X"F6",X"A4",X"26",X"E2",X"10",X"8E",X"F6",X"CC",X"AE",X"A4",X"BF",X"BF",X"06",X"A6",X"24",
		X"A7",X"84",X"7C",X"BF",X"06",X"C6",X"39",X"F7",X"CB",X"FF",X"BE",X"BF",X"06",X"AC",X"22",X"26",
		X"EF",X"31",X"25",X"10",X"8C",X"F7",X"08",X"26",X"E0",X"10",X"8E",X"F7",X"08",X"AE",X"A4",X"A6",
		X"24",X"A7",X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"AC",X"22",X"26",X"F5",X"31",X"25",X"10",X"8C",
		X"F7",X"1C",X"26",X"E9",X"86",X"21",X"B7",X"43",X"7E",X"86",X"20",X"B7",X"93",X"7E",X"8E",X"4B",
		X"0A",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",
		X"6D",X"26",X"EE",X"8E",X"4B",X"90",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",
		X"FF",X"A7",X"80",X"8C",X"4B",X"F3",X"26",X"EE",X"8E",X"0B",X"18",X"BF",X"BF",X"06",X"BE",X"BF",
		X"06",X"A6",X"84",X"84",X"F0",X"8A",X"01",X"A7",X"84",X"F6",X"BF",X"07",X"CB",X"22",X"25",X"05",
		X"F7",X"BF",X"07",X"20",X"E9",X"C6",X"18",X"F7",X"BF",X"07",X"F6",X"BF",X"06",X"CB",X"10",X"F7",
		X"BF",X"06",X"C1",X"9B",X"26",X"D8",X"C6",X"01",X"F7",X"BF",X"FF",X"F7",X"C9",X"00",X"C6",X"39",
		X"F7",X"CB",X"FF",X"39",X"04",X"07",X"94",X"07",X"04",X"29",X"94",X"29",X"04",X"4B",X"94",X"4B",
		X"04",X"6D",X"94",X"6D",X"04",X"8F",X"94",X"8F",X"04",X"B1",X"94",X"B1",X"04",X"D3",X"94",X"D3",
		X"04",X"F5",X"94",X"F5",X"03",X"07",X"03",X"F5",X"13",X"07",X"13",X"F5",X"23",X"07",X"23",X"F5",
		X"33",X"07",X"33",X"F5",X"43",X"07",X"43",X"F5",X"53",X"07",X"53",X"F5",X"63",X"07",X"63",X"F5",
		X"73",X"07",X"73",X"F5",X"83",X"07",X"83",X"F5",X"93",X"07",X"93",X"F5",X"45",X"05",X"52",X"05",
		X"44",X"45",X"06",X"52",X"06",X"44",X"45",X"07",X"52",X"07",X"00",X"45",X"08",X"52",X"08",X"33",
		X"45",X"09",X"52",X"09",X"33",X"45",X"F3",X"52",X"F3",X"33",X"45",X"F4",X"52",X"F4",X"33",X"45",
		X"F5",X"52",X"F5",X"00",X"45",X"F6",X"52",X"F6",X"44",X"45",X"F7",X"52",X"F7",X"44",X"04",X"7E",
		X"43",X"7E",X"22",X"54",X"7E",X"93",X"7E",X"22",X"02",X"6F",X"02",X"8E",X"04",X"03",X"6F",X"03",
		X"8E",X"30",X"93",X"6F",X"93",X"8E",X"00",X"94",X"6F",X"94",X"8E",X"34",X"BD",X"32",X"45",X"86",
		X"05",X"BD",X"E2",X"12",X"86",X"80",X"B7",X"BF",X"1F",X"4F",X"BD",X"F9",X"97",X"BD",X"F9",X"8A",
		X"25",X"33",X"7A",X"BF",X"1F",X"26",X"F2",X"B6",X"F7",X"95",X"8D",X"71",X"8D",X"28",X"8E",X"F7",
		X"95",X"A6",X"80",X"BF",X"BF",X"06",X"8D",X"65",X"86",X"80",X"B7",X"BF",X"1F",X"4F",X"BD",X"F9",
		X"97",X"BD",X"F9",X"8A",X"25",X"0F",X"7A",X"BF",X"1F",X"26",X"F2",X"BE",X"BF",X"06",X"8C",X"F7",
		X"9D",X"25",X"DE",X"20",X"D9",X"39",X"8E",X"00",X"00",X"10",X"8E",X"F7",X"9D",X"BF",X"BF",X"06",
		X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"C6",X"39",X"F7",X"CB",X"FF",X"BC",
		X"BF",X"06",X"26",X"F2",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"10",X"8C",
		X"F7",X"AD",X"26",X"D9",X"39",X"02",X"03",X"04",X"10",X"18",X"20",X"40",X"80",X"00",X"FF",X"11",
		X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",X"8E",X"C0",X"00",
		X"A7",X"80",X"8C",X"C0",X"10",X"25",X"F9",X"39",X"86",X"0A",X"B7",X"BF",X"06",X"BD",X"32",X"45",
		X"86",X"06",X"BD",X"E2",X"12",X"C6",X"39",X"F7",X"CB",X"FF",X"CE",X"BF",X"1F",X"6F",X"C0",X"11",
		X"83",X"BF",X"28",X"23",X"F8",X"CE",X"F8",X"99",X"8D",X"29",X"86",X"34",X"B7",X"C8",X"07",X"C6",
		X"39",X"F7",X"CB",X"FF",X"8D",X"1D",X"86",X"3C",X"B7",X"C8",X"07",X"8D",X"26",X"BD",X"F9",X"8A",
		X"24",X"0A",X"C6",X"39",X"F7",X"CB",X"FF",X"7A",X"BF",X"06",X"27",X"06",X"4F",X"BD",X"F9",X"97",
		X"20",X"D3",X"39",X"AE",X"C1",X"27",X"0B",X"10",X"AE",X"C1",X"A6",X"84",X"A8",X"A4",X"A7",X"21",
		X"20",X"F1",X"39",X"CE",X"F8",X"B1",X"10",X"8E",X"BF",X"1F",X"C6",X"01",X"E5",X"21",X"27",X"02",
		X"8D",X"15",X"33",X"43",X"58",X"24",X"F5",X"C6",X"39",X"F7",X"CB",X"FF",X"31",X"22",X"10",X"8C",
		X"BF",X"28",X"22",X"02",X"20",X"E4",X"39",X"34",X"14",X"86",X"3F",X"B7",X"C8",X"0E",X"E8",X"A4",
		X"E7",X"A4",X"E6",X"E4",X"E5",X"A4",X"26",X"2A",X"A6",X"42",X"27",X"4B",X"C6",X"60",X"1F",X"01",
		X"C6",X"39",X"F7",X"CB",X"FF",X"CC",X"07",X"84",X"FD",X"CA",X"06",X"BF",X"CA",X"04",X"BF",X"CA",
		X"04",X"C6",X"00",X"F7",X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",X"C6",X"39",X"F7",X"CB",X"FF",
		X"35",X"94",X"A6",X"42",X"27",X"21",X"C6",X"60",X"1F",X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",
		X"BB",X"A6",X"C4",X"BD",X"E2",X"0C",X"A6",X"41",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"BD",
		X"E2",X"0F",X"86",X"38",X"B7",X"C8",X"0E",X"35",X"94",X"C8",X"0C",X"BF",X"1F",X"C8",X"04",X"BF",
		X"21",X"C8",X"06",X"BF",X"23",X"00",X"00",X"C8",X"04",X"BF",X"25",X"C8",X"06",X"BF",X"27",X"00",
		X"00",X"11",X"FF",X"74",X"12",X"FF",X"71",X"13",X"FF",X"6E",X"14",X"FF",X"6B",X"15",X"FF",X"68",
		X"16",X"FF",X"65",X"17",X"FF",X"62",X"00",X"00",X"00",X"1A",X"F2",X"3B",X"1B",X"F2",X"38",X"1C",
		X"F2",X"35",X"1D",X"F2",X"32",X"1E",X"F2",X"2F",X"1F",X"F2",X"2C",X"20",X"F2",X"29",X"21",X"F2",
		X"26",X"22",X"F2",X"23",X"23",X"F2",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"FF",X"41",
		X"19",X"FF",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"F1",X"5F",X"1B",X"F1",X"5C",X"1C",
		X"F1",X"59",X"1D",X"F1",X"56",X"1E",X"F1",X"53",X"1F",X"F1",X"50",X"20",X"F1",X"4D",X"21",X"F1",
		X"4A",X"22",X"F1",X"47",X"23",X"F1",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F4",X"01",X"20",X"03",X"CE",X"F3",
		X"DD",X"10",X"CE",X"BF",X"00",X"10",X"8E",X"F9",X"3E",X"86",X"01",X"7E",X"F1",X"FD",X"B6",X"C8",
		X"0C",X"85",X"02",X"26",X"F0",X"10",X"8E",X"F9",X"4E",X"86",X"01",X"7E",X"F1",X"FD",X"B6",X"C8",
		X"0C",X"85",X"02",X"27",X"F0",X"10",X"8E",X"F9",X"5E",X"86",X"01",X"7E",X"F1",X"FD",X"B6",X"C8",
		X"0C",X"85",X"02",X"26",X"F0",X"6E",X"C4",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"06",X"86",X"01",
		X"8D",X"25",X"20",X"F3",X"7F",X"C0",X"00",X"BD",X"32",X"45",X"20",X"07",X"B6",X"C8",X"0C",X"85",
		X"02",X"27",X"06",X"86",X"01",X"8D",X"10",X"20",X"F3",X"39",X"B6",X"C8",X"0C",X"85",X"02",X"27",
		X"03",X"1A",X"01",X"39",X"1C",X"FE",X"39",X"C6",X"39",X"8E",X"03",X"00",X"F7",X"CB",X"FF",X"30",
		X"1F",X"26",X"F9",X"4A",X"2A",X"F1",X"39",X"86",X"BF",X"1F",X"8B",X"BD",X"F4",X"90",X"8D",X"DA",
		X"24",X"02",X"8D",X"B3",X"86",X"07",X"BD",X"E2",X"12",X"CE",X"CD",X"02",X"8E",X"6F",X"18",X"86",
		X"26",X"34",X"12",X"C6",X"88",X"BD",X"E2",X"03",X"1E",X"31",X"BD",X"4A",X"70",X"C5",X"F0",X"26",
		X"08",X"CA",X"F0",X"C5",X"0F",X"26",X"02",X"CA",X"0F",X"1F",X"98",X"43",X"34",X"06",X"BD",X"4A",
		X"6E",X"6D",X"E0",X"26",X"12",X"85",X"F0",X"26",X"0E",X"8A",X"F0",X"85",X"0F",X"26",X"08",X"8A",
		X"0F",X"C5",X"F0",X"26",X"02",X"CA",X"F0",X"1F",X"02",X"1E",X"31",X"1F",X"10",X"C6",X"B8",X"1F",
		X"01",X"35",X"02",X"C6",X"88",X"BD",X"E2",X"06",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"20",X"34",
		X"04",X"C6",X"88",X"BD",X"E2",X"06",X"35",X"02",X"BD",X"E2",X"06",X"86",X"39",X"B7",X"CB",X"FF",
		X"35",X"12",X"30",X"89",X"F6",X"00",X"4C",X"11",X"83",X"CD",X"2C",X"23",X"94",X"86",X"2E",X"C6",
		X"88",X"BD",X"E2",X"03",X"1F",X"10",X"C6",X"C2",X"1F",X"01",X"1E",X"31",X"8E",X"CD",X"20",X"BD",
		X"4A",X"70",X"F7",X"BF",X"10",X"BD",X"4A",X"6E",X"FD",X"BF",X"11",X"8E",X"CD",X"2C",X"BD",X"4A",
		X"70",X"F7",X"BF",X"13",X"BD",X"4A",X"6E",X"FD",X"BF",X"14",X"1E",X"31",X"8D",X"21",X"C6",X"88",
		X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",X"E2",X"06",X"86",X"32",X"BD",X"E2",X"00",X"B6",X"BF",
		X"12",X"BD",X"E2",X"06",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"F9",X"67",X"7E",X"FB",X"80",X"34",
		X"30",X"8D",X"7A",X"FC",X"BF",X"10",X"27",X"0F",X"86",X"99",X"34",X"02",X"B7",X"BF",X"12",X"7F",
		X"BF",X"11",X"7F",X"BF",X"10",X"20",X"4C",X"B6",X"BF",X"12",X"34",X"02",X"FC",X"BF",X"0D",X"FD",
		X"BF",X"10",X"B6",X"BF",X"0F",X"B7",X"BF",X"12",X"CC",X"00",X"00",X"FD",X"BF",X"0D",X"B7",X"BF",
		X"0F",X"86",X"04",X"78",X"BF",X"12",X"79",X"BF",X"11",X"79",X"BF",X"10",X"79",X"BF",X"0F",X"4A",
		X"26",X"F1",X"8E",X"BF",X"13",X"10",X"8E",X"BF",X"13",X"CE",X"BF",X"13",X"8D",X"17",X"FC",X"BF",
		X"0F",X"FD",X"BF",X"16",X"FC",X"BF",X"11",X"FD",X"BF",X"18",X"8E",X"BF",X"1A",X"8D",X"06",X"8D",
		X"04",X"8D",X"23",X"35",X"B2",X"34",X"70",X"C6",X"04",X"20",X"04",X"34",X"70",X"C6",X"03",X"1C",
		X"FE",X"A6",X"82",X"A9",X"A2",X"19",X"A7",X"C2",X"5A",X"26",X"F6",X"35",X"F0",X"CC",X"00",X"00",
		X"FD",X"BF",X"0D",X"B7",X"BF",X"0F",X"FC",X"BF",X"13",X"26",X"0F",X"B6",X"BF",X"15",X"26",X"0A",
		X"CC",X"00",X"00",X"FD",X"BF",X"10",X"B7",X"BF",X"12",X"39",X"86",X"07",X"B7",X"BF",X"16",X"8E",
		X"BF",X"10",X"10",X"8E",X"BF",X"16",X"CE",X"BF",X"1A",X"8D",X"35",X"7A",X"BF",X"16",X"26",X"02",
		X"20",X"2E",X"86",X"04",X"78",X"BF",X"12",X"79",X"BF",X"11",X"79",X"BF",X"10",X"79",X"BF",X"0F",
		X"79",X"BF",X"0E",X"79",X"BF",X"0D",X"4A",X"26",X"EB",X"8D",X"A0",X"25",X"02",X"20",X"DC",X"FC",
		X"BF",X"17",X"FD",X"BF",X"0D",X"B6",X"BF",X"19",X"B7",X"BF",X"0F",X"7C",X"BF",X"12",X"20",X"E9",
		X"34",X"20",X"C6",X"03",X"86",X"99",X"A0",X"A2",X"A7",X"A4",X"5A",X"26",X"F7",X"10",X"AE",X"E4",
		X"C6",X"03",X"1A",X"01",X"A6",X"3F",X"89",X"00",X"19",X"A7",X"A2",X"5A",X"26",X"F6",X"35",X"A0",
		X"8E",X"CC",X"1A",X"6F",X"80",X"8C",X"CC",X"24",X"25",X"F9",X"BD",X"32",X"45",X"BD",X"F9",X"8A",
		X"24",X"03",X"BD",X"F9",X"67",X"86",X"08",X"BD",X"E2",X"12",X"CE",X"CC",X"00",X"8E",X"78",X"20",
		X"86",X"30",X"34",X"12",X"C6",X"22",X"BD",X"E2",X"0C",X"F7",X"BF",X"1A",X"F7",X"BF",X"0D",X"1F",
		X"12",X"BD",X"FD",X"60",X"33",X"42",X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"12",X"30",X"89",X"FB",
		X"00",X"4C",X"11",X"83",X"CC",X"24",X"2D",X"DA",X"86",X"09",X"BD",X"E2",X"15",X"7F",X"BF",X"0D",
		X"B6",X"CC",X"0D",X"84",X"0F",X"81",X"09",X"26",X"0B",X"86",X"4C",X"F6",X"BF",X"1A",X"8E",X"5A",
		X"98",X"BD",X"E2",X"0C",X"10",X"8E",X"78",X"18",X"CE",X"CC",X"00",X"1F",X"21",X"86",X"30",X"C6",
		X"33",X"FD",X"BF",X"1F",X"BD",X"E2",X"09",X"86",X"39",X"B7",X"CB",X"FF",X"C6",X"34",X"F7",X"C8",
		X"07",X"BD",X"48",X"F3",X"84",X"03",X"27",X"02",X"8D",X"1A",X"BD",X"48",X"F3",X"84",X"30",X"27",
		X"03",X"BD",X"FC",X"BD",X"C6",X"3C",X"F7",X"C8",X"07",X"BD",X"F9",X"8A",X"24",X"D9",X"BD",X"F9",
		X"67",X"7E",X"49",X"4C",X"B7",X"BF",X"23",X"B1",X"BF",X"21",X"27",X"15",X"7F",X"BF",X"22",X"B6",
		X"BF",X"23",X"B7",X"BF",X"21",X"86",X"02",X"BD",X"F9",X"97",X"BD",X"48",X"F3",X"84",X"03",X"26",
		X"1D",X"C6",X"05",X"F7",X"BF",X"24",X"BD",X"48",X"F3",X"84",X"03",X"26",X"04",X"7F",X"BF",X"21",
		X"39",X"86",X"02",X"BD",X"F9",X"97",X"7A",X"BF",X"24",X"26",X"EB",X"BD",X"48",X"F3",X"85",X"02",
		X"26",X"25",X"85",X"01",X"27",X"48",X"10",X"8C",X"78",X"18",X"27",X"42",X"8D",X"45",X"31",X"A9",
		X"05",X"00",X"33",X"5E",X"11",X"83",X"CC",X"18",X"26",X"0B",X"7D",X"BF",X"0A",X"27",X"06",X"31",
		X"A9",X"1E",X"00",X"33",X"54",X"20",X"1F",X"10",X"8C",X"23",X"18",X"27",X"21",X"8D",X"24",X"31",
		X"A9",X"FB",X"00",X"33",X"42",X"11",X"83",X"CC",X"0E",X"26",X"0B",X"7D",X"BF",X"0A",X"27",X"06",
		X"31",X"A9",X"E2",X"00",X"33",X"4C",X"1F",X"21",X"FC",X"BF",X"1F",X"BD",X"E2",X"09",X"4F",X"BD",
		X"F9",X"97",X"39",X"1F",X"21",X"B6",X"BF",X"1F",X"5F",X"BD",X"E2",X"09",X"39",X"B7",X"BF",X"23",
		X"B1",X"BF",X"25",X"27",X"15",X"7F",X"BF",X"26",X"B6",X"BF",X"23",X"B7",X"BF",X"25",X"86",X"02",
		X"BD",X"F9",X"97",X"BD",X"48",X"F3",X"84",X"30",X"26",X"1E",X"C6",X"08",X"F7",X"BF",X"28",X"BD",
		X"48",X"F3",X"84",X"30",X"26",X"04",X"7F",X"BF",X"26",X"39",X"4F",X"BD",X"F9",X"97",X"7A",X"BF",
		X"28",X"26",X"EC",X"BD",X"48",X"F3",X"84",X"30",X"34",X"02",X"1F",X"31",X"BD",X"4A",X"5F",X"34",
		X"02",X"7F",X"BF",X"1A",X"8D",X"5A",X"C6",X"39",X"F7",X"CB",X"FF",X"8E",X"FD",X"3C",X"1F",X"30",
		X"30",X"85",X"35",X"06",X"C5",X"10",X"26",X"0C",X"C5",X"20",X"27",X"14",X"A1",X"84",X"27",X"10",
		X"8B",X"99",X"20",X"06",X"A1",X"01",X"27",X"08",X"8B",X"01",X"19",X"1F",X"31",X"BD",X"4A",X"78",
		X"C6",X"22",X"F7",X"BF",X"1A",X"BD",X"FD",X"60",X"4F",X"7E",X"F9",X"97",X"01",X"99",X"00",X"99",
		X"01",X"99",X"00",X"09",X"00",X"01",X"00",X"01",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"99",
		X"01",X"99",X"00",X"99",X"00",X"99",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",
		X"1F",X"30",X"54",X"8E",X"FD",X"C1",X"30",X"85",X"6D",X"84",X"2B",X"2C",X"1F",X"31",X"BD",X"4A",
		X"5F",X"11",X"83",X"CC",X"0C",X"26",X"0A",X"B7",X"BF",X"0A",X"7D",X"BF",X"0D",X"26",X"02",X"8D",
		X"52",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"34",X"02",X"1F",X"20",X"C6",X"C4",X"1F",X"01",X"35",
		X"02",X"F6",X"BF",X"1A",X"BD",X"E2",X"0F",X"39",X"A6",X"84",X"85",X"01",X"26",X"1C",X"1F",X"31",
		X"BD",X"4A",X"70",X"86",X"08",X"5D",X"27",X"02",X"86",X"44",X"34",X"02",X"1F",X"20",X"C6",X"C4",
		X"1F",X"01",X"35",X"02",X"F6",X"BF",X"1A",X"7E",X"E2",X"0C",X"8D",X"B0",X"86",X"2F",X"7E",X"E2",
		X"09",X"81",X"81",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"80",X"80",X"80",X"34",X"76",X"8E",X"FE",X"30",X"81",X"09",X"26",X"0F",X"34",X"12",X"86",X"4C",
		X"F6",X"BF",X"1A",X"8E",X"5A",X"98",X"BD",X"E2",X"0C",X"35",X"12",X"1F",X"89",X"58",X"34",X"04",
		X"58",X"EB",X"E0",X"3A",X"33",X"42",X"1E",X"31",X"8C",X"CC",X"1A",X"27",X"31",X"A6",X"C0",X"BD",
		X"4A",X"78",X"C6",X"39",X"F7",X"CB",X"FF",X"1E",X"31",X"31",X"A9",X"FB",X"00",X"34",X"10",X"30",
		X"5E",X"BD",X"4A",X"5F",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"34",X"02",X"1F",X"20",X"C6",X"C4",
		X"1F",X"01",X"35",X"02",X"F6",X"BF",X"1A",X"BD",X"E2",X"0F",X"35",X"10",X"20",X"C8",X"35",X"F6",
		X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",
		X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",
		X"01",X"02",X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",
		X"01",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"32",X"45",X"CC",
		X"FE",X"01",X"FD",X"BF",X"20",X"39",X"34",X"10",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",
		X"F9",X"97",X"4F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"97",X"86",X"3F",X"B7",X"C8",X"0E",
		X"86",X"03",X"BD",X"F9",X"97",X"FC",X"BF",X"20",X"84",X"3F",X"B7",X"C8",X"0E",X"C6",X"99",X"8E",
		X"4C",X"54",X"86",X"24",X"BD",X"E2",X"03",X"AF",X"E4",X"B6",X"BF",X"21",X"8A",X"F0",X"C6",X"99",
		X"BD",X"E2",X"06",X"86",X"40",X"B7",X"BF",X"1F",X"86",X"01",X"BD",X"F9",X"97",X"BD",X"F9",X"8A",
		X"25",X"05",X"7A",X"BF",X"1F",X"26",X"F1",X"B6",X"BF",X"08",X"26",X"06",X"B6",X"C8",X"0C",X"46",
		X"24",X"1C",X"AE",X"E4",X"B6",X"BF",X"21",X"8A",X"F0",X"C6",X"00",X"BD",X"E2",X"06",X"FC",X"BF",
		X"20",X"1A",X"01",X"49",X"7E",X"FF",X"D0",X"25",X"02",X"8D",X"84",X"FD",X"BF",X"20",X"35",X"90",
		X"8E",X"CC",X"00",X"10",X"8E",X"9C",X"00",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",
		X"C6",X"06",X"FE",X"BF",X"0B",X"10",X"BE",X"BF",X"0A",X"8E",X"CC",X"00",X"BD",X"FF",X"57",X"A7",
		X"80",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"F1",X"10",X"BF",X"BF",X"0A",X"FF",
		X"BF",X"0B",X"8E",X"CC",X"00",X"BD",X"FF",X"57",X"A8",X"80",X"84",X"0F",X"26",X"24",X"86",X"39",
		X"B7",X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"ED",X"5A",X"26",X"C7",X"8D",X"03",X"1C",X"FE",X"39",
		X"CE",X"9C",X"00",X"10",X"8E",X"CC",X"00",X"A6",X"C0",X"A7",X"A0",X"10",X"8C",X"D0",X"00",X"26",
		X"F6",X"39",X"8D",X"EC",X"1A",X"01",X"39",X"34",X"04",X"F6",X"BF",X"0A",X"86",X"03",X"3D",X"CB",
		X"11",X"B6",X"BF",X"0C",X"44",X"44",X"44",X"B8",X"BF",X"0C",X"44",X"76",X"BF",X"0B",X"76",X"BF",
		X"0C",X"FB",X"BF",X"0C",X"F9",X"BF",X"0B",X"F7",X"BF",X"0A",X"B6",X"BF",X"0A",X"35",X"84",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"20",X"57",X"49",
		X"34",X"10",X"BD",X"46",X"DB",X"FF",X"A1",X"05",X"A1",X"6D",X"6F",X"04",X"35",X"10",X"7E",X"7C",
		X"6D",X"6A",X"24",X"26",X"02",X"0F",X"95",X"EC",X"3E",X"DD",X"42",X"39",X"00",X"00",X"00",X"00",
		X"CC",X"38",X"7A",X"ED",X"25",X"E7",X"27",X"6F",X"A8",X"10",X"6E",X"B8",X"1A",X"00",X"00",X"00",
		X"7F",X"C0",X"00",X"7F",X"CA",X"01",X"BD",X"32",X"45",X"7E",X"F0",X"82",X"00",X"00",X"00",X"00",
		X"5C",X"C1",X"03",X"26",X"03",X"7E",X"FE",X"E1",X"C1",X"06",X"7E",X"FE",X"E7",X"00",X"00",X"DA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"1F",X"F0",X"1F",X"F0",X"1F",X"F0",X"1F",X"E0",X"0B",X"F0",X"1F",X"F0",X"1F",X"F0",X"1F",
		X"00",X"00",X"7E",X"2E",X"45",X"00",X"FF",X"06",X"09",X"01",X"07",X"01",X"3D",X"05",X"04",X"06",
		X"09",X"01",X"4F",X"01",X"85",X"05",X"04",X"06",X"0A",X"01",X"97",X"01",X"D3",X"05",X"04",X"06",
		X"0A",X"01",X"E7",X"02",X"23",X"05",X"05",X"06",X"0A",X"02",X"37",X"02",X"73",X"05",X"04",X"05",
		X"0B",X"02",X"87",X"02",X"BE",X"05",X"04",X"06",X"0B",X"02",X"D4",X"03",X"16",X"05",X"04",X"05",
		X"0B",X"03",X"2C",X"03",X"63",X"04",X"03",X"05",X"0B",X"03",X"79",X"03",X"B0",X"04",X"03",X"05",
		X"0B",X"03",X"C6",X"03",X"FD",X"04",X"03",X"06",X"0B",X"04",X"13",X"04",X"55",X"04",X"03",X"05",
		X"0A",X"04",X"6B",X"04",X"9D",X"03",X"03",X"06",X"0A",X"04",X"B1",X"04",X"ED",X"04",X"03",X"06",
		X"09",X"05",X"01",X"05",X"37",X"04",X"03",X"06",X"0A",X"05",X"49",X"05",X"85",X"05",X"03",X"06",
		X"0A",X"05",X"99",X"05",X"D5",X"05",X"03",X"06",X"09",X"05",X"E7",X"06",X"1D",X"05",X"03",X"06",
		X"09",X"06",X"2F",X"06",X"65",X"05",X"03",X"06",X"0A",X"06",X"77",X"06",X"B3",X"05",X"03",X"06",
		X"09",X"06",X"C7",X"06",X"FD",X"05",X"02",X"06",X"0A",X"07",X"0F",X"07",X"4B",X"04",X"03",X"05",
		X"0B",X"07",X"5F",X"07",X"96",X"03",X"04",X"06",X"0B",X"07",X"AC",X"07",X"EE",X"04",X"04",X"05",
		X"0A",X"08",X"04",X"08",X"36",X"04",X"04",X"05",X"0B",X"08",X"4A",X"08",X"81",X"04",X"04",X"05",
		X"0B",X"08",X"97",X"08",X"CE",X"04",X"04",X"06",X"0B",X"08",X"E4",X"09",X"26",X"06",X"04",X"06",
		X"0B",X"09",X"3C",X"09",X"7E",X"06",X"04",X"06",X"0A",X"09",X"94",X"09",X"D0",X"05",X"03",X"06",
		X"0A",X"09",X"E4",X"0A",X"20",X"05",X"02",X"06",X"0B",X"0A",X"34",X"0A",X"76",X"05",X"03",X"06",
		X"09",X"0A",X"8C",X"0A",X"C2",X"05",X"03",X"0A",X"55",X"A0",X"00",X"00",X"00",X"0A",X"41",X"2A",
		X"00",X"00",X"00",X"0A",X"42",X"12",X"A0",X"00",X"00",X"A5",X"54",X"21",X"14",X"A0",X"00",X"65",
		X"11",X"11",X"22",X"44",X"A0",X"A6",X"55",X"55",X"55",X"A0",X"00",X"0A",X"66",X"55",X"A0",X"00",
		X"00",X"0A",X"54",X"5A",X"00",X"00",X"00",X"0A",X"56",X"A0",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"01",X"01",X"01",X"05",X"06",X"07",X"09",X"0A",X"09",X"07",X"06",X"05",X"00",
		X"A5",X"A0",X"00",X"00",X"00",X"00",X"A4",X"1A",X"00",X"00",X"00",X"00",X"A4",X"21",X"A0",X"00",
		X"00",X"0A",X"45",X"42",X"1A",X"00",X"00",X"A4",X"42",X"11",X"22",X"4A",X"00",X"06",X"44",X"22",
		X"21",X"14",X"60",X"0A",X"65",X"54",X"45",X"AA",X"A0",X"0A",X"54",X"45",X"A0",X"00",X"00",X"06",
		X"56",X"A0",X"00",X"00",X"00",X"02",X"02",X"02",X"01",X"00",X"01",X"01",X"01",X"01",X"05",X"06",
		X"07",X"08",X"0A",X"0B",X"0B",X"07",X"05",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"06",X"64",
		X"A0",X"00",X"00",X"00",X"A6",X"54",X"4A",X"00",X"00",X"06",X"54",X"45",X"46",X"00",X"00",X"06",
		X"44",X"22",X"25",X"A0",X"00",X"0A",X"44",X"41",X"22",X"4A",X"00",X"0A",X"66",X"44",X"41",X"15",
		X"00",X"0A",X"56",X"66",X"55",X"54",X"60",X"A6",X"54",X"66",X"A0",X"00",X"00",X"0A",X"AA",X"A0",
		X"00",X"00",X"00",X"03",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"05",X"07",X"08",
		X"08",X"09",X"0A",X"0A",X"0B",X"07",X"05",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"A6",
		X"A0",X"00",X"00",X"00",X"AA",X"A5",X"4A",X"00",X"00",X"0A",X"64",X"45",X"46",X"00",X"00",X"0A",
		X"52",X"24",X"46",X"A0",X"00",X"0A",X"54",X"12",X"24",X"A0",X"00",X"0A",X"65",X"41",X"22",X"60",
		X"00",X"A6",X"56",X"65",X"41",X"5A",X"00",X"A5",X"44",X"56",X"66",X"46",X"00",X"0A",X"AA",X"A0",
		X"00",X"0A",X"A0",X"05",X"04",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"06",X"07",X"08",
		X"08",X"09",X"09",X"09",X"0A",X"0A",X"0B",X"00",X"00",X"0A",X"60",X"00",X"00",X"00",X"AA",X"A5",
		X"56",X"00",X"00",X"0A",X"64",X"42",X"25",X"00",X"00",X"0A",X"51",X"24",X"25",X"A0",X"00",X"06",
		X"54",X"12",X"44",X"A0",X"00",X"A5",X"65",X"41",X"24",X"A0",X"00",X"65",X"56",X"54",X"12",X"60",
		X"00",X"06",X"65",X"55",X"41",X"50",X"00",X"00",X"00",X"AA",X"65",X"1A",X"00",X"00",X"00",X"00",
		X"00",X"A6",X"00",X"05",X"02",X"01",X"01",X"01",X"00",X"00",X"01",X"04",X"08",X"07",X"08",X"08",
		X"09",X"09",X"09",X"09",X"09",X"0A",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"A6",X"6A",X"55",
		X"A0",X"00",X"64",X"44",X"42",X"00",X"0A",X"54",X"14",X"42",X"A0",X"AA",X"65",X"12",X"44",X"A0",
		X"64",X"65",X"41",X"24",X"A0",X"A6",X"66",X"44",X"25",X"00",X"00",X"A6",X"64",X"14",X"00",X"00",
		X"00",X"A6",X"64",X"A0",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",X"00",X"00",X"A0",X"06",X"02",
		X"02",X"01",X"00",X"00",X"00",X"02",X"04",X"06",X"08",X"08",X"09",X"08",X"09",X"09",X"09",X"08",
		X"08",X"09",X"09",X"09",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"06",X"6A",X"A6",X"6A",X"00",
		X"00",X"A5",X"24",X"65",X"4A",X"00",X"0A",X"A5",X"22",X"42",X"4A",X"00",X"A6",X"55",X"41",X"24",
		X"5A",X"00",X"05",X"55",X"42",X"24",X"60",X"00",X"0A",X"65",X"54",X"15",X"A0",X"00",X"00",X"A6",
		X"54",X"25",X"00",X"00",X"00",X"00",X"A6",X"46",X"00",X"00",X"00",X"00",X"00",X"65",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"08",X"03",X"02",X"01",X"00",X"01",X"01",X"02",X"04",X"06",
		X"07",X"09",X"0A",X"0A",X"0A",X"0A",X"09",X"09",X"08",X"08",X"08",X"08",X"00",X"00",X"6A",X"00",
		X"00",X"00",X"0A",X"44",X"AA",X"60",X"AA",X"A5",X"42",X"51",X"10",X"65",X"56",X"21",X"41",X"20",
		X"64",X"46",X"21",X"21",X"A0",X"A6",X"55",X"42",X"44",X"00",X"00",X"A5",X"52",X"4A",X"00",X"00",
		X"0A",X"54",X"50",X"00",X"00",X"00",X"64",X"A0",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"04",X"03",X"00",X"00",X"00",X"00",X"02",X"03",X"04",X"05",X"05",X"06",X"09",
		X"09",X"09",X"09",X"08",X"08",X"07",X"07",X"06",X"06",X"00",X"0A",X"6A",X"00",X"00",X"AA",X"A5",
		X"26",X"AA",X"A0",X"55",X"65",X"12",X"21",X"40",X"64",X"65",X"12",X"22",X"50",X"A5",X"55",X"14",
		X"44",X"A0",X"0A",X"55",X"14",X"4A",X"00",X"00",X"A5",X"25",X"A0",X"00",X"00",X"05",X"45",X"00",
		X"00",X"00",X"0A",X"5A",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"03",X"04",X"04",X"06",X"09",X"09",X"09",X"09",
		X"08",X"07",X"06",X"06",X"05",X"05",X"00",X"0A",X"60",X"00",X"00",X"6A",X"A5",X"1A",X"00",X"00",
		X"52",X"54",X"14",X"AA",X"A0",X"54",X"54",X"14",X"12",X"60",X"A5",X"52",X"24",X"24",X"A0",X"05",
		X"52",X"24",X"4A",X"00",X"0A",X"62",X"45",X"A0",X"00",X"00",X"64",X"56",X"00",X"00",X"00",X"A4",
		X"60",X"00",X"00",X"00",X"A5",X"A0",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"02",X"05",X"06",X"09",X"09",X"09",X"08",X"07",X"06",
		X"05",X"05",X"04",X"0A",X"00",X"00",X"00",X"00",X"00",X"06",X"AA",X"A6",X"6A",X"00",X"00",X"A2",
		X"26",X"24",X"5A",X"00",X"00",X"A4",X"24",X"21",X"46",X"AA",X"00",X"A4",X"44",X"12",X"45",X"6A",
		X"00",X"06",X"44",X"14",X"44",X"50",X"00",X"0A",X"64",X"44",X"46",X"A0",X"00",X"00",X"54",X"55",
		X"6A",X"00",X"00",X"00",X"64",X"6A",X"00",X"00",X"00",X"00",X"56",X"A0",X"00",X"00",X"00",X"00",
		X"6A",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"02",
		X"02",X"08",X"08",X"0A",X"0A",X"09",X"09",X"08",X"06",X"05",X"04",X"0A",X"A0",X"00",X"00",X"00",
		X"A5",X"6A",X"66",X"A0",X"00",X"A2",X"55",X"41",X"6A",X"00",X"A2",X"54",X"22",X"4A",X"00",X"A4",
		X"44",X"14",X"46",X"A0",X"A6",X"52",X"44",X"42",X"60",X"06",X"44",X"54",X"46",X"00",X"06",X"45",
		X"6A",X"A0",X"00",X"04",X"6A",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"03",X"07",X"08",X"08",X"09",X"09",X"08",X"07",X"04",
		X"03",X"00",X"06",X"A0",X"00",X"00",X"00",X"00",X"64",X"6A",X"AA",X"00",X"00",X"00",X"54",X"44",
		X"46",X"A0",X"00",X"0A",X"54",X"42",X"12",X"A0",X"00",X"0A",X"54",X"21",X"24",X"A0",X"00",X"0A",
		X"54",X"12",X"44",X"6A",X"00",X"06",X"52",X"44",X"54",X"47",X"00",X"06",X"45",X"55",X"55",X"60",
		X"00",X"A5",X"66",X"AA",X"A0",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"02",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"05",X"08",X"09",X"09",X"09",X"0A",X"0A",X"09",X"07",
		X"02",X"00",X"00",X"6A",X"00",X"00",X"00",X"00",X"06",X"26",X"AA",X"00",X"00",X"00",X"A4",X"44",
		X"46",X"A0",X"00",X"00",X"A4",X"44",X"21",X"60",X"00",X"00",X"65",X"31",X"23",X"60",X"00",X"0A",
		X"54",X"23",X"35",X"A0",X"00",X"A6",X"33",X"53",X"55",X"6A",X"00",X"63",X"66",X"63",X"22",X"5A",
		X"00",X"A0",X"00",X"AA",X"AA",X"A0",X"00",X"04",X"03",X"02",X"02",X"02",X"01",X"00",X"00",X"00",
		X"06",X"08",X"09",X"09",X"09",X"09",X"0A",X"0A",X"09",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"A5",X"6A",X"00",X"00",X"00",X"0A",X"64",X"56",X"AA",X"00",X"00",X"06",X"44",X"44",X"56",
		X"00",X"00",X"A5",X"44",X"21",X"46",X"00",X"0A",X"65",X"41",X"12",X"2A",X"00",X"A6",X"44",X"44",
		X"44",X"6A",X"00",X"65",X"65",X"54",X"42",X"2A",X"00",X"00",X"00",X"A6",X"54",X"26",X"00",X"00",
		X"00",X"00",X"AA",X"A0",X"00",X"06",X"04",X"03",X"03",X"02",X"01",X"00",X"00",X"04",X"06",X"08",
		X"08",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"09",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",
		X"00",X"06",X"44",X"A0",X"00",X"00",X"00",X"64",X"44",X"A0",X"00",X"00",X"A6",X"55",X"44",X"2A",
		X"00",X"0A",X"65",X"54",X"11",X"11",X"60",X"65",X"44",X"55",X"55",X"56",X"A0",X"AA",X"A6",X"66",
		X"55",X"5A",X"00",X"00",X"00",X"A5",X"54",X"4A",X"00",X"00",X"00",X"00",X"A5",X"56",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"05",X"04",X"02",X"01",X"00",X"00",X"04",X"06",X"09",X"09",
		X"09",X"0A",X"0B",X"0B",X"0A",X"0A",X"0A",X"00",X"00",X"00",X"A5",X"4A",X"00",X"00",X"00",X"0A",
		X"42",X"1A",X"00",X"00",X"00",X"A4",X"42",X"2A",X"00",X"00",X"A5",X"54",X"42",X"25",X"A0",X"A5",
		X"54",X"21",X"11",X"12",X"60",X"00",X"A5",X"55",X"55",X"55",X"A0",X"00",X"00",X"A5",X"56",X"6A",
		X"00",X"00",X"00",X"0A",X"54",X"5A",X"00",X"00",X"00",X"00",X"A6",X"5A",X"00",X"06",X"05",X"04",
		X"02",X"00",X"02",X"04",X"05",X"06",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0A",X"0A",X"0A",X"00",
		X"00",X"00",X"A2",X"16",X"00",X"00",X"00",X"A4",X"11",X"1A",X"00",X"00",X"A5",X"44",X"24",X"5A",
		X"00",X"65",X"44",X"22",X"11",X"24",X"A0",X"00",X"65",X"54",X"22",X"44",X"60",X"00",X"0A",X"55",
		X"66",X"5A",X"00",X"00",X"00",X"A5",X"45",X"A0",X"00",X"00",X"00",X"06",X"45",X"A0",X"00",X"00",
		X"00",X"0A",X"66",X"A0",X"00",X"06",X"04",X"02",X"00",X"02",X"03",X"04",X"05",X"05",X"0A",X"0A",
		X"0A",X"0B",X"0B",X"0A",X"09",X"09",X"09",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"A6",
		X"44",X"46",X"A0",X"65",X"65",X"54",X"42",X"56",X"00",X"06",X"42",X"12",X"24",X"6A",X"00",X"00",
		X"64",X"22",X"12",X"4A",X"00",X"00",X"A5",X"54",X"44",X"26",X"00",X"00",X"06",X"55",X"55",X"56",
		X"00",X"00",X"0A",X"65",X"5A",X"A0",X"00",X"00",X"00",X"A5",X"6A",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"06",X"04",X"00",X"01",X"02",X"02",X"03",X"03",X"04",X"06",X"0A",X"0B",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"09",X"08",X"07",X"AA",X"A0",X"0A",X"AA",X"6A",X"00",X"06",X"44",X"54",
		X"42",X"25",X"A0",X"0A",X"51",X"22",X"44",X"45",X"A0",X"00",X"64",X"41",X"24",X"4A",X"00",X"00",
		X"A6",X"44",X"11",X"46",X"00",X"00",X"06",X"65",X"54",X"46",X"00",X"00",X"0A",X"66",X"65",X"6A",
		X"00",X"00",X"00",X"65",X"AA",X"00",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",X"00",X"01",X"01",
		X"02",X"02",X"03",X"03",X"04",X"04",X"0A",X"0B",X"0B",X"0A",X"0A",X"0A",X"0A",X"08",X"07",X"6A",
		X"00",X"00",X"00",X"00",X"00",X"A1",X"56",X"AA",X"A0",X"00",X"00",X"05",X"12",X"44",X"55",X"60",
		X"00",X"06",X"41",X"24",X"22",X"56",X"00",X"06",X"54",X"12",X"42",X"5A",X"00",X"0A",X"55",X"41",
		X"24",X"A0",X"00",X"0A",X"56",X"54",X"14",X"A0",X"00",X"0A",X"65",X"65",X"56",X"A0",X"00",X"00",
		X"65",X"56",X"AA",X"00",X"00",X"00",X"06",X"A0",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"01",X"01",X"01",X"02",X"03",X"02",X"07",X"09",X"0A",X"0A",X"09",X"09",X"09",X"08",X"05",X"A0",
		X"00",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",X"00",X"04",X"56",X"A0",X"00",X"00",X"06",X"12",
		X"45",X"60",X"00",X"06",X"42",X"25",X"44",X"00",X"06",X"51",X"24",X"55",X"60",X"A5",X"64",X"12",
		X"4A",X"A0",X"A4",X"65",X"42",X"4A",X"00",X"A4",X"56",X"55",X"6A",X"00",X"A5",X"6A",X"A6",X"A0",
		X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"05",X"07",X"08",X"09",X"09",X"08",X"08",X"07",X"03",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"45",X"A0",X"00",X"00",X"00",X"00",X"51",X"4A",X"00",X"00",X"00",X"00",X"51",
		X"25",X"6A",X"00",X"00",X"0A",X"54",X"22",X"44",X"A0",X"00",X"06",X"64",X"12",X"54",X"40",X"00",
		X"A6",X"64",X"42",X"45",X"6A",X"00",X"A4",X"66",X"44",X"46",X"6A",X"00",X"A5",X"56",X"44",X"5A",
		X"00",X"00",X"A6",X"AA",X"A6",X"60",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"05",X"06",X"08",X"09",X"09",X"0A",
		X"0A",X"08",X"07",X"02",X"00",X"A6",X"00",X"00",X"00",X"00",X"A4",X"A0",X"00",X"00",X"00",X"A1",
		X"40",X"00",X"00",X"00",X"51",X"2A",X"00",X"00",X"0A",X"42",X"21",X"A0",X"00",X"05",X"42",X"12",
		X"1A",X"00",X"A4",X"52",X"14",X"21",X"A0",X"64",X"54",X"25",X"44",X"50",X"55",X"64",X"44",X"AA",
		X"A0",X"6A",X"A6",X"4A",X"00",X"00",X"02",X"02",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",
		X"04",X"05",X"05",X"06",X"07",X"08",X"09",X"09",X"09",X"06",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"0A",X"4A",X"00",X"00",X"00",X"05",X"24",X"00",X"00",X"00",X"A5",
		X"21",X"A0",X"00",X"0A",X"55",X"11",X"2A",X"00",X"A5",X"55",X"12",X"12",X"A0",X"64",X"65",X"14",
		X"21",X"50",X"55",X"65",X"15",X"44",X"50",X"AA",X"A6",X"55",X"AA",X"A0",X"00",X"0A",X"6A",X"00",
		X"00",X"04",X"04",X"03",X"03",X"02",X"01",X"00",X"00",X"00",X"00",X"03",X"05",X"05",X"06",X"06",
		X"07",X"08",X"09",X"09",X"09",X"09",X"06",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"A2",X"A0",
		X"00",X"00",X"00",X"51",X"A0",X"00",X"00",X"0A",X"41",X"40",X"00",X"00",X"A5",X"22",X"4A",X"00",
		X"0A",X"54",X"22",X"15",X"00",X"A4",X"45",X"22",X"21",X"A0",X"65",X"65",X"24",X"42",X"60",X"AA",
		X"A5",X"45",X"54",X"40",X"00",X"0A",X"46",X"AA",X"60",X"00",X"00",X"A0",X"00",X"00",X"05",X"04",
		X"04",X"03",X"02",X"01",X"00",X"00",X"00",X"03",X"04",X"06",X"07",X"07",X"07",X"08",X"08",X"09",
		X"09",X"09",X"09",X"05",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"06",X"50",X"00",
		X"00",X"00",X"0A",X"51",X"50",X"00",X"00",X"0A",X"A5",X"41",X"40",X"00",X"00",X"A6",X"42",X"21",
		X"5A",X"00",X"0A",X"64",X"52",X"12",X"46",X"00",X"AA",X"66",X"42",X"14",X"56",X"00",X"0A",X"A6",
		X"44",X"44",X"54",X"A0",X"00",X"0A",X"65",X"46",X"55",X"A0",X"00",X"0A",X"66",X"AA",X"A6",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"08",X"07",X"05",X"03",X"02",X"01",X"00",X"01",X"03",X"03",
		X"08",X"09",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0B",X"0B",X"0A",X"0A",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"0A",X"6A",X"00",X"00",X"00",X"0A",X"65",X"4A",X"00",X"00",X"AA",
		X"65",X"41",X"40",X"00",X"0A",X"62",X"44",X"22",X"50",X"00",X"A6",X"44",X"42",X"14",X"6A",X"00",
		X"0A",X"A5",X"41",X"24",X"4A",X"00",X"00",X"A5",X"44",X"45",X"4A",X"00",X"00",X"A6",X"55",X"56",
		X"2A",X"00",X"00",X"0A",X"66",X"A6",X"6A",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"09",X"07",
		X"05",X"02",X"01",X"00",X"01",X"02",X"02",X"03",X"07",X"0A",X"0A",X"0A",X"09",X"09",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"09",X"00",X"00",X"00",X"00",X"A6",X"00",X"00",X"0A",X"AA",X"65",X"1A",X"00",
		X"06",X"65",X"45",X"21",X"50",X"00",X"65",X"54",X"42",X"12",X"60",X"00",X"A6",X"54",X"21",X"25",
		X"60",X"00",X"0A",X"52",X"12",X"44",X"A0",X"00",X"0A",X"51",X"24",X"45",X"A0",X"00",X"0A",X"65",
		X"55",X"56",X"A0",X"00",X"00",X"AA",X"A6",X"56",X"00",X"00",X"00",X"00",X"0A",X"60",X"00",X"00",
		X"08",X"03",X"01",X"00",X"00",X"01",X"01",X"01",X"02",X"05",X"0A",X"0A",X"09",X"09",X"09",X"09",
		X"09",X"09",X"08",X"07",X"0A",X"AA",X"A0",X"00",X"AA",X"A0",X"A6",X"24",X"46",X"54",X"46",X"00",
		X"A6",X"65",X"44",X"21",X"5A",X"00",X"0A",X"54",X"21",X"24",X"60",X"00",X"06",X"54",X"12",X"45",
		X"A0",X"00",X"06",X"54",X"44",X"46",X"00",X"00",X"0A",X"65",X"54",X"2A",X"00",X"00",X"00",X"AA",
		X"A4",X"6A",X"00",X"00",X"00",X"00",X"A6",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"04",X"05",X"0B",X"0A",X"0A",X"09",X"09",X"08",
		X"08",X"08",X"07",X"06",X"00",X"AA",X"00",X"00",X"00",X"00",X"A6",X"66",X"66",X"A0",X"00",X"00",
		X"AA",X"55",X"54",X"54",X"55",X"60",X"0A",X"64",X"42",X"11",X"16",X"00",X"0A",X"44",X"11",X"24",
		X"50",X"00",X"06",X"54",X"22",X"25",X"A0",X"00",X"06",X"64",X"45",X"4A",X"00",X"00",X"0A",X"A6",
		X"64",X"6A",X"00",X"00",X"00",X"0A",X"66",X"A0",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"03",
		X"04",X"04",X"07",X"0B",X"0A",X"09",X"09",X"08",X"08",X"07",X"06",X"05",X"06",X"46",X"A0",X"00",
		X"00",X"00",X"0A",X"42",X"15",X"A0",X"00",X"00",X"0A",X"54",X"21",X"44",X"AA",X"00",X"06",X"54",
		X"22",X"21",X"12",X"60",X"A4",X"42",X"22",X"24",X"5A",X"00",X"0A",X"55",X"54",X"5A",X"00",X"00",
		X"00",X"A6",X"45",X"A0",X"00",X"00",X"00",X"A5",X"4A",X"00",X"00",X"00",X"00",X"A6",X"A0",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"01",X"02",X"02",X"02",X"05",X"07",X"0A",X"0B",X"0A",
		X"08",X"07",X"06",X"05",X"03",X"05",X"0A",X"F6",X"0A",X"EC",X"02",X"02",X"03",X"05",X"0B",X"05",
		X"0A",X"EC",X"02",X"02",X"03",X"05",X"0B",X"14",X"0A",X"EC",X"02",X"02",X"01",X"00",X"00",X"00",
		X"01",X"04",X"05",X"05",X"05",X"04",X"09",X"92",X"00",X"29",X"B9",X"90",X"9B",X"BB",X"90",X"99",
		X"B9",X"20",X"02",X"99",X"00",X"09",X"29",X"00",X"99",X"D9",X"90",X"2D",X"DD",X"20",X"99",X"D9",
		X"90",X"09",X"29",X"00",X"02",X"99",X"00",X"99",X"F9",X"20",X"9F",X"1F",X"90",X"29",X"F9",X"90",
		X"09",X"92",X"00",X"0E",X"1A",X"0B",X"2B",X"0C",X"97",X"0D",X"0D",X"00",X"00",X"00",X"00",X"0A",
		X"AA",X"65",X"45",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"5A",X"AA",X"6A",X"54",
		X"55",X"44",X"60",X"00",X"00",X"00",X"00",X"00",X"A6",X"55",X"45",X"45",X"4A",X"65",X"56",X"62",
		X"5A",X"00",X"00",X"00",X"00",X"00",X"55",X"66",X"66",X"55",X"56",X"A6",X"5A",X"65",X"4A",X"66",
		X"00",X"00",X"00",X"0A",X"64",X"54",X"55",X"54",X"44",X"6A",X"BA",X"65",X"46",X"54",X"56",X"00",
		X"00",X"0A",X"64",X"45",X"44",X"55",X"54",X"44",X"AB",X"45",X"55",X"44",X"45",X"00",X"00",X"0A",
		X"A6",X"55",X"45",X"66",X"55",X"55",X"5A",X"66",X"54",X"55",X"44",X"60",X"00",X"0A",X"A5",X"65",
		X"56",X"A6",X"65",X"55",X"45",X"A6",X"55",X"65",X"52",X"46",X"00",X"AB",X"AA",X"A6",X"66",X"AB",
		X"66",X"65",X"54",X"A6",X"66",X"65",X"54",X"46",X"00",X"AA",X"AA",X"AA",X"AB",X"AA",X"AA",X"A6",
		X"55",X"4A",X"65",X"66",X"54",X"4A",X"00",X"AB",X"AB",X"AA",X"AA",X"65",X"56",X"A6",X"54",X"44",
		X"45",X"65",X"54",X"6A",X"00",X"AA",X"AA",X"66",X"66",X"44",X"45",X"A6",X"55",X"55",X"54",X"65",
		X"55",X"6A",X"00",X"AA",X"BA",X"AA",X"55",X"45",X"45",X"AB",X"65",X"66",X"55",X"64",X"56",X"56",
		X"00",X"AA",X"AA",X"AA",X"65",X"56",X"54",X"AA",X"65",X"65",X"66",X"55",X"56",X"55",X"00",X"0A",
		X"AB",X"AA",X"A6",X"56",X"45",X"5A",X"66",X"55",X"44",X"45",X"66",X"45",X"00",X"0A",X"AA",X"AA",
		X"AA",X"BA",X"65",X"4A",X"AA",X"66",X"55",X"54",X"56",X"54",X"00",X"0A",X"AB",X"AA",X"AA",X"AA",
		X"A6",X"56",X"AA",X"A6",X"66",X"66",X"64",X"46",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",
		X"AA",X"AA",X"BA",X"B6",X"55",X"60",X"00",X"00",X"AA",X"BA",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",
		X"AA",X"65",X"44",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AB",X"AA",X"AA",X"AB",X"AA",X"64",
		X"56",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"BA",X"AA",X"66",X"60",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"AB",X"AA",X"AA",X"AB",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AB",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",
		X"AA",X"0A",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"04",X"02",X"02",X"01",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"05",X"06",X"07",
		X"09",X"11",X"13",X"14",X"16",X"18",X"18",X"19",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"1A",X"1A",X"19",X"18",X"18",X"17",X"16",X"15",X"13",X"12",X"0B",X"0D",X"18",X"0C",X"D3",X"0E",
		X"0B",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"56",X"44",X"66",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"A6",X"66",X"54",X"44",X"45",X"46",X"A0",X"00",X"00",X"00",X"00",X"0A",X"A5",X"44",X"46",
		X"55",X"45",X"56",X"54",X"46",X"A0",X"00",X"00",X"00",X"65",X"55",X"65",X"44",X"66",X"56",X"45",
		X"54",X"42",X"60",X"00",X"00",X"0A",X"55",X"65",X"66",X"54",X"6A",X"A6",X"54",X"65",X"54",X"4A",
		X"00",X"00",X"06",X"55",X"AB",X"AB",X"64",X"A6",X"55",X"44",X"56",X"A6",X"46",X"00",X"0A",X"6A",
		X"AB",X"AA",X"A6",X"A6",X"55",X"44",X"45",X"6A",X"64",X"46",X"00",X"06",X"AA",X"BA",X"AA",X"AA",
		X"55",X"45",X"44",X"56",X"56",X"54",X"55",X"00",X"0A",X"AA",X"AA",X"AA",X"A5",X"66",X"AA",X"65",
		X"44",X"5A",X"54",X"55",X"00",X"AA",X"AA",X"AA",X"AA",X"56",X"AA",X"AA",X"BA",X"64",X"6A",X"55",
		X"66",X"00",X"AA",X"AA",X"AA",X"AA",X"6B",X"AA",X"AA",X"AA",X"B5",X"A6",X"54",X"5A",X"00",X"AA",
		X"AA",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"65",X"54",X"6A",X"00",X"AA",X"BA",X"AA",X"BA",
		X"AA",X"AA",X"AA",X"AA",X"B5",X"55",X"44",X"5A",X"00",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AB",X"AA",X"65",X"64",X"5A",X"00",X"0A",X"AA",X"AA",X"BA",X"AA",X"AA",X"AB",X"AA",X"AA",X"56",
		X"66",X"60",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"60",X"00",
		X"0A",X"AA",X"AB",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"40",X"00",X"00",X"00",X"0A",X"AA",X"BA",X"AA",X"AA",
		X"AA",X"BA",X"AA",X"AA",X"50",X"00",X"00",X"00",X"00",X"00",X"AB",X"AA",X"AA",X"AA",X"AA",X"BA",
		X"B6",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"AB",X"AB",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0A",X"07",X"05",X"04",
		X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"03",X"06",
		X"06",X"07",X"0A",X"10",X"13",X"15",X"17",X"17",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",
		X"18",X"18",X"17",X"17",X"17",X"15",X"15",X"14",X"12",X"10",X"0E",X"0A",X"12",X"0E",X"43",X"0E",
		X"F7",X"09",X"09",X"00",X"00",X"0A",X"65",X"55",X"44",X"6A",X"00",X"00",X"00",X"00",X"A6",X"55",
		X"56",X"66",X"45",X"55",X"44",X"6A",X"00",X"00",X"55",X"56",X"65",X"45",X"65",X"66",X"54",X"44",
		X"00",X"05",X"56",X"65",X"44",X"45",X"56",X"65",X"54",X"55",X"00",X"06",X"66",X"AA",X"B4",X"6A",
		X"66",X"44",X"46",X"45",X"00",X"A6",X"6A",X"AB",X"A6",X"AA",X"A4",X"24",X"56",X"5A",X"00",X"A6",
		X"AA",X"AA",X"6A",X"AA",X"AA",X"44",X"5A",X"5A",X"00",X"AB",X"AA",X"A6",X"AA",X"AA",X"AA",X"54",
		X"56",X"5A",X"00",X"AA",X"AA",X"AB",X"AA",X"AA",X"AA",X"65",X"64",X"50",X"00",X"0A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"55",X"A4",X"60",X"00",X"0A",X"AA",X"AA",X"BA",X"AA",X"AA",X"6A",X"64",X"50",
		X"00",X"0A",X"AA",X"AA",X"AA",X"BA",X"AB",X"AA",X"45",X"60",X"00",X"00",X"AA",X"AA",X"AA",X"AA",
		X"BA",X"54",X"44",X"A0",X"00",X"00",X"AB",X"AA",X"AA",X"AA",X"AA",X"65",X"54",X"00",X"00",X"00",
		X"AA",X"BA",X"AA",X"AA",X"AA",X"A6",X"64",X"00",X"00",X"00",X"0A",X"AA",X"BA",X"BA",X"AA",X"AA",
		X"66",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AB",X"AA",X"AB",X"6A",X"00",X"00",X"00",X"00",X"00",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"05",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"02",X"02",X"02",X"03",X"04",X"06",X"0E",X"12",X"12",X"12",X"12",X"12",X"12",
		X"12",X"11",X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"10",X"0E",X"0C",X"1B",X"0F",X"23",X"10",
		X"67",X"0B",X"0D",X"00",X"00",X"A5",X"46",X"54",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"64",X"44",X"65",X"54",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"A6",X"54",X"A6",
		X"44",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"A6",X"64",X"A6",X"54",X"25",X"50",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"AA",X"65",X"A6",X"54",X"44",X"44",X"A0",X"00",X"00",X"00",X"0A",
		X"AA",X"BA",X"6B",X"A6",X"54",X"56",X"44",X"64",X"40",X"00",X"00",X"0A",X"AA",X"A6",X"6A",X"A6",
		X"55",X"65",X"54",X"65",X"46",X"00",X"00",X"0A",X"AA",X"A6",X"AB",X"66",X"54",X"65",X"45",X"A5",
		X"44",X"A0",X"00",X"AA",X"AA",X"AA",X"BA",X"A6",X"56",X"A5",X"56",X"A6",X"52",X"4A",X"00",X"AA",
		X"AA",X"BA",X"AA",X"66",X"66",X"A4",X"56",X"A6",X"45",X"4A",X"00",X"AA",X"AB",X"AA",X"AA",X"65",
		X"6A",X"A5",X"46",X"AA",X"55",X"5A",X"00",X"AA",X"AA",X"AA",X"AA",X"A6",X"AA",X"65",X"6A",X"BA",
		X"64",X"60",X"00",X"0A",X"AA",X"AA",X"AA",X"6A",X"AA",X"66",X"6A",X"AA",X"64",X"A0",X"00",X"0A",
		X"AA",X"AA",X"AA",X"AB",X"AA",X"66",X"AB",X"AA",X"65",X"A0",X"00",X"0A",X"AA",X"AA",X"AA",X"BA",
		X"A6",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"AA",
		X"56",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"AA",X"4A",X"00",X"00",X"00",
		X"0A",X"AA",X"BA",X"AA",X"AA",X"AB",X"AA",X"AA",X"5A",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",
		X"AB",X"AA",X"AA",X"A6",X"A0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"BA",X"AA",X"AA",X"A6",
		X"A0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"BA",X"AA",X"AA",X"AA",X"66",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"66",X"4A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A5",X"5A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"AA",X"66",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"AA",X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"02",X"02",X"02",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"03",X"03",X"04",X"04",X"05",X"06",X"07",X"08",
		X"09",X"0B",X"0C",X"0D",X"0E",X"0F",X"11",X"13",X"14",X"15",X"16",X"16",X"16",X"15",X"15",X"15",
		X"14",X"14",X"14",X"14",X"13",X"13",X"12",X"12",X"11",X"10",X"10",X"0F",X"0E",X"10",X"1C",X"10",
		X"A5",X"12",X"65",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"06",X"65",
		X"66",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"66",X"A0",X"00",X"AA",X"66",X"45",
		X"24",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A6",X"44",X"60",X"0A",X"66",X"64",X"54",
		X"44",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A6",X"52",X"60",X"AA",X"66",X"54",X"45",
		X"42",X"6A",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"65",X"64",X"4A",X"A6",X"55",X"54",X"54",
		X"46",X"6A",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"45",X"45",X"2A",X"55",X"55",X"65",X"45",
		X"24",X"6A",X"AA",X"00",X"00",X"00",X"00",X"A6",X"65",X"54",X"64",X"46",X"55",X"65",X"55",X"55",
		X"45",X"46",X"66",X"6A",X"00",X"00",X"0A",X"65",X"45",X"64",X"46",X"5A",X"66",X"66",X"55",X"55",
		X"56",X"54",X"42",X"66",X"00",X"0A",X"A6",X"64",X"42",X"65",X"46",X"45",X"AA",X"A6",X"66",X"AA",
		X"64",X"54",X"56",X"45",X"00",X"A6",X"55",X"55",X"54",X"46",X"66",X"64",X"42",X"4A",X"AA",X"4B",
		X"A6",X"65",X"55",X"4A",X"00",X"AA",X"55",X"66",X"65",X"44",X"6A",X"65",X"44",X"64",X"44",X"26",
		X"AA",X"A6",X"66",X"5A",X"00",X"AB",X"65",X"66",X"46",X"65",X"4A",X"66",X"55",X"55",X"55",X"44",
		X"26",X"AA",X"A5",X"6A",X"00",X"AA",X"AA",X"6A",X"64",X"65",X"5A",X"66",X"55",X"56",X"65",X"55",
		X"42",X"5A",X"A6",X"A0",X"00",X"0A",X"AA",X"AA",X"A5",X"46",X"46",X"AA",X"66",X"66",X"65",X"55",
		X"44",X"5A",X"AA",X"00",X"00",X"0A",X"AA",X"AA",X"A6",X"5A",X"54",X"5A",X"AA",X"AA",X"66",X"65",
		X"56",X"6A",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"6A",X"64",X"44",X"44",X"6B",X"AA",X"66",
		X"66",X"A0",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"BA",X"65",X"56",X"66",X"4A",X"AA",X"AA",
		X"A6",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"AA",X"44",X"A0",X"AA",
		X"A0",X"00",X"00",X"00",X"00",X"0A",X"AB",X"AA",X"AA",X"BA",X"AA",X"AB",X"A5",X"64",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"BA",X"AA",X"AB",X"AA",X"AA",X"BA",X"AA",X"65",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"BA",X"BA",X"AA",X"AA",X"AA",X"AA",X"A6",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",X"AA",X"6A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"BA",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"AA",X"AA",X"A6",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"AA",X"A6",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"13",X"0A",X"09",X"08",X"07",X"07",X"05",X"04",X"03",X"01",X"00",
		X"00",X"00",X"00",X"01",X"01",X"02",X"02",X"02",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",
		X"06",X"18",X"19",X"1A",X"1A",X"1A",X"1A",X"1C",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1D",X"1C",
		X"1A",X"19",X"18",X"17",X"13",X"13",X"12",X"12",X"11",X"0D",X"0C",X"0B",X"09",X"06",X"0A",X"13",
		X"1D",X"13",X"59",X"04",X"04",X"07",X"0C",X"13",X"6D",X"13",X"C1",X"06",X"05",X"08",X"0D",X"13",
		X"D9",X"14",X"41",X"06",X"05",X"07",X"0D",X"14",X"5B",X"14",X"B6",X"05",X"06",X"06",X"0A",X"14",
		X"D0",X"15",X"0C",X"05",X"04",X"07",X"0D",X"15",X"20",X"15",X"7B",X"05",X"06",X"07",X"0E",X"15",
		X"95",X"15",X"F7",X"06",X"06",X"07",X"0C",X"16",X"13",X"16",X"67",X"05",X"05",X"06",X"0A",X"16",
		X"7F",X"16",X"BB",X"04",X"04",X"07",X"0C",X"16",X"CF",X"17",X"23",X"05",X"05",X"08",X"0D",X"17",
		X"3B",X"17",X"A3",X"06",X"06",X"07",X"0D",X"17",X"BD",X"18",X"18",X"05",X"05",X"06",X"0A",X"18",
		X"32",X"18",X"6E",X"04",X"04",X"07",X"0D",X"18",X"82",X"18",X"DD",X"05",X"05",X"07",X"0E",X"18",
		X"F7",X"19",X"59",X"05",X"06",X"07",X"0C",X"19",X"75",X"19",X"C9",X"06",X"05",X"00",X"00",X"00",
		X"CC",X"DC",X"00",X"9D",X"DC",X"CD",X"DD",X"0D",X"00",X"9C",X"CC",X"DD",X"D0",X"00",X"00",X"00",
		X"0D",X"DD",X"DF",X"DC",X"00",X"00",X"DD",X"DD",X"DD",X"D0",X"00",X"00",X"CD",X"DD",X"DD",X"D0",
		X"00",X"00",X"0C",X"DD",X"DF",X"DC",X"00",X"9D",X"CC",X"CC",X"D0",X"00",X"00",X"9C",X"CC",X"CC",
		X"DD",X"0D",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"06",X"00",X"00",X"03",X"02",X"02",X"03",
		X"00",X"00",X"06",X"0A",X"0A",X"07",X"0A",X"09",X"09",X"0A",X"07",X"0A",X"0A",X"00",X"09",X"90",
		X"00",X"00",X"00",X"00",X"00",X"09",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DC",
		X"DD",X"00",X"00",X"00",X"0C",X"DD",X"DC",X"CC",X"D0",X"00",X"00",X"CD",X"DD",X"D0",X"00",X"C0",
		X"00",X"00",X"DD",X"DD",X"DF",X"C0",X"00",X"09",X"00",X"CD",X"DD",X"DD",X"CC",X"00",X"99",X"DD",
		X"CC",X"DD",X"DD",X"00",X"00",X"00",X"CD",X"CC",X"CC",X"FD",X"C0",X"00",X"00",X"00",X"CC",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"0C",X"00",X"00",X"00",X"00",X"00",X"0D",X"DC",X"00",
		X"00",X"03",X"03",X"04",X"05",X"04",X"04",X"01",X"00",X"02",X"04",X"06",X"07",X"05",X"06",X"0C",
		X"0D",X"0D",X"0B",X"0C",X"0A",X"0B",X"07",X"0A",X"0A",X"00",X"00",X"09",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"CC",X"DD",X"C0",X"00",X"00",X"09",X"00",X"CD",X"DD",X"DD",X"DD",X"C0",
		X"00",X"99",X"D0",X"CD",X"DD",X"DD",X"DD",X"CC",X"00",X"0C",X"CD",X"CD",X"DD",X"DF",X"00",X"0D",
		X"00",X"00",X"CC",X"CC",X"DD",X"CD",X"D0",X"0C",X"00",X"00",X"0C",X"CC",X"CD",X"D0",X"00",X"00",
		X"00",X"00",X"00",X"CD",X"0F",X"D0",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"D0",X"00",X"00",
		X"00",X"05",X"05",X"06",X"06",X"01",X"00",X"01",X"02",X"03",X"04",X"05",X"05",X"06",X"07",X"08",
		X"09",X"0B",X"0D",X"0E",X"0E",X"0E",X"09",X"09",X"07",X"07",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"9D",X"C0",X"00",X"00",X"09",X"00",X"00",X"CC",X"D0",X"00",X"00",
		X"99",X"90",X"CC",X"0C",X"DC",X"00",X"00",X"0C",X"D0",X"CC",X"CD",X"DD",X"00",X"00",X"0C",X"DC",
		X"CD",X"DD",X"DD",X"C0",X"00",X"0C",X"CC",X"DD",X"DD",X"DD",X"DC",X"00",X"00",X"CC",X"DD",X"DD",
		X"D0",X"CD",X"00",X"00",X"CC",X"CD",X"DC",X"F0",X"0D",X"00",X"00",X"CC",X"0F",X"CD",X"DD",X"0C",
		X"00",X"00",X"CD",X"00",X"DD",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"DC",X"00",X"00",X"00",X"00",X"06",X"06",X"01",X"00",X"01",X"01",X"01",X"02",X"02",X"02",
		X"02",X"03",X"03",X"08",X"09",X"09",X"0A",X"0A",X"0B",X"0C",X"0C",X"0C",X"0C",X"08",X"04",X"06",
		X"09",X"90",X"00",X"09",X"90",X"00",X"0D",X"D0",X"00",X"0D",X"D0",X"00",X"0C",X"D0",X"CD",X"0C",
		X"D0",X"00",X"0C",X"CC",X"DD",X"DD",X"C0",X"00",X"0C",X"CD",X"DD",X"DD",X"D0",X"00",X"0C",X"CD",
		X"DD",X"DD",X"D0",X"00",X"CC",X"CC",X"DD",X"DD",X"DC",X"00",X"DC",X"0F",X"CD",X"F0",X"CD",X"00",
		X"C0",X"0C",X"CD",X"C0",X"0D",X"00",X"CD",X"0C",X"00",X"C0",X"DC",X"00",X"01",X"01",X"01",X"01",
		X"01",X"01",X"00",X"00",X"00",X"00",X"09",X"09",X"09",X"09",X"09",X"09",X"0A",X"0A",X"0A",X"0A",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"0D",X"C0",X"CC",X"00",X"99",X"00",X"00",X"CC",X"CC",X"DD",
		X"0D",X"D9",X"00",X"00",X"CC",X"DD",X"DD",X"DD",X"C0",X"00",X"0C",X"CC",X"DD",X"DD",X"DD",X"00",
		X"00",X"CC",X"0C",X"DD",X"DD",X"DD",X"00",X"00",X"D0",X"0F",X"CD",X"DD",X"DC",X"00",X"00",X"CC",
		X"0C",X"CC",X"F0",X"CC",X"00",X"00",X"00",X"0D",X"0C",X"D0",X"CD",X"00",X"00",X"00",X"00",X"0C",
		X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"0C",X"C0",X"00",X"00",X"04",X"04",X"03",X"03",X"02",
		X"02",X"01",X"00",X"00",X"00",X"03",X"05",X"07",X"05",X"06",X"05",X"0C",X"0C",X"0B",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"0A",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",
		X"90",X"00",X"00",X"00",X"00",X"0C",X"DD",X"00",X"00",X"00",X"00",X"00",X"CC",X"D0",X"00",X"00",
		X"00",X"00",X"0C",X"CC",X"DC",X"D0",X"00",X"00",X"0C",X"CC",X"CD",X"DD",X"D0",X"09",X"90",X"CC",
		X"C0",X"CD",X"DD",X"DD",X"CD",X"90",X"C0",X"0F",X"CD",X"DD",X"DD",X"DD",X"00",X"C0",X"0D",X"CD",
		X"DD",X"DD",X"C0",X"00",X"00",X"00",X"0C",X"FD",X"DC",X"00",X"00",X"00",X"00",X"0C",X"0C",X"DC",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"0C",X"D0",X"00",X"00",
		X"00",X"00",X"0C",X"DC",X"00",X"00",X"00",X"07",X"06",X"05",X"04",X"03",X"01",X"00",X"00",X"00",
		X"05",X"05",X"07",X"07",X"05",X"08",X"09",X"08",X"07",X"09",X"0D",X"0D",X"0C",X"0B",X"0A",X"0A",
		X"09",X"09",X"08",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"0C",X"D9",X"90",
		X"00",X"00",X"CC",X"DD",X"CD",X"DD",X"00",X"00",X"CD",X"CD",X"DD",X"DD",X"00",X"00",X"00",X"C0",
		X"00",X"CD",X"DD",X"DD",X"00",X"00",X"00",X"0F",X"DD",X"DD",X"DC",X"00",X"00",X"00",X"DD",X"DD",
		X"DD",X"D0",X"09",X"90",X"00",X"0C",X"DD",X"DD",X"DC",X"DD",X"90",X"00",X"0D",X"FC",X"CD",X"DD",
		X"DC",X"00",X"00",X"00",X"00",X"CD",X"CC",X"00",X"00",X"00",X"00",X"0C",X"DD",X"00",X"00",X"00",
		X"00",X"0C",X"DD",X"D0",X"00",X"00",X"00",X"09",X"07",X"02",X"00",X"00",X"03",X"02",X"03",X"03",
		X"06",X"05",X"03",X"0A",X"0B",X"0A",X"08",X"0A",X"0A",X"0D",X"0D",X"0C",X"0A",X"08",X"07",X"CC",
		X"DC",X"00",X"00",X"00",X"00",X"C0",X"CD",X"CD",X"DD",X"D9",X"00",X"00",X"0D",X"DD",X"DC",X"D9",
		X"00",X"CC",X"FC",X"DD",X"D0",X"00",X"00",X"0C",X"CD",X"DD",X"DD",X"00",X"00",X"0C",X"CD",X"DD",
		X"DC",X"00",X"00",X"CC",X"FC",X"DD",X"C0",X"00",X"00",X"00",X"0C",X"CC",X"DD",X"D9",X"00",X"C0",
		X"CC",X"CC",X"CC",X"D9",X"00",X"CD",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",
		X"01",X"00",X"03",X"00",X"00",X"04",X"0A",X"0A",X"07",X"08",X"08",X"07",X"0A",X"0A",X"04",X"00",
		X"0C",X"DD",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"C0",X"00",X"00",X"00",X"DC",X"FD",X"DD",X"DD",X"D0",X"00",X"00",X"0D",X"DD",X"DD",X"DC",
		X"D9",X"90",X"0C",X"CD",X"DD",X"DD",X"D0",X"09",X"00",X"00",X"CF",X"DD",X"DD",X"DD",X"00",X"00",
		X"C0",X"00",X"CD",X"DD",X"CC",X"00",X"00",X"CD",X"CD",X"CC",X"CC",X"00",X"00",X"00",X"0C",X"DC",
		X"CC",X"CD",X"D0",X"00",X"00",X"00",X"00",X"00",X"0C",X"D9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"03",X"03",X"06",X"02",X"03",X"01",X"02",X"00",X"00",X"01",X"07",X"08",X"06",
		X"07",X"09",X"0B",X"0D",X"0C",X"0A",X"0A",X"08",X"09",X"0A",X"0A",X"00",X"00",X"0C",X"CD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"0D",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"0D",X"C0",X"DD",X"00",X"00",X"00",X"00",X"00",X"0C",X"FD",X"DD",
		X"D0",X"00",X"00",X"0D",X"0D",X"DD",X"DD",X"DD",X"DD",X"00",X"00",X"D0",X"00",X"FD",X"DD",X"DD",
		X"DD",X"D0",X"00",X"CD",X"DC",X"DD",X"DD",X"DD",X"0C",X"99",X"00",X"0C",X"CC",X"CC",X"DD",X"DD",
		X"00",X"90",X"00",X"00",X"0C",X"CD",X"DC",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"90",
		X"00",X"00",X"00",X"05",X"05",X"07",X"05",X"05",X"01",X"00",X"00",X"01",X"03",X"05",X"06",X"07",
		X"08",X"09",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0D",X"08",X"08",X"09",X"09",X"00",X"00",X"00",
		X"CD",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"0D",X"00",X"DD",
		X"00",X"00",X"C0",X"CD",X"DD",X"F0",X"CD",X"00",X"00",X"D0",X"0D",X"DD",X"DD",X"DD",X"00",X"00",
		X"DC",X"0F",X"DD",X"DD",X"DD",X"00",X"00",X"CD",X"CC",X"DD",X"DD",X"DD",X"C0",X"00",X"0C",X"CC",
		X"CD",X"DD",X"CC",X"D0",X"00",X"00",X"CC",X"CC",X"CD",X"0C",X"D0",X"00",X"00",X"CD",X"D0",X"CC",
		X"0C",X"99",X"00",X"00",X"0C",X"DC",X"00",X"00",X"90",X"00",X"00",X"0C",X"D9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"06",X"08",X"05",X"00",X"00",X"00",X"00",X"01",
		X"02",X"02",X"03",X"03",X"04",X"09",X"09",X"0A",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0C",X"0B",
		X"06",X"06",X"CC",X"0D",X"00",X"D0",X"DC",X"00",X"D0",X"0C",X"DD",X"D0",X"0D",X"00",X"CD",X"0F",
		X"DD",X"F0",X"CD",X"00",X"CC",X"DC",X"DD",X"DD",X"DC",X"00",X"0C",X"CD",X"DD",X"DD",X"D0",X"00",
		X"0C",X"CD",X"DD",X"DD",X"D0",X"00",X"0C",X"CC",X"DD",X"DC",X"D0",X"00",X"0C",X"D0",X"DD",X"0D",
		X"D0",X"00",X"0C",X"D0",X"00",X"0C",X"D0",X"00",X"09",X"90",X"00",X"09",X"90",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"0A",X"0A",X"0A",X"0A",X"09",X"09",X"09",X"09",
		X"09",X"09",X"00",X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"CD",X"00",X"C0",X"00",X"00",X"00",
		X"00",X"CD",X"0C",X"D0",X"D0",X"00",X"00",X"00",X"CD",X"0F",X"DD",X"D0",X"CC",X"00",X"00",X"CD",
		X"DD",X"DD",X"F0",X"0D",X"00",X"00",X"CD",X"DD",X"DD",X"D0",X"DD",X"00",X"00",X"CC",X"DD",X"DD",
		X"DD",X"D0",X"00",X"0C",X"CC",X"CD",X"DD",X"DD",X"C0",X"00",X"9D",X"D0",X"CC",X"CD",X"DC",X"00",
		X"00",X"99",X"00",X"CC",X"0C",X"D0",X"00",X"00",X"00",X"00",X"00",X"0D",X"D0",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"03",X"02",X"02",
		X"02",X"02",X"02",X"02",X"01",X"00",X"00",X"07",X"06",X"07",X"05",X"07",X"09",X"0C",X"0C",X"0C",
		X"0B",X"0B",X"0A",X"09",X"09",X"08",X"08",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"0D",X"00",X"00",X"00",X"00",X"00",X"CD",X"00",X"00",X"00",X"00",X"00",X"0C",X"DC",X"0D",
		X"00",X"00",X"00",X"00",X"0D",X"DD",X"FD",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"DD",X"0C",
		X"C0",X"0D",X"DD",X"DD",X"DD",X"FC",X"00",X"D0",X"9D",X"DC",X"DD",X"DD",X"D0",X"CD",X"C0",X"99",
		X"00",X"CD",X"DD",X"DD",X"DC",X"00",X"00",X"00",X"CC",X"CC",X"CD",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"C0",X"00",X"00",X"00",X"00",X"0D",X"DC",X"00",X"00",X"00",X"00",X"00",X"99",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"05",X"04",X"04",X"03",X"03",X"02",X"01",
		X"00",X"00",X"04",X"06",X"05",X"04",X"05",X"08",X"08",X"06",X"08",X"08",X"0D",X"0D",X"0D",X"0C",
		X"0A",X"09",X"08",X"07",X"06",X"00",X"00",X"00",X"CC",X"DD",X"00",X"00",X"00",X"00",X"0C",X"DC",
		X"00",X"00",X"00",X"00",X"0C",X"DD",X"D0",X"00",X"00",X"00",X"0C",X"DC",X"DD",X"DF",X"DD",X"00",
		X"00",X"9C",X"CC",X"DD",X"DD",X"DC",X"00",X"00",X"99",X"00",X"DD",X"DD",X"DD",X"D0",X"00",X"00",
		X"00",X"DD",X"DD",X"DF",X"00",X"00",X"00",X"00",X"CD",X"DD",X"D0",X"00",X"D0",X"00",X"00",X"0C",
		X"CD",X"CD",X"CD",X"C0",X"00",X"0C",X"CC",X"CC",X"CC",X"C0",X"00",X"00",X"99",X"DC",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"06",X"05",X"03",X"01",X"00",X"00",X"04",
		X"04",X"05",X"03",X"02",X"03",X"0A",X"08",X"07",X"0A",X"0A",X"0B",X"0A",X"0D",X"0D",X"0B",X"06",
		X"04",X"08",X"11",X"19",X"E9",X"1A",X"71",X"07",X"08",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AB",X"AA",X"A0",X"00",X"00",X"00",X"0A",X"AA",X"BD",X"BA",X"AA",X"00",
		X"00",X"00",X"BC",X"BA",X"BB",X"BA",X"BD",X"B0",X"00",X"0A",X"CC",X"AA",X"AB",X"AA",X"AD",X"DA",
		X"00",X"AA",X"BA",X"BA",X"BB",X"BA",X"BA",X"BA",X"A0",X"AA",X"AA",X"AA",X"44",X"4A",X"AA",X"AA",
		X"A0",X"0A",X"BA",X"B4",X"54",X"24",X"BA",X"BA",X"00",X"0C",X"BB",X"B5",X"6D",X"54",X"BB",X"BD",
		X"00",X"0A",X"BA",X"B5",X"56",X"54",X"BA",X"BA",X"00",X"AA",X"AA",X"AA",X"55",X"5A",X"AA",X"AA",
		X"A0",X"AA",X"BA",X"BA",X"BB",X"BA",X"BA",X"BA",X"A0",X"0A",X"CC",X"AA",X"AB",X"AA",X"AC",X"CA",
		X"00",X"00",X"BC",X"BA",X"BB",X"BA",X"BC",X"B0",X"00",X"00",X"0A",X"AA",X"BC",X"BA",X"AA",X"00",
		X"00",X"00",X"00",X"AA",X"AB",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",
		X"00",X"05",X"04",X"03",X"02",X"01",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"01",X"02",X"03",
		X"04",X"05",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"0F",X"0E",X"0E",X"0E",X"0F",X"0F",X"0E",X"0D",
		X"0C",X"0B",X"0A",X"05",X"05",X"1A",X"D4",X"00",X"00",X"02",X"02",X"04",X"07",X"1A",X"ED",X"00",
		X"00",X"02",X"02",X"03",X"09",X"1B",X"09",X"00",X"00",X"02",X"02",X"04",X"07",X"1B",X"24",X"00",
		X"00",X"04",X"02",X"05",X"05",X"1B",X"40",X"00",X"00",X"06",X"02",X"04",X"07",X"1B",X"59",X"00",
		X"00",X"04",X"04",X"03",X"09",X"1B",X"75",X"00",X"00",X"02",X"06",X"04",X"07",X"1B",X"90",X"00",
		X"00",X"02",X"04",X"00",X"04",X"44",X"00",X"00",X"00",X"45",X"42",X"40",X"00",X"00",X"56",X"D5",
		X"44",X"42",X"20",X"55",X"65",X"40",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"04",X"44",X"00",
		X"00",X"45",X"42",X"40",X"00",X"56",X"D5",X"40",X"00",X"55",X"65",X"40",X"00",X"05",X"55",X"20",
		X"00",X"00",X"00",X"52",X"00",X"00",X"00",X"06",X"20",X"04",X"44",X"00",X"45",X"42",X"40",X"56",
		X"D5",X"40",X"55",X"65",X"40",X"05",X"55",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",
		X"00",X"00",X"20",X"00",X"00",X"04",X"44",X"00",X"00",X"45",X"42",X"40",X"00",X"56",X"D5",X"40",
		X"00",X"55",X"65",X"40",X"06",X"25",X"55",X"00",X"62",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"00",X"04",X"44",X"00",X"00",X"00",X"45",X"42",X"40",X"22",X"24",X"46",X"D5",X"40",X"00",
		X"00",X"55",X"65",X"40",X"00",X"00",X"05",X"55",X"00",X"20",X"00",X"00",X"00",X"62",X"00",X"00",
		X"00",X"06",X"24",X"44",X"00",X"00",X"45",X"42",X"40",X"00",X"56",X"D5",X"40",X"00",X"55",X"65",
		X"40",X"00",X"05",X"55",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",X"00",X"00",X"20",
		X"00",X"04",X"44",X"00",X"45",X"42",X"40",X"56",X"D5",X"40",X"55",X"65",X"40",X"05",X"55",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"52",X"00",X"04",X"44",X"20",X"00",X"45",X"42",X"40",X"00",
		X"56",X"D5",X"40",X"00",X"55",X"65",X"40",X"00",X"05",X"55",X"00",X"00",X"06",X"0D",X"1B",X"BC",
		X"1C",X"0A",X"06",X"06",X"06",X"0D",X"1C",X"04",X"1C",X"16",X"06",X"06",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"02",X"33",X"00",X"00",X"00",X"00",X"23",X"44",X"40",X"02",X"00",X"02",X"44",
		X"55",X"55",X"23",X"30",X"24",X"45",X"66",X"63",X"33",X"00",X"00",X"00",X"12",X"42",X"20",X"00",
		X"00",X"00",X"23",X"32",X"00",X"00",X"00",X"00",X"23",X"22",X"00",X"00",X"00",X"04",X"33",X"22",
		X"00",X"00",X"00",X"04",X"43",X"21",X"00",X"00",X"00",X"05",X"54",X"42",X"00",X"00",X"00",X"00",
		X"05",X"65",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"04",X"03",X"02",X"01",X"00",X"04",
		X"04",X"04",X"03",X"03",X"03",X"05",X"06",X"05",X"06",X"0A",X"0B",X"0A",X"09",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"07",X"07",X"1C",X"2C",X"1C",X"5D",X"07",X"03",X"05",X"56",X"22",X"11",
		X"22",X"20",X"00",X"05",X"56",X"52",X"22",X"23",X"35",X"00",X"BA",X"AA",X"51",X"23",X"34",X"4A",
		X"00",X"BB",X"BA",X"61",X"22",X"34",X"4A",X"00",X"BA",X"AA",X"51",X"23",X"34",X"4A",X"00",X"05",
		X"56",X"52",X"22",X"23",X"35",X"00",X"05",X"56",X"22",X"11",X"22",X"20",X"00",X"01",X"01",X"00",
		X"00",X"00",X"01",X"01",X"0B",X"0C",X"0C",X"0C",X"0C",X"0C",X"0B",X"0A",X"12",X"1C",X"7B",X"1D",
		X"2F",X"0A",X"09",X"0A",X"12",X"1D",X"25",X"1D",X"40",X"0A",X"09",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"34",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"23",X"44",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"02",X"23",X"55",X"61",X"22",
		X"00",X"00",X"00",X"00",X"53",X"22",X"35",X"56",X"22",X"33",X"20",X"00",X"00",X"05",X"54",X"44",
		X"45",X"52",X"23",X"33",X"43",X"00",X"00",X"65",X"36",X"BB",X"35",X"22",X"33",X"33",X"44",X"34",
		X"00",X"54",X"3B",X"0A",X"A2",X"23",X"33",X"44",X"30",X"00",X"00",X"54",X"30",X"00",X"42",X"23",
		X"44",X"45",X"50",X"00",X"00",X"44",X"3C",X"0A",X"21",X"34",X"45",X"54",X"45",X"00",X"00",X"54",
		X"60",X"03",X"13",X"34",X"55",X"45",X"54",X"50",X"00",X"55",X"A0",X"51",X"23",X"45",X"54",X"54",
		X"55",X"40",X"00",X"56",X"A5",X"22",X"34",X"54",X"43",X"45",X"54",X"50",X"00",X"00",X"02",X"23",
		X"45",X"42",X"34",X"55",X"55",X"54",X"00",X"00",X"32",X"34",X"54",X"23",X"44",X"55",X"55",X"45",
		X"00",X"00",X"23",X"45",X"56",X"66",X"55",X"55",X"55",X"54",X"00",X"00",X"02",X"04",X"00",X"23",
		X"00",X"55",X"50",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"08",
		X"07",X"06",X"05",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",X"02",X"03",
		X"0D",X"09",X"0A",X"0D",X"0E",X"0F",X"10",X"12",X"0F",X"0F",X"10",X"11",X"11",X"11",X"12",X"12",
		X"12",X"12",X"0E",X"08",X"08",X"1D",X"63",X"1D",X"A3",X"08",X"04",X"08",X"08",X"1D",X"9B",X"1D",
		X"AA",X"08",X"04",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",
		X"55",X"56",X"00",X"00",X"00",X"00",X"03",X"42",X"22",X"22",X"00",X"00",X"00",X"00",X"45",X"22",
		X"34",X"54",X"00",X"00",X"00",X"05",X"52",X"23",X"34",X"50",X"00",X"00",X"03",X"56",X"22",X"33",
		X"45",X"40",X"00",X"00",X"35",X"65",X"33",X"34",X"5A",X"00",X"00",X"33",X"55",X"63",X"33",X"52",
		X"00",X"00",X"00",X"09",X"08",X"07",X"06",X"05",X"03",X"02",X"00",X"0A",X"0E",X"0E",X"0E",X"0D",
		X"0D",X"0C",X"0A",X"06",X"0B",X"1D",X"BB",X"1D",X"FD",X"06",X"05",X"00",X"30",X"00",X"00",X"00",
		X"00",X"11",X"23",X"30",X"00",X"00",X"00",X"02",X"34",X"44",X"00",X"00",X"00",X"00",X"24",X"54",
		X"44",X"54",X"50",X"0A",X"23",X"5A",X"05",X"45",X"00",X"0A",X"23",X"45",X"A0",X"B5",X"00",X"00",
		X"23",X"5A",X"05",X"45",X"00",X"00",X"24",X"54",X"44",X"54",X"50",X"02",X"34",X"44",X"00",X"00",
		X"00",X"11",X"23",X"30",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"02",X"00",X"01",
		X"02",X"01",X"01",X"02",X"02",X"01",X"00",X"02",X"03",X"05",X"06",X"0B",X"0A",X"0A",X"0A",X"0B",
		X"06",X"05",X"03",X"07",X"0F",X"1E",X"23",X"1E",X"8C",X"07",X"07",X"07",X"0F",X"1E",X"85",X"1E",
		X"9A",X"07",X"07",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"A5",X"AB",X"00",X"00",X"00",X"00",
		X"0A",X"A5",X"5A",X"B0",X"00",X"00",X"65",X"5A",X"AB",X"BB",X"B0",X"00",X"00",X"A6",X"64",X"43",
		X"45",X"5B",X"AA",X"00",X"06",X"55",X"43",X"45",X"6B",X"AA",X"00",X"00",X"65",X"53",X"45",X"5B",
		X"AA",X"00",X"00",X"65",X"53",X"45",X"6B",X"AA",X"00",X"00",X"56",X"54",X"55",X"5B",X"AA",X"00",
		X"00",X"06",X"54",X"55",X"6B",X"AA",X"00",X"00",X"0A",X"AB",X"BA",X"A0",X"00",X"00",X"00",X"0A",
		X"AB",X"BB",X"A0",X"00",X"00",X"00",X"0A",X"0B",X"0A",X"00",X"00",X"00",X"05",X"05",X"04",X"04",
		X"03",X"00",X"00",X"01",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"07",X"07",X"08",X"08",X"09",
		X"09",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"09",X"09",X"08",X"06",X"0B",X"1E",X"BA",X"1E",X"FC",
		X"06",X"05",X"06",X"0B",X"1E",X"F6",X"1F",X"06",X"06",X"05",X"A0",X"00",X"00",X"00",X"05",X"30",
		X"CC",X"00",X"00",X"05",X"43",X"A0",X"CC",X"C0",X"05",X"44",X"45",X"A0",X"DC",X"C4",X"34",X"44",
		X"4A",X"00",X"D2",X"22",X"33",X"34",X"5A",X"00",X"24",X"42",X"22",X"34",X"A0",X"00",X"55",X"44",
		X"32",X"34",X"00",X"00",X"65",X"54",X"42",X"30",X"00",X"00",X"06",X"55",X"44",X"40",X"00",X"00",
		X"00",X"65",X"54",X"00",X"00",X"00",X"00",X"06",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"02",X"03",X"0B",X"0B",X"0B",X"0A",X"0A",X"09",X"08",X"07",X"07",
		X"06",X"06",X"08",X"0D",X"1F",X"22",X"1F",X"8A",X"08",X"06",X"08",X"0D",X"1F",X"82",X"1F",X"96",
		X"08",X"06",X"00",X"0A",X"AA",X"AA",X"20",X"00",X"00",X"00",X"00",X"06",X"BB",X"B2",X"40",X"00",
		X"00",X"00",X"0A",X"A4",X"55",X"62",X"4A",X"BA",X"00",X"00",X"AA",X"A3",X"46",X"23",X"4A",X"5B",
		X"BA",X"00",X"0B",X"A3",X"44",X"23",X"46",X"55",X"5B",X"00",X"BB",X"B2",X"42",X"33",X"4A",X"34",
		X"55",X"00",X"0B",X"B3",X"52",X"33",X"4B",X"53",X"45",X"00",X"BB",X"B5",X"33",X"44",X"5B",X"65",
		X"34",X"00",X"0B",X"B5",X"34",X"44",X"5B",X"B6",X"55",X"00",X"BB",X"53",X"44",X"55",X"50",X"5B",
		X"63",X"00",X"0B",X"53",X"45",X"65",X"00",X"05",X"63",X"00",X"0A",X"05",X"56",X"50",X"00",X"00",
		X"60",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"01",X"04",X"09",X"09",X"0C",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0D",X"06",X"07",X"0D",X"1F",X"B4",X"20",X"0F",X"07",X"06",X"07",X"0D",X"20",X"08",
		X"20",X"1B",X"07",X"06",X"00",X"00",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"00",X"6B",X"BB",X"B0",
		X"00",X"00",X"0A",X"BB",X"46",X"66",X"5A",X"A0",X"00",X"B5",X"45",X"25",X"55",X"5A",X"AA",X"00",
		X"53",X"32",X"23",X"43",X"3A",X"B0",X"00",X"44",X"43",X"23",X"22",X"2B",X"BB",X"00",X"45",X"43",
		X"12",X"33",X"3B",X"B0",X"00",X"55",X"54",X"13",X"44",X"3B",X"BB",X"00",X"55",X"55",X"14",X"35",
		X"5B",X"B0",X"00",X"55",X"55",X"23",X"06",X"5B",X"B5",X"00",X"45",X"56",X"50",X"00",X"6B",X"B0",
		X"00",X"45",X"56",X"00",X"00",X"0A",X"A0",X"00",X"34",X"60",X"00",X"00",X"00",X"00",X"00",X"04",
		X"04",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",X"0B",X"0C",
		X"0B",X"0C",X"0B",X"0C",X"0B",X"0C",X"0B",X"0B",X"03",X"07",X"0D",X"20",X"39",X"20",X"94",X"07",
		X"06",X"07",X"0D",X"20",X"8D",X"20",X"A0",X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"CC",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"00",X"00",X"00",
		X"00",X"0C",X"CC",X"CC",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CD",X"00",X"00",X"00",X"0B",X"CC",
		X"CC",X"DD",X"00",X"00",X"00",X"BC",X"CC",X"CD",X"DD",X"00",X"00",X"AB",X"35",X"54",X"33",X"33",
		X"00",X"00",X"A6",X"45",X"43",X"32",X"32",X"00",X"0A",X"B3",X"54",X"32",X"22",X"23",X"30",X"0A",
		X"54",X"43",X"22",X"12",X"22",X"00",X"AB",X"34",X"32",X"21",X"11",X"20",X"00",X"AB",X"65",X"44",
		X"33",X"33",X"00",X"00",X"0B",X"09",X"08",X"07",X"06",X"05",X"04",X"02",X"02",X"01",X"01",X"00",
		X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0D",X"0C",X"0B",X"0A",X"06",X"09",
		X"20",X"BE",X"20",X"F4",X"06",X"04",X"06",X"09",X"20",X"EE",X"20",X"FC",X"06",X"04",X"A6",X"54",
		X"12",X"23",X"33",X"40",X"A5",X"44",X"12",X"33",X"30",X"00",X"A6",X"41",X"23",X"33",X"00",X"00",
		X"A5",X"41",X"23",X"00",X"00",X"00",X"A6",X"12",X"33",X"50",X"00",X"00",X"A5",X"12",X"33",X"40",
		X"00",X"00",X"00",X"AB",X"BB",X"00",X"00",X"00",X"00",X"AB",X"BB",X"00",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"03",X"0B",X"09",X"08",
		X"06",X"07",X"07",X"06",X"06",X"06",X"0A",X"19",X"21",X"0A",X"00",X"00",X"00",X"55",X"61",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"56",X"22",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"52",X"23",X"30",X"40",X"00",X"00",X"00",X"30",X"00",X"05",X"22",X"33",X"33",X"40",X"00",
		X"00",X"00",X"3B",X"E0",X"A2",X"23",X"33",X"44",X"36",X"50",X"00",X"00",X"3E",X"EE",X"42",X"23",
		X"44",X"45",X"5A",X"00",X"00",X"00",X"3C",X"EA",X"21",X"34",X"45",X"54",X"45",X"60",X"00",X"00",
		X"0E",X"E3",X"13",X"34",X"55",X"45",X"50",X"00",X"00",X"00",X"AE",X"51",X"23",X"45",X"54",X"54",
		X"50",X"00",X"00",X"00",X"05",X"22",X"34",X"54",X"43",X"45",X"50",X"00",X"00",X"00",X"02",X"23",
		X"45",X"42",X"34",X"55",X"50",X"00",X"00",X"00",X"32",X"34",X"54",X"23",X"44",X"55",X"55",X"45",
		X"AA",X"00",X"23",X"45",X"56",X"66",X"55",X"55",X"55",X"54",X"AA",X"00",X"0A",X"19",X"21",X"90",
		X"00",X"00",X"00",X"45",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"55",X"62",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"22",X"30",X"30",X"00",X"00",X"00",X"30",X"00",
		X"03",X"52",X"23",X"34",X"40",X"00",X"00",X"00",X"4B",X"E0",X"B4",X"52",X"33",X"44",X"44",X"50",
		X"00",X"00",X"4E",X"EE",X"B5",X"22",X"33",X"44",X"55",X"00",X"00",X"00",X"4D",X"EA",X"B2",X"13",
		X"34",X"45",X"56",X"A0",X"00",X"00",X"0E",X"EB",X"51",X"34",X"44",X"55",X"50",X"00",X"00",X"00",
		X"BE",X"B5",X"22",X"34",X"45",X"54",X"50",X"00",X"00",X"00",X"0B",X"45",X"23",X"44",X"54",X"45",
		X"50",X"00",X"00",X"00",X"04",X"62",X"33",X"45",X"43",X"45",X"50",X"00",X"00",X"00",X"45",X"52",
		X"34",X"54",X"34",X"55",X"55",X"45",X"AA",X"00",X"56",X"23",X"34",X"66",X"55",X"55",X"55",X"54",
		X"AA",X"00",X"0A",X"19",X"22",X"16",X"00",X"00",X"00",X"45",X"56",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"55",X"64",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"55",X"52",X"20",
		X"40",X"00",X"00",X"00",X"40",X"00",X"03",X"44",X"52",X"33",X"40",X"00",X"00",X"00",X"4A",X"E0",
		X"B4",X"45",X"22",X"34",X"44",X"40",X"00",X"00",X"4E",X"EE",X"B4",X"52",X"23",X"34",X"44",X"00",
		X"00",X"00",X"4D",X"BA",X"B5",X"51",X"33",X"44",X"46",X"A0",X"00",X"00",X"0E",X"EB",X"45",X"22",
		X"34",X"44",X"50",X"00",X"00",X"00",X"AE",X"B4",X"55",X"23",X"34",X"45",X"50",X"00",X"00",X"00",
		X"0B",X"44",X"52",X"23",X"44",X"55",X"50",X"00",X"00",X"00",X"04",X"56",X"22",X"34",X"45",X"45",
		X"50",X"00",X"00",X"00",X"45",X"55",X"23",X"44",X"54",X"55",X"55",X"45",X"AB",X"00",X"55",X"62",
		X"23",X"45",X"66",X"55",X"55",X"54",X"AA",X"00",X"08",X"19",X"22",X"9C",X"00",X"00",X"00",X"00",
		X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"35",X"55",X"56",X"00",X"00",X"00",X"00",X"03",X"42",X"22",X"22",X"00",X"00",X"00",X"00",X"45",
		X"22",X"34",X"54",X"00",X"00",X"00",X"05",X"52",X"23",X"34",X"54",X"00",X"00",X"03",X"56",X"22",
		X"33",X"45",X"40",X"00",X"00",X"35",X"65",X"33",X"34",X"5A",X"00",X"00",X"33",X"55",X"63",X"33",
		X"52",X"10",X"00",X"00",X"05",X"56",X"22",X"11",X"22",X"22",X"00",X"00",X"05",X"56",X"52",X"22",
		X"23",X"35",X"20",X"00",X"BA",X"AA",X"51",X"23",X"34",X"4A",X"20",X"00",X"BB",X"BA",X"61",X"22",
		X"34",X"4A",X"20",X"00",X"08",X"19",X"23",X"08",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"55",X"66",X"00",
		X"00",X"00",X"00",X"05",X"44",X"22",X"23",X"00",X"00",X"00",X"00",X"53",X"BC",X"CB",X"B5",X"00",
		X"00",X"00",X"05",X"25",X"BE",X"EC",X"B3",X"00",X"00",X"04",X"52",X"4B",X"EE",X"EE",X"50",X"00",
		X"00",X"45",X"24",X"BC",X"EE",X"E4",X"00",X"00",X"45",X"63",X"2B",X"BC",X"EA",X"20",X"00",X"00",
		X"04",X"33",X"22",X"3A",X"BE",X"E5",X"00",X"00",X"0A",X"23",X"5A",X"CB",X"BA",X"EA",X"30",X"00",
		X"AA",X"32",X"35",X"CC",X"CB",X"EA",X"20",X"00",X"AA",X"51",X"25",X"BB",X"CC",X"BA",X"20",X"00",
		X"08",X"19",X"23",X"74",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"55",X"66",X"00",X"00",X"00",X"00",X"05",
		X"32",X"22",X"22",X"00",X"00",X"00",X"00",X"45",X"23",X"CB",X"A5",X"00",X"00",X"00",X"05",X"52",
		X"24",X"AC",X"B4",X"00",X"00",X"04",X"55",X"22",X"5E",X"EE",X"50",X"00",X"00",X"45",X"62",X"25",
		X"CE",X"E4",X"00",X"00",X"45",X"56",X"22",X"35",X"EA",X"20",X"00",X"00",X"06",X"42",X"12",X"23",
		X"4A",X"E5",X"00",X"00",X"06",X"A5",X"33",X"45",X"BA",X"EA",X"30",X"00",X"BA",X"A5",X"22",X"35",
		X"CB",X"EA",X"20",X"00",X"BA",X"A6",X"12",X"25",X"CC",X"BA",X"20",X"00",X"07",X"0C",X"23",X"E4",
		X"00",X"00",X"06",X"05",X"00",X"0A",X"66",X"AB",X"BB",X"A0",X"00",X"00",X"06",X"55",X"6B",X"CB",
		X"B0",X"00",X"00",X"A6",X"44",X"56",X"D5",X"46",X"00",X"0A",X"61",X"15",X"45",X"44",X"56",X"00",
		X"A6",X"65",X"23",X"31",X"35",X"6A",X"00",X"63",X"22",X"54",X"41",X"23",X"56",X"00",X"65",X"45",
		X"35",X"62",X"44",X"66",X"00",X"A6",X"56",X"44",X"54",X"46",X"6A",X"00",X"0B",X"66",X"55",X"24",
		X"55",X"6A",X"00",X"0A",X"BB",X"42",X"13",X"66",X"6A",X"00",X"06",X"42",X"43",X"56",X"6A",X"A0",
		X"00",X"0A",X"55",X"56",X"6A",X"A0",X"00",X"00",X"05",X"01",X"24",X"B8",X"24",X"BD",X"04",X"00",
		X"05",X"03",X"24",X"BF",X"24",X"CE",X"04",X"01",X"04",X"05",X"24",X"D4",X"24",X"E8",X"03",X"02",
		X"04",X"05",X"24",X"F2",X"25",X"06",X"03",X"02",X"04",X"07",X"25",X"10",X"25",X"2C",X"03",X"03",
		X"03",X"07",X"25",X"3A",X"25",X"4F",X"02",X"03",X"03",X"07",X"25",X"5D",X"25",X"72",X"02",X"03",
		X"02",X"09",X"25",X"80",X"25",X"92",X"01",X"04",X"01",X"09",X"25",X"A4",X"25",X"AD",X"00",X"04",
		X"02",X"09",X"25",X"BF",X"25",X"D1",X"01",X"04",X"03",X"07",X"25",X"E3",X"25",X"F8",X"02",X"03",
		X"03",X"07",X"26",X"06",X"26",X"1B",X"02",X"03",X"04",X"07",X"26",X"29",X"26",X"45",X"03",X"03",
		X"04",X"05",X"26",X"53",X"26",X"67",X"03",X"02",X"04",X"05",X"26",X"71",X"26",X"85",X"03",X"02",
		X"05",X"03",X"26",X"8F",X"26",X"9E",X"04",X"01",X"51",X"11",X"11",X"11",X"50",X"00",X"09",X"A5",
		X"50",X"00",X"00",X"00",X"05",X"51",X"11",X"55",X"00",X"00",X"00",X"00",X"55",X"A0",X"00",X"01",
		X"06",X"03",X"08",X"09",X"A0",X"00",X"00",X"00",X"11",X"50",X"00",X"00",X"00",X"51",X"50",X"00",
		X"00",X"00",X"51",X"10",X"00",X"00",X"00",X"A0",X"00",X"00",X"02",X"04",X"06",X"01",X"03",X"05",
		X"07",X"07",X"15",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"51",X"50",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"05",X"10",X"00",X"01",X"02",X"04",X"05",X"02",X"03",X"05",X"06",X"07",
		X"AA",X"00",X"00",X"00",X"A1",X"A0",X"00",X"00",X"0A",X"1A",X"00",X"00",X"00",X"A1",X"A0",X"00",
		X"00",X"0A",X"1A",X"00",X"00",X"00",X"A1",X"A0",X"00",X"00",X"0A",X"A0",X"00",X"00",X"01",X"02",
		X"03",X"04",X"05",X"02",X"03",X"04",X"05",X"06",X"07",X"07",X"10",X"00",X"00",X"51",X"00",X"00",
		X"01",X"50",X"00",X"00",X"10",X"00",X"00",X"51",X"00",X"00",X"01",X"50",X"00",X"00",X"10",X"00",
		X"00",X"01",X"02",X"02",X"03",X"04",X"01",X"02",X"03",X"03",X"04",X"05",X"05",X"A1",X"00",X"00",
		X"01",X"00",X"00",X"05",X"50",X"00",X"00",X"10",X"00",X"00",X"55",X"00",X"00",X"01",X"00",X"00",
		X"01",X"A0",X"00",X"01",X"01",X"02",X"02",X"03",X"03",X"02",X"02",X"03",X"03",X"04",X"04",X"05",
		X"A0",X"00",X"55",X"00",X"55",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"05",X"50",X"05",X"50",
		X"00",X"A0",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"02",X"02",X"02",
		X"02",X"03",X"03",X"03",X"50",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"A0",X"05",X"50",X"05",X"50",X"01",X"00",X"01",X"00",X"01",X"00",X"55",X"00",X"55",X"00",X"A0",
		X"00",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"03",X"03",X"03",X"02",X"02",X"02",
		X"02",X"02",X"01",X"00",X"01",X"A0",X"00",X"01",X"00",X"00",X"55",X"00",X"00",X"10",X"00",X"05",
		X"50",X"00",X"01",X"00",X"00",X"A1",X"00",X"00",X"03",X"03",X"02",X"02",X"01",X"01",X"00",X"05",
		X"04",X"04",X"03",X"03",X"02",X"02",X"00",X"00",X"10",X"00",X"01",X"50",X"00",X"51",X"00",X"00",
		X"10",X"00",X"01",X"50",X"00",X"51",X"00",X"00",X"10",X"00",X"00",X"04",X"03",X"02",X"02",X"01",
		X"00",X"00",X"05",X"05",X"04",X"03",X"03",X"02",X"01",X"00",X"00",X"0A",X"A0",X"00",X"00",X"A1",
		X"A0",X"00",X"0A",X"1A",X"00",X"00",X"A1",X"A0",X"00",X"0A",X"1A",X"00",X"00",X"A1",X"A0",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"05",X"04",X"03",X"02",X"01",X"00",X"00",X"07",X"07",X"06",X"05",
		X"04",X"03",X"02",X"00",X"00",X"05",X"10",X"00",X"00",X"11",X"00",X"00",X"51",X"50",X"00",X"01",
		X"10",X"00",X"00",X"15",X"00",X"00",X"00",X"05",X"04",X"02",X"01",X"00",X"07",X"06",X"05",X"03",
		X"02",X"00",X"00",X"00",X"A0",X"00",X"00",X"51",X"10",X"00",X"51",X"50",X"00",X"11",X"50",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"06",X"04",X"02",X"00",X"00",X"07",X"07",X"05",X"03",X"01",X"00",
		X"00",X"00",X"55",X"A0",X"05",X"51",X"11",X"55",X"00",X"A5",X"50",X"00",X"00",X"00",X"06",X"01",
		X"00",X"02",X"02",X"26",X"A9",X"26",X"AD",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"02",
		X"02",X"03",X"04",X"26",X"B9",X"26",X"C5",X"01",X"01",X"A1",X"1A",X"00",X"1F",X"F1",X"00",X"1F",
		X"F1",X"00",X"A1",X"1A",X"00",X"01",X"00",X"00",X"01",X"03",X"04",X"04",X"03",X"05",X"0B",X"27",
		X"0E",X"00",X"00",X"05",X"06",X"05",X"0B",X"27",X"45",X"00",X"00",X"05",X"06",X"05",X"08",X"27",
		X"7C",X"00",X"00",X"05",X"04",X"06",X"0B",X"27",X"A4",X"00",X"00",X"06",X"06",X"06",X"09",X"27",
		X"E6",X"00",X"00",X"06",X"05",X"04",X"07",X"28",X"1C",X"00",X"00",X"04",X"04",X"06",X"09",X"28",
		X"38",X"00",X"00",X"06",X"05",X"06",X"0B",X"28",X"6E",X"00",X"00",X"06",X"06",X"00",X"00",X"0A",
		X"65",X"5A",X"00",X"0A",X"66",X"43",X"45",X"00",X"0A",X"36",X"45",X"45",X"00",X"AA",X"65",X"64",
		X"54",X"00",X"AA",X"66",X"6A",X"45",X"50",X"AA",X"A6",X"AA",X"65",X"40",X"0A",X"AA",X"AA",X"A5",
		X"50",X"0A",X"AA",X"AA",X"56",X"60",X"0A",X"AB",X"AA",X"36",X"A0",X"00",X"AA",X"AA",X"AA",X"00",
		X"00",X"0A",X"AA",X"00",X"00",X"00",X"0A",X"55",X"A0",X"00",X"00",X"A4",X"65",X"4A",X"00",X"0A",
		X"AA",X"A4",X"54",X"A0",X"0A",X"AA",X"A5",X"55",X"40",X"AA",X"65",X"AA",X"54",X"40",X"AA",X"A6",
		X"4A",X"55",X"A0",X"AB",X"AA",X"54",X"AA",X"00",X"0A",X"AA",X"34",X"50",X"00",X"0A",X"AA",X"66",
		X"A0",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"0A",X"A0",X"00",X"00",X"00",X"A5",X"44",X"50",
		X"00",X"0A",X"56",X"65",X"54",X"00",X"AA",X"AA",X"A6",X"31",X"50",X"AA",X"AA",X"AA",X"63",X"40",
		X"AB",X"AA",X"AA",X"64",X"50",X"0A",X"AA",X"AA",X"45",X"00",X"00",X"AA",X"A6",X"3A",X"00",X"00",
		X"0A",X"AA",X"A0",X"00",X"00",X"00",X"A4",X"46",X"00",X"00",X"00",X"00",X"A4",X"44",X"A0",X"00",
		X"00",X"0A",X"65",X"A3",X"4A",X"00",X"00",X"0A",X"AA",X"A5",X"5A",X"00",X"0A",X"5A",X"55",X"4A",
		X"6A",X"00",X"A5",X"43",X"5A",X"44",X"A0",X"00",X"A6",X"34",X"AA",X"53",X"40",X"00",X"AA",X"6A",
		X"6A",X"A6",X"A0",X"00",X"AA",X"AA",X"36",X"AA",X"00",X"00",X"AB",X"AA",X"6A",X"00",X"00",X"00",
		X"0A",X"AA",X"A0",X"00",X"00",X"00",X"00",X"0A",X"55",X"A0",X"00",X"00",X"00",X"AA",X"A5",X"44",
		X"00",X"00",X"0A",X"AB",X"A6",X"54",X"4A",X"00",X"AB",X"AA",X"AA",X"65",X"45",X"00",X"AA",X"AA",
		X"AA",X"A6",X"44",X"00",X"AB",X"AB",X"AA",X"A6",X"55",X"00",X"0A",X"AA",X"AA",X"A4",X"5A",X"00",
		X"00",X"AA",X"AA",X"65",X"A0",X"00",X"00",X"0A",X"A6",X"AA",X"00",X"00",X"00",X"05",X"4A",X"00",
		X"00",X"AA",X"44",X"50",X"0A",X"5A",X"44",X"60",X"A5",X"5A",X"55",X"A0",X"A6",X"4A",X"AA",X"00",
		X"0A",X"64",X"A0",X"00",X"00",X"AA",X"00",X"00",X"0A",X"45",X"A0",X"00",X"00",X"00",X"0A",X"45",
		X"5A",X"A0",X"00",X"00",X"A6",X"5A",X"A5",X"45",X"A0",X"00",X"A6",X"AA",X"AA",X"44",X"4A",X"00",
		X"AA",X"AA",X"A6",X"36",X"45",X"A0",X"0A",X"AA",X"A6",X"63",X"55",X"A0",X"0A",X"AA",X"AA",X"A6",
		X"56",X"A0",X"00",X"AA",X"AB",X"AA",X"AA",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",X"00",X"00",
		X"54",X"5A",X"00",X"00",X"00",X"A6",X"55",X"45",X"45",X"00",X"0A",X"65",X"66",X"66",X"53",X"50",
		X"0A",X"64",X"54",X"56",X"54",X"60",X"A6",X"66",X"45",X"44",X"55",X"60",X"A6",X"A6",X"66",X"43",
		X"6A",X"60",X"AB",X"AA",X"A6",X"56",X"AA",X"A0",X"0A",X"AB",X"AA",X"AA",X"AA",X"00",X"00",X"AA",
		X"AA",X"AA",X"AA",X"00",X"00",X"0A",X"AA",X"AA",X"A0",X"00",X"00",X"00",X"AA",X"AA",X"00",X"00",
		X"03",X"03",X"28",X"D0",X"28",X"D9",X"02",X"01",X"03",X"04",X"28",X"DF",X"28",X"EB",X"02",X"02",
		X"02",X"05",X"28",X"F3",X"28",X"FD",X"01",X"02",X"03",X"04",X"29",X"07",X"29",X"13",X"02",X"02",
		X"00",X"D0",X"00",X"CD",X"FD",X"C0",X"00",X"D0",X"00",X"02",X"00",X"02",X"03",X"05",X"03",X"C0",
		X"00",X"00",X"0D",X"F0",X"00",X"0D",X"D0",X"00",X"00",X"0C",X"00",X"00",X"01",X"01",X"03",X"01",
		X"03",X"03",X"04",X"0C",X"00",X"0D",X"00",X"DF",X"D0",X"0D",X"00",X"0C",X"00",X"01",X"01",X"00",
		X"01",X"01",X"02",X"02",X"03",X"02",X"02",X"00",X"0C",X"00",X"0D",X"D0",X"00",X"0D",X"F0",X"00",
		X"C0",X"00",X"00",X"03",X"01",X"01",X"00",X"04",X"03",X"03",X"01",X"04",X"03",X"29",X"3C",X"00",
		X"00",X"03",X"01",X"03",X"04",X"29",X"48",X"00",X"00",X"02",X"02",X"04",X"03",X"29",X"54",X"00",
		X"00",X"03",X"01",X"03",X"04",X"29",X"60",X"00",X"00",X"02",X"02",X"00",X"A1",X"14",X"00",X"00",
		X"0A",X"22",X"14",X"00",X"A4",X"45",X"00",X"00",X"2A",X"0A",X"A0",X"24",X"44",X"A0",X"12",X"4A",
		X"00",X"14",X"A0",X"00",X"A2",X"12",X"26",X"00",X"24",X"12",X"12",X"20",X"A2",X"54",X"46",X"00",
		X"14",X"A0",X"00",X"12",X"2A",X"00",X"11",X"24",X"A0",X"4A",X"0A",X"A0",X"0C",X"13",X"29",X"8C",
		X"00",X"00",X"0C",X"0A",X"0D",X"13",X"2A",X"70",X"00",X"00",X"0D",X"0A",X"0D",X"14",X"2B",X"67",
		X"00",X"00",X"0D",X"0A",X"0D",X"14",X"2C",X"6B",X"00",X"00",X"0D",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"CF",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"DD",X"DD",X"2D",X"DD",X"0D",X"00",X"00",X"00",
		X"00",X"00",X"FD",X"DD",X"DF",X"DF",X"F2",X"FD",X"DD",X"F0",X"00",X"00",X"C0",X"00",X"0C",X"DF",
		X"F2",X"F2",X"22",X"FF",X"2D",X"00",X"D0",X"00",X"00",X"00",X"0D",X"DF",X"F2",X"21",X"12",X"22",
		X"FF",X"DD",X"00",X"00",X"0D",X"0D",X"0D",X"FF",X"22",X"12",X"11",X"12",X"2F",X"D0",X"CF",X"00",
		X"00",X"00",X"CD",X"F2",X"22",X"11",X"11",X"11",X"F2",X"FD",X"D0",X"00",X"00",X"0C",X"DF",X"F2",
		X"11",X"11",X"11",X"11",X"22",X"FF",X"D0",X"00",X"00",X"DD",X"F2",X"21",X"11",X"11",X"11",X"11",
		X"12",X"2F",X"FC",X"D0",X"00",X"0C",X"DF",X"F2",X"11",X"11",X"11",X"11",X"22",X"FF",X"DC",X"00",
		X"00",X"0C",X"DD",X"F2",X"F1",X"11",X"11",X"12",X"2F",X"DD",X"D0",X"00",X"00",X"00",X"DC",X"DF",
		X"2F",X"11",X"11",X"1F",X"2F",X"DD",X"0C",X"00",X"00",X"0D",X"00",X"D2",X"F2",X"21",X"11",X"22",
		X"FD",X"CF",X"00",X"00",X"00",X"00",X"00",X"DD",X"DF",X"22",X"12",X"2F",X"2D",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"DD",X"FF",X"2F",X"FD",X"DF",X"F0",X"00",X"00",X"00",X"00",X"0C",X"FC",
		X"0D",X"DD",X"FF",X"DD",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0C",X"DD",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"C0",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"BC",X"DC",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"BC",X"CC",
		X"DD",X"BC",X"00",X"0B",X"00",X"00",X"00",X"00",X"0D",X"CD",X"CC",X"CC",X"DD",X"FD",X"CC",X"CB",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"0C",X"DB",X"CD",X"DD",X"2D",X"DD",X"DC",X"00",X"D0",X"00",
		X"00",X"C0",X"00",X"0B",X"CC",X"DD",X"DF",X"22",X"FD",X"DC",X"CB",X"00",X"0C",X"00",X"00",X"0D",
		X"0D",X"CD",X"DD",X"22",X"22",X"2F",X"D2",X"C0",X"BB",X"00",X"00",X"00",X"00",X"BC",X"DD",X"22",
		X"22",X"2F",X"22",X"2D",X"CB",X"D0",X"00",X"00",X"00",X"0B",X"BC",X"DD",X"DF",X"2F",X"FF",X"22",
		X"DD",X"DD",X"B0",X"00",X"00",X"0C",X"0D",X"CD",X"D2",X"22",X"2F",X"DF",X"F2",X"22",X"FD",X"DB",
		X"DB",X"00",X"00",X"0C",X"BC",X"DD",X"DF",X"2F",X"FF",X"22",X"2F",X"DC",X"BB",X"00",X"00",X"00",
		X"0B",X"CD",X"CD",X"22",X"F2",X"F2",X"22",X"DD",X"DB",X"D0",X"00",X"00",X"00",X"00",X"DB",X"CD",
		X"DD",X"22",X"22",X"2F",X"DC",X"BB",X"0B",X"00",X"00",X"00",X"00",X"00",X"CC",X"D2",X"F2",X"2F",
		X"22",X"DD",X"B0",X"C0",X"00",X"00",X"00",X"00",X"00",X"DD",X"DD",X"DD",X"2D",X"FD",X"CD",X"C0",
		X"00",X"00",X"00",X"0C",X"00",X"00",X"0C",X"CC",X"CD",X"DD",X"DC",X"DD",X"B0",X"0C",X"00",X"00",
		X"00",X"00",X"BB",X"0B",X"0C",X"DD",X"DC",X"CB",X"B0",X"0D",X"00",X"00",X"00",X"00",X"00",X"BD",
		X"0B",X"0D",X"0B",X"DC",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
		X"BB",X"C0",X"B0",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0B",X"CB",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"0B",X"BC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"BC",X"BC",X"CC",X"DC",X"BC",X"00",X"CB",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"CC",X"CC",X"CD",X"DC",X"CC",X"CB",X"B0",X"0C",X"00",X"00",X"00",X"00",X"0C",X"DB",X"CD",
		X"DD",X"FD",X"CC",X"DC",X"00",X"B0",X"00",X"A0",X"A0",X"00",X"0B",X"CC",X"DD",X"DD",X"FF",X"DD",
		X"CC",X"CB",X"00",X"00",X"00",X"00",X"C0",X"0C",X"CC",X"DD",X"CF",X"00",X"FF",X"DC",X"C0",X"BB",
		X"00",X"00",X"00",X"00",X"BC",X"CD",X"DD",X"FF",X"00",X"0F",X"DD",X"CB",X"B0",X"00",X"00",X"00",
		X"0B",X"BC",X"CD",X"DD",X"F0",X"00",X"00",X"FC",X"CC",X"B0",X"00",X"00",X"0B",X"C0",X"CD",X"DD",
		X"DF",X"00",X"00",X"0F",X"DD",X"DD",X"DB",X"CB",X"00",X"00",X"0C",X"BC",X"CD",X"DD",X"F0",X"00",
		X"0F",X"DD",X"DC",X"BB",X"00",X"00",X"00",X"0B",X"CC",X"CD",X"DF",X"F0",X"00",X"FF",X"DD",X"CB",
		X"C0",X"00",X"00",X"00",X"00",X"0B",X"CC",X"DD",X"DF",X"0F",X"FD",X"DC",X"BB",X"0B",X"00",X"00",
		X"00",X"0C",X"00",X"CC",X"DD",X"DD",X"FD",X"DD",X"DC",X"B0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"CC",X"DD",X"DD",X"DC",X"CD",X"C0",X"00",X"00",X"00",X"A0",X"00",X"0C",X"0C",X"CC",X"CC",
		X"DD",X"CC",X"CB",X"B0",X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"0C",X"DC",X"DC",X"CB",X"B0",
		X"CB",X"00",X"A0",X"00",X"00",X"00",X"B0",X"0B",X"00",X"0B",X"CC",X"00",X"00",X"00",X"C0",X"00",
		X"00",X"00",X"00",X"C0",X"00",X"0C",X"00",X"BB",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"B0",X"0B",X"00",X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",
		X"0A",X"BA",X"00",X"00",X"0A",X"00",X"0A",X"00",X"00",X"0A",X"00",X"00",X"0B",X"0B",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"B0",X"00",X"00",X"BB",X"0B",X"0B",X"00",
		X"A0",X"00",X"00",X"00",X"AB",X"00",X"00",X"D0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"B0",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0B",X"0A",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"0A",X"B0",X"00",X"00",X"00",X"00",X"00",X"0B",X"0B",X"00",X"00",X"A0",X"00",
		X"0B",X"00",X"0C",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"0B",
		X"B0",X"00",X"0B",X"00",X"BB",X"00",X"A0",X"00",X"00",X"00",X"A0",X"0B",X"00",X"0A",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"0A",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"90",X"00",
		X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",
		X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",
		X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",
		X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",
		X"00",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"90",X"0A",X"50",X"00",X"0A",X"22",X"00",X"05",
		X"11",X"24",X"0A",X"65",X"00",X"0A",X"60",X"00",X"09",X"22",X"90",X"02",X"99",X"20",X"02",X"99",
		X"20",X"09",X"22",X"90",X"00",X"00",X"00",X"01",X"10",X"01",X"10",X"BD",X"65",X"03",X"7D",X"A1",
		X"BB",X"27",X"07",X"BD",X"68",X"CC",X"25",X"02",X"4F",X"5F",X"39",X"49",X"4C",X"4C",X"49",X"41",
		X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",
		X"49",X"4E",X"43",X"2E",X"E1",X"95",X"E1",X"95",X"E1",X"95",X"E1",X"95",X"6C",X"83",X"2E",X"E3",
		X"6C",X"8A",X"2F",X"0D",X"E1",X"95",X"E1",X"95",X"E1",X"95",X"E1",X"95",X"6D",X"7D",X"6C",X"F6",
		X"6C",X"CA",X"6C",X"BA",X"39",X"10",X"CE",X"BF",X"00",X"86",X"98",X"1F",X"8B",X"4F",X"5F",X"97",
		X"39",X"B7",X"CA",X"01",X"97",X"54",X"97",X"57",X"B7",X"DC",X"77",X"B7",X"DC",X"79",X"97",X"5A",
		X"FD",X"9F",X"F6",X"FD",X"9F",X"F8",X"FD",X"9F",X"FA",X"97",X"8A",X"B7",X"BF",X"1C",X"7E",X"8E",
		X"49",X"8E",X"C8",X"00",X"A7",X"05",X"A7",X"07",X"A7",X"0D",X"A7",X"0F",X"C6",X"34",X"E7",X"05",
		X"E7",X"07",X"86",X"3F",X"ED",X"0E",X"CC",X"80",X"05",X"ED",X"0C",X"A7",X"0C",X"39",X"C8",X"06",
		X"97",X"58",X"B6",X"C8",X"0C",X"97",X"59",X"CC",X"45",X"66",X"DD",X"76",X"CC",X"50",X"23",X"DD",
		X"7D",X"CC",X"F1",X"F0",X"DD",X"5B",X"8E",X"CD",X"00",X"BD",X"4A",X"5F",X"81",X"20",X"23",X"01",
		X"4F",X"B7",X"BF",X"1B",X"30",X"1E",X"BD",X"4A",X"78",X"86",X"FF",X"8E",X"CD",X"22",X"BD",X"4A",
		X"70",X"DD",X"30",X"BD",X"4A",X"70",X"DD",X"2E",X"86",X"30",X"97",X"80",X"BD",X"52",X"A4",X"BD",
		X"31",X"49",X"0F",X"96",X"BD",X"31",X"49",X"BD",X"51",X"4F",X"10",X"CE",X"BF",X"00",X"1C",X"EF",
		X"7E",X"34",X"5E",X"8E",X"CC",X"0C",X"BD",X"4A",X"5F",X"81",X"09",X"27",X"08",X"B6",X"BF",X"1B",
		X"81",X"02",X"24",X"01",X"39",X"0F",X"96",X"BD",X"32",X"45",X"86",X"02",X"97",X"8A",X"86",X"13",
		X"BD",X"30",X"AC",X"BD",X"33",X"45",X"86",X"B4",X"BD",X"30",X"AC",X"20",X"1E",X"8E",X"CC",X"0C",
		X"BD",X"4A",X"5F",X"81",X"09",X"27",X"06",X"B6",X"BF",X"1B",X"26",X"01",X"39",X"0F",X"96",X"BD",
		X"32",X"45",X"86",X"01",X"97",X"8A",X"86",X"13",X"BD",X"30",X"AC",X"4F",X"5F",X"97",X"80",X"CC",
		X"FC",X"7A",X"DD",X"69",X"DD",X"67",X"86",X"01",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"86",X"05",
		X"B7",X"CA",X"06",X"86",X"01",X"97",X"00",X"BD",X"32",X"FA",X"96",X"00",X"8B",X"09",X"81",X"35",
		X"25",X"F3",X"7F",X"CA",X"01",X"86",X"05",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"BD",X"32",X"0F",
		X"BD",X"51",X"45",X"B6",X"9F",X"FC",X"C6",X"02",X"BD",X"3C",X"0C",X"BD",X"3C",X"74",X"BD",X"31",
		X"49",X"BD",X"46",X"DB",X"2F",X"7C",X"08",X"A1",X"5F",X"7E",X"2E",X"DA",X"96",X"8A",X"4A",X"27",
		X"36",X"B6",X"9F",X"FC",X"26",X"27",X"BD",X"32",X"0C",X"B6",X"A0",X"99",X"27",X"2E",X"BD",X"31",
		X"D8",X"34",X"20",X"8E",X"49",X"60",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"4D",X"BD",X"E2",X"03",
		X"86",X"4E",X"BD",X"E2",X"03",X"35",X"20",X"CC",X"00",X"B4",X"BD",X"34",X"19",X"B6",X"A0",X"99",
		X"27",X"3F",X"BD",X"33",X"45",X"20",X"3A",X"B6",X"9F",X"FC",X"26",X"35",X"B6",X"A0",X"0A",X"2A",
		X"03",X"BD",X"33",X"45",X"34",X"20",X"BD",X"38",X"91",X"4D",X"F2",X"8E",X"49",X"60",X"BD",X"2E",
		X"44",X"C6",X"DD",X"86",X"4D",X"BD",X"E2",X"03",X"86",X"4E",X"BD",X"E2",X"03",X"86",X"30",X"97",
		X"80",X"7E",X"87",X"84",X"33",X"8E",X"35",X"20",X"CC",X"01",X"2C",X"BD",X"34",X"19",X"7E",X"2E",
		X"D4",X"34",X"20",X"BD",X"32",X"0F",X"BD",X"31",X"D8",X"7E",X"85",X"60",X"BD",X"32",X"0F",X"4F",
		X"5F",X"DD",X"44",X"DD",X"46",X"97",X"48",X"DD",X"49",X"97",X"4B",X"DD",X"4C",X"DD",X"4E",X"97",
		X"61",X"FD",X"A1",X"3E",X"FD",X"A1",X"40",X"97",X"7F",X"97",X"95",X"97",X"85",X"97",X"86",X"8E",
		X"9F",X"60",X"CE",X"4F",X"A0",X"86",X"00",X"BD",X"48",X"02",X"34",X"02",X"CC",X"02",X"74",X"BD",
		X"47",X"FA",X"35",X"04",X"ED",X"84",X"A6",X"C0",X"A7",X"02",X"6F",X"03",X"30",X"04",X"8C",X"9F",
		X"88",X"25",X"E2",X"BD",X"46",X"BB",X"3C",X"65",X"A1",X"74",X"CC",X"4B",X"C3",X"FD",X"A1",X"3C",
		X"BD",X"43",X"22",X"BF",X"A1",X"42",X"CC",X"27",X"7A",X"ED",X"05",X"E7",X"07",X"4F",X"5F",X"ED",
		X"0C",X"ED",X"0E",X"97",X"50",X"BD",X"43",X"5E",X"CC",X"A1",X"38",X"ED",X"88",X"1C",X"FD",X"A1",
		X"36",X"FD",X"A1",X"38",X"BD",X"46",X"DB",X"3F",X"74",X"06",X"A1",X"74",X"DC",X"48",X"F0",X"99",
		X"05",X"82",X"00",X"47",X"56",X"E7",X"04",X"DC",X"4B",X"F0",X"99",X"07",X"82",X"00",X"47",X"56",
		X"47",X"56",X"E7",X"05",X"BD",X"32",X"7E",X"BD",X"33",X"B4",X"BD",X"51",X"89",X"86",X"0F",X"0D",
		X"96",X"27",X"02",X"86",X"38",X"97",X"80",X"35",X"20",X"7E",X"47",X"55",X"B7",X"A0",X"0A",X"4F",
		X"5F",X"B7",X"A0",X"13",X"FD",X"9F",X"FD",X"FD",X"9F",X"FF",X"FD",X"A0",X"06",X"FD",X"A0",X"08",
		X"B7",X"A0",X"12",X"FD",X"A0",X"01",X"B7",X"A0",X"05",X"FD",X"A0",X"0C",X"8E",X"CC",X"00",X"BD",
		X"4A",X"5F",X"5F",X"BD",X"48",X"EA",X"FD",X"A0",X"0E",X"FD",X"A0",X"03",X"BD",X"4A",X"5F",X"5F",
		X"BD",X"48",X"EA",X"FD",X"A0",X"10",X"BD",X"4A",X"70",X"BD",X"4B",X"89",X"1F",X"98",X"B7",X"9F",
		X"FC",X"C6",X"02",X"BD",X"3C",X"0C",X"4A",X"26",X"FA",X"86",X"FF",X"B7",X"A0",X"09",X"BD",X"3C",
		X"74",X"86",X"81",X"F6",X"A0",X"0A",X"1F",X"01",X"C6",X"99",X"86",X"4F",X"BD",X"E2",X"0C",X"86",
		X"50",X"BD",X"E2",X"0C",X"BD",X"3B",X"C0",X"CC",X"50",X"02",X"FD",X"A0",X"16",X"CC",X"4F",X"B2",
		X"FD",X"A0",X"14",X"96",X"96",X"26",X"1E",X"8E",X"CC",X"0C",X"BD",X"4A",X"5F",X"81",X"09",X"27",
		X"14",X"B6",X"BF",X"1B",X"8B",X"99",X"19",X"B7",X"BF",X"1B",X"8E",X"CD",X"00",X"BD",X"4A",X"78",
		X"C6",X"08",X"BD",X"4A",X"8E",X"BD",X"52",X"9D",X"39",X"34",X"01",X"1A",X"10",X"97",X"3F",X"8E",
		X"98",X"1E",X"EC",X"89",X"B8",X"AD",X"ED",X"81",X"8C",X"98",X"2E",X"25",X"F5",X"8E",X"99",X"00",
		X"9F",X"3D",X"30",X"88",X"22",X"AF",X"88",X"DE",X"8C",X"9F",X"3E",X"26",X"F5",X"4F",X"5F",X"ED",
		X"84",X"8E",X"A2",X"25",X"9F",X"3B",X"30",X"02",X"AF",X"1E",X"8C",X"A5",X"23",X"25",X"F7",X"4F",
		X"5F",X"ED",X"84",X"DD",X"33",X"DD",X"88",X"97",X"32",X"CC",X"A5",X"25",X"DD",X"6B",X"CC",X"BE",
		X"C0",X"DD",X"6D",X"86",X"FF",X"97",X"71",X"86",X"30",X"97",X"75",X"CC",X"18",X"8B",X"DD",X"73",
		X"8E",X"A1",X"5F",X"CC",X"46",X"7B",X"ED",X"84",X"AF",X"02",X"33",X"02",X"EF",X"04",X"6F",X"06",
		X"30",X"07",X"8C",X"A1",X"9E",X"26",X"EF",X"CC",X"46",X"9E",X"ED",X"84",X"AF",X"02",X"33",X"02",
		X"EF",X"04",X"86",X"01",X"A7",X"06",X"CC",X"A1",X"9E",X"DD",X"40",X"CC",X"A1",X"A0",X"DD",X"42",
		X"BD",X"E2",X"22",X"12",X"12",X"12",X"35",X"81",X"34",X"36",X"96",X"8A",X"4A",X"27",X"2B",X"B6",
		X"A0",X"0A",X"2B",X"14",X"8E",X"60",X"66",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"51",X"BD",X"E2",
		X"03",X"86",X"52",X"BD",X"E2",X"03",X"20",X"12",X"8E",X"60",X"66",X"BD",X"2E",X"44",X"C6",X"DD",
		X"86",X"51",X"BD",X"E2",X"03",X"86",X"53",X"BD",X"E2",X"03",X"35",X"B6",X"7E",X"8C",X"74",X"34",
		X"06",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"CC",X"1C",
		X"35",X"FD",X"CA",X"06",X"CC",X"75",X"68",X"FD",X"CA",X"02",X"FD",X"CA",X"04",X"C6",X"12",X"F7",
		X"CA",X"00",X"86",X"05",X"B7",X"CA",X"06",X"86",X"8D",X"B7",X"CA",X"04",X"86",X"52",X"B7",X"CA",
		X"00",X"86",X"73",X"20",X"11",X"34",X"06",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"86",X"97",X"C6",X"05",X"F7",X"CA",X"06",X"C6",X"FB",X"F7",X"CA",X"07",
		X"7F",X"CA",X"05",X"B7",X"CA",X"04",X"C6",X"12",X"F7",X"CA",X"00",X"C6",X"39",X"F7",X"CB",X"FF",
		X"80",X"01",X"24",X"EF",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"86",X"34",X"16",
		X"CC",X"D7",X"7C",X"FD",X"CA",X"02",X"FD",X"CA",X"04",X"CC",X"1E",X"35",X"FD",X"CA",X"06",X"B6",
		X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"86",X"10",X"B7",X"CA",
		X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"8E",X"9F",X"94",X"86",X"4B",X"C6",X"31",
		X"BD",X"32",X"F0",X"40",X"BD",X"32",X"F0",X"FC",X"A0",X"14",X"34",X"06",X"FC",X"A0",X"16",X"10",
		X"83",X"4F",X"E2",X"26",X"15",X"FD",X"A0",X"14",X"8E",X"50",X"02",X"BF",X"A0",X"16",X"BD",X"3D",
		X"4E",X"10",X"B3",X"A0",X"14",X"25",X"F7",X"FD",X"A0",X"16",X"8E",X"4F",X"B2",X"BD",X"3D",X"7E",
		X"AC",X"E4",X"27",X"08",X"BD",X"3D",X"4E",X"BE",X"A0",X"14",X"20",X"F4",X"32",X"62",X"35",X"96",
		X"3A",X"34",X"14",X"A7",X"82",X"5A",X"26",X"FB",X"35",X"94",X"CC",X"14",X"66",X"8D",X"09",X"96",
		X"00",X"8B",X"03",X"97",X"00",X"CC",X"11",X"AA",X"F7",X"CA",X"01",X"8D",X"04",X"4A",X"26",X"FB",
		X"39",X"34",X"02",X"81",X"11",X"23",X"02",X"86",X"11",X"34",X"02",X"48",X"8B",X"35",X"88",X"04",
		X"B7",X"CA",X"07",X"C6",X"66",X"E0",X"E0",X"A6",X"E4",X"9B",X"00",X"46",X"34",X"01",X"8B",X"74",
		X"81",X"98",X"23",X"01",X"4F",X"FD",X"CA",X"04",X"86",X"52",X"35",X"01",X"24",X"02",X"86",X"92",
		X"B7",X"CA",X"00",X"35",X"82",X"34",X"72",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"8E",X"05",X"99",X"BF",X"CA",X"06",X"8E",X"A0",X"99",X"BF",X"CA",X"02",
		X"10",X"8E",X"D7",X"7C",X"10",X"BF",X"CA",X"04",X"86",X"04",X"B7",X"CA",X"00",X"CE",X"9F",X"FC",
		X"FF",X"CA",X"02",X"BF",X"CA",X"04",X"B7",X"CA",X"00",X"12",X"10",X"BF",X"CA",X"02",X"FF",X"CA",
		X"04",X"7F",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"F2",X"34",X"16",
		X"96",X"8A",X"26",X"1E",X"7D",X"BF",X"1B",X"27",X"19",X"8E",X"10",X"6D",X"BD",X"2E",X"44",X"C6",
		X"11",X"86",X"54",X"BD",X"E2",X"0C",X"B6",X"BF",X"1B",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",
		X"E2",X"0F",X"35",X"96",X"34",X"06",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",
		X"B7",X"C9",X"00",X"CC",X"05",X"FB",X"FD",X"CA",X"06",X"CC",X"74",X"00",X"FD",X"CA",X"04",X"B6",
		X"A0",X"18",X"B7",X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",X"C6",X"31",X"F7",X"CA",X"07",X"CC",
		X"8E",X"66",X"FD",X"CA",X"04",X"C6",X"52",X"F7",X"CA",X"00",X"86",X"8D",X"B7",X"CA",X"04",X"C6",
		X"92",X"F7",X"CA",X"00",X"CC",X"1D",X"06",X"FD",X"CA",X"06",X"86",X"75",X"B7",X"CA",X"04",X"C6",
		X"12",X"F7",X"CA",X"00",X"86",X"99",X"B7",X"CA",X"05",X"F7",X"CA",X"00",X"35",X"02",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"7F",X"CA",X"01",X"35",X"86",X"ED",X"24",X"35",X"06",X"ED",X"26",X"CC",
		X"34",X"29",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"EC",X"24",X"83",X"00",X"01",X"ED",X"24",
		X"26",X"ED",X"6E",X"B8",X"06",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",
		X"39",X"38",X"33",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",
		X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"0A",X"32",
		X"2F",X"03",X"7E",X"37",X"F0",X"2A",X"0E",X"AE",X"9F",X"98",X"42",X"10",X"AE",X"94",X"AD",X"B8",
		X"02",X"96",X"32",X"2B",X"F2",X"BD",X"35",X"3E",X"10",X"9E",X"33",X"26",X"32",X"20",X"DF",X"AE",
		X"22",X"27",X"27",X"A6",X"26",X"A1",X"06",X"24",X"21",X"EE",X"A4",X"DF",X"00",X"EF",X"84",X"AF",
		X"42",X"AE",X"02",X"A1",X"06",X"25",X"FA",X"EE",X"84",X"10",X"AF",X"84",X"AF",X"22",X"EF",X"A4",
		X"10",X"AF",X"42",X"10",X"9E",X"00",X"26",X"07",X"20",X"B4",X"10",X"AE",X"A4",X"27",X"AF",X"E6",
		X"26",X"EB",X"2B",X"24",X"02",X"C6",X"FF",X"D7",X"3A",X"A6",X"B8",X"12",X"2B",X"32",X"AE",X"A4",
		X"E1",X"06",X"23",X"2C",X"A6",X"A8",X"11",X"A1",X"05",X"2F",X"1F",X"A6",X"25",X"A1",X"88",X"11",
		X"2C",X"18",X"EE",X"88",X"12",X"EC",X"42",X"A4",X"B8",X"12",X"26",X"09",X"D7",X"00",X"EC",X"B8",
		X"12",X"D4",X"00",X"27",X"03",X"BD",X"39",X"8E",X"D6",X"3A",X"AE",X"84",X"E1",X"06",X"22",X"D4",
		X"96",X"32",X"2E",X"47",X"96",X"3A",X"8B",X"20",X"25",X"2D",X"B1",X"CB",X"00",X"25",X"3C",X"10",
		X"9F",X"1C",X"AE",X"9F",X"98",X"42",X"10",X"AE",X"94",X"AD",X"B8",X"02",X"96",X"32",X"2E",X"28",
		X"96",X"3A",X"8B",X"20",X"25",X"14",X"B1",X"CB",X"00",X"25",X"1D",X"AE",X"9F",X"98",X"42",X"10",
		X"AE",X"94",X"AD",X"B8",X"02",X"20",X"E5",X"10",X"9F",X"1C",X"AE",X"9F",X"98",X"42",X"10",X"AE",
		X"94",X"AD",X"B8",X"02",X"96",X"32",X"2F",X"F2",X"10",X"9E",X"1C",X"6E",X"B8",X"18",X"DE",X"40",
		X"DC",X"42",X"ED",X"44",X"0C",X"3F",X"27",X"1F",X"8E",X"A1",X"5F",X"C6",X"07",X"96",X"3F",X"3A",
		X"44",X"24",X"FC",X"A6",X"06",X"4C",X"26",X"01",X"3F",X"A7",X"06",X"A1",X"46",X"25",X"08",X"26",
		X"04",X"9C",X"40",X"24",X"02",X"33",X"84",X"B6",X"A1",X"65",X"4C",X"26",X"01",X"3F",X"B7",X"A1",
		X"65",X"A1",X"46",X"25",X"03",X"CE",X"A1",X"5F",X"DF",X"40",X"EC",X"44",X"DD",X"42",X"BD",X"38",
		X"07",X"96",X"54",X"27",X"09",X"0A",X"54",X"26",X"05",X"DE",X"55",X"BD",X"38",X"BA",X"86",X"00",
		X"BD",X"48",X"08",X"86",X"02",X"BD",X"48",X"02",X"84",X"06",X"8E",X"4F",X"98",X"EC",X"86",X"DD",
		X"76",X"BD",X"37",X"DA",X"96",X"8A",X"26",X"01",X"39",X"0F",X"53",X"CC",X"22",X"22",X"FD",X"81",
		X"80",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"CC",X"03",
		X"0A",X"FD",X"CA",X"06",X"CC",X"2D",X"77",X"FD",X"CA",X"02",X"DC",X"67",X"10",X"93",X"69",X"27",
		X"17",X"DD",X"00",X"DC",X"69",X"8B",X"03",X"46",X"FD",X"CA",X"04",X"86",X"1A",X"24",X"02",X"8A",
		X"20",X"B7",X"CA",X"00",X"DC",X"00",X"DD",X"69",X"8B",X"03",X"46",X"FD",X"CA",X"04",X"86",X"1A",
		X"24",X"02",X"8A",X"20",X"F6",X"A0",X"18",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"02",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"7F",X"CA",X"01",X"BD",X"51",X"08",X"10",X"8E",X"99",X"00",X"96",
		X"80",X"85",X"04",X"10",X"27",X"00",X"AC",X"8E",X"4E",X"01",X"B6",X"C8",X"04",X"84",X"70",X"44",
		X"44",X"44",X"44",X"E6",X"86",X"58",X"58",X"D7",X"00",X"B6",X"C8",X"04",X"84",X"07",X"E6",X"86",
		X"DA",X"00",X"10",X"27",X"00",X"8D",X"8E",X"4E",X"09",X"EC",X"85",X"97",X"53",X"B6",X"C8",X"04",
		X"2B",X"01",X"50",X"85",X"08",X"26",X"03",X"50",X"CB",X"80",X"D0",X"50",X"96",X"53",X"D7",X"00",
		X"3D",X"2A",X"02",X"90",X"53",X"C3",X"00",X"80",X"1F",X"89",X"9B",X"50",X"97",X"50",X"BD",X"47",
		X"DA",X"DD",X"51",X"D6",X"00",X"CB",X"20",X"C1",X"40",X"24",X"58",X"D6",X"52",X"1D",X"58",X"49",
		X"58",X"49",X"A3",X"2E",X"97",X"00",X"96",X"53",X"3D",X"97",X"02",X"96",X"53",X"D6",X"00",X"3D",
		X"2A",X"02",X"90",X"53",X"DB",X"02",X"89",X"00",X"47",X"56",X"47",X"56",X"47",X"56",X"C9",X"00",
		X"89",X"00",X"E3",X"2E",X"ED",X"2E",X"D6",X"51",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"A3",
		X"2C",X"97",X"00",X"96",X"53",X"3D",X"97",X"02",X"96",X"53",X"D6",X"00",X"3D",X"2A",X"02",X"90",
		X"53",X"DB",X"02",X"89",X"00",X"47",X"56",X"47",X"56",X"47",X"56",X"C9",X"00",X"89",X"00",X"E3",
		X"2C",X"ED",X"2C",X"96",X"80",X"85",X"08",X"26",X"01",X"39",X"A6",X"25",X"E6",X"26",X"E3",X"2E",
		X"D3",X"44",X"81",X"08",X"25",X"04",X"81",X"6C",X"25",X"08",X"EC",X"2E",X"43",X"50",X"82",X"FF",
		X"DD",X"44",X"EC",X"2C",X"D3",X"46",X"E3",X"27",X"81",X"10",X"25",X"04",X"81",X"F0",X"25",X"08",
		X"EC",X"2C",X"43",X"50",X"82",X"FF",X"DD",X"46",X"DC",X"51",X"47",X"47",X"47",X"57",X"57",X"57",
		X"DD",X"00",X"C6",X"7B",X"E0",X"27",X"57",X"D0",X"00",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",
		X"A3",X"2C",X"93",X"46",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"34",X"06",
		X"47",X"56",X"E3",X"E1",X"D3",X"46",X"DD",X"46",X"C6",X"38",X"E0",X"25",X"D0",X"01",X"1D",X"58",
		X"49",X"58",X"49",X"58",X"49",X"A3",X"2E",X"93",X"44",X"47",X"56",X"47",X"56",X"47",X"56",X"47",
		X"56",X"47",X"56",X"34",X"06",X"47",X"56",X"E3",X"E1",X"D3",X"44",X"DD",X"44",X"DC",X"44",X"2A",
		X"08",X"D3",X"49",X"25",X"0A",X"0A",X"48",X"20",X"06",X"D3",X"49",X"24",X"02",X"0C",X"48",X"DD",
		X"49",X"DC",X"46",X"2A",X"08",X"D3",X"4C",X"25",X"0A",X"0A",X"4B",X"20",X"06",X"D3",X"4C",X"24",
		X"02",X"0C",X"4B",X"DD",X"4C",X"D6",X"50",X"CB",X"04",X"C4",X"F8",X"8E",X"00",X"07",X"3A",X"AC",
		X"A8",X"14",X"27",X"09",X"AF",X"A8",X"16",X"8E",X"43",X"B8",X"AF",X"A8",X"18",X"A6",X"25",X"44",
		X"40",X"97",X"65",X"8B",X"3A",X"97",X"63",X"A6",X"27",X"44",X"44",X"40",X"97",X"66",X"8B",X"3F",
		X"97",X"64",X"0A",X"85",X"2A",X"05",X"CC",X"1D",X"12",X"20",X"07",X"0A",X"85",X"2A",X"0B",X"CC",
		X"1C",X"02",X"97",X"85",X"B6",X"9F",X"FC",X"BD",X"3C",X"0C",X"96",X"86",X"27",X"1B",X"0A",X"86",
		X"26",X"17",X"BD",X"39",X"1D",X"8E",X"CC",X"08",X"BD",X"4A",X"5F",X"27",X"0C",X"96",X"87",X"81",
		X"0A",X"24",X"04",X"8B",X"00",X"97",X"87",X"97",X"86",X"39",X"B6",X"C8",X"06",X"97",X"00",X"98",
		X"58",X"94",X"80",X"26",X"01",X"39",X"D6",X"00",X"D7",X"58",X"8E",X"2E",X"24",X"7E",X"E1",X"46",
		X"86",X"FF",X"12",X"12",X"0A",X"32",X"7E",X"34",X"5E",X"9F",X"00",X"8D",X"0A",X"9E",X"00",X"DE",
		X"88",X"4F",X"5F",X"DD",X"88",X"6E",X"C4",X"9E",X"6D",X"8C",X"BE",X"C0",X"25",X"19",X"9E",X"71",
		X"8C",X"BE",X"C0",X"24",X"6D",X"30",X"1C",X"9F",X"6D",X"EC",X"84",X"33",X"8B",X"DF",X"6F",X"D3",
		X"73",X"DD",X"73",X"86",X"FF",X"97",X"71",X"BF",X"CA",X"04",X"DE",X"6F",X"11",X"93",X"6B",X"24",
		X"0E",X"A6",X"42",X"26",X"13",X"EC",X"C4",X"33",X"CB",X"D3",X"73",X"DD",X"73",X"20",X"ED",X"9F",
		X"6B",X"CC",X"BE",X"C0",X"DD",X"6D",X"20",X"3A",X"FF",X"CA",X"02",X"DC",X"6D",X"C3",X"00",X"04",
		X"ED",X"D8",X"02",X"EC",X"C4",X"30",X"8B",X"9F",X"6D",X"33",X"CB",X"DF",X"6F",X"4D",X"27",X"01",
		X"3F",X"86",X"05",X"C8",X"04",X"FD",X"CA",X"06",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"C6",X"04",X"F7",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"96",X"73",X"2A",X"0A",X"9E",X"71",X"8C",X"BE",X"C0",X"10",X"25",X"FF",X"78",X"3F",
		X"39",X"34",X"56",X"AE",X"66",X"EE",X"81",X"AF",X"66",X"96",X"96",X"27",X"06",X"11",X"83",X"4D",
		X"FC",X"26",X"15",X"A6",X"C0",X"91",X"57",X"23",X"0F",X"4F",X"B7",X"9F",X"88",X"B7",X"9F",X"8B",
		X"B7",X"9F",X"8E",X"B7",X"9F",X"91",X"8D",X"02",X"35",X"D6",X"A6",X"C4",X"85",X"C0",X"26",X"3E",
		X"4D",X"26",X"0D",X"0F",X"57",X"86",X"FF",X"B7",X"C8",X"0E",X"86",X"01",X"B7",X"C8",X"0E",X"39",
		X"8E",X"9F",X"88",X"11",X"A3",X"84",X"27",X"16",X"30",X"03",X"8C",X"9F",X"94",X"26",X"F4",X"8E",
		X"9F",X"88",X"E6",X"84",X"27",X"04",X"30",X"03",X"20",X"F8",X"EF",X"84",X"A7",X"02",X"6A",X"02",
		X"27",X"06",X"A6",X"41",X"33",X"C6",X"20",X"C2",X"6F",X"84",X"33",X"42",X"20",X"BC",X"2A",X"10",
		X"C6",X"FF",X"F7",X"C8",X"0E",X"B7",X"C8",X"0E",X"33",X"41",X"85",X"40",X"27",X"AC",X"20",X"06",
		X"A6",X"C0",X"84",X"3F",X"97",X"57",X"A6",X"C0",X"97",X"54",X"DF",X"55",X"39",X"BD",X"38",X"91",
		X"4D",X"AE",X"96",X"75",X"27",X"67",X"BD",X"43",X"4F",X"CC",X"4D",X"11",X"ED",X"88",X"12",X"D6",
		X"50",X"CB",X"04",X"C4",X"78",X"4F",X"C3",X"24",X"38",X"1F",X"03",X"BD",X"43",X"32",X"96",X"50",
		X"BD",X"47",X"DA",X"34",X"02",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"F3",X"99",X"0E",X"ED",
		X"0E",X"35",X"04",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"F3",X"99",X"0C",X"ED",
		X"0C",X"10",X"BE",X"99",X"14",X"A6",X"26",X"A0",X"46",X"5F",X"47",X"56",X"34",X"06",X"FC",X"99",
		X"07",X"AB",X"27",X"A0",X"47",X"ED",X"07",X"A7",X"06",X"35",X"06",X"F9",X"99",X"04",X"B9",X"99",
		X"05",X"A7",X"05",X"E7",X"04",X"AB",X"C4",X"A7",X"88",X"11",X"BD",X"43",X"5E",X"39",X"EC",X"05",
		X"CA",X"7F",X"A3",X"25",X"58",X"49",X"97",X"00",X"D6",X"3A",X"E0",X"06",X"E1",X"0B",X"25",X"02",
		X"E6",X"0B",X"D7",X"01",X"A6",X"06",X"A0",X"26",X"9F",X"5D",X"EE",X"88",X"14",X"E6",X"88",X"10",
		X"2A",X"09",X"E6",X"41",X"E0",X"0B",X"AE",X"44",X"3A",X"20",X"02",X"AE",X"44",X"10",X"9F",X"5F",
		X"EE",X"A8",X"14",X"E6",X"A8",X"10",X"2A",X"0B",X"E6",X"41",X"E0",X"2B",X"10",X"AE",X"44",X"31",
		X"A5",X"20",X"03",X"10",X"AE",X"44",X"31",X"A6",X"A6",X"A4",X"10",X"8C",X"9F",X"94",X"25",X"08",
		X"1E",X"12",X"8D",X"69",X"1E",X"12",X"96",X"02",X"90",X"00",X"8C",X"9F",X"94",X"25",X"06",X"8D",
		X"5C",X"91",X"02",X"20",X"02",X"A1",X"84",X"2E",X"04",X"DE",X"5F",X"20",X"06",X"DE",X"5D",X"1E",
		X"12",X"00",X"00",X"EC",X"D8",X"14",X"31",X"A5",X"D6",X"01",X"A6",X"A0",X"90",X"00",X"A1",X"80",
		X"2E",X"09",X"5A",X"26",X"F5",X"9E",X"5D",X"10",X"9E",X"5F",X"39",X"9E",X"5D",X"EE",X"88",X"12",
		X"A6",X"44",X"97",X"00",X"10",X"9E",X"5F",X"EE",X"A8",X"12",X"A6",X"44",X"91",X"00",X"24",X"09",
		X"1E",X"12",X"97",X"00",X"EE",X"A8",X"12",X"A6",X"44",X"E6",X"44",X"5C",X"3D",X"C3",X"50",X"47",
		X"1F",X"03",X"96",X"00",X"48",X"AD",X"D6",X"9E",X"5D",X"10",X"9E",X"5F",X"39",X"34",X"10",X"D6",
		X"01",X"3A",X"C6",X"FF",X"E1",X"82",X"23",X"02",X"E6",X"84",X"AC",X"E4",X"22",X"F6",X"D7",X"02",
		X"35",X"90",X"A6",X"88",X"10",X"85",X"03",X"27",X"09",X"A6",X"A8",X"10",X"85",X"03",X"10",X"26",
		X"00",X"92",X"EE",X"88",X"12",X"A6",X"49",X"97",X"02",X"EE",X"A8",X"12",X"A6",X"49",X"97",X"03",
		X"9B",X"02",X"24",X"03",X"46",X"20",X"05",X"81",X"20",X"25",X"07",X"44",X"04",X"02",X"04",X"03",
		X"20",X"F5",X"CE",X"4E",X"28",X"33",X"C6",X"A6",X"C4",X"D6",X"02",X"26",X"08",X"EC",X"2E",X"DD",
		X"04",X"EC",X"2C",X"20",X"34",X"3D",X"D7",X"08",X"A6",X"C4",X"D6",X"03",X"26",X"08",X"EC",X"0E",
		X"DD",X"04",X"EC",X"0C",X"20",X"23",X"3D",X"D7",X"09",X"CE",X"98",X"08",X"EC",X"0E",X"8D",X"55",
		X"DD",X"04",X"EC",X"0C",X"8D",X"4F",X"DD",X"06",X"CE",X"98",X"09",X"EC",X"2E",X"8D",X"46",X"D3",
		X"04",X"DD",X"04",X"EC",X"2C",X"8D",X"3E",X"D3",X"06",X"58",X"49",X"C9",X"00",X"89",X"00",X"DD",
		X"06",X"A3",X"0C",X"ED",X"0C",X"DC",X"06",X"A3",X"2C",X"ED",X"2C",X"DC",X"04",X"58",X"49",X"C9",
		X"00",X"89",X"00",X"DD",X"04",X"A3",X"0E",X"ED",X"0E",X"DC",X"04",X"A3",X"2E",X"ED",X"2E",X"BD",
		X"38",X"91",X"4D",X"A9",X"A6",X"88",X"10",X"8A",X"02",X"A7",X"88",X"10",X"A6",X"A8",X"10",X"8A",
		X"02",X"A7",X"A8",X"10",X"39",X"97",X"00",X"A6",X"C4",X"3D",X"97",X"01",X"A6",X"C4",X"D6",X"00",
		X"3D",X"2A",X"02",X"A0",X"C4",X"DB",X"01",X"89",X"00",X"39",X"34",X"56",X"7C",X"A0",X"0B",X"CE",
		X"A0",X"02",X"8E",X"9F",X"FD",X"8D",X"59",X"24",X"05",X"7F",X"A0",X"12",X"20",X"0C",X"8E",X"9F",
		X"FD",X"8D",X"6D",X"25",X"49",X"B6",X"A0",X"12",X"26",X"44",X"8E",X"A0",X"0C",X"FC",X"A0",X"10",
		X"8D",X"3E",X"A6",X"01",X"27",X"07",X"6F",X"01",X"CC",X"FF",X"FF",X"ED",X"02",X"FC",X"A0",X"0E",
		X"30",X"5F",X"8D",X"2C",X"A6",X"84",X"27",X"05",X"B7",X"A0",X"12",X"6F",X"84",X"8D",X"51",X"BD",
		X"38",X"91",X"4D",X"DF",X"B6",X"9F",X"FC",X"C6",X"02",X"BD",X"3C",X"0C",X"4C",X"27",X"BF",X"B7",
		X"9F",X"FC",X"C6",X"05",X"BD",X"4A",X"8E",X"C6",X"02",X"BD",X"3C",X"0C",X"20",X"B0",X"35",X"D6",
		X"34",X"16",X"A6",X"03",X"AB",X"61",X"19",X"A7",X"03",X"A6",X"02",X"A9",X"E4",X"19",X"A7",X"02",
		X"A6",X"01",X"89",X"00",X"19",X"A7",X"01",X"A6",X"84",X"89",X"00",X"19",X"A7",X"84",X"35",X"96",
		X"34",X"06",X"EC",X"84",X"10",X"A3",X"C4",X"26",X"05",X"EC",X"02",X"10",X"A3",X"42",X"35",X"86",
		X"34",X"56",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"CC",
		X"07",X"1B",X"FD",X"CA",X"06",X"86",X"81",X"F6",X"A0",X"0A",X"CB",X"22",X"1F",X"01",X"BF",X"CA",
		X"04",X"86",X"12",X"B7",X"CA",X"00",X"C6",X"99",X"CE",X"A0",X"02",X"A6",X"C0",X"27",X"FC",X"85",
		X"F0",X"26",X"06",X"8A",X"F0",X"20",X"02",X"A6",X"C0",X"BD",X"E2",X"0F",X"11",X"83",X"A0",X"06",
		X"25",X"F5",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"D6",X"34",X"06",X"4A",X"81",
		X"09",X"22",X"50",X"C6",X"06",X"3D",X"FB",X"A0",X"0A",X"86",X"7D",X"FD",X"CA",X"04",X"CC",X"2D",
		X"D9",X"20",X"1D",X"34",X"06",X"4A",X"C6",X"89",X"81",X"0A",X"2D",X"04",X"80",X"0A",X"CB",X"03",
		X"34",X"04",X"C6",X"06",X"3D",X"FB",X"A0",X"0A",X"35",X"02",X"FD",X"CA",X"04",X"CC",X"2D",X"E8",
		X"FD",X"CA",X"02",X"CC",X"07",X"01",X"FD",X"CA",X"06",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",
		X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"A6",X"62",X"B7",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",
		X"B7",X"C9",X"00",X"35",X"86",X"B6",X"A0",X"0B",X"27",X"05",X"8D",X"08",X"7F",X"A0",X"0B",X"EC",
		X"3E",X"DD",X"42",X"39",X"34",X"56",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",
		X"B7",X"C9",X"00",X"CC",X"85",X"03",X"FB",X"A0",X"0A",X"1F",X"01",X"CE",X"9F",X"FD",X"A6",X"C4",
		X"A1",X"49",X"27",X"0C",X"86",X"0F",X"8D",X"1F",X"86",X"F0",X"8D",X"1B",X"A6",X"C4",X"A7",X"49",
		X"30",X"0E",X"33",X"41",X"11",X"83",X"A0",X"01",X"25",X"E4",X"7F",X"CA",X"01",X"35",X"02",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"35",X"D6",X"97",X"00",X"A6",X"C4",X"9A",X"00",X"97",X"01",X"A6",
		X"49",X"9A",X"00",X"91",X"01",X"27",X"11",X"5F",X"BD",X"E2",X"06",X"30",X"12",X"A6",X"C4",X"9A",
		X"00",X"C6",X"DD",X"BD",X"E2",X"06",X"30",X"12",X"39",X"34",X"56",X"BE",X"A0",X"14",X"8C",X"4F",
		X"B2",X"26",X"0C",X"BE",X"A0",X"16",X"8C",X"4F",X"E2",X"26",X"5E",X"8D",X"5E",X"20",X"5A",X"30",
		X"1C",X"CC",X"FF",X"18",X"BD",X"3D",X"C1",X"BD",X"3D",X"7E",X"EE",X"9F",X"98",X"78",X"EE",X"4A",
		X"27",X"19",X"EC",X"02",X"44",X"AB",X"45",X"EB",X"47",X"FD",X"CA",X"04",X"EC",X"94",X"4C",X"88",
		X"04",X"C8",X"04",X"FD",X"CA",X"06",X"86",X"12",X"B7",X"CA",X"00",X"AE",X"9F",X"98",X"78",X"EC",
		X"08",X"6D",X"0A",X"27",X"04",X"9B",X"8D",X"DB",X"8E",X"BD",X"3F",X"B1",X"4D",X"6E",X"FE",X"A0",
		X"14",X"EE",X"0A",X"27",X"10",X"96",X"8D",X"5F",X"47",X"56",X"47",X"56",X"ED",X"4E",X"96",X"8E",
		X"5F",X"47",X"56",X"ED",X"4C",X"DC",X"8D",X"ED",X"06",X"35",X"D6",X"12",X"12",X"39",X"34",X"16",
		X"BE",X"A0",X"14",X"BC",X"A0",X"16",X"27",X"21",X"CC",X"FF",X"08",X"8D",X"64",X"30",X"04",X"BC",
		X"A0",X"16",X"26",X"15",X"8C",X"50",X"02",X"26",X"10",X"8E",X"4F",X"E2",X"BF",X"A0",X"14",X"BF",
		X"A0",X"16",X"CC",X"50",X"02",X"DD",X"7A",X"20",X"03",X"BD",X"3D",X"7E",X"35",X"96",X"34",X"56",
		X"BF",X"A0",X"14",X"EC",X"02",X"47",X"97",X"91",X"49",X"EE",X"84",X"E3",X"46",X"80",X"17",X"47",
		X"47",X"97",X"8D",X"D7",X"92",X"C0",X"16",X"57",X"57",X"D7",X"8E",X"FC",X"A0",X"16",X"10",X"83",
		X"4F",X"E2",X"26",X"03",X"8E",X"50",X"02",X"EC",X"1E",X"EE",X"1C",X"E3",X"46",X"47",X"97",X"8F",
		X"49",X"80",X"17",X"47",X"47",X"97",X"8B",X"D7",X"90",X"C0",X"16",X"57",X"57",X"D7",X"8C",X"35",
		X"D6",X"34",X"76",X"32",X"E8",X"E8",X"A6",X"03",X"A7",X"62",X"C6",X"1A",X"3D",X"10",X"8E",X"D7",
		X"7C",X"31",X"AB",X"E6",X"02",X"E7",X"63",X"54",X"A6",X"E8",X"19",X"24",X"02",X"8A",X"20",X"A7",
		X"E4",X"31",X"A5",X"EE",X"84",X"86",X"05",X"B7",X"CA",X"07",X"A6",X"41",X"A7",X"61",X"A7",X"66",
		X"E6",X"C4",X"C8",X"04",X"F7",X"CA",X"06",X"C8",X"04",X"86",X"19",X"A0",X"62",X"81",X"03",X"2E",
		X"02",X"4F",X"50",X"8C",X"50",X"02",X"24",X"01",X"4F",X"A7",X"67",X"AE",X"44",X"AF",X"64",X"AE",
		X"42",X"33",X"68",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",
		X"10",X"BF",X"CA",X"02",X"FF",X"CA",X"04",X"7F",X"CA",X"00",X"A6",X"61",X"BF",X"CA",X"02",X"B7",
		X"CA",X"00",X"86",X"04",X"FF",X"CA",X"02",X"10",X"BF",X"CA",X"04",X"B7",X"CA",X"00",X"31",X"A8",
		X"1A",X"6A",X"68",X"26",X"01",X"50",X"30",X"85",X"6A",X"62",X"26",X"D4",X"35",X"02",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"A6",X"E8",X"18",X"10",X"27",X"00",X"81",X"1D",X"8A",X"01",X"A7",X"61",
		X"8E",X"9F",X"94",X"E6",X"62",X"3A",X"A6",X"E4",X"85",X"10",X"26",X"29",X"EE",X"64",X"A6",X"66",
		X"31",X"C6",X"E6",X"C4",X"EB",X"63",X"E1",X"84",X"2C",X"02",X"E7",X"84",X"E6",X"A4",X"EB",X"63",
		X"E1",X"88",X"31",X"2F",X"03",X"E7",X"88",X"31",X"E6",X"61",X"33",X"C5",X"31",X"A5",X"30",X"01",
		X"4A",X"26",X"DF",X"20",X"47",X"86",X"1A",X"3D",X"C3",X"D7",X"7C",X"1F",X"03",X"A6",X"88",X"31",
		X"44",X"34",X"02",X"E6",X"84",X"54",X"A6",X"C5",X"26",X"0E",X"5C",X"E1",X"E4",X"23",X"F7",X"32",
		X"61",X"C6",X"4B",X"E7",X"84",X"50",X"20",X"18",X"58",X"85",X"F0",X"26",X"01",X"5C",X"E7",X"84",
		X"35",X"04",X"A6",X"C5",X"26",X"03",X"5A",X"20",X"F9",X"5C",X"58",X"85",X"0F",X"26",X"01",X"5A",
		X"E7",X"88",X"31",X"33",X"C8",X"1A",X"30",X"01",X"6A",X"66",X"26",X"C1",X"32",X"E8",X"18",X"35",
		X"F6",X"34",X"76",X"EE",X"88",X"12",X"A6",X"C8",X"1E",X"D6",X"75",X"3D",X"4D",X"10",X"27",X"00",
		X"81",X"34",X"06",X"1F",X"12",X"AE",X"A8",X"14",X"EC",X"06",X"E3",X"25",X"34",X"06",X"EE",X"A8",
		X"12",X"EE",X"C8",X"1F",X"BD",X"43",X"4F",X"CC",X"4D",X"9B",X"ED",X"88",X"12",X"1F",X"30",X"BD",
		X"43",X"32",X"CC",X"00",X"55",X"BD",X"47",X"FA",X"8B",X"55",X"AB",X"63",X"A7",X"63",X"BD",X"47",
		X"DA",X"34",X"06",X"CC",X"02",X"09",X"BD",X"47",X"FA",X"8B",X"03",X"10",X"8C",X"99",X"00",X"26",
		X"01",X"44",X"35",X"04",X"34",X"02",X"BD",X"47",X"BE",X"E3",X"2C",X"ED",X"0C",X"35",X"06",X"BD",
		X"47",X"BE",X"47",X"56",X"E3",X"2E",X"ED",X"0E",X"EC",X"E4",X"A3",X"46",X"A1",X"25",X"24",X"02",
		X"A6",X"25",X"E1",X"26",X"24",X"02",X"E6",X"26",X"ED",X"05",X"E7",X"07",X"AB",X"C4",X"A7",X"88",
		X"11",X"BD",X"43",X"5E",X"6A",X"62",X"27",X"08",X"33",X"48",X"A6",X"C4",X"26",X"96",X"20",X"8E",
		X"32",X"64",X"35",X"F6",X"DC",X"48",X"F0",X"99",X"05",X"82",X"00",X"47",X"56",X"E0",X"24",X"D7",
		X"61",X"EB",X"24",X"E7",X"24",X"DC",X"4B",X"F0",X"99",X"07",X"82",X"00",X"47",X"56",X"47",X"56",
		X"E0",X"25",X"D7",X"62",X"EB",X"25",X"E7",X"25",X"B6",X"99",X"05",X"C6",X"18",X"3D",X"43",X"97",
		X"67",X"B6",X"99",X"07",X"C6",X"0C",X"3D",X"40",X"8B",X"7F",X"97",X"68",X"EC",X"3E",X"DD",X"42",
		X"39",X"34",X"46",X"AE",X"64",X"EE",X"81",X"AF",X"64",X"6C",X"D8",X"12",X"E6",X"C8",X"14",X"4F",
		X"BD",X"46",X"FB",X"CC",X"41",X"07",X"6D",X"C8",X"17",X"26",X"03",X"CC",X"41",X"12",X"ED",X"02",
		X"EF",X"04",X"4F",X"5F",X"ED",X"0A",X"EC",X"9F",X"98",X"7D",X"ED",X"06",X"DC",X"7D",X"C3",X"00",
		X"02",X"10",X"83",X"50",X"35",X"25",X"03",X"CC",X"50",X"23",X"DD",X"7D",X"EC",X"E4",X"ED",X"08",
		X"10",X"83",X"80",X"80",X"10",X"26",X"00",X"82",X"86",X"00",X"BD",X"48",X"08",X"ED",X"08",X"0D",
		X"7F",X"10",X"27",X"00",X"C1",X"86",X"02",X"BD",X"48",X"08",X"C4",X"07",X"84",X"07",X"C0",X"04",
		X"80",X"04",X"DB",X"62",X"9B",X"61",X"34",X"06",X"2A",X"01",X"40",X"34",X"02",X"5D",X"2A",X"01",
		X"50",X"EB",X"E4",X"86",X"00",X"BD",X"48",X"02",X"3D",X"A1",X"E0",X"22",X"09",X"E6",X"E4",X"1D",
		X"8B",X"80",X"A7",X"08",X"20",X"07",X"E6",X"61",X"1D",X"8B",X"80",X"A7",X"09",X"32",X"62",X"EC",
		X"06",X"9B",X"61",X"26",X"12",X"34",X"02",X"96",X"31",X"2B",X"06",X"6C",X"06",X"6C",X"E4",X"20",
		X"04",X"6A",X"06",X"6A",X"E4",X"35",X"02",X"AB",X"08",X"28",X"02",X"63",X"08",X"DB",X"62",X"26",
		X"11",X"34",X"02",X"96",X"31",X"48",X"2B",X"05",X"6C",X"07",X"5C",X"20",X"03",X"6A",X"07",X"5A",
		X"35",X"02",X"EB",X"09",X"28",X"50",X"63",X"09",X"20",X"4C",X"0D",X"75",X"27",X"48",X"A3",X"C8",
		X"15",X"91",X"63",X"2C",X"41",X"D1",X"64",X"2C",X"3D",X"EC",X"08",X"E3",X"C8",X"15",X"91",X"65",
		X"2F",X"34",X"D1",X"66",X"2F",X"30",X"34",X"20",X"1F",X"12",X"1F",X"30",X"BD",X"43",X"22",X"A6",
		X"28",X"90",X"65",X"48",X"A7",X"05",X"A6",X"29",X"90",X"66",X"2A",X"01",X"4F",X"48",X"48",X"A7",
		X"07",X"A7",X"06",X"AB",X"98",X"14",X"24",X"07",X"A6",X"0B",X"40",X"A7",X"07",X"A7",X"06",X"BD",
		X"42",X"7B",X"1F",X"21",X"35",X"20",X"CE",X"A1",X"74",X"EC",X"C4",X"ED",X"84",X"EC",X"1E",X"ED",
		X"C4",X"35",X"C6",X"EE",X"24",X"EC",X"26",X"9B",X"61",X"AB",X"28",X"29",X"06",X"DB",X"62",X"EB",
		X"29",X"28",X"03",X"6E",X"D8",X"10",X"ED",X"28",X"A3",X"C8",X"15",X"91",X"63",X"2C",X"17",X"D1",
		X"64",X"2C",X"13",X"EC",X"28",X"E3",X"C8",X"15",X"91",X"65",X"2F",X"0A",X"D1",X"66",X"2F",X"06",
		X"96",X"75",X"10",X"26",X"00",X"BD",X"39",X"8D",X"10",X"8D",X"C8",X"8D",X"61",X"EC",X"3E",X"DD",
		X"42",X"39",X"8D",X"BF",X"EC",X"3E",X"DD",X"42",X"39",X"86",X"30",X"E6",X"28",X"3D",X"2A",X"02",
		X"80",X"30",X"47",X"34",X"01",X"8B",X"81",X"97",X"00",X"86",X"30",X"E6",X"29",X"3D",X"2A",X"02",
		X"80",X"30",X"8B",X"80",X"97",X"01",X"35",X"01",X"25",X"08",X"CC",X"00",X"00",X"ED",X"9F",X"98",
		X"00",X"39",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"CC",
		X"06",X"06",X"FD",X"CA",X"06",X"DC",X"00",X"FD",X"CA",X"04",X"CC",X"2D",X"F7",X"FD",X"CA",X"02",
		X"86",X"1A",X"B7",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"39",X"86",X"30",
		X"E6",X"28",X"3D",X"2A",X"02",X"80",X"30",X"47",X"34",X"01",X"8B",X"81",X"97",X"00",X"86",X"30",
		X"E6",X"29",X"3D",X"2A",X"02",X"80",X"30",X"8B",X"80",X"97",X"01",X"35",X"01",X"25",X"08",X"EC",
		X"C8",X"17",X"ED",X"9F",X"98",X"00",X"39",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"CC",X"06",X"06",X"FD",X"CA",X"06",X"DC",X"00",X"FD",X"CA",X"04",X"30",
		X"C8",X"19",X"BF",X"CA",X"02",X"86",X"0A",X"B7",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"39",X"DC",X"63",X"E3",X"C8",X"15",X"A0",X"28",X"97",X"00",X"8E",X"50",X"37",X"E0",
		X"29",X"D1",X"00",X"2C",X"05",X"D7",X"00",X"8E",X"50",X"3B",X"EC",X"28",X"E3",X"C8",X"15",X"90",
		X"65",X"91",X"00",X"2C",X"05",X"97",X"00",X"8E",X"50",X"39",X"D0",X"66",X"D1",X"00",X"2C",X"03",
		X"8E",X"50",X"3D",X"11",X"83",X"4D",X"2D",X"26",X"02",X"30",X"08",X"EC",X"84",X"DD",X"01",X"1F",
		X"30",X"BD",X"43",X"22",X"6E",X"9F",X"98",X"01",X"CC",X"FF",X"73",X"ED",X"04",X"20",X"06",X"A6",
		X"98",X"14",X"40",X"A7",X"05",X"6F",X"88",X"10",X"A6",X"29",X"A0",X"C8",X"16",X"90",X"66",X"2B",
		X"14",X"48",X"48",X"A7",X"07",X"A7",X"06",X"AB",X"0B",X"24",X"50",X"86",X"FF",X"A7",X"07",X"A7",
		X"06",X"86",X"40",X"20",X"09",X"6F",X"06",X"A6",X"0B",X"40",X"A7",X"07",X"86",X"80",X"A7",X"88",
		X"10",X"A6",X"28",X"A0",X"C8",X"15",X"90",X"65",X"48",X"A7",X"05",X"20",X"2E",X"CC",X"FF",X"73",
		X"ED",X"04",X"20",X"02",X"6F",X"05",X"A6",X"29",X"90",X"66",X"2B",X"14",X"48",X"48",X"A7",X"07",
		X"A7",X"06",X"AB",X"98",X"14",X"24",X"14",X"A6",X"0B",X"40",X"A7",X"07",X"A7",X"06",X"20",X"04",
		X"6F",X"06",X"6F",X"07",X"A6",X"28",X"90",X"65",X"48",X"A7",X"05",X"A6",X"05",X"AB",X"98",X"14",
		X"A7",X"88",X"11",X"EC",X"3E",X"ED",X"88",X"1C",X"A6",X"26",X"5F",X"47",X"56",X"47",X"56",X"ED",
		X"0E",X"A6",X"27",X"5F",X"47",X"56",X"ED",X"0C",X"AF",X"2A",X"BD",X"43",X"5E",X"6E",X"D8",X"0E",
		X"CC",X"45",X"47",X"ED",X"88",X"1A",X"CC",X"42",X"AC",X"ED",X"22",X"39",X"8D",X"1E",X"EC",X"3E",
		X"DD",X"42",X"39",X"CC",X"45",X"47",X"ED",X"88",X"1A",X"CC",X"42",X"BF",X"ED",X"22",X"39",X"BD",
		X"41",X"19",X"8D",X"08",X"BD",X"41",X"6E",X"EC",X"3E",X"DD",X"42",X"39",X"EE",X"24",X"AE",X"2A",
		X"F6",X"99",X"07",X"54",X"54",X"D7",X"00",X"E6",X"07",X"54",X"54",X"A6",X"88",X"10",X"2A",X"02",
		X"CB",X"C0",X"D0",X"00",X"B6",X"99",X"05",X"44",X"97",X"00",X"A6",X"05",X"8B",X"50",X"44",X"80",
		X"28",X"90",X"00",X"AB",X"C8",X"15",X"ED",X"28",X"39",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",
		X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",X"49",X"4E",
		X"43",X"2E",X"34",X"06",X"8D",X"29",X"EC",X"E4",X"ED",X"88",X"12",X"C3",X"00",X"0A",X"ED",X"E4",
		X"EC",X"F1",X"34",X"46",X"EE",X"E4",X"EF",X"88",X"14",X"EC",X"42",X"ED",X"09",X"A6",X"41",X"A7",
		X"0B",X"CC",X"44",X"22",X"ED",X"88",X"18",X"CC",X"45",X"EA",X"ED",X"88",X"1A",X"35",X"C6",X"0A",
		X"75",X"9E",X"3D",X"26",X"01",X"3F",X"EC",X"84",X"DD",X"3D",X"6F",X"88",X"10",X"39",X"34",X"62",
		X"A6",X"06",X"CE",X"98",X"33",X"31",X"C4",X"EE",X"C4",X"27",X"04",X"A1",X"46",X"22",X"F6",X"EE",
		X"A4",X"EF",X"84",X"AF",X"A4",X"10",X"AF",X"02",X"AF",X"42",X"A6",X"05",X"EE",X"88",X"14",X"AB",
		X"C4",X"A7",X"88",X"11",X"35",X"E2",X"CC",X"43",X"93",X"ED",X"88",X"18",X"CC",X"4B",X"B5",X"ED",
		X"88",X"12",X"39",X"AE",X"A8",X"14",X"A6",X"84",X"E6",X"2B",X"88",X"04",X"C8",X"04",X"FD",X"CA",
		X"06",X"EC",X"25",X"FD",X"CA",X"04",X"EC",X"29",X"FD",X"CA",X"02",X"E6",X"24",X"1D",X"84",X"20",
		X"8A",X"1A",X"B7",X"CA",X"00",X"7E",X"46",X"65",X"AE",X"A8",X"14",X"A6",X"84",X"E6",X"2B",X"88",
		X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"25",X"FD",X"CA",X"04",X"EC",X"29",X"FD",X"CA",X"02",
		X"E6",X"24",X"1D",X"84",X"20",X"8A",X"1A",X"B7",X"CA",X"00",X"EC",X"06",X"AE",X"A8",X"16",X"AF",
		X"A8",X"14",X"A0",X"06",X"E0",X"07",X"D7",X"01",X"EB",X"2C",X"E7",X"2C",X"5F",X"47",X"56",X"DD",
		X"02",X"E3",X"2E",X"ED",X"2E",X"EC",X"02",X"ED",X"29",X"FD",X"CA",X"02",X"EC",X"84",X"E7",X"2B",
		X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"A8",X"1A",X"DD",X"04",X"CC",X"45",X"2D",X"ED",
		X"A8",X"1A",X"A6",X"A8",X"10",X"2A",X"2D",X"A6",X"27",X"AB",X"01",X"25",X"27",X"7E",X"45",X"27",
		X"20",X"22",X"AE",X"A8",X"14",X"A6",X"84",X"E6",X"2B",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",
		X"EC",X"25",X"FD",X"CA",X"04",X"EC",X"29",X"FD",X"CA",X"02",X"E6",X"24",X"1D",X"84",X"20",X"8A",
		X"1A",X"B7",X"CA",X"00",X"AE",X"A8",X"14",X"EC",X"2C",X"D3",X"46",X"2A",X"31",X"E3",X"27",X"ED",
		X"27",X"25",X"17",X"E6",X"A8",X"10",X"CA",X"80",X"E7",X"A8",X"10",X"5F",X"E7",X"26",X"F7",X"CA",
		X"05",X"97",X"00",X"AB",X"01",X"25",X"6E",X"7E",X"45",X"27",X"E6",X"A8",X"10",X"2B",X"F2",X"A7",
		X"26",X"B7",X"CA",X"05",X"C5",X"40",X"27",X"71",X"AB",X"01",X"25",X"1F",X"20",X"43",X"E3",X"27",
		X"ED",X"27",X"25",X"25",X"E6",X"A8",X"10",X"2B",X"48",X"A7",X"26",X"B7",X"CA",X"05",X"C5",X"40",
		X"26",X"09",X"AB",X"01",X"24",X"53",X"CA",X"40",X"E7",X"A8",X"10",X"A6",X"27",X"43",X"2F",X"0E",
		X"A7",X"2B",X"88",X"04",X"B7",X"CA",X"07",X"20",X"40",X"E6",X"A8",X"10",X"2B",X"07",X"86",X"FF",
		X"A7",X"27",X"7E",X"45",X"27",X"A7",X"26",X"B7",X"CA",X"05",X"EC",X"02",X"ED",X"29",X"FD",X"CA",
		X"02",X"C4",X"3F",X"E7",X"A8",X"10",X"A6",X"01",X"A7",X"2B",X"88",X"04",X"B7",X"CA",X"07",X"20",
		X"18",X"97",X"00",X"AB",X"01",X"A7",X"2B",X"88",X"04",X"B7",X"CA",X"07",X"96",X"00",X"40",X"E6",
		X"84",X"3D",X"E3",X"02",X"ED",X"29",X"FD",X"CA",X"02",X"E6",X"24",X"A6",X"25",X"2B",X"0C",X"E3",
		X"2E",X"D3",X"44",X"2B",X"0C",X"81",X"74",X"25",X"13",X"20",X"2C",X"E3",X"2E",X"D3",X"44",X"2A",
		X"0B",X"A7",X"25",X"B7",X"CA",X"04",X"AB",X"84",X"25",X"0D",X"20",X"1B",X"A7",X"25",X"B7",X"CA",
		X"04",X"AB",X"84",X"2A",X"02",X"86",X"7F",X"A7",X"A8",X"11",X"E7",X"24",X"1D",X"84",X"20",X"8A",
		X"0A",X"B7",X"CA",X"00",X"6E",X"B8",X"1A",X"AE",X"A8",X"12",X"6E",X"98",X"0C",X"A6",X"2C",X"90",
		X"01",X"A7",X"2C",X"EC",X"2E",X"93",X"02",X"ED",X"2E",X"CC",X"44",X"22",X"ED",X"A8",X"18",X"DC",
		X"04",X"ED",X"A8",X"1A",X"6E",X"B8",X"1A",X"A6",X"A8",X"10",X"85",X"C0",X"26",X"15",X"A6",X"24",
		X"48",X"EC",X"25",X"49",X"E3",X"06",X"81",X"E8",X"24",X"09",X"44",X"06",X"00",X"1F",X"01",X"6E",
		X"9F",X"98",X"76",X"7E",X"45",X"EA",X"96",X"7C",X"A7",X"A8",X"1E",X"A6",X"A8",X"21",X"A7",X"A8",
		X"1F",X"A7",X"A8",X"20",X"20",X"30",X"96",X"7C",X"A7",X"A8",X"1F",X"A6",X"A8",X"20",X"A7",X"A8",
		X"1E",X"A7",X"A8",X"21",X"20",X"20",X"96",X"7C",X"A7",X"A8",X"20",X"A6",X"A8",X"1F",X"A7",X"A8",
		X"1E",X"A7",X"A8",X"21",X"20",X"10",X"96",X"7C",X"A7",X"A8",X"21",X"A6",X"A8",X"1E",X"A7",X"A8",
		X"1F",X"A7",X"A8",X"20",X"20",X"00",X"A6",X"A8",X"1E",X"48",X"48",X"48",X"48",X"AA",X"A8",X"1F",
		X"E6",X"A8",X"20",X"58",X"58",X"58",X"58",X"EA",X"A8",X"21",X"0D",X"00",X"2B",X"04",X"ED",X"84",
		X"20",X"1A",X"B7",X"DC",X"76",X"F7",X"DC",X"78",X"CC",X"06",X"06",X"FD",X"CA",X"06",X"CC",X"DC",
		X"76",X"FD",X"CA",X"02",X"BF",X"CA",X"04",X"86",X"2A",X"B7",X"CA",X"00",X"8E",X"4F",X"AA",X"86",
		X"00",X"BD",X"48",X"08",X"C4",X"07",X"A6",X"85",X"97",X"7C",X"A6",X"A8",X"10",X"85",X"03",X"10",
		X"27",X"EE",X"8C",X"6A",X"A8",X"10",X"7E",X"34",X"7F",X"A6",X"A8",X"10",X"85",X"C0",X"26",X"28",
		X"EE",X"A8",X"1E",X"EC",X"C4",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"42",X"FD",X"CA",
		X"02",X"A6",X"24",X"48",X"EC",X"25",X"49",X"E3",X"06",X"A3",X"46",X"44",X"FD",X"CA",X"04",X"86",
		X"0A",X"24",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"7E",X"45",X"EA",X"AE",X"A8",X"12",X"CC",X"41",
		X"07",X"6D",X"88",X"17",X"26",X"03",X"CC",X"41",X"12",X"AE",X"B8",X"1C",X"ED",X"02",X"EC",X"2E",
		X"C3",X"00",X"20",X"58",X"49",X"58",X"49",X"A7",X"06",X"EC",X"2C",X"C3",X"00",X"20",X"58",X"49",
		X"A7",X"07",X"34",X"20",X"1F",X"12",X"BD",X"41",X"19",X"BD",X"42",X"CC",X"BD",X"41",X"6E",X"4F",
		X"5F",X"ED",X"2A",X"35",X"20",X"AE",X"A4",X"DC",X"3D",X"ED",X"A4",X"10",X"9F",X"3D",X"10",X"AE",
		X"22",X"AF",X"A4",X"10",X"AF",X"02",X"0C",X"75",X"7E",X"34",X"AA",X"46",X"7B",X"46",X"7F",X"9E",
		X"40",X"33",X"02",X"EF",X"04",X"6A",X"06",X"4F",X"A1",X"06",X"24",X"04",X"33",X"84",X"A6",X"06",
		X"30",X"07",X"8C",X"A1",X"A5",X"26",X"F1",X"DF",X"40",X"EC",X"44",X"DD",X"42",X"39",X"46",X"9E",
		X"46",X"A2",X"CC",X"A1",X"A0",X"DD",X"42",X"39",X"35",X"06",X"ED",X"22",X"EC",X"A4",X"DE",X"42",
		X"ED",X"D4",X"EC",X"84",X"ED",X"A4",X"EC",X"3E",X"ED",X"84",X"39",X"34",X"66",X"CC",X"00",X"04",
		X"8D",X"39",X"10",X"AE",X"66",X"EC",X"A4",X"31",X"24",X"10",X"AF",X"66",X"ED",X"02",X"10",X"AE",
		X"3E",X"EC",X"A4",X"ED",X"84",X"EC",X"1E",X"ED",X"A4",X"35",X"E6",X"34",X"66",X"10",X"AE",X"66",
		X"EE",X"A4",X"31",X"25",X"10",X"AF",X"66",X"E6",X"3D",X"4F",X"8D",X"0F",X"EF",X"02",X"10",X"AE",
		X"3E",X"EC",X"A4",X"ED",X"84",X"EC",X"1E",X"ED",X"A4",X"35",X"E6",X"34",X"40",X"DE",X"3B",X"26",
		X"01",X"3F",X"AE",X"C4",X"9F",X"3B",X"C3",X"00",X"04",X"9E",X"6B",X"30",X"8B",X"8C",X"BE",X"C0",
		X"22",X"0A",X"9E",X"6B",X"ED",X"84",X"D3",X"6B",X"DD",X"6B",X"20",X"11",X"9E",X"6D",X"30",X"8B",
		X"9C",X"6F",X"25",X"01",X"3F",X"9E",X"6D",X"ED",X"84",X"D3",X"6D",X"DD",X"6D",X"DC",X"73",X"A3",
		X"81",X"DD",X"73",X"24",X"12",X"DC",X"88",X"27",X"01",X"3F",X"FC",X"BE",X"FE",X"DD",X"88",X"CC",
		X"37",X"F9",X"FD",X"BE",X"FE",X"DC",X"73",X"EF",X"81",X"AF",X"C4",X"35",X"C0",X"BD",X"41",X"19",
		X"EE",X"24",X"6A",X"D8",X"12",X"EC",X"A4",X"AE",X"9F",X"98",X"42",X"20",X"02",X"AE",X"94",X"10",
		X"AC",X"94",X"26",X"F9",X"ED",X"84",X"30",X"A4",X"34",X"46",X"9C",X"6D",X"24",X"06",X"9C",X"71",
		X"24",X"02",X"9F",X"71",X"EE",X"1E",X"DC",X"3B",X"ED",X"C4",X"DF",X"3B",X"4F",X"5F",X"ED",X"1E",
		X"35",X"C6",X"34",X"14",X"ED",X"E3",X"2A",X"01",X"40",X"5D",X"2A",X"01",X"50",X"85",X"F0",X"27",
		X"06",X"44",X"54",X"85",X"F0",X"26",X"F6",X"C5",X"F0",X"27",X"06",X"44",X"54",X"C5",X"F0",X"26",
		X"F6",X"A7",X"E2",X"58",X"58",X"58",X"58",X"EB",X"E0",X"30",X"8D",X"06",X"EB",X"3A",X"A6",X"84",
		X"E6",X"E0",X"2A",X"03",X"40",X"8B",X"80",X"E6",X"E0",X"2A",X"01",X"40",X"35",X"94",X"34",X"06",
		X"4D",X"2A",X"01",X"40",X"5D",X"2A",X"01",X"50",X"3D",X"6D",X"E0",X"2A",X"04",X"43",X"50",X"82",
		X"FF",X"6D",X"E0",X"2A",X"04",X"43",X"50",X"82",X"FF",X"39",X"34",X"52",X"84",X"C0",X"44",X"44",
		X"44",X"44",X"CE",X"4E",X"89",X"33",X"C6",X"8E",X"4E",X"49",X"35",X"02",X"A8",X"C4",X"E6",X"86",
		X"E8",X"41",X"88",X"3F",X"A6",X"86",X"A8",X"42",X"35",X"D0",X"34",X"04",X"8D",X"0A",X"35",X"04",
		X"3D",X"39",X"34",X"04",X"8D",X"02",X"35",X"84",X"34",X"10",X"8E",X"98",X"2E",X"30",X"86",X"A6",
		X"84",X"48",X"A8",X"84",X"48",X"48",X"EC",X"84",X"59",X"49",X"ED",X"84",X"26",X"01",X"3F",X"35",
		X"90",X"34",X"56",X"5F",X"20",X"02",X"34",X"56",X"AE",X"66",X"EE",X"94",X"30",X"1F",X"A3",X"C4",
		X"2C",X"04",X"8D",X"68",X"20",X"02",X"8D",X"20",X"30",X"03",X"AF",X"66",X"35",X"D6",X"34",X"56",
		X"5F",X"20",X"02",X"34",X"56",X"AE",X"66",X"30",X"1F",X"4D",X"2A",X"04",X"8D",X"4E",X"20",X"02",
		X"8D",X"06",X"30",X"03",X"AF",X"66",X"35",X"D6",X"34",X"10",X"AE",X"01",X"EE",X"84",X"EB",X"41",
		X"E7",X"41",X"89",X"00",X"27",X"34",X"34",X"02",X"AB",X"C4",X"A1",X"C4",X"2C",X"0B",X"CC",X"7F",
		X"FF",X"A0",X"C4",X"32",X"61",X"35",X"10",X"20",X"DF",X"A7",X"C4",X"30",X"02",X"A6",X"E4",X"E6",
		X"84",X"27",X"15",X"3D",X"2A",X"0A",X"A0",X"E4",X"58",X"49",X"8D",X"10",X"30",X"03",X"20",X"ED",
		X"58",X"49",X"8D",X"C4",X"30",X"03",X"20",X"E5",X"32",X"61",X"35",X"90",X"34",X"10",X"AE",X"01",
		X"EE",X"84",X"EB",X"41",X"E7",X"41",X"89",X"00",X"27",X"38",X"34",X"02",X"AB",X"C4",X"A1",X"C4",
		X"2F",X"0B",X"CC",X"80",X"00",X"A0",X"C4",X"32",X"61",X"35",X"10",X"20",X"DF",X"A7",X"C4",X"30",
		X"02",X"A6",X"E4",X"E6",X"84",X"27",X"19",X"3D",X"2A",X"0C",X"A0",X"E4",X"A0",X"84",X"58",X"49",
		X"8D",X"86",X"30",X"03",X"20",X"EB",X"A0",X"84",X"58",X"49",X"8D",X"C0",X"30",X"03",X"20",X"E1",
		X"32",X"61",X"35",X"90",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",
		X"47",X"56",X"39",X"34",X"04",X"B6",X"C8",X"06",X"84",X"03",X"48",X"48",X"48",X"48",X"F6",X"C8",
		X"04",X"C5",X"20",X"26",X"08",X"8A",X"08",X"C5",X"80",X"26",X"02",X"88",X"0C",X"C5",X"02",X"26",
		X"08",X"8A",X"01",X"C5",X"08",X"26",X"02",X"88",X"03",X"35",X"84",X"34",X"02",X"A6",X"80",X"1E",
		X"12",X"BD",X"4A",X"78",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",X"34",X"36",X"8E",X"49",X"3A",
		X"10",X"8E",X"CC",X"00",X"C6",X"12",X"8D",X"E3",X"35",X"B6",X"30",X"30",X"03",X"05",X"01",X"01",
		X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"49",X"B8",X"BD",
		X"32",X"45",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1D",X"84",X"0F",X"27",X"11",
		X"7F",X"CC",X"1D",X"BD",X"49",X"B8",X"BD",X"32",X"45",X"BD",X"4A",X"4F",X"86",X"28",X"BD",X"F0",
		X"09",X"B6",X"CC",X"1F",X"84",X"0F",X"27",X"0C",X"7F",X"CC",X"1F",X"8D",X"3B",X"8D",X"45",X"86",
		X"40",X"BD",X"F0",X"09",X"B6",X"CC",X"23",X"84",X"0F",X"27",X"07",X"7F",X"CC",X"23",X"8D",X"28",
		X"8D",X"35",X"B6",X"CC",X"21",X"84",X"0F",X"27",X"0A",X"7F",X"CC",X"21",X"8D",X"1A",X"8D",X"07",
		X"7E",X"F0",X"06",X"8D",X"02",X"20",X"52",X"B6",X"CC",X"1B",X"84",X"0F",X"27",X"09",X"7C",X"CC",
		X"28",X"7C",X"CC",X"28",X"7F",X"CC",X"1B",X"39",X"34",X"12",X"8D",X"0E",X"8E",X"CC",X"28",X"BD",
		X"4A",X"78",X"35",X"92",X"7E",X"8B",X"64",X"7E",X"89",X"8E",X"34",X"34",X"8E",X"CC",X"00",X"10",
		X"8E",X"CC",X"24",X"8D",X"02",X"35",X"B4",X"10",X"BF",X"BF",X"06",X"4F",X"E6",X"80",X"C4",X"0F",
		X"34",X"04",X"AB",X"E0",X"BC",X"BF",X"06",X"26",X"F3",X"8B",X"37",X"39",X"8D",X"DC",X"34",X"02",
		X"8E",X"CC",X"28",X"BD",X"4A",X"5F",X"A1",X"E0",X"39",X"8D",X"F1",X"27",X"36",X"86",X"39",X"B7",
		X"CB",X"FF",X"BD",X"49",X"2B",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"AC",X"86",X"39",X"B7",X"CB",
		X"FF",X"BD",X"32",X"45",X"86",X"39",X"B7",X"CB",X"FF",X"8D",X"1E",X"8D",X"CF",X"27",X"16",X"86",
		X"0A",X"BD",X"E2",X"12",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F4",
		X"7E",X"2E",X"45",X"20",X"FB",X"86",X"0B",X"20",X"E8",X"8E",X"CD",X"02",X"C6",X"04",X"A6",X"80",
		X"84",X"0F",X"81",X"09",X"23",X"03",X"5A",X"27",X"06",X"8C",X"CD",X"32",X"26",X"F0",X"39",X"86",
		X"0C",X"BD",X"E2",X"12",X"8E",X"CD",X"02",X"6F",X"80",X"8C",X"CD",X"32",X"26",X"F9",X"39",X"A6",
		X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",X"8D",X"EF",
		X"34",X"02",X"8D",X"EB",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",
		X"A7",X"81",X"35",X"82",X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",X"34",X"16",
		X"86",X"01",X"20",X"02",X"34",X"16",X"0D",X"96",X"26",X"35",X"C4",X"0F",X"58",X"34",X"04",X"58",
		X"EB",X"E0",X"8E",X"CC",X"FC",X"3A",X"8D",X"C8",X"34",X"04",X"8D",X"C4",X"34",X"04",X"8D",X"C0",
		X"34",X"04",X"AB",X"E4",X"19",X"A7",X"E4",X"A6",X"61",X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",
		X"89",X"00",X"19",X"30",X"1A",X"8D",X"B1",X"35",X"04",X"35",X"02",X"8D",X"B7",X"35",X"02",X"35",
		X"96",X"34",X"12",X"BB",X"BF",X"1B",X"19",X"24",X"02",X"86",X"99",X"B7",X"BF",X"1B",X"8E",X"CD",
		X"00",X"BD",X"4A",X"78",X"8E",X"10",X"6D",X"86",X"02",X"C6",X"26",X"6F",X"8B",X"5A",X"2A",X"FB",
		X"4A",X"2A",X"F6",X"35",X"92",X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",
		X"04",X"34",X"16",X"C6",X"01",X"96",X"96",X"34",X"02",X"0F",X"96",X"BD",X"38",X"91",X"4D",X"FC",
		X"BD",X"4A",X"8E",X"58",X"8E",X"CC",X"0C",X"3A",X"BD",X"4A",X"70",X"8D",X"6C",X"B6",X"BF",X"1D",
		X"34",X"04",X"AB",X"E4",X"B7",X"BF",X"1D",X"B6",X"BF",X"1C",X"AB",X"E0",X"B7",X"BF",X"1C",X"8E",
		X"CC",X"18",X"BD",X"4A",X"70",X"8D",X"52",X"34",X"04",X"A1",X"E0",X"25",X"30",X"8E",X"CC",X"14",
		X"BD",X"4A",X"70",X"8D",X"44",X"8D",X"2C",X"34",X"02",X"F7",X"BF",X"1C",X"8E",X"CC",X"16",X"BD",
		X"4A",X"70",X"B6",X"BF",X"1D",X"8D",X"32",X"8D",X"1A",X"4D",X"27",X"06",X"7F",X"BF",X"1C",X"7F",
		X"BF",X"1D",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"4A",X"94",X"BD",X"4A",X"D1",X"35",X"02",X"97",
		X"96",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",
		X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",X"4F",X"C1",X"10",X"25",X"06",
		X"8B",X"0A",X"C0",X"10",X"20",X"F6",X"34",X"04",X"AB",X"E0",X"1F",X"89",X"35",X"82",X"34",X"04",
		X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",
		X"AB",X"E0",X"19",X"35",X"84",X"80",X"00",X"00",X"00",X"00",X"E1",X"96",X"E1",X"96",X"00",X"00",
		X"00",X"46",X"65",X"2F",X"A0",X"40",X"00",X"00",X"75",X"5F",X"72",X"19",X"05",X"00",X"07",X"FF",
		X"B0",X"42",X"B9",X"E1",X"96",X"A0",X"39",X"19",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"40",X"29",X"1B",X"00",X"7F",X"E0",X"20",X"00",X"01",X"74",X"A1",X"71",X"C7",X"60",X"0B",
		X"23",X"6F",X"A2",X"42",X"B9",X"5D",X"26",X"A0",X"21",X"16",X"03",X"03",X"AA",X"AA",X"0A",X"A0",
		X"0A",X"A0",X"00",X"42",X"26",X"CD",X"0D",X"7F",X"E0",X"20",X"00",X"01",X"74",X"AA",X"71",X"CE",
		X"50",X"0C",X"CB",X"6F",X"A2",X"42",X"B9",X"5D",X"26",X"A0",X"24",X"16",X"03",X"03",X"AA",X"AA",
		X"0A",X"A0",X"0A",X"A0",X"00",X"37",X"26",X"CD",X"0D",X"7F",X"E0",X"20",X"00",X"01",X"74",X"B3",
		X"71",X"D5",X"20",X"0E",X"3B",X"6F",X"A2",X"42",X"B9",X"5D",X"26",X"A0",X"27",X"16",X"02",X"02",
		X"AA",X"AA",X"0A",X"A0",X"0A",X"A0",X"00",X"16",X"26",X"CD",X"0D",X"7F",X"E0",X"20",X"00",X"01",
		X"74",X"BC",X"71",X"DC",X"50",X"0F",X"1B",X"6F",X"A2",X"42",X"B9",X"5D",X"26",X"A0",X"2A",X"16",
		X"03",X"03",X"AA",X"AA",X"0A",X"A0",X"0A",X"A0",X"00",X"37",X"26",X"CD",X"0D",X"7F",X"E0",X"20",
		X"00",X"01",X"74",X"C5",X"71",X"E3",X"90",X"10",X"9D",X"6F",X"A2",X"42",X"B9",X"5D",X"26",X"A0",
		X"2D",X"22",X"04",X"03",X"AA",X"AA",X"0A",X"A0",X"0A",X"A0",X"00",X"63",X"26",X"CD",X"19",X"27",
		X"A0",X"10",X"00",X"02",X"75",X"0C",X"72",X"06",X"01",X"DC",X"7D",X"46",X"2B",X"42",X"B9",X"5D",
		X"2F",X"98",X"95",X"19",X"00",X"00",X"99",X"99",X"09",X"90",X"09",X"90",X"06",X"00",X"2D",X"6F",
		X"00",X"7F",X"F0",X"04",X"00",X"04",X"74",X"83",X"6C",X"73",X"01",X"12",X"9D",X"46",X"2B",X"42",
		X"B9",X"5D",X"26",X"A0",X"1B",X"27",X"01",X"01",X"CC",X"CC",X"0C",X"C0",X"0C",X"C0",X"0A",X"00",
		X"7F",X"D0",X"01",X"00",X"06",X"74",X"8C",X"71",X"91",X"02",X"19",X"E1",X"6A",X"2E",X"69",X"F8",
		X"5D",X"26",X"A0",X"1E",X"27",X"02",X"02",X"BB",X"BB",X"0B",X"B0",X"0B",X"B0",X"0C",X"00",X"7D",
		X"80",X"00",X"80",X"07",X"75",X"34",X"59",X"B0",X"FF",X"50",X"1A",X"6F",X"A2",X"42",X"B9",X"5D",
		X"BE",X"A0",X"36",X"22",X"06",X"06",X"FF",X"FF",X"0F",X"F0",X"0F",X"F0",X"04",X"00",X"2D",X"6F",
		X"19",X"27",X"20",X"00",X"40",X"08",X"E1",X"96",X"E1",X"96",X"00",X"24",X"38",X"46",X"65",X"76",
		X"50",X"00",X"20",X"09",X"E1",X"96",X"E1",X"96",X"00",X"24",X"38",X"46",X"65",X"6F",X"80",X"08",
		X"00",X"03",X"74",X"E9",X"6C",X"70",X"01",X"26",X"A1",X"46",X"2B",X"42",X"A0",X"5D",X"26",X"A0",
		X"33",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"2D",X"6F",X"00",X"7F",
		X"70",X"02",X"00",X"05",X"74",X"95",X"71",X"95",X"02",X"12",X"9D",X"46",X"2B",X"42",X"B3",X"5D",
		X"6A",X"A0",X"1B",X"27",X"01",X"01",X"CC",X"CC",X"0C",X"C0",X"0C",X"C0",X"0A",X"00",X"07",X"20",
		X"00",X"10",X"0A",X"E1",X"96",X"72",X"1D",X"00",X"23",X"DC",X"E1",X"96",X"7A",X"76",X"5D",X"26",
		X"00",X"00",X"0D",X"01",X"01",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"E1",X"96",X"E1",X"96",X"00",X"00",X"00",X"7A",X"66",X"07",X"20",X"00",X"10",X"0A",
		X"E1",X"96",X"E1",X"96",X"00",X"24",X"38",X"46",X"65",X"10",X"AB",X"42",X"03",X"00",X"13",X"AE",
		X"52",X"10",X"00",X"28",X"B3",X"60",X"10",X"58",X"20",X"00",X"21",X"AD",X"50",X"10",X"48",X"10",
		X"00",X"38",X"B8",X"79",X"0C",X"B7",X"79",X"80",X"00",X"21",X"AA",X"5A",X"20",X"00",X"21",X"A6",
		X"60",X"09",X"00",X"24",X"AF",X"60",X"10",X"52",X"FF",X"00",X"21",X"A3",X"58",X"20",X"00",X"38",
		X"BC",X"70",X"20",X"58",X"20",X"00",X"21",X"BE",X"60",X"30",X"00",X"38",X"A4",X"70",X"30",X"58",
		X"88",X"00",X"38",X"A6",X"70",X"FF",X"00",X"12",X"A7",X"50",X"40",X"00",X"3F",X"B0",X"7E",X"60",
		X"00",X"06",X"04",X"00",X"02",X"04",X"00",X"02",X"00",X"00",X"00",X"0D",X"00",X"32",X"00",X"72",
		X"00",X"0D",X"40",X"19",X"20",X"3F",X"13",X"7F",X"0D",X"32",X"40",X"3F",X"2D",X"66",X"20",X"7F",
		X"18",X"72",X"40",X"7F",X"33",X"7F",X"28",X"7F",X"20",X"FF",X"80",X"55",X"40",X"33",X"2B",X"25",
		X"20",X"1C",X"1A",X"17",X"15",X"14",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"0D",X"0C",X"0C",X"0B",
		X"0B",X"0A",X"0A",X"0A",X"09",X"09",X"09",X"08",X"08",X"00",X"03",X"06",X"09",X"0C",X"0F",X"12",
		X"15",X"18",X"1B",X"1E",X"21",X"24",X"27",X"2A",X"2D",X"30",X"33",X"36",X"39",X"3B",X"3E",X"41",
		X"43",X"46",X"49",X"4B",X"4E",X"50",X"52",X"55",X"57",X"59",X"5B",X"5E",X"60",X"62",X"64",X"66",
		X"67",X"69",X"6B",X"6C",X"6E",X"70",X"71",X"72",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"3F",X"00",X"00",X"00",X"40",X"FF",X"00",
		X"00",X"BF",X"FF",X"FF",X"00",X"C0",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"12",X"0E",X"0A",X"08",X"06",X"04",
		X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"40",X"2E",X"20",X"1A",X"12",X"0E",X"0E",X"0A",
		X"0A",X"08",X"08",X"06",X"06",X"06",X"04",X"04",X"40",X"32",X"26",X"20",X"1C",X"18",X"12",X"10",
		X"0E",X"0E",X"0A",X"0A",X"0A",X"08",X"08",X"08",X"40",X"36",X"2E",X"24",X"20",X"1C",X"1A",X"16",
		X"12",X"10",X"0E",X"0E",X"0E",X"0E",X"0A",X"0A",X"40",X"38",X"32",X"28",X"24",X"20",X"1E",X"1A",
		X"18",X"16",X"12",X"10",X"10",X"0E",X"0E",X"0E",X"40",X"3A",X"32",X"2E",X"26",X"22",X"20",X"1E",
		X"1C",X"1A",X"18",X"16",X"12",X"10",X"10",X"0E",X"40",X"3C",X"36",X"30",X"2A",X"26",X"22",X"20",
		X"1E",X"1C",X"1A",X"18",X"18",X"16",X"12",X"12",X"40",X"3C",X"36",X"32",X"2E",X"28",X"24",X"22",
		X"20",X"20",X"1C",X"1A",X"1A",X"18",X"16",X"16",X"40",X"3C",X"38",X"32",X"30",X"2A",X"26",X"24",
		X"20",X"20",X"20",X"1E",X"1C",X"1A",X"18",X"18",X"40",X"3E",X"38",X"36",X"32",X"2E",X"28",X"26",
		X"24",X"20",X"20",X"20",X"1E",X"1C",X"1A",X"1A",X"40",X"3E",X"3A",X"36",X"32",X"30",X"2A",X"28",
		X"26",X"22",X"20",X"20",X"20",X"1E",X"1C",X"1C",X"40",X"3E",X"3A",X"36",X"32",X"30",X"2E",X"28",
		X"26",X"24",X"22",X"20",X"20",X"20",X"1E",X"1C",X"40",X"3E",X"3A",X"38",X"32",X"32",X"30",X"2A",
		X"28",X"26",X"24",X"22",X"20",X"20",X"20",X"1E",X"40",X"3E",X"3C",X"38",X"36",X"32",X"30",X"2E",
		X"2A",X"28",X"26",X"24",X"22",X"20",X"20",X"20",X"40",X"3E",X"3C",X"38",X"36",X"32",X"32",X"2E",
		X"2A",X"28",X"26",X"24",X"24",X"22",X"20",X"20",X"45",X"66",X"45",X"76",X"45",X"86",X"45",X"96",
		X"CC",X"66",X"99",X"55",X"DD",X"CC",X"66",X"99",X"55",X"DD",X"01",X"02",X"03",X"04",X"05",X"09",
		X"0D",X"0F",X"1E",X"13",X"27",X"0B",X"1E",X"1B",X"27",X"17",X"1E",X"AA",X"25",X"04",X"1F",X"12",
		X"17",X"00",X"1E",X"B2",X"25",X"22",X"1F",X"1A",X"17",X"24",X"1F",X"AC",X"0E",X"24",X"1F",X"A4",
		X"0E",X"00",X"20",X"29",X"02",X"04",X"20",X"AE",X"00",X"11",X"20",X"B6",X"00",X"17",X"20",X"31",
		X"02",X"20",X"1D",X"5B",X"06",X"1C",X"1B",X"AC",X"10",X"09",X"1C",X"24",X"06",X"15",X"1D",X"53",
		X"06",X"0D",X"1C",X"6B",X"18",X"09",X"1B",X"B4",X"10",X"1B",X"1C",X"73",X"18",X"16",X"1D",X"B3",
		X"10",X"13",X"22",X"98",X"06",X"0C",X"21",X"06",X"1A",X"0C",X"23",X"04",X"06",X"0C",X"21",X"8C",
		X"1A",X"0C",X"23",X"70",X"06",X"0C",X"22",X"12",X"1A",X"0C",X"1A",X"31",X"D7",X"7C",X"9F",X"94",
		X"19",X"18",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"01",X"01",X"FF",X"01",X"01",X"FF",
		X"01",X"FF",X"FF",X"01",X"00",X"A1",X"38",X"42",X"08",X"42",X"0F",X"42",X"2B",X"42",X"35",X"42",
		X"4D",X"42",X"54",X"42",X"67",X"42",X"70",X"E1",X"96",X"57",X"1C",X"57",X"33",X"E1",X"96",X"57",
		X"56",X"E1",X"96",X"56",X"6C",X"57",X"2A",X"E1",X"96",X"55",X"EB",X"55",X"E4",X"57",X"2A",X"57",
		X"6F",X"56",X"FE",X"55",X"EB",X"55",X"E4",X"57",X"2A",X"57",X"6F",X"55",X"EB",X"55",X"EB",X"55",
		X"EB",X"55",X"E4",X"57",X"2A",X"57",X"8E",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",X"EB",X"55",
		X"EE",X"57",X"4B",X"57",X"C7",X"57",X"28",X"57",X"28",X"E1",X"96",X"57",X"28",X"57",X"33",X"E1",
		X"96",X"57",X"50",X"E1",X"96",X"E1",X"96",X"56",X"D5",X"56",X"D5",X"57",X"FC",X"E1",X"96",X"E1",
		X"96",X"56",X"EE",X"57",X"50",X"57",X"E9",X"E1",X"96",X"56",X"D5",X"56",X"D5",X"E1",X"96",X"E1",
		X"96",X"58",X"1E",X"E1",X"96",X"E1",X"96",X"E1",X"96",X"E1",X"96",X"E1",X"96",X"58",X"18",X"58",
		X"18",X"58",X"18",X"E1",X"96",X"E1",X"96",X"58",X"15",X"E1",X"96",X"00",X"FF",X"BF",X"AE",X"AD",
		X"A4",X"9A",X"00",X"00",X"C9",X"50",X"4B",X"05",X"07",X"00",X"37",X"00",X"DD",X"BB",X"66",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"BD",X"51",X"0F",X"BD",X"54",X"33",X"39",X"12",
		X"12",X"12",X"7D",X"A1",X"B8",X"26",X"01",X"39",X"8E",X"DC",X"7A",X"6C",X"80",X"2F",X"05",X"6F",
		X"1F",X"6A",X"1F",X"39",X"10",X"AE",X"84",X"31",X"28",X"10",X"8C",X"0A",X"EC",X"2D",X"04",X"10",
		X"8E",X"0A",X"D4",X"10",X"AF",X"81",X"30",X"08",X"10",X"AE",X"22",X"C6",X"0F",X"A6",X"A0",X"A7",
		X"80",X"5A",X"2E",X"F9",X"39",X"12",X"12",X"12",X"BD",X"59",X"56",X"FD",X"A1",X"A9",X"39",X"BD",
		X"7C",X"58",X"0D",X"96",X"27",X"14",X"7E",X"8E",X"31",X"BD",X"46",X"DB",X"51",X"6D",X"08",X"A1",
		X"5F",X"4F",X"5F",X"ED",X"04",X"ED",X"06",X"39",X"2E",X"DA",X"0C",X"96",X"39",X"8E",X"99",X"00",
		X"EC",X"0E",X"E3",X"24",X"47",X"56",X"ED",X"0E",X"ED",X"24",X"EC",X"0C",X"E3",X"26",X"47",X"56",
		X"ED",X"0C",X"ED",X"26",X"EC",X"3E",X"DD",X"42",X"39",X"BD",X"51",X"ED",X"7F",X"A1",X"B9",X"86",
		X"FF",X"B7",X"A1",X"BC",X"7F",X"A1",X"BA",X"7F",X"A1",X"BB",X"0F",X"86",X"BD",X"46",X"BB",X"51",
		X"A4",X"A1",X"97",X"39",X"96",X"2E",X"B7",X"A1",X"B6",X"B7",X"A1",X"B7",X"CC",X"51",X"B6",X"ED",
		X"22",X"EC",X"3E",X"DD",X"42",X"39",X"CC",X"51",X"C0",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",
		X"CC",X"51",X"CA",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"96",X"2E",X"B7",X"A1",X"B6",X"CC",
		X"51",X"D9",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"CC",X"51",X"E3",X"ED",X"22",X"EC",X"3E",
		X"DD",X"42",X"39",X"CC",X"51",X"A4",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"BD",X"74",X"15",
		X"8E",X"DC",X"7D",X"10",X"8E",X"0A",X"D4",X"EE",X"A4",X"EF",X"81",X"CE",X"DC",X"85",X"EF",X"81",
		X"EE",X"24",X"EF",X"81",X"EE",X"26",X"EF",X"81",X"8E",X"DC",X"7B",X"BD",X"51",X"33",X"BD",X"55",
		X"A0",X"0F",X"94",X"7F",X"A1",X"B2",X"7F",X"A1",X"B8",X"0F",X"93",X"0A",X"93",X"BD",X"46",X"BB",
		X"55",X"D4",X"A1",X"89",X"7F",X"A1",X"AC",X"7F",X"A1",X"AB",X"8E",X"55",X"50",X"BF",X"A1",X"A9",
		X"7D",X"A1",X"B3",X"2A",X"11",X"BD",X"46",X"BB",X"52",X"3E",X"A1",X"5F",X"20",X"08",X"BD",X"3C",
		X"D9",X"EC",X"3E",X"DD",X"42",X"39",X"0D",X"96",X"27",X"37",X"B6",X"9F",X"FC",X"27",X"0A",X"C6",
		X"12",X"BD",X"3C",X"0C",X"7A",X"9F",X"FC",X"20",X"F1",X"BD",X"56",X"7E",X"4C",X"81",X"05",X"2D",
		X"F8",X"BD",X"46",X"DB",X"52",X"82",X"08",X"A1",X"5F",X"BD",X"46",X"BB",X"52",X"8F",X"A1",X"5F",
		X"BD",X"46",X"DB",X"6C",X"59",X"08",X"A1",X"66",X"CC",X"03",X"DE",X"ED",X"04",X"4F",X"BD",X"8E",
		X"37",X"39",X"86",X"3B",X"97",X"80",X"CC",X"0E",X"10",X"BD",X"34",X"19",X"7E",X"58",X"32",X"96",
		X"8A",X"0F",X"8A",X"BD",X"33",X"8E",X"97",X"8A",X"EC",X"3E",X"DD",X"42",X"39",X"BD",X"74",X"0B",
		X"BD",X"52",X"F5",X"39",X"BD",X"80",X"57",X"4F",X"97",X"96",X"4F",X"5F",X"FD",X"A1",X"A9",X"34",
		X"50",X"8E",X"00",X"00",X"CC",X"00",X"EF",X"B7",X"A1",X"B3",X"30",X"02",X"8B",X"10",X"2B",X"1C",
		X"EE",X"8B",X"11",X"A3",X"89",X"52",X"E1",X"1A",X"0A",X"1C",X"DE",X"26",X"02",X"1A",X"0B",X"7D",
		X"A1",X"B3",X"25",X"E6",X"2E",X"E4",X"5C",X"F7",X"A1",X"B3",X"24",X"DE",X"35",X"50",X"39",X"52",
		X"69",X"63",X"68",X"6A",X"00",X"00",X"00",X"0C",X"4A",X"15",X"91",X"45",X"43",X"01",X"50",X"35",
		X"02",X"57",X"69",X"74",X"74",X"7D",X"A0",X"13",X"26",X"12",X"34",X"37",X"86",X"8A",X"F6",X"A0",
		X"0A",X"1F",X"01",X"C6",X"FF",X"86",X"55",X"BD",X"E2",X"03",X"35",X"37",X"39",X"34",X"36",X"86",
		X"8A",X"F6",X"A0",X"0A",X"1F",X"01",X"C6",X"00",X"86",X"55",X"BD",X"E2",X"03",X"35",X"36",X"7D",
		X"A1",X"B3",X"10",X"2C",X"DB",X"1E",X"34",X"36",X"34",X"16",X"AE",X"9F",X"98",X"78",X"A6",X"0A",
		X"27",X"32",X"BE",X"A0",X"16",X"8C",X"4F",X"E2",X"26",X"2A",X"9E",X"7A",X"31",X"89",X"AF",X"FE",
		X"1F",X"20",X"47",X"56",X"47",X"56",X"47",X"56",X"1F",X"02",X"A6",X"A9",X"53",X"69",X"97",X"2C",
		X"CC",X"00",X"08",X"30",X"04",X"BD",X"3D",X"C1",X"30",X"04",X"8C",X"50",X"1A",X"25",X"03",X"8E",
		X"50",X"02",X"9F",X"7A",X"35",X"16",X"35",X"36",X"39",X"07",X"03",X"00",X"34",X"12",X"BE",X"A0",
		X"16",X"8C",X"4F",X"E2",X"26",X"2B",X"A6",X"F8",X"03",X"81",X"0B",X"27",X"15",X"7D",X"A1",X"AB",
		X"27",X"08",X"81",X"08",X"27",X"04",X"81",X"09",X"26",X"17",X"81",X"02",X"27",X"04",X"0D",X"94",
		X"26",X"0F",X"8E",X"53",X"AA",X"48",X"AD",X"96",X"7C",X"A1",X"AB",X"BF",X"A1",X"A9",X"7F",X"A1",
		X"AC",X"AE",X"63",X"30",X"01",X"AF",X"63",X"35",X"12",X"39",X"2E",X"44",X"53",X"C2",X"53",X"CB",
		X"53",X"D4",X"53",X"DD",X"53",X"E6",X"53",X"EF",X"53",X"F8",X"54",X"01",X"54",X"0D",X"54",X"19",
		X"54",X"22",X"BD",X"38",X"91",X"55",X"56",X"8E",X"54",X"88",X"39",X"BD",X"38",X"91",X"55",X"5B",
		X"8E",X"54",X"A2",X"39",X"BD",X"38",X"91",X"55",X"60",X"8E",X"54",X"C0",X"39",X"BD",X"38",X"91",
		X"55",X"65",X"8E",X"54",X"CE",X"39",X"BD",X"38",X"91",X"55",X"6A",X"8E",X"54",X"EC",X"39",X"BD",
		X"38",X"91",X"55",X"6F",X"8E",X"55",X"04",X"39",X"BD",X"38",X"91",X"55",X"74",X"8E",X"55",X"20",
		X"39",X"BD",X"38",X"91",X"55",X"79",X"7F",X"A1",X"AB",X"8E",X"55",X"3A",X"39",X"BD",X"38",X"91",
		X"55",X"7E",X"7F",X"A1",X"AB",X"8E",X"55",X"46",X"39",X"BD",X"38",X"91",X"54",X"2E",X"8E",X"55",
		X"50",X"39",X"BD",X"38",X"91",X"55",X"5B",X"7F",X"A1",X"AB",X"8E",X"54",X"A2",X"39",X"3F",X"A0",
		X"41",X"01",X"00",X"34",X"76",X"7A",X"A1",X"AC",X"2C",X"3F",X"BE",X"A1",X"A9",X"27",X"2E",X"EC",
		X"84",X"81",X"FF",X"27",X"28",X"30",X"02",X"BF",X"A1",X"A9",X"5A",X"2D",X"ED",X"F7",X"A1",X"AC",
		X"AE",X"9F",X"98",X"78",X"AE",X"0A",X"27",X"21",X"BE",X"A0",X"16",X"8C",X"4F",X"E2",X"26",X"19",
		X"8E",X"54",X"7C",X"30",X"86",X"CC",X"00",X"08",X"BD",X"3D",X"C1",X"20",X"0C",X"8E",X"55",X"54",
		X"7F",X"A1",X"AB",X"BF",X"A1",X"A9",X"7F",X"A1",X"AC",X"35",X"76",X"39",X"22",X"98",X"06",X"0C",
		X"23",X"70",X"06",X"0C",X"23",X"04",X"06",X"0C",X"00",X"01",X"08",X"0E",X"04",X"08",X"08",X"06",
		X"00",X"14",X"04",X"0C",X"00",X"01",X"04",X"0A",X"00",X"03",X"08",X"19",X"04",X"03",X"00",X"01",
		X"FF",X"06",X"00",X"01",X"08",X"02",X"04",X"10",X"00",X"05",X"04",X"03",X"08",X"07",X"04",X"0E",
		X"00",X"0D",X"08",X"0C",X"04",X"08",X"08",X"07",X"00",X"03",X"04",X"0F",X"00",X"01",X"FF",X"06",
		X"00",X"01",X"08",X"05",X"04",X"0B",X"08",X"0C",X"04",X"18",X"00",X"01",X"FF",X"06",X"00",X"01",
		X"08",X"02",X"04",X"10",X"00",X"07",X"04",X"03",X"08",X"05",X"04",X"0E",X"00",X"0D",X"04",X"08",
		X"00",X"06",X"04",X"03",X"08",X"05",X"04",X"0D",X"00",X"0D",X"FF",X"06",X"00",X"01",X"04",X"04",
		X"08",X"0E",X"04",X"06",X"00",X"0D",X"04",X"08",X"00",X"06",X"04",X"03",X"08",X"05",X"04",X"0D",
		X"00",X"0D",X"FF",X"06",X"00",X"01",X"04",X"04",X"08",X"0E",X"04",X"06",X"00",X"0D",X"04",X"04",
		X"08",X"0E",X"04",X"06",X"00",X"0D",X"04",X"04",X"08",X"0E",X"04",X"06",X"00",X"0D",X"FF",X"06",
		X"00",X"01",X"08",X"05",X"04",X"0B",X"08",X"0C",X"04",X"18",X"00",X"0D",X"04",X"08",X"00",X"06",
		X"04",X"03",X"08",X"05",X"04",X"0D",X"00",X"0D",X"FF",X"06",X"00",X"01",X"04",X"14",X"08",X"7E",
		X"04",X"02",X"00",X"01",X"FF",X"06",X"00",X"01",X"04",X"14",X"08",X"7E",X"04",X"02",X"FF",X"06",
		X"00",X"01",X"FF",X"00",X"FF",X"00",X"3C",X"B2",X"7B",X"80",X"00",X"3C",X"B1",X"7B",X"80",X"00",
		X"3A",X"B0",X"7B",X"60",X"00",X"3A",X"AC",X"7B",X"80",X"00",X"3A",X"B4",X"7B",X"80",X"00",X"3A",
		X"A2",X"7B",X"80",X"00",X"3A",X"B9",X"7B",X"80",X"00",X"3A",X"BD",X"7B",X"A0",X"00",X"3C",X"BD",
		X"7B",X"A0",X"00",X"34",X"12",X"86",X"04",X"97",X"93",X"A6",X"62",X"BB",X"A0",X"0A",X"A7",X"62",
		X"35",X"12",X"39",X"91",X"57",X"23",X"09",X"0F",X"57",X"BD",X"38",X"91",X"4D",X"E6",X"97",X"57",
		X"34",X"16",X"86",X"FF",X"97",X"93",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",
		X"B7",X"C9",X"00",X"CC",X"03",X"45",X"FD",X"CA",X"06",X"F6",X"A0",X"0A",X"86",X"76",X"FD",X"CA",
		X"02",X"FD",X"CA",X"04",X"86",X"12",X"B7",X"CA",X"00",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",
		X"00",X"35",X"16",X"39",X"0D",X"93",X"2D",X"07",X"0A",X"93",X"2C",X"03",X"BD",X"55",X"A0",X"EC",
		X"3E",X"DD",X"42",X"39",X"7D",X"A1",X"B2",X"10",X"26",X"D8",X"59",X"7E",X"3A",X"62",X"7D",X"A1",
		X"B2",X"10",X"26",X"D8",X"4F",X"FC",X"A0",X"16",X"10",X"83",X"4F",X"E2",X"10",X"26",X"01",X"28",
		X"7D",X"A1",X"BB",X"10",X"27",X"00",X"01",X"39",X"4F",X"5F",X"ED",X"2E",X"ED",X"2C",X"FD",X"99",
		X"0E",X"FD",X"99",X"0C",X"86",X"08",X"97",X"80",X"0F",X"86",X"CC",X"4B",X"B5",X"FD",X"99",X"12",
		X"7F",X"A1",X"AB",X"BD",X"53",X"6C",X"09",X"BD",X"46",X"DB",X"56",X"34",X"05",X"A1",X"5F",X"86",
		X"92",X"A7",X"04",X"39",X"B6",X"A1",X"BB",X"26",X"2C",X"96",X"2E",X"97",X"50",X"7F",X"A1",X"B9",
		X"AE",X"9F",X"98",X"78",X"A6",X"0C",X"84",X"F0",X"A7",X"0C",X"6A",X"24",X"27",X"05",X"EC",X"3E",
		X"DD",X"42",X"39",X"7F",X"A1",X"AB",X"BD",X"53",X"6C",X"0A",X"CC",X"4B",X"C3",X"FD",X"99",X"12",
		X"BD",X"58",X"32",X"20",X"04",X"86",X"0F",X"97",X"80",X"7E",X"47",X"55",X"BD",X"56",X"7E",X"AE",
		X"B8",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"CC",X"02",X"00",X"BD",X"3B",X"2A",X"39",X"34",X"36",
		X"B6",X"A0",X"13",X"26",X"03",X"BD",X"53",X"0D",X"4C",X"81",X"14",X"2F",X"33",X"BD",X"38",X"91",
		X"56",X"D0",X"86",X"10",X"BD",X"55",X"93",X"8E",X"7A",X"00",X"BD",X"55",X"83",X"C6",X"AA",X"86",
		X"56",X"BD",X"E2",X"0C",X"86",X"57",X"BD",X"E2",X"0C",X"8E",X"76",X"00",X"BD",X"55",X"83",X"86",
		X"58",X"BD",X"E2",X"0C",X"86",X"59",X"BD",X"E2",X"0C",X"86",X"5A",X"BD",X"E2",X"0C",X"20",X"0D",
		X"BD",X"38",X"91",X"4D",X"DA",X"B7",X"A0",X"13",X"C6",X"02",X"BD",X"3C",X"23",X"35",X"36",X"39",
		X"21",X"A8",X"5A",X"0C",X"00",X"BD",X"38",X"91",X"4D",X"B3",X"AE",X"98",X"1C",X"EE",X"04",X"AD",
		X"D8",X"07",X"30",X"A4",X"BD",X"43",X"86",X"CC",X"01",X"50",X"BD",X"3B",X"2A",X"39",X"7D",X"A1",
		X"B2",X"10",X"26",X"D7",X"4F",X"30",X"A4",X"BD",X"43",X"86",X"BD",X"58",X"32",X"39",X"EE",X"B8",
		X"1C",X"EC",X"88",X"1C",X"10",X"A3",X"C8",X"11",X"27",X"01",X"39",X"BD",X"38",X"91",X"4D",X"C9",
		X"AE",X"98",X"1C",X"BD",X"6C",X"70",X"AE",X"B8",X"1C",X"7E",X"6C",X"64",X"7D",X"A1",X"B2",X"10",
		X"26",X"D7",X"21",X"86",X"01",X"B7",X"A1",X"B4",X"1E",X"12",X"BD",X"6C",X"79",X"BD",X"3A",X"62",
		X"7E",X"6C",X"76",X"34",X"10",X"30",X"A4",X"BD",X"6C",X"79",X"35",X"10",X"BD",X"6C",X"79",X"BD",
		X"3A",X"62",X"BD",X"6C",X"76",X"30",X"A4",X"BD",X"6C",X"76",X"39",X"BD",X"6C",X"56",X"20",X"E3",
		X"BD",X"6C",X"56",X"7E",X"58",X"18",X"BD",X"38",X"91",X"4D",X"B3",X"AE",X"98",X"1C",X"EE",X"04",
		X"AD",X"D8",X"07",X"AE",X"B8",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"BD",X"57",X"A9",X"39",X"BD",
		X"38",X"91",X"4D",X"B3",X"AE",X"98",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"AE",X"B8",X"1C",X"EE",
		X"04",X"AD",X"D8",X"07",X"CC",X"01",X"50",X"BD",X"3B",X"2A",X"BD",X"57",X"A9",X"39",X"BD",X"38",
		X"91",X"4D",X"B3",X"AE",X"98",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"AE",X"B8",X"1C",X"EE",X"04",
		X"AD",X"D8",X"07",X"CC",X"05",X"00",X"BD",X"3B",X"2A",X"86",X"20",X"BD",X"55",X"93",X"8E",X"7A",
		X"00",X"BD",X"55",X"83",X"C6",X"FF",X"86",X"5B",X"BD",X"E2",X"0C",X"8E",X"76",X"00",X"BD",X"55",
		X"83",X"86",X"5C",X"BD",X"E2",X"0C",X"39",X"BD",X"38",X"91",X"4D",X"B3",X"34",X"10",X"30",X"A4",
		X"BD",X"6C",X"56",X"35",X"10",X"AE",X"98",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"BD",X"58",X"B9",
		X"B6",X"A1",X"B9",X"8B",X"02",X"B7",X"A1",X"B9",X"39",X"BD",X"38",X"91",X"4D",X"B3",X"AE",X"98",
		X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"30",X"A4",X"BD",X"43",X"86",X"39",X"BD",X"38",X"91",X"4D",
		X"B3",X"AE",X"98",X"1C",X"EE",X"04",X"AD",X"D8",X"07",X"30",X"A4",X"BD",X"43",X"86",X"CC",X"05",
		X"00",X"BD",X"3B",X"2A",X"39",X"BD",X"43",X"86",X"30",X"A4",X"BD",X"43",X"86",X"39",X"BD",X"38",
		X"91",X"4D",X"B3",X"BD",X"43",X"86",X"30",X"A4",X"BD",X"43",X"86",X"CC",X"01",X"00",X"BD",X"3B",
		X"2A",X"39",X"96",X"96",X"27",X"07",X"0F",X"96",X"0F",X"8A",X"7E",X"8C",X"F0",X"BD",X"38",X"91",
		X"4D",X"C1",X"86",X"FF",X"97",X"1E",X"4F",X"5F",X"FD",X"99",X"0E",X"FD",X"99",X"0C",X"DD",X"44",
		X"DD",X"46",X"0F",X"80",X"B6",X"9F",X"FC",X"C6",X"12",X"BD",X"3C",X"0C",X"7A",X"9F",X"FC",X"C6",
		X"07",X"BD",X"4A",X"8E",X"7C",X"A1",X"BA",X"8E",X"99",X"00",X"BD",X"6C",X"61",X"CC",X"4B",X"B5",
		X"FD",X"99",X"12",X"BD",X"46",X"DB",X"58",X"7C",X"08",X"A1",X"5F",X"39",X"96",X"95",X"BA",X"A1",
		X"AB",X"27",X"05",X"EC",X"3E",X"DD",X"42",X"39",X"CC",X"00",X"3C",X"BD",X"34",X"19",X"AE",X"9F",
		X"98",X"78",X"AE",X"0A",X"26",X"0A",X"BD",X"53",X"6C",X"01",X"CC",X"00",X"3C",X"BD",X"34",X"19",
		X"BD",X"55",X"A0",X"CC",X"58",X"AD",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"7D",X"A1",X"AB",
		X"10",X"27",X"D6",X"AF",X"EC",X"3E",X"DD",X"42",X"39",X"34",X"36",X"FC",X"A0",X"14",X"10",X"83",
		X"4F",X"B2",X"26",X"24",X"FC",X"A0",X"16",X"10",X"83",X"4F",X"E2",X"10",X"26",X"00",X"84",X"7D",
		X"A1",X"BB",X"26",X"7F",X"7C",X"A1",X"BB",X"BD",X"6C",X"6D",X"CC",X"70",X"00",X"BD",X"3B",X"2A",
		X"CC",X"80",X"00",X"BD",X"3B",X"2A",X"20",X"6B",X"BD",X"3C",X"D9",X"BD",X"53",X"6C",X"08",X"10",
		X"AE",X"9F",X"98",X"78",X"4F",X"AE",X"2A",X"27",X"0C",X"EC",X"0E",X"47",X"56",X"ED",X"0E",X"EC",
		X"0C",X"47",X"56",X"ED",X"0C",X"A6",X"26",X"47",X"A7",X"26",X"E6",X"27",X"57",X"E7",X"27",X"A6",
		X"A8",X"18",X"E6",X"A8",X"19",X"47",X"57",X"8A",X"01",X"CA",X"01",X"3D",X"47",X"47",X"47",X"47",
		X"47",X"26",X"01",X"4C",X"97",X"1E",X"86",X"10",X"BD",X"55",X"93",X"8E",X"7A",X"00",X"BD",X"55",
		X"83",X"C6",X"AA",X"86",X"5B",X"BD",X"E2",X"0C",X"86",X"5D",X"BD",X"E2",X"0C",X"8E",X"76",X"00",
		X"BD",X"55",X"83",X"86",X"5E",X"BD",X"E2",X"0C",X"86",X"5F",X"BD",X"E2",X"0C",X"CC",X"05",X"00",
		X"BD",X"3B",X"2A",X"35",X"36",X"39",X"C3",X"D6",X"D7",X"E8",X"D9",X"C9",X"C7",X"C8",X"E3",X"40",
		X"4D",X"C3",X"5D",X"40",X"F1",X"F9",X"F8",X"F2",X"40",X"E6",X"C9",X"D3",X"D3",X"C9",X"C1",X"D4",
		X"E2",X"40",X"C5",X"D3",X"C5",X"C3",X"E3",X"D9",X"D6",X"D5",X"C9",X"C3",X"E2",X"6B",X"40",X"C9",
		X"D5",X"C3",X"4B",X"00",X"39",X"A0",X"19",X"06",X"59",X"A4",X"14",X"59",X"A7",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"A0",X"1C",X"00",X"A0",X"1F",X"00",X"A0",X"2E",X"00",X"A0",X"3C",X"00",
		X"34",X"36",X"7C",X"A1",X"B2",X"CC",X"50",X"02",X"FD",X"A0",X"16",X"7C",X"A0",X"3E",X"28",X"03",
		X"7A",X"A0",X"3E",X"7E",X"8E",X"65",X"26",X"0C",X"86",X"07",X"97",X"1E",X"BD",X"46",X"DB",X"59",
		X"D7",X"0C",X"A1",X"5F",X"35",X"36",X"39",X"BD",X"46",X"BB",X"5C",X"8B",X"A1",X"9E",X"AE",X"1E",
		X"AF",X"28",X"BD",X"46",X"BB",X"5C",X"8B",X"A1",X"6D",X"AE",X"1E",X"AF",X"2A",X"86",X"FF",X"B7",
		X"A1",X"BC",X"BD",X"46",X"BB",X"5B",X"06",X"A1",X"5F",X"CC",X"5A",X"03",X"ED",X"22",X"EC",X"3E",
		X"DD",X"42",X"39",X"AE",X"9F",X"98",X"78",X"AE",X"0A",X"26",X"05",X"EC",X"3E",X"DD",X"42",X"39",
		X"CC",X"00",X"5A",X"BD",X"34",X"19",X"7F",X"A1",X"BC",X"BD",X"32",X"0F",X"AE",X"B8",X"08",X"CC",
		X"5C",X"ED",X"ED",X"02",X"AE",X"B8",X"0A",X"CC",X"5C",X"ED",X"ED",X"02",X"CC",X"00",X"B4",X"BD",
		X"34",X"19",X"7C",X"A1",X"BC",X"BD",X"32",X"0F",X"AE",X"B8",X"08",X"CC",X"5C",X"B8",X"ED",X"02",
		X"AE",X"B8",X"0A",X"CC",X"5C",X"B8",X"ED",X"02",X"34",X"36",X"B6",X"A1",X"AD",X"BD",X"47",X"DA",
		X"34",X"02",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"FD",X"A1",X"AE",X"35",X"04",
		X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"FD",X"A1",X"B0",X"BD",X"46",
		X"BB",X"5B",X"68",X"A1",X"5F",X"35",X"36",X"CC",X"00",X"78",X"BD",X"34",X"19",X"BD",X"32",X"0F",
		X"AE",X"B8",X"08",X"CC",X"5C",X"ED",X"ED",X"02",X"AE",X"B8",X"0A",X"CC",X"5C",X"ED",X"ED",X"02",
		X"CC",X"00",X"B4",X"BD",X"34",X"19",X"34",X"36",X"BD",X"46",X"BB",X"5B",X"AE",X"A1",X"6D",X"BD",
		X"6C",X"7C",X"AE",X"B8",X"08",X"CC",X"5C",X"06",X"ED",X"02",X"AE",X"B8",X"0A",X"CC",X"5C",X"06",
		X"ED",X"02",X"35",X"36",X"CC",X"00",X"78",X"BD",X"34",X"19",X"34",X"36",X"BD",X"32",X"0F",X"AE",
		X"B8",X"08",X"CC",X"47",X"55",X"ED",X"02",X"AE",X"B8",X"0A",X"CC",X"47",X"55",X"ED",X"02",X"86",
		X"FF",X"B7",X"A1",X"BC",X"4F",X"5F",X"10",X"AE",X"9F",X"98",X"78",X"AE",X"2A",X"27",X"04",X"ED",
		X"0E",X"ED",X"0C",X"A7",X"26",X"A7",X"27",X"B6",X"A1",X"AD",X"BD",X"47",X"DA",X"34",X"02",X"1D",
		X"58",X"49",X"DD",X"81",X"35",X"04",X"1D",X"58",X"49",X"DD",X"83",X"7F",X"A1",X"B2",X"7F",X"A1",
		X"BB",X"35",X"36",X"7E",X"8E",X"88",X"7D",X"A1",X"BC",X"2F",X"03",X"7E",X"47",X"55",X"34",X"36",
		X"0C",X"96",X"10",X"AE",X"9F",X"50",X"35",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"38",X"BD",X"64",
		X"DD",X"8B",X"80",X"97",X"50",X"86",X"01",X"F6",X"A1",X"B7",X"34",X"16",X"BD",X"63",X"38",X"8E",
		X"5C",X"F6",X"BD",X"65",X"03",X"BD",X"65",X"40",X"FC",X"99",X"0E",X"43",X"50",X"82",X"FF",X"DD",
		X"44",X"35",X"16",X"BD",X"63",X"49",X"8E",X"5C",X"F6",X"BD",X"65",X"03",X"BD",X"65",X"69",X"FC",
		X"99",X"0C",X"43",X"50",X"82",X"FF",X"DD",X"46",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"79",X"0A",
		X"96",X"35",X"36",X"EC",X"3E",X"DD",X"42",X"39",X"34",X"36",X"FC",X"A1",X"B0",X"4D",X"2C",X"04",
		X"43",X"50",X"82",X"FF",X"10",X"83",X"02",X"00",X"24",X"10",X"FC",X"A1",X"AE",X"4D",X"2C",X"04",
		X"43",X"50",X"82",X"FF",X"10",X"83",X"01",X"00",X"25",X"1F",X"FC",X"A1",X"AE",X"FD",X"99",X"0E",
		X"43",X"50",X"82",X"FF",X"DD",X"44",X"FC",X"A1",X"B0",X"FD",X"99",X"0C",X"43",X"50",X"82",X"FF",
		X"DD",X"46",X"35",X"36",X"EC",X"3E",X"DD",X"42",X"39",X"35",X"36",X"7E",X"47",X"55",X"34",X"36",
		X"FC",X"A1",X"B0",X"4D",X"2C",X"04",X"43",X"50",X"82",X"FF",X"10",X"83",X"02",X"00",X"24",X"10",
		X"FC",X"A1",X"AE",X"4D",X"2C",X"04",X"43",X"50",X"82",X"FF",X"10",X"83",X"01",X"00",X"25",X"31",
		X"FC",X"A1",X"AE",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"43",X"50",X"82",X"FF",X"F3",
		X"A1",X"AE",X"FD",X"A1",X"AE",X"FC",X"A1",X"B0",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",
		X"43",X"50",X"82",X"FF",X"F3",X"A1",X"B0",X"FD",X"A1",X"B0",X"35",X"36",X"EC",X"3E",X"DD",X"42",
		X"39",X"35",X"36",X"7E",X"47",X"55",X"34",X"36",X"B6",X"A0",X"3E",X"84",X"03",X"26",X"16",X"8E",
		X"4E",X"43",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"60",X"BD",X"E2",X"03",X"C6",X"99",X"86",X"61",
		X"BD",X"E2",X"03",X"20",X"46",X"4A",X"26",X"16",X"8E",X"4E",X"39",X"BD",X"2E",X"44",X"C6",X"DD",
		X"86",X"60",X"BD",X"E2",X"03",X"C6",X"99",X"86",X"62",X"BD",X"E2",X"03",X"20",X"2D",X"4A",X"26",
		X"16",X"8E",X"4E",X"38",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"60",X"BD",X"E2",X"03",X"C6",X"99",
		X"86",X"63",X"BD",X"E2",X"03",X"20",X"14",X"8E",X"4E",X"2B",X"BD",X"2E",X"44",X"C6",X"DD",X"86",
		X"60",X"BD",X"E2",X"03",X"C6",X"99",X"86",X"64",X"BD",X"E2",X"03",X"C6",X"DD",X"86",X"65",X"BD",
		X"E2",X"03",X"8E",X"3A",X"40",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"66",X"BD",X"E2",X"03",X"86",
		X"58",X"BD",X"E2",X"03",X"86",X"67",X"BD",X"E2",X"03",X"20",X"64",X"34",X"36",X"8E",X"4E",X"4E",
		X"BD",X"2E",X"44",X"C6",X"99",X"86",X"68",X"BD",X"E2",X"03",X"8E",X"2E",X"2B",X"BD",X"2E",X"44",
		X"C6",X"99",X"86",X"69",X"BD",X"E2",X"03",X"86",X"6A",X"BD",X"E2",X"03",X"86",X"6B",X"BD",X"E2",
		X"03",X"86",X"6C",X"BD",X"E2",X"03",X"20",X"37",X"34",X"36",X"8E",X"4E",X"36",X"BD",X"2E",X"44",
		X"C6",X"FF",X"86",X"6B",X"BD",X"E2",X"03",X"86",X"67",X"BD",X"E2",X"03",X"86",X"6D",X"BD",X"E2",
		X"03",X"86",X"6E",X"BD",X"E2",X"03",X"8E",X"46",X"3A",X"BD",X"2E",X"44",X"86",X"6F",X"BD",X"E2",
		X"03",X"86",X"59",X"BD",X"E2",X"03",X"86",X"5A",X"BD",X"E2",X"03",X"20",X"02",X"34",X"36",X"35",
		X"36",X"EC",X"3E",X"DD",X"42",X"39",X"7F",X"FF",X"1F",X"FF",X"48",X"EC",X"00",X"FA",X"01",X"00",
		X"48",X"E8",X"00",X"64",X"00",X"70",X"48",X"EE",X"00",X"40",X"00",X"70",X"48",X"EE",X"00",X"30",
		X"00",X"60",X"48",X"EE",X"00",X"20",X"00",X"40",X"48",X"EE",X"00",X"10",X"00",X"20",X"48",X"F0",
		X"00",X"00",X"00",X"00",X"48",X"F2",X"34",X"10",X"30",X"A4",X"AD",X"D8",X"07",X"35",X"90",X"34",
		X"36",X"0D",X"94",X"26",X"08",X"BE",X"A0",X"14",X"8C",X"4F",X"B2",X"26",X"2A",X"30",X"A4",X"AD",
		X"D8",X"07",X"86",X"00",X"BD",X"48",X"02",X"4D",X"2B",X"1D",X"86",X"20",X"BD",X"55",X"93",X"8E",
		X"7A",X"00",X"BD",X"55",X"83",X"C6",X"FF",X"86",X"5B",X"BD",X"E2",X"0C",X"8E",X"76",X"00",X"BD",
		X"55",X"83",X"86",X"5C",X"BD",X"E2",X"0C",X"35",X"36",X"39",X"0D",X"94",X"27",X"03",X"BD",X"5D",
		X"7B",X"34",X"10",X"30",X"A4",X"AD",X"D8",X"07",X"35",X"10",X"39",X"34",X"06",X"FC",X"A0",X"14",
		X"10",X"B3",X"A0",X"16",X"27",X"19",X"7D",X"A1",X"B2",X"26",X"14",X"BD",X"3D",X"4E",X"BD",X"38",
		X"91",X"4D",X"CE",X"FC",X"A0",X"14",X"10",X"B3",X"A0",X"16",X"26",X"03",X"BD",X"5D",X"A2",X"35",
		X"06",X"39",X"BD",X"53",X"6C",X"02",X"34",X"22",X"10",X"AE",X"9F",X"98",X"78",X"86",X"00",X"BD",
		X"48",X"02",X"B7",X"A1",X"B5",X"84",X"F0",X"8A",X"0C",X"A7",X"2C",X"35",X"22",X"39",X"7E",X"E1",
		X"B7",X"32",X"62",X"EC",X"28",X"34",X"02",X"1D",X"DD",X"83",X"35",X"04",X"1D",X"DD",X"81",X"0A",
		X"94",X"BD",X"55",X"A0",X"CC",X"5D",X"D9",X"ED",X"22",X"E6",X"26",X"DB",X"61",X"1D",X"D3",X"81",
		X"DD",X"81",X"E6",X"27",X"DB",X"62",X"1D",X"D3",X"83",X"DD",X"83",X"C3",X"00",X"80",X"4D",X"26",
		X"08",X"DC",X"81",X"C3",X"00",X"80",X"4D",X"27",X"51",X"9E",X"83",X"DC",X"81",X"34",X"16",X"2A",
		X"01",X"40",X"D6",X"83",X"2A",X"01",X"50",X"64",X"E4",X"66",X"61",X"64",X"62",X"66",X"63",X"4D",
		X"26",X"03",X"5D",X"27",X"04",X"44",X"54",X"20",X"EE",X"A6",X"61",X"E6",X"63",X"32",X"64",X"BD",
		X"47",X"82",X"8B",X"20",X"C6",X"80",X"48",X"25",X"0E",X"48",X"24",X"06",X"43",X"8B",X"80",X"5A",
		X"20",X"11",X"8B",X"80",X"5A",X"20",X"0A",X"48",X"24",X"04",X"8B",X"80",X"20",X"05",X"43",X"8B",
		X"80",X"1E",X"89",X"ED",X"28",X"EC",X"3E",X"DD",X"42",X"39",X"0F",X"94",X"34",X"20",X"86",X"30",
		X"BD",X"55",X"93",X"8E",X"7A",X"00",X"BD",X"55",X"83",X"C6",X"DD",X"86",X"6C",X"BD",X"E2",X"0C",
		X"86",X"6E",X"BD",X"E2",X"0C",X"86",X"70",X"BD",X"E2",X"0C",X"8E",X"76",X"00",X"BD",X"55",X"83",
		X"86",X"71",X"BD",X"E2",X"0C",X"86",X"72",X"BD",X"E2",X"0C",X"86",X"73",X"BD",X"E2",X"0C",X"35",
		X"20",X"BD",X"6C",X"80",X"CC",X"41",X"07",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"0F",X"A0",
		X"7F",X"FF",X"48",X"EC",X"02",X"00",X"11",X"00",X"48",X"EA",X"00",X"80",X"06",X"00",X"48",X"EC",
		X"00",X"40",X"04",X"00",X"48",X"EC",X"00",X"20",X"02",X"00",X"48",X"EC",X"00",X"10",X"01",X"00",
		X"48",X"EE",X"00",X"08",X"00",X"C0",X"48",X"F0",X"00",X"00",X"00",X"40",X"48",X"F2",X"7F",X"FF",
		X"07",X"FF",X"48",X"E8",X"0F",X"A0",X"10",X"00",X"48",X"EA",X"04",X"00",X"00",X"80",X"48",X"F0",
		X"02",X"58",X"01",X"40",X"48",X"E8",X"00",X"50",X"01",X"00",X"48",X"EC",X"00",X"40",X"00",X"C0",
		X"48",X"EA",X"00",X"20",X"00",X"80",X"48",X"EA",X"00",X"10",X"00",X"60",X"48",X"EC",X"00",X"00",
		X"00",X"40",X"48",X"EE",X"7F",X"FF",X"1F",X"FF",X"48",X"EC",X"00",X"64",X"02",X"00",X"48",X"EA",
		X"00",X"30",X"01",X"C0",X"48",X"EC",X"00",X"28",X"01",X"70",X"48",X"EC",X"00",X"20",X"01",X"48",
		X"48",X"EC",X"00",X"18",X"00",X"F8",X"48",X"EE",X"00",X"10",X"00",X"80",X"48",X"EE",X"00",X"08",
		X"00",X"30",X"48",X"F0",X"00",X"04",X"00",X"00",X"48",X"F0",X"00",X"00",X"00",X"00",X"48",X"F2",
		X"04",X"00",X"0F",X"FF",X"48",X"EA",X"01",X"28",X"03",X"00",X"48",X"EA",X"00",X"88",X"02",X"00",
		X"48",X"EA",X"00",X"40",X"01",X"00",X"48",X"EC",X"00",X"28",X"00",X"80",X"48",X"EC",X"00",X"18",
		X"00",X"00",X"48",X"EE",X"00",X"08",X"00",X"00",X"48",X"F0",X"00",X"00",X"FF",X"F0",X"48",X"EA",
		X"06",X"00",X"04",X"10",X"48",X"EC",X"00",X"00",X"03",X"00",X"48",X"EA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"A0",
		X"0F",X"FF",X"48",X"EE",X"00",X"50",X"03",X"00",X"48",X"EC",X"00",X"40",X"02",X"C0",X"48",X"EC",
		X"00",X"30",X"02",X"40",X"48",X"EE",X"00",X"20",X"02",X"00",X"48",X"EE",X"00",X"10",X"01",X"00",
		X"48",X"F0",X"00",X"08",X"00",X"80",X"48",X"F0",X"00",X"00",X"00",X"00",X"48",X"F2",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"0F",X"FF",X"48",X"EC",
		X"02",X"00",X"04",X"50",X"48",X"EA",X"01",X"00",X"03",X"C5",X"48",X"EA",X"00",X"80",X"03",X"20",
		X"48",X"EC",X"00",X"40",X"02",X"00",X"48",X"EC",X"00",X"20",X"01",X"80",X"48",X"EE",X"00",X"10",
		X"00",X"E0",X"48",X"EE",X"00",X"00",X"00",X"90",X"48",X"F0",X"18",X"00",X"04",X"10",X"48",X"EC",
		X"0C",X"80",X"02",X"A0",X"48",X"EE",X"06",X"00",X"01",X"90",X"48",X"F0",X"05",X"00",X"01",X"80",
		X"48",X"F0",X"04",X"00",X"01",X"60",X"48",X"F0",X"03",X"00",X"01",X"20",X"48",X"F0",X"02",X"00",
		X"00",X"C0",X"48",X"F0",X"01",X"00",X"00",X"70",X"48",X"EC",X"00",X"00",X"00",X"30",X"48",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",
		X"31",X"39",X"38",X"33",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",
		X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"06",
		X"00",X"04",X"10",X"48",X"EC",X"00",X"50",X"03",X"00",X"48",X"EA",X"00",X"40",X"02",X"C0",X"48",
		X"EA",X"00",X"30",X"02",X"40",X"48",X"EC",X"00",X"20",X"02",X"00",X"48",X"EC",X"00",X"08",X"01",
		X"00",X"48",X"EE",X"00",X"00",X"00",X"C0",X"48",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"06",
		X"00",X"04",X"10",X"48",X"EC",X"00",X"30",X"02",X"40",X"48",X"EA",X"00",X"20",X"02",X"00",X"48",
		X"EC",X"00",X"08",X"01",X"00",X"48",X"EE",X"00",X"00",X"00",X"80",X"48",X"F0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"1F",X"FF",X"48",X"EC",X"00",X"64",X"00",X"E8",X"48",
		X"EE",X"00",X"40",X"00",X"A0",X"48",X"F2",X"00",X"20",X"00",X"70",X"48",X"F2",X"00",X"10",X"00",
		X"40",X"48",X"F0",X"00",X"00",X"00",X"00",X"48",X"EE",X"5F",X"60",X"5F",X"BA",X"60",X"E1",X"5F",
		X"30",X"7D",X"00",X"08",X"C0",X"48",X"EA",X"06",X"00",X"02",X"30",X"48",X"EA",X"05",X"00",X"01",
		X"E0",X"48",X"EA",X"04",X"00",X"01",X"A0",X"48",X"EA",X"03",X"00",X"01",X"50",X"48",X"EC",X"02",
		X"00",X"00",X"B0",X"48",X"EE",X"00",X"00",X"00",X"40",X"48",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7D",X"00",X"07",
		X"D0",X"48",X"EA",X"0C",X"80",X"02",X"10",X"48",X"EC",X"06",X"00",X"01",X"C0",X"48",X"EE",X"05",
		X"00",X"01",X"70",X"48",X"EE",X"04",X"00",X"01",X"48",X"48",X"EE",X"03",X"00",X"00",X"F8",X"48",
		X"EE",X"02",X"00",X"00",X"80",X"48",X"F0",X"01",X"00",X"00",X"30",X"48",X"F0",X"00",X"00",X"00",
		X"00",X"48",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"61",X"61",X"61",X"62",X"61",X"64",X"61",
		X"67",X"80",X"80",X"C0",X"80",X"C0",X"A0",X"80",X"40",X"80",X"40",X"34",X"36",X"10",X"AE",X"B8",
		X"04",X"4F",X"E6",X"A8",X"1D",X"8E",X"61",X"81",X"AD",X"95",X"35",X"36",X"EC",X"3E",X"DD",X"42",
		X"39",X"61",X"8D",X"61",X"A6",X"62",X"00",X"62",X"37",X"62",X"B7",X"FF",X"FF",X"34",X"76",X"AE",
		X"B8",X"11",X"A6",X"A8",X"1A",X"8B",X"10",X"A7",X"A8",X"1A",X"86",X"02",X"BD",X"69",X"DA",X"10",
		X"24",X"00",X"14",X"35",X"76",X"39",X"34",X"76",X"AE",X"B8",X"11",X"BD",X"69",X"DA",X"10",X"25",
		X"00",X"4B",X"BD",X"64",X"96",X"86",X"08",X"34",X"10",X"BD",X"64",X"D2",X"F6",X"A1",X"B6",X"34",
		X"02",X"34",X"04",X"BD",X"63",X"5A",X"34",X"06",X"8E",X"5F",X"EA",X"BD",X"65",X"03",X"BD",X"65",
		X"40",X"AE",X"64",X"A6",X"63",X"E6",X"62",X"BD",X"63",X"96",X"34",X"06",X"8E",X"5F",X"EA",X"BD",
		X"65",X"03",X"BD",X"65",X"69",X"35",X"06",X"58",X"49",X"58",X"49",X"34",X"02",X"EC",X"61",X"58",
		X"49",X"58",X"49",X"35",X"04",X"BD",X"47",X"82",X"BD",X"62",X"C8",X"32",X"66",X"35",X"76",X"39",
		X"34",X"76",X"AE",X"B8",X"11",X"BD",X"64",X"D2",X"A6",X"A8",X"1A",X"BD",X"62",X"C8",X"BD",X"69",
		X"DA",X"10",X"25",X"00",X"1F",X"BD",X"64",X"96",X"34",X"10",X"BD",X"63",X"38",X"8E",X"60",X"4F",
		X"BD",X"65",X"03",X"BD",X"65",X"40",X"35",X"10",X"BD",X"63",X"49",X"8E",X"60",X"4F",X"BD",X"65",
		X"03",X"BD",X"65",X"69",X"35",X"76",X"39",X"34",X"76",X"AE",X"B8",X"11",X"BD",X"69",X"DA",X"10",
		X"25",X"00",X"71",X"BD",X"63",X"F7",X"BD",X"64",X"96",X"7D",X"A1",X"BB",X"26",X"17",X"FC",X"A0",
		X"14",X"10",X"B3",X"A0",X"16",X"27",X"0E",X"7D",X"A0",X"3E",X"26",X"15",X"FC",X"A0",X"16",X"10",
		X"83",X"4F",X"E2",X"26",X"0C",X"BD",X"62",X"6A",X"20",X"43",X"34",X"76",X"86",X"20",X"7E",X"61",
		X"B7",X"BD",X"64",X"D2",X"BD",X"63",X"38",X"8E",X"60",X"7F",X"BD",X"65",X"03",X"BD",X"65",X"40",
		X"AE",X"9F",X"98",X"78",X"BD",X"63",X"49",X"8E",X"60",X"7F",X"BD",X"65",X"03",X"BD",X"65",X"69",
		X"A6",X"A8",X"1A",X"BD",X"62",X"C8",X"A6",X"A8",X"18",X"AA",X"A8",X"19",X"85",X"FC",X"26",X"0D",
		X"BD",X"5D",X"7B",X"EC",X"3E",X"ED",X"A8",X"11",X"1F",X"21",X"BD",X"6C",X"73",X"AE",X"9F",X"98",
		X"78",X"BD",X"64",X"79",X"35",X"76",X"39",X"34",X"76",X"BD",X"69",X"DA",X"25",X"07",X"AE",X"9F",
		X"50",X"35",X"7E",X"61",X"B5",X"35",X"76",X"39",X"34",X"26",X"10",X"AE",X"2A",X"27",X"19",X"A6",
		X"E4",X"8B",X"08",X"47",X"47",X"47",X"47",X"8B",X"08",X"C6",X"08",X"3D",X"C3",X"12",X"9D",X"ED",
		X"A8",X"16",X"CC",X"43",X"B8",X"ED",X"A8",X"18",X"35",X"26",X"39",X"34",X"60",X"EE",X"0A",X"27",
		X"1A",X"10",X"AE",X"9F",X"50",X"35",X"10",X"AE",X"2A",X"4F",X"E6",X"25",X"58",X"89",X"00",X"34",
		X"06",X"4F",X"E6",X"45",X"58",X"89",X"00",X"A3",X"E1",X"20",X"07",X"E6",X"08",X"1D",X"58",X"49",
		X"58",X"49",X"35",X"60",X"39",X"34",X"60",X"EE",X"0A",X"27",X"13",X"10",X"AE",X"9F",X"50",X"35",
		X"10",X"AE",X"2A",X"E6",X"27",X"4F",X"34",X"06",X"E6",X"47",X"A3",X"E1",X"20",X"07",X"E6",X"09",
		X"1D",X"58",X"49",X"58",X"49",X"35",X"60",X"39",X"34",X"10",X"BD",X"62",X"EB",X"34",X"06",X"30",
		X"A4",X"BD",X"62",X"EB",X"A3",X"E1",X"35",X"10",X"39",X"34",X"10",X"BD",X"63",X"15",X"34",X"06",
		X"30",X"A4",X"BD",X"63",X"15",X"A3",X"E1",X"35",X"10",X"39",X"34",X"32",X"A6",X"08",X"5F",X"BD",
		X"48",X"EE",X"34",X"06",X"BD",X"64",X"DD",X"BD",X"47",X"DA",X"E6",X"62",X"50",X"BD",X"47",X"BE",
		X"E3",X"E4",X"ED",X"E4",X"E6",X"06",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"58",
		X"49",X"58",X"49",X"58",X"49",X"E3",X"E4",X"ED",X"E4",X"5F",X"A6",X"28",X"BD",X"48",X"EE",X"A3",
		X"E1",X"32",X"61",X"35",X"30",X"39",X"34",X"32",X"A6",X"09",X"5F",X"BD",X"48",X"EE",X"34",X"06",
		X"BD",X"64",X"DD",X"BD",X"47",X"DA",X"A6",X"62",X"BD",X"47",X"BE",X"E3",X"E4",X"ED",X"E4",X"E6",
		X"06",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",
		X"E3",X"E4",X"ED",X"E4",X"5F",X"A6",X"29",X"BD",X"48",X"EE",X"A3",X"E1",X"32",X"61",X"35",X"30",
		X"39",X"34",X"40",X"EE",X"0A",X"27",X"04",X"EC",X"4E",X"20",X"06",X"12",X"A6",X"06",X"5F",X"47",
		X"56",X"35",X"40",X"39",X"34",X"40",X"EE",X"0A",X"27",X"04",X"EC",X"4E",X"20",X"06",X"12",X"A6",
		X"07",X"5F",X"47",X"56",X"35",X"40",X"39",X"34",X"46",X"A6",X"08",X"E6",X"09",X"DD",X"02",X"9B",
		X"8D",X"29",X"02",X"A7",X"08",X"DB",X"8E",X"29",X"02",X"E7",X"09",X"EE",X"0A",X"27",X"26",X"A6",
		X"45",X"E6",X"47",X"DD",X"00",X"34",X"04",X"9B",X"91",X"81",X"C0",X"25",X"01",X"4F",X"A7",X"45",
		X"E6",X"C8",X"10",X"1D",X"35",X"04",X"DB",X"92",X"89",X"00",X"27",X"07",X"2B",X"04",X"C6",X"FF",
		X"20",X"01",X"5F",X"E7",X"47",X"35",X"46",X"39",X"34",X"46",X"A6",X"08",X"E6",X"09",X"DD",X"02",
		X"9B",X"8B",X"29",X"02",X"A7",X"08",X"DB",X"8C",X"29",X"02",X"E7",X"09",X"EE",X"0A",X"27",X"26",
		X"A6",X"45",X"E6",X"47",X"DD",X"00",X"34",X"04",X"9B",X"8F",X"81",X"C0",X"25",X"01",X"4F",X"A7",
		X"45",X"E6",X"C8",X"10",X"1D",X"35",X"04",X"DB",X"90",X"89",X"00",X"27",X"07",X"2B",X"04",X"C6",
		X"FF",X"20",X"01",X"5F",X"E7",X"47",X"35",X"46",X"39",X"34",X"46",X"DC",X"02",X"A7",X"08",X"E7",
		X"09",X"EE",X"0A",X"27",X"06",X"DC",X"00",X"A7",X"45",X"E7",X"47",X"35",X"46",X"39",X"34",X"16",
		X"AE",X"9F",X"50",X"35",X"20",X"05",X"34",X"16",X"AE",X"B8",X"11",X"4F",X"9C",X"78",X"26",X"04",
		X"A6",X"89",X"98",X"8D",X"AB",X"08",X"A1",X"28",X"2D",X"04",X"A0",X"28",X"20",X"04",X"A6",X"28",
		X"A0",X"08",X"A7",X"A8",X"18",X"4F",X"9C",X"78",X"26",X"04",X"A6",X"89",X"98",X"8E",X"AB",X"09",
		X"A1",X"29",X"2D",X"04",X"A0",X"29",X"20",X"04",X"A6",X"29",X"A0",X"09",X"A7",X"A8",X"19",X"35",
		X"16",X"39",X"34",X"02",X"BD",X"64",X"DD",X"A7",X"A8",X"1A",X"35",X"02",X"39",X"34",X"04",X"A6",
		X"28",X"A0",X"08",X"28",X"09",X"34",X"01",X"86",X"7F",X"35",X"01",X"2E",X"01",X"43",X"E6",X"29",
		X"E0",X"09",X"28",X"09",X"34",X"01",X"C6",X"7F",X"35",X"01",X"2E",X"01",X"53",X"BD",X"47",X"82",
		X"35",X"04",X"39",X"34",X"12",X"6F",X"E4",X"6A",X"E4",X"4D",X"2C",X"06",X"60",X"E4",X"43",X"50",
		X"82",X"FF",X"10",X"A3",X"84",X"2C",X"04",X"30",X"06",X"20",X"F7",X"EC",X"02",X"6D",X"E0",X"2C",
		X"04",X"43",X"50",X"82",X"FF",X"35",X"10",X"1F",X"13",X"34",X"06",X"4D",X"2C",X"04",X"43",X"50",
		X"82",X"FF",X"10",X"A3",X"42",X"2C",X"04",X"33",X"46",X"20",X"F7",X"EE",X"44",X"35",X"06",X"39",
		X"34",X"26",X"BD",X"65",X"EE",X"34",X"06",X"E6",X"26",X"4F",X"BD",X"48",X"F0",X"93",X"44",X"1F",
		X"02",X"35",X"06",X"BD",X"65",X"B9",X"10",X"AE",X"62",X"10",X"AE",X"2A",X"26",X"07",X"10",X"AE",
		X"62",X"31",X"26",X"20",X"29",X"31",X"2E",X"20",X"41",X"34",X"26",X"58",X"49",X"BD",X"65",X"EE",
		X"34",X"06",X"E6",X"27",X"4F",X"BD",X"48",X"F0",X"93",X"46",X"1F",X"02",X"35",X"06",X"BD",X"65",
		X"B9",X"10",X"AE",X"62",X"10",X"AE",X"2A",X"26",X"1E",X"10",X"AE",X"62",X"31",X"27",X"BD",X"48",
		X"E6",X"E0",X"A4",X"27",X"10",X"1D",X"AD",X"C4",X"5D",X"2B",X"04",X"CA",X"01",X"20",X"02",X"C4",
		X"FE",X"EB",X"A4",X"E7",X"A4",X"20",X"0F",X"31",X"2C",X"12",X"A3",X"A4",X"27",X"08",X"AD",X"C4",
		X"CA",X"01",X"E3",X"A4",X"ED",X"A4",X"35",X"26",X"39",X"34",X"26",X"1F",X"20",X"4D",X"2D",X"0F",
		X"6D",X"E4",X"2D",X"25",X"E3",X"E1",X"10",X"A3",X"02",X"2F",X"20",X"EC",X"02",X"20",X"1C",X"6D",
		X"E4",X"2C",X"16",X"E3",X"E1",X"34",X"06",X"4D",X"2C",X"04",X"43",X"50",X"82",X"FF",X"10",X"A3",
		X"02",X"2F",X"06",X"4F",X"5F",X"A3",X"02",X"ED",X"E4",X"35",X"06",X"35",X"20",X"39",X"34",X"40",
		X"EE",X"24",X"11",X"83",X"4C",X"8F",X"27",X"0C",X"11",X"83",X"4C",X"EF",X"27",X"0D",X"10",X"AE",
		X"B8",X"11",X"35",X"C0",X"10",X"AE",X"9F",X"98",X"78",X"35",X"C0",X"10",X"AE",X"9F",X"50",X"35",
		X"35",X"C0",X"34",X"36",X"10",X"AE",X"B8",X"04",X"BD",X"64",X"96",X"E6",X"A8",X"1D",X"8E",X"66",
		X"57",X"EE",X"2A",X"27",X"29",X"A6",X"45",X"81",X"08",X"23",X"23",X"81",X"6C",X"24",X"1F",X"A6",
		X"47",X"81",X"10",X"23",X"19",X"81",X"F0",X"24",X"15",X"34",X"04",X"A6",X"2C",X"1F",X"89",X"C4",
		X"0F",X"27",X"09",X"5A",X"34",X"04",X"84",X"F0",X"AA",X"E0",X"A7",X"2C",X"35",X"04",X"AD",X"95",
		X"35",X"36",X"EC",X"3E",X"DD",X"42",X"39",X"66",X"65",X"66",X"8D",X"66",X"F3",X"67",X"71",X"67",
		X"A7",X"67",X"DC",X"FF",X"FF",X"34",X"76",X"AE",X"9F",X"50",X"35",X"BD",X"66",X"78",X"BD",X"69",
		X"DA",X"10",X"24",X"00",X"6A",X"35",X"76",X"39",X"34",X"02",X"A6",X"A8",X"1A",X"34",X"02",X"BD",
		X"64",X"D2",X"35",X"02",X"BD",X"68",X"36",X"BD",X"68",X"4C",X"35",X"02",X"39",X"34",X"76",X"AE",
		X"B8",X"11",X"BD",X"66",X"78",X"BD",X"69",X"DA",X"24",X"09",X"35",X"76",X"7D",X"A1",X"B3",X"10",
		X"2C",X"C7",X"A1",X"1F",X"21",X"EC",X"88",X"16",X"10",X"83",X"00",X"00",X"26",X"06",X"AE",X"B8",
		X"11",X"7E",X"67",X"16",X"86",X"06",X"F6",X"A1",X"B7",X"AE",X"B8",X"11",X"BD",X"63",X"5A",X"8E",
		X"5F",X"EA",X"BD",X"65",X"03",X"BD",X"65",X"40",X"AE",X"B8",X"11",X"86",X"06",X"F6",X"A1",X"B7",
		X"BD",X"63",X"96",X"8E",X"5F",X"EA",X"BD",X"65",X"03",X"BD",X"65",X"69",X"7E",X"66",X"DF",X"BD",
		X"68",X"CC",X"25",X"0C",X"AE",X"9F",X"50",X"35",X"BD",X"6A",X"57",X"25",X"03",X"BD",X"68",X"DD",
		X"35",X"76",X"39",X"34",X"76",X"AE",X"B8",X"11",X"A6",X"A8",X"1A",X"34",X"02",X"BD",X"64",X"D2",
		X"35",X"02",X"BD",X"68",X"36",X"BD",X"68",X"4C",X"BD",X"69",X"DA",X"24",X"09",X"35",X"76",X"7D",
		X"A1",X"B3",X"10",X"2C",X"C7",X"2E",X"BD",X"63",X"38",X"34",X"06",X"8E",X"5F",X"30",X"BD",X"65",
		X"03",X"BD",X"65",X"40",X"AE",X"B8",X"11",X"BD",X"63",X"49",X"34",X"06",X"8E",X"5F",X"30",X"BD",
		X"65",X"03",X"BD",X"65",X"69",X"AE",X"B8",X"11",X"EC",X"E4",X"2C",X"04",X"43",X"50",X"82",X"FF",
		X"10",X"83",X"00",X"50",X"2E",X"26",X"EC",X"62",X"2C",X"04",X"43",X"50",X"82",X"FF",X"10",X"83",
		X"00",X"50",X"2E",X"18",X"CC",X"02",X"02",X"BD",X"47",X"FA",X"4D",X"26",X"0F",X"A6",X"A8",X"1D",
		X"81",X"04",X"27",X"05",X"32",X"64",X"7E",X"66",X"DF",X"BD",X"68",X"DD",X"32",X"64",X"35",X"76",
		X"39",X"BD",X"69",X"DA",X"24",X"01",X"39",X"34",X"76",X"AE",X"9F",X"50",X"35",X"BD",X"66",X"78",
		X"86",X"08",X"F6",X"A1",X"B7",X"AE",X"B8",X"11",X"34",X"16",X"BD",X"63",X"5A",X"8E",X"61",X"1D",
		X"BD",X"65",X"03",X"BD",X"65",X"40",X"35",X"16",X"BD",X"63",X"96",X"8E",X"61",X"1D",X"BD",X"65",
		X"03",X"BD",X"65",X"69",X"7E",X"66",X"DF",X"34",X"76",X"AE",X"B8",X"11",X"BD",X"66",X"78",X"BD",
		X"69",X"DA",X"24",X"03",X"35",X"76",X"39",X"BD",X"63",X"38",X"8E",X"5F",X"BA",X"BD",X"65",X"03",
		X"BD",X"65",X"40",X"AE",X"B8",X"11",X"BD",X"63",X"49",X"8E",X"5F",X"BA",X"BD",X"65",X"03",X"BD",
		X"65",X"69",X"0D",X"96",X"26",X"DE",X"AE",X"B8",X"11",X"7E",X"66",X"DF",X"34",X"76",X"BD",X"69",
		X"DA",X"25",X"50",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"38",X"BD",X"66",X"78",X"86",X"06",X"F6",
		X"A1",X"B7",X"1F",X"21",X"BD",X"65",X"EE",X"1E",X"12",X"34",X"16",X"BD",X"63",X"5A",X"8E",X"60",
		X"B5",X"BD",X"65",X"03",X"BD",X"65",X"40",X"35",X"16",X"BD",X"63",X"96",X"8E",X"60",X"B5",X"BD",
		X"65",X"03",X"BD",X"65",X"69",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"79",X"CC",X"02",X"08",X"BD",
		X"47",X"FA",X"8B",X"FF",X"25",X"0D",X"B6",X"A0",X"13",X"27",X"08",X"BD",X"E1",X"F1",X"27",X"03",
		X"BD",X"6C",X"5E",X"35",X"76",X"39",X"34",X"02",X"A6",X"A8",X"1A",X"A0",X"E0",X"AB",X"A8",X"20",
		X"47",X"4C",X"84",X"FE",X"A7",X"A8",X"20",X"48",X"AB",X"A8",X"1A",X"39",X"34",X"36",X"10",X"8C",
		X"A1",X"38",X"27",X"51",X"AE",X"2A",X"27",X"4A",X"E6",X"2C",X"C4",X"7F",X"A0",X"A8",X"1F",X"2A",
		X"01",X"40",X"81",X"20",X"2E",X"05",X"A6",X"A8",X"1F",X"20",X"02",X"A6",X"E4",X"8B",X"10",X"84",
		X"E0",X"A0",X"A8",X"1F",X"81",X"20",X"2F",X"04",X"86",X"20",X"CA",X"80",X"81",X"E0",X"2C",X"04",
		X"86",X"E0",X"CA",X"80",X"AB",X"A8",X"1F",X"E7",X"2C",X"A7",X"A8",X"1F",X"47",X"47",X"47",X"47",
		X"47",X"8B",X"04",X"C6",X"08",X"3D",X"C3",X"1A",X"93",X"ED",X"88",X"1E",X"CC",X"45",X"F9",X"ED",
		X"88",X"1A",X"35",X"36",X"39",X"8B",X"80",X"97",X"50",X"20",X"F7",X"34",X"70",X"10",X"AE",X"B8",
		X"0D",X"EE",X"24",X"DF",X"04",X"AE",X"98",X"0D",X"EE",X"04",X"EF",X"24",X"35",X"70",X"39",X"34",
		X"60",X"10",X"AE",X"B8",X"0D",X"DE",X"04",X"EF",X"24",X"35",X"60",X"39",X"34",X"06",X"4F",X"5F",
		X"10",X"A3",X"2A",X"35",X"06",X"27",X"03",X"1C",X"FE",X"39",X"1A",X"01",X"39",X"34",X"76",X"EE",
		X"0A",X"10",X"27",X"00",X"ED",X"EE",X"2A",X"10",X"27",X"00",X"E7",X"96",X"75",X"10",X"27",X"00",
		X"E1",X"A6",X"45",X"81",X"08",X"10",X"23",X"00",X"D9",X"81",X"6C",X"10",X"24",X"00",X"D3",X"A6",
		X"47",X"81",X"10",X"10",X"23",X"00",X"CB",X"81",X"F0",X"10",X"24",X"00",X"C5",X"A6",X"A8",X"1D",
		X"81",X"04",X"27",X"08",X"A6",X"2C",X"84",X"0F",X"10",X"26",X"00",X"B6",X"10",X"8C",X"A1",X"38",
		X"10",X"27",X"00",X"B1",X"BD",X"64",X"DD",X"34",X"02",X"A6",X"A8",X"1F",X"8B",X"80",X"8B",X"10",
		X"84",X"E0",X"1F",X"89",X"E0",X"E0",X"2C",X"01",X"50",X"C1",X"10",X"2F",X"00",X"E6",X"2C",X"C5",
		X"80",X"10",X"26",X"00",X"8D",X"34",X"02",X"BD",X"38",X"91",X"4D",X"BA",X"BD",X"43",X"4F",X"10",
		X"8E",X"4D",X"1F",X"10",X"AF",X"88",X"12",X"E6",X"E4",X"C4",X"60",X"57",X"57",X"57",X"57",X"57",
		X"86",X"08",X"3D",X"C3",X"28",X"B0",X"1F",X"03",X"BD",X"43",X"32",X"A6",X"E4",X"BD",X"47",X"DA",
		X"1E",X"89",X"34",X"02",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"10",X"AE",X"66",X"10",X"AE",
		X"2A",X"E3",X"2C",X"ED",X"0C",X"35",X"04",X"1D",X"58",X"49",X"58",X"49",X"10",X"AE",X"65",X"10",
		X"AE",X"2A",X"E3",X"2E",X"ED",X"0E",X"10",X"AE",X"65",X"35",X"02",X"10",X"AE",X"2A",X"34",X"20",
		X"10",X"AE",X"A8",X"14",X"A6",X"26",X"A0",X"46",X"5F",X"BD",X"48",X"F0",X"34",X"06",X"A6",X"27",
		X"A0",X"47",X"5F",X"10",X"AE",X"62",X"EB",X"28",X"A9",X"27",X"A7",X"07",X"E7",X"08",X"A7",X"06",
		X"35",X"06",X"35",X"20",X"EB",X"24",X"A9",X"25",X"A7",X"05",X"E7",X"04",X"6F",X"88",X"10",X"BD",
		X"43",X"5E",X"35",X"76",X"39",X"BD",X"39",X"1D",X"20",X"F8",X"34",X"42",X"A6",X"2C",X"EE",X"2A",
		X"26",X"04",X"85",X"20",X"26",X"09",X"8A",X"20",X"A7",X"2C",X"35",X"42",X"1C",X"FE",X"39",X"84",
		X"DF",X"A7",X"2C",X"35",X"42",X"1A",X"01",X"39",X"34",X"36",X"E6",X"A8",X"1D",X"C4",X"FE",X"2D",
		X"09",X"C1",X"0C",X"2C",X"05",X"8E",X"6A",X"0E",X"6E",X"95",X"C6",X"00",X"20",X"F7",X"6A",X"18",
		X"6A",X"1D",X"6A",X"1D",X"6A",X"1D",X"6A",X"1D",X"8E",X"A1",X"38",X"20",X"03",X"AE",X"B8",X"11",
		X"BD",X"64",X"D2",X"A6",X"A8",X"1A",X"A7",X"A8",X"1F",X"35",X"36",X"7E",X"42",X"B9",X"34",X"20",
		X"10",X"AE",X"B8",X"1C",X"BD",X"6A",X"3C",X"35",X"20",X"7E",X"46",X"2B",X"34",X"02",X"86",X"04",
		X"34",X"02",X"B6",X"A0",X"3C",X"43",X"6C",X"E4",X"8B",X"28",X"28",X"FA",X"A6",X"2C",X"84",X"F0",
		X"AA",X"E0",X"A7",X"2C",X"35",X"02",X"39",X"34",X"06",X"CC",X"00",X"A0",X"BD",X"47",X"FA",X"34",
		X"02",X"B6",X"A0",X"3C",X"8B",X"20",X"A1",X"E0",X"35",X"06",X"39",X"FA",X"8B",X"FF",X"35",X"06",
		X"39",X"34",X"76",X"10",X"AE",X"B8",X"04",X"BD",X"69",X"DA",X"10",X"25",X"00",X"83",X"EE",X"2A",
		X"26",X"0C",X"EE",X"B8",X"13",X"BD",X"6B",X"0E",X"EE",X"B8",X"15",X"BD",X"6B",X"0E",X"BE",X"A0",
		X"16",X"8C",X"4F",X"E2",X"27",X"09",X"FC",X"A0",X"14",X"10",X"83",X"4F",X"B2",X"27",X"62",X"AE",
		X"9F",X"98",X"78",X"BD",X"64",X"38",X"BD",X"63",X"38",X"34",X"06",X"8E",X"5E",X"8E",X"BD",X"65",
		X"03",X"BD",X"65",X"40",X"AE",X"9F",X"98",X"78",X"BD",X"63",X"49",X"34",X"06",X"BD",X"64",X"79",
		X"8E",X"5E",X"8E",X"BD",X"65",X"03",X"BD",X"65",X"69",X"EE",X"2A",X"26",X"3B",X"0D",X"94",X"26",
		X"37",X"AE",X"9F",X"98",X"78",X"EE",X"0A",X"26",X"2F",X"EC",X"62",X"4D",X"2C",X"04",X"43",X"50",
		X"82",X"FF",X"ED",X"62",X"35",X"06",X"4D",X"2C",X"04",X"43",X"50",X"82",X"FF",X"AA",X"E0",X"EA",
		X"E0",X"10",X"83",X"00",X"50",X"2E",X"0A",X"1F",X"21",X"EE",X"04",X"AD",X"D8",X"07",X"BD",X"58",
		X"B9",X"35",X"76",X"EC",X"3E",X"DD",X"42",X"39",X"35",X"06",X"35",X"06",X"20",X"F3",X"34",X"76",
		X"34",X"03",X"6F",X"61",X"6C",X"61",X"35",X"01",X"27",X"23",X"CC",X"00",X"14",X"A1",X"C8",X"18",
		X"25",X"16",X"E1",X"C8",X"19",X"25",X"11",X"EC",X"4A",X"26",X"0D",X"34",X"40",X"1F",X"31",X"EE",
		X"04",X"AD",X"D8",X"07",X"35",X"40",X"6F",X"E4",X"EE",X"D8",X"16",X"20",X"DB",X"6D",X"E0",X"26",
		X"24",X"1F",X"21",X"EE",X"04",X"AD",X"D8",X"07",X"86",X"20",X"BD",X"55",X"93",X"8E",X"7A",X"00",
		X"BD",X"55",X"83",X"C6",X"FF",X"86",X"5B",X"BD",X"E2",X"0C",X"8E",X"76",X"00",X"BD",X"55",X"83",
		X"86",X"5C",X"BD",X"E2",X"0C",X"35",X"76",X"39",X"34",X"76",X"FC",X"A0",X"16",X"10",X"83",X"4F",
		X"E2",X"10",X"26",X"00",X"6E",X"10",X"AE",X"9F",X"98",X"78",X"BD",X"69",X"DA",X"10",X"25",X"00",
		X"62",X"BD",X"64",X"8E",X"BD",X"53",X"26",X"E6",X"2C",X"A6",X"2C",X"C4",X"0F",X"27",X"0A",X"C1",
		X"09",X"2E",X"05",X"BD",X"68",X"CC",X"25",X"01",X"5A",X"34",X"04",X"84",X"F0",X"AA",X"E0",X"A7",
		X"2C",X"7D",X"A1",X"B9",X"27",X"03",X"7A",X"A1",X"B9",X"BD",X"6C",X"24",X"25",X"35",X"AE",X"9F",
		X"98",X"78",X"DC",X"8F",X"34",X"06",X"CC",X"04",X"12",X"DD",X"8F",X"BD",X"64",X"38",X"AE",X"9F",
		X"50",X"35",X"BD",X"6B",X"EA",X"BD",X"2D",X"FB",X"BD",X"65",X"40",X"AE",X"9F",X"50",X"35",X"BD",
		X"6C",X"07",X"BD",X"2D",X"FB",X"BD",X"65",X"69",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"79",X"35",
		X"06",X"DD",X"8F",X"35",X"76",X"EC",X"3E",X"DD",X"42",X"39",X"A6",X"2C",X"84",X"0F",X"27",X"10",
		X"F6",X"A1",X"B5",X"81",X"0C",X"2F",X"02",X"86",X"0C",X"BD",X"63",X"5A",X"8E",X"5E",X"F4",X"39",
		X"BD",X"63",X"38",X"8E",X"5E",X"BE",X"39",X"A6",X"2C",X"84",X"0F",X"27",X"10",X"F6",X"A1",X"B5",
		X"81",X"0C",X"2F",X"02",X"86",X"0C",X"BD",X"63",X"96",X"8E",X"5E",X"F4",X"39",X"BD",X"63",X"49",
		X"8E",X"5E",X"BE",X"39",X"34",X"20",X"7D",X"A1",X"B9",X"26",X"17",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"0D",X"96",X"27",X"05",X"BD",X"68",X"CC",X"24",X"04",X"1C",X"FE",
		X"20",X"11",X"6F",X"26",X"6F",X"27",X"10",X"AE",X"2A",X"27",X"06",X"4F",X"5F",X"ED",X"2E",X"ED",
		X"2C",X"1A",X"01",X"35",X"20",X"39",X"7E",X"6F",X"4C",X"7E",X"8C",X"8C",X"42",X"39",X"7E",X"6D",
		X"30",X"7E",X"73",X"5F",X"7E",X"6F",X"B0",X"7E",X"76",X"02",X"7E",X"75",X"B6",X"7E",X"7F",X"4B",
		X"7E",X"71",X"F6",X"7E",X"71",X"8D",X"7E",X"6F",X"30",X"7E",X"6F",X"14",X"7E",X"7B",X"B0",X"39",
		X"7E",X"79",X"EF",X"7C",X"A1",X"B4",X"7C",X"A1",X"B4",X"39",X"86",X"C3",X"B1",X"A1",X"B4",X"10",
		X"26",X"C1",X"B1",X"34",X"36",X"8E",X"43",X"51",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"74",X"BD",
		X"E2",X"03",X"30",X"1A",X"86",X"75",X"BD",X"E2",X"0C",X"30",X"0B",X"86",X"76",X"BD",X"E2",X"03",
		X"30",X"1A",X"86",X"77",X"BD",X"E2",X"0C",X"35",X"36",X"39",X"0D",X"96",X"26",X"08",X"86",X"01",
		X"97",X"86",X"86",X"08",X"97",X"87",X"78",X"A1",X"B4",X"39",X"0F",X"86",X"7D",X"A1",X"BD",X"10",
		X"26",X"C1",X"71",X"0D",X"8A",X"27",X"08",X"0D",X"96",X"10",X"27",X"C1",X"67",X"0F",X"8A",X"0F",
		X"96",X"7E",X"2E",X"D4",X"0F",X"86",X"0D",X"8A",X"26",X"05",X"0F",X"96",X"7E",X"2E",X"D4",X"0D",
		X"96",X"10",X"26",X"EB",X"3D",X"39",X"0D",X"96",X"10",X"26",X"C1",X"48",X"B6",X"A0",X"13",X"10",
		X"26",X"FF",X"5B",X"86",X"10",X"BD",X"55",X"93",X"8E",X"7A",X"00",X"BD",X"55",X"83",X"C6",X"AA",
		X"86",X"78",X"BD",X"E2",X"0C",X"86",X"56",X"BD",X"E2",X"0C",X"86",X"79",X"BD",X"E2",X"0C",X"8E",
		X"76",X"00",X"BD",X"55",X"83",X"86",X"7A",X"BD",X"E2",X"0C",X"86",X"5B",X"BD",X"E2",X"0C",X"39",
		X"34",X"36",X"C6",X"12",X"BD",X"3C",X"23",X"7C",X"A1",X"B8",X"7A",X"A0",X"13",X"26",X"03",X"BD",
		X"52",X"F5",X"BD",X"38",X"91",X"4D",X"D3",X"CC",X"00",X"00",X"8E",X"4C",X"8F",X"AD",X"98",X"05",
		X"31",X"84",X"AE",X"9F",X"98",X"78",X"BD",X"64",X"38",X"BD",X"64",X"DD",X"8B",X"80",X"BD",X"64",
		X"79",X"BD",X"47",X"DA",X"34",X"06",X"35",X"04",X"1D",X"58",X"49",X"F3",X"99",X"0C",X"AE",X"2A",
		X"ED",X"0C",X"35",X"04",X"1D",X"F3",X"99",X"0E",X"ED",X"0E",X"35",X"36",X"39",X"8E",X"BF",X"1B",
		X"BD",X"4A",X"5F",X"4D",X"26",X"03",X"77",X"A1",X"B4",X"86",X"C3",X"B1",X"A1",X"B4",X"26",X"19",
		X"8E",X"BF",X"1B",X"BD",X"4A",X"5F",X"81",X"30",X"26",X"0F",X"BD",X"46",X"DB",X"6D",X"AA",X"05",
		X"A1",X"6D",X"86",X"F0",X"A7",X"04",X"7F",X"A1",X"B4",X"39",X"6A",X"24",X"26",X"06",X"BD",X"32",
		X"0F",X"7E",X"47",X"55",X"BD",X"6C",X"93",X"34",X"36",X"8E",X"57",X"66",X"BD",X"2E",X"44",X"C6",
		X"FF",X"86",X"7B",X"BD",X"E2",X"0C",X"8E",X"57",X"87",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"7C",
		X"BD",X"E2",X"0C",X"8E",X"5F",X"6A",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"7D",X"BD",X"E2",X"0C",
		X"8E",X"5B",X"6A",X"BD",X"2E",X"44",X"86",X"7E",X"BD",X"E2",X"0C",X"8E",X"57",X"6A",X"BD",X"2E",
		X"44",X"86",X"7F",X"BD",X"E2",X"0C",X"8E",X"53",X"6A",X"BD",X"2E",X"44",X"86",X"80",X"BD",X"E2",
		X"0C",X"8E",X"47",X"6A",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"81",X"BD",X"E2",X"0C",X"8E",X"43",
		X"6A",X"BD",X"2E",X"44",X"86",X"7F",X"BD",X"E2",X"0C",X"8E",X"3F",X"6A",X"BD",X"2E",X"44",X"86",
		X"82",X"BD",X"E2",X"0C",X"8E",X"3B",X"6A",X"BD",X"2E",X"44",X"86",X"83",X"BD",X"E2",X"0C",X"8E",
		X"37",X"6A",X"BD",X"2E",X"44",X"86",X"84",X"BD",X"E2",X"0C",X"8E",X"33",X"6A",X"BD",X"2E",X"44",
		X"86",X"76",X"BD",X"E2",X"0C",X"8E",X"2F",X"6A",X"BD",X"2E",X"44",X"86",X"85",X"BD",X"E2",X"0C",
		X"8E",X"2B",X"6A",X"BD",X"2E",X"44",X"86",X"7D",X"BD",X"E2",X"0C",X"8E",X"2F",X"66",X"BD",X"2E",
		X"44",X"C6",X"FF",X"86",X"86",X"BD",X"E2",X"0C",X"8E",X"2F",X"8B",X"BD",X"2E",X"44",X"C6",X"FF",
		X"86",X"7F",X"BD",X"E2",X"0C",X"8E",X"2F",X"95",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"87",X"BD",
		X"E2",X"0C",X"8E",X"57",X"9B",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"88",X"BD",X"E2",X"0C",X"8E",
		X"53",X"9B",X"BD",X"2E",X"44",X"86",X"7E",X"BD",X"E2",X"0C",X"8E",X"4F",X"9B",X"BD",X"2E",X"44",
		X"86",X"89",X"BD",X"E2",X"0C",X"8E",X"4B",X"9B",X"BD",X"2E",X"44",X"86",X"76",X"BD",X"E2",X"0C",
		X"8E",X"47",X"9B",X"BD",X"2E",X"44",X"86",X"88",X"BD",X"E2",X"0C",X"8E",X"43",X"9B",X"BD",X"2E",
		X"44",X"86",X"84",X"BD",X"E2",X"0C",X"8E",X"3B",X"9B",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"8A",
		X"BD",X"E2",X"0C",X"8E",X"33",X"9B",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"8B",X"BD",X"E2",X"0C",
		X"8E",X"2F",X"9B",X"BD",X"2E",X"44",X"86",X"85",X"BD",X"E2",X"0C",X"8E",X"2B",X"9B",X"BD",X"2E",
		X"44",X"86",X"8C",X"BD",X"E2",X"0C",X"8E",X"27",X"9B",X"BD",X"2E",X"44",X"86",X"7F",X"BD",X"E2",
		X"0C",X"8E",X"23",X"9B",X"BD",X"2E",X"44",X"86",X"82",X"BD",X"E2",X"0C",X"35",X"36",X"EC",X"3E",
		X"DD",X"42",X"39",X"39",X"34",X"06",X"AE",X"98",X"1C",X"EE",X"04",X"A6",X"C8",X"21",X"33",X"86",
		X"AE",X"0A",X"EC",X"0E",X"A3",X"42",X"ED",X"0E",X"EC",X"0C",X"A3",X"44",X"ED",X"0C",X"35",X"86",
		X"34",X"46",X"AE",X"98",X"1C",X"EE",X"04",X"A6",X"C8",X"21",X"33",X"86",X"AE",X"0A",X"EC",X"0E",
		X"E3",X"42",X"ED",X"0E",X"EC",X"0C",X"E3",X"44",X"ED",X"0C",X"35",X"C6",X"34",X"76",X"EE",X"88",
		X"12",X"10",X"AE",X"98",X"1C",X"10",X"9C",X"78",X"26",X"07",X"86",X"30",X"97",X"00",X"7E",X"6F",
		X"78",X"E6",X"2C",X"54",X"54",X"54",X"54",X"26",X"01",X"5C",X"4F",X"C3",X"4E",X"28",X"DD",X"00",
		X"A6",X"9F",X"98",X"00",X"44",X"44",X"97",X"00",X"A6",X"C8",X"21",X"EE",X"98",X"1C",X"33",X"C6",
		X"EC",X"C4",X"26",X"11",X"EC",X"88",X"1C",X"BD",X"46",X"DB",X"6F",X"DF",X"08",X"A1",X"6D",X"ED",
		X"04",X"AE",X"1E",X"AF",X"C4",X"A6",X"46",X"81",X"60",X"2C",X"04",X"9B",X"00",X"A7",X"46",X"35",
		X"76",X"39",X"30",X"A4",X"BD",X"6C",X"79",X"4F",X"5F",X"ED",X"42",X"ED",X"44",X"7E",X"46",X"2B",
		X"34",X"06",X"EC",X"0A",X"27",X"12",X"34",X"10",X"AE",X"0A",X"CC",X"45",X"47",X"ED",X"88",X"1A",
		X"CC",X"4D",X"4F",X"ED",X"88",X"12",X"35",X"10",X"CC",X"4D",X"4F",X"ED",X"04",X"DC",X"78",X"ED",
		X"88",X"11",X"86",X"06",X"A7",X"88",X"1D",X"86",X"FF",X"A7",X"88",X"13",X"35",X"06",X"39",X"34",
		X"20",X"BD",X"70",X"8D",X"27",X"7A",X"BD",X"70",X"9B",X"35",X"20",X"CC",X"6F",X"F5",X"ED",X"22",
		X"EC",X"3E",X"DD",X"42",X"39",X"34",X"20",X"BD",X"70",X"8D",X"27",X"64",X"BD",X"70",X"BF",X"35",
		X"20",X"CC",X"70",X"0B",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"34",X"20",X"BD",X"70",X"8D",
		X"27",X"4E",X"BD",X"71",X"1E",X"BD",X"70",X"DE",X"EC",X"88",X"1C",X"10",X"93",X"78",X"27",X"1C",
		X"A6",X"46",X"80",X"02",X"A7",X"46",X"81",X"60",X"2D",X"23",X"BD",X"70",X"74",X"4F",X"5F",X"ED",
		X"C4",X"6F",X"46",X"ED",X"42",X"ED",X"44",X"35",X"20",X"7E",X"47",X"55",X"A6",X"46",X"80",X"04",
		X"28",X"01",X"4F",X"A7",X"46",X"81",X"60",X"2D",X"04",X"86",X"60",X"A7",X"46",X"A6",X"46",X"2A",
		X"95",X"6F",X"46",X"4F",X"5F",X"ED",X"C4",X"ED",X"42",X"ED",X"44",X"35",X"20",X"7E",X"47",X"55",
		X"A6",X"46",X"80",X"02",X"A7",X"46",X"2B",X"E9",X"35",X"20",X"CC",X"6F",X"DF",X"ED",X"22",X"EC",
		X"3E",X"DD",X"42",X"39",X"34",X"56",X"BD",X"38",X"91",X"4D",X"B3",X"CC",X"00",X"05",X"BD",X"3B",
		X"2A",X"EE",X"88",X"12",X"AE",X"98",X"1C",X"AD",X"D8",X"07",X"35",X"56",X"39",X"AE",X"B8",X"04",
		X"10",X"AE",X"04",X"A6",X"A8",X"21",X"33",X"86",X"AE",X"0A",X"39",X"E6",X"46",X"4F",X"58",X"49",
		X"58",X"49",X"34",X"06",X"BD",X"70",X"F3",X"BD",X"71",X"0A",X"ED",X"42",X"E3",X"0E",X"ED",X"0E",
		X"35",X"06",X"BD",X"70",X"F3",X"BD",X"71",X"0A",X"ED",X"44",X"E3",X"0C",X"ED",X"0C",X"39",X"EC",
		X"42",X"43",X"53",X"C3",X"00",X"01",X"ED",X"42",X"E3",X"42",X"E3",X"0E",X"ED",X"0E",X"EC",X"44",
		X"43",X"53",X"C3",X"00",X"01",X"ED",X"44",X"E3",X"44",X"E3",X"0C",X"ED",X"0C",X"39",X"EC",X"0E",
		X"A3",X"42",X"ED",X"0E",X"6F",X"42",X"6F",X"43",X"EC",X"0C",X"A3",X"44",X"ED",X"0C",X"6F",X"44",
		X"6F",X"45",X"39",X"34",X"02",X"86",X"00",X"BD",X"48",X"02",X"4C",X"2B",X"05",X"35",X"02",X"7E",
		X"71",X"09",X"35",X"02",X"43",X"53",X"C3",X"00",X"01",X"39",X"34",X"02",X"86",X"00",X"BD",X"48",
		X"02",X"4C",X"2B",X"05",X"35",X"02",X"7E",X"71",X"1D",X"35",X"02",X"47",X"56",X"39",X"34",X"36",
		X"CC",X"4C",X"EF",X"10",X"A3",X"88",X"12",X"27",X"5E",X"A6",X"46",X"80",X"10",X"23",X"58",X"34",
		X"02",X"86",X"00",X"BD",X"48",X"02",X"A1",X"E0",X"22",X"4D",X"34",X"10",X"10",X"AE",X"98",X"1C",
		X"A6",X"2C",X"80",X"08",X"24",X"01",X"4F",X"A7",X"2C",X"EC",X"28",X"C3",X"01",X"01",X"10",X"8E",
		X"4D",X"2D",X"AD",X"B8",X"05",X"35",X"20",X"AE",X"0A",X"27",X"24",X"EC",X"2E",X"A3",X"42",X"ED",
		X"0E",X"86",X"00",X"BD",X"48",X"02",X"1F",X"89",X"1D",X"E3",X"0E",X"ED",X"0E",X"EC",X"2C",X"A3",
		X"44",X"ED",X"0C",X"86",X"02",X"BD",X"48",X"02",X"1F",X"89",X"1D",X"E3",X"0C",X"ED",X"0C",X"A6",
		X"46",X"44",X"A7",X"46",X"7E",X"71",X"8A",X"BD",X"E1",X"95",X"35",X"36",X"39",X"BD",X"72",X"35",
		X"39",X"BD",X"72",X"3C",X"39",X"34",X"46",X"EC",X"1E",X"ED",X"88",X"11",X"EE",X"0A",X"27",X"08",
		X"EC",X"4E",X"DD",X"00",X"EC",X"4C",X"DD",X"02",X"EE",X"08",X"BD",X"72",X"35",X"1F",X"30",X"C3",
		X"01",X"01",X"CE",X"4D",X"2D",X"AD",X"D8",X"05",X"EE",X"0A",X"27",X"08",X"DC",X"00",X"ED",X"4E",
		X"DC",X"02",X"ED",X"4C",X"35",X"46",X"39",X"BD",X"72",X"21",X"BD",X"73",X"32",X"39",X"BD",X"72",
		X"21",X"BD",X"73",X"32",X"39",X"BD",X"72",X"21",X"BD",X"73",X"32",X"39",X"BD",X"72",X"21",X"BD",
		X"73",X"32",X"39",X"34",X"46",X"EE",X"98",X"0F",X"CC",X"47",X"55",X"ED",X"42",X"BD",X"72",X"21",
		X"BD",X"72",X"B0",X"35",X"46",X"39",X"34",X"46",X"EE",X"98",X"0F",X"CC",X"47",X"55",X"ED",X"42",
		X"BD",X"72",X"B0",X"35",X"46",X"39",X"34",X"46",X"EE",X"98",X"0F",X"CC",X"47",X"55",X"ED",X"42",
		X"BD",X"72",X"B0",X"7A",X"A1",X"B8",X"35",X"46",X"39",X"BD",X"72",X"B0",X"39",X"BD",X"73",X"32",
		X"39",X"34",X"36",X"10",X"AE",X"04",X"A6",X"A8",X"21",X"10",X"AE",X"96",X"27",X"05",X"CC",X"47",
		X"55",X"ED",X"22",X"35",X"B6",X"34",X"66",X"86",X"00",X"7E",X"72",X"40",X"34",X"66",X"86",X"01",
		X"34",X"02",X"EC",X"0A",X"27",X"0F",X"34",X"10",X"1F",X"01",X"BD",X"6C",X"61",X"CC",X"45",X"EA",
		X"ED",X"88",X"1A",X"35",X"10",X"10",X"AE",X"98",X"0D",X"CC",X"47",X"55",X"ED",X"22",X"10",X"AE",
		X"1E",X"10",X"AC",X"88",X"11",X"27",X"23",X"EE",X"98",X"11",X"A6",X"E4",X"31",X"C8",X"11",X"6A",
		X"A6",X"48",X"8B",X"13",X"10",X"AE",X"1E",X"10",X"AC",X"C6",X"27",X"07",X"EE",X"D6",X"86",X"16",
		X"BD",X"73",X"42",X"10",X"AE",X"88",X"16",X"10",X"AF",X"C6",X"A6",X"E4",X"48",X"CE",X"A1",X"A5",
		X"10",X"AE",X"1E",X"10",X"AC",X"C6",X"27",X"07",X"EE",X"D6",X"86",X"14",X"BD",X"73",X"42",X"10",
		X"AE",X"88",X"14",X"10",X"AF",X"C6",X"1F",X"12",X"BD",X"73",X"4D",X"32",X"61",X"35",X"66",X"39",
		X"34",X"66",X"EE",X"04",X"A6",X"C8",X"21",X"27",X"0C",X"34",X"10",X"10",X"AE",X"96",X"CC",X"47",
		X"55",X"ED",X"22",X"35",X"10",X"EC",X"0A",X"27",X"18",X"34",X"10",X"AE",X"0A",X"EC",X"88",X"12",
		X"10",X"83",X"4D",X"2D",X"27",X"06",X"BD",X"6C",X"61",X"7E",X"72",X"DF",X"BD",X"43",X"86",X"35",
		X"10",X"86",X"08",X"EE",X"98",X"13",X"BD",X"73",X"02",X"86",X"00",X"EE",X"98",X"15",X"BD",X"73",
		X"02",X"10",X"AE",X"98",X"0D",X"CC",X"47",X"55",X"ED",X"22",X"1F",X"12",X"BD",X"73",X"4D",X"35",
		X"66",X"39",X"34",X"02",X"27",X"29",X"A6",X"E4",X"A7",X"C8",X"1D",X"CC",X"FF",X"FF",X"ED",X"C8",
		X"18",X"86",X"01",X"A7",X"C8",X"1C",X"86",X"01",X"A7",X"C8",X"13",X"EC",X"5E",X"ED",X"C8",X"11",
		X"10",X"AE",X"C8",X"16",X"CC",X"00",X"00",X"ED",X"C8",X"16",X"EE",X"A4",X"7E",X"73",X"04",X"35",
		X"02",X"39",X"34",X"16",X"CC",X"47",X"4D",X"ED",X"02",X"AE",X"0A",X"27",X"03",X"BD",X"6C",X"61",
		X"35",X"96",X"10",X"AC",X"C6",X"27",X"05",X"EE",X"D6",X"7E",X"73",X"42",X"39",X"34",X"06",X"CC",
		X"47",X"4D",X"ED",X"22",X"35",X"86",X"34",X"76",X"10",X"8E",X"FF",X"FF",X"7E",X"73",X"65",X"34",
		X"76",X"10",X"8E",X"00",X"00",X"BD",X"3E",X"E1",X"8C",X"99",X"00",X"26",X"05",X"BD",X"7C",X"6A",
		X"20",X"0C",X"EC",X"88",X"12",X"10",X"83",X"4C",X"D0",X"26",X"03",X"BD",X"7C",X"67",X"CC",X"4D",
		X"8D",X"ED",X"88",X"12",X"33",X"84",X"10",X"8C",X"00",X"00",X"27",X"0B",X"BD",X"46",X"DB",X"73",
		X"B9",X"07",X"A1",X"74",X"7E",X"73",X"AB",X"BD",X"46",X"DB",X"73",X"B9",X"07",X"A1",X"5F",X"CC",
		X"2D",X"6F",X"ED",X"C8",X"16",X"CC",X"43",X"B8",X"ED",X"C8",X"18",X"EF",X"04",X"6F",X"06",X"6A",
		X"06",X"AE",X"1E",X"AF",X"C8",X"1C",X"35",X"76",X"39",X"CC",X"73",X"C3",X"ED",X"22",X"EC",X"3E",
		X"DD",X"42",X"39",X"8E",X"A1",X"6D",X"CC",X"73",X"CC",X"7E",X"46",X"AA",X"34",X"36",X"AE",X"24",
		X"A6",X"26",X"4C",X"81",X"04",X"2C",X"18",X"A7",X"26",X"C6",X"08",X"3D",X"C3",X"29",X"6C",X"ED",
		X"88",X"16",X"CC",X"43",X"B8",X"ED",X"88",X"18",X"35",X"36",X"EC",X"3E",X"DD",X"42",X"39",X"8C",
		X"99",X"00",X"26",X"0F",X"CC",X"2D",X"6F",X"ED",X"88",X"16",X"CC",X"43",X"B8",X"ED",X"88",X"18",
		X"7E",X"74",X"06",X"BD",X"43",X"86",X"35",X"36",X"7E",X"47",X"55",X"BD",X"85",X"59",X"7F",X"A0",
		X"3E",X"BD",X"6C",X"7C",X"39",X"BD",X"82",X"F1",X"CE",X"A0",X"1B",X"6F",X"C4",X"33",X"43",X"11",
		X"83",X"A0",X"3C",X"2D",X"F6",X"8E",X"00",X"00",X"BF",X"A1",X"A5",X"BF",X"A1",X"A7",X"10",X"8E",
		X"80",X"80",X"4F",X"97",X"7F",X"BD",X"79",X"00",X"CE",X"4B",X"C3",X"AD",X"D8",X"05",X"86",X"FF",
		X"97",X"7F",X"CC",X"80",X"80",X"CE",X"4C",X"EF",X"AD",X"D8",X"05",X"BD",X"46",X"BB",X"7A",X"3C",
		X"A1",X"97",X"BD",X"46",X"BB",X"78",X"EC",X"A1",X"9E",X"BD",X"46",X"BB",X"79",X"BB",X"A1",X"89",
		X"B6",X"A0",X"3E",X"27",X"04",X"84",X"03",X"27",X"07",X"BD",X"46",X"BB",X"79",X"65",X"A1",X"97",
		X"12",X"86",X"00",X"CE",X"4D",X"4F",X"97",X"00",X"0A",X"00",X"2B",X"06",X"AD",X"D8",X"05",X"7E",
		X"74",X"78",X"39",X"BD",X"3F",X"B1",X"4C",X"B1",X"BD",X"75",X"74",X"39",X"BD",X"3F",X"B1",X"4C",
		X"D0",X"BD",X"6C",X"6A",X"39",X"BD",X"3F",X"B1",X"4D",X"4F",X"BD",X"75",X"74",X"BD",X"6C",X"64",
		X"39",X"BD",X"3F",X"B1",X"4B",X"E5",X"BD",X"76",X"35",X"39",X"BD",X"3F",X"B1",X"4C",X"07",X"BD",
		X"76",X"35",X"39",X"BD",X"3F",X"B1",X"4C",X"29",X"BD",X"76",X"35",X"39",X"BD",X"3F",X"B1",X"4C",
		X"4B",X"BD",X"76",X"35",X"39",X"34",X"40",X"BD",X"3F",X"B1",X"4C",X"6D",X"34",X"10",X"BD",X"76",
		X"35",X"BD",X"6C",X"67",X"BD",X"46",X"DB",X"78",X"99",X"08",X"A1",X"89",X"EE",X"E4",X"EC",X"5E",
		X"ED",X"04",X"EC",X"1E",X"ED",X"4F",X"35",X"50",X"39",X"34",X"40",X"BD",X"3F",X"B1",X"4D",X"2D",
		X"34",X"10",X"BD",X"6C",X"67",X"BD",X"46",X"DB",X"77",X"EC",X"07",X"A1",X"89",X"EE",X"E4",X"EC",
		X"5E",X"ED",X"04",X"EC",X"1E",X"ED",X"4F",X"6F",X"06",X"35",X"50",X"39",X"34",X"40",X"BD",X"3F",
		X"B1",X"4C",X"8F",X"34",X"10",X"86",X"00",X"BD",X"48",X"02",X"A7",X"0C",X"BD",X"6C",X"67",X"BD",
		X"46",X"DB",X"6A",X"71",X"08",X"A1",X"74",X"EE",X"E4",X"EC",X"5E",X"ED",X"04",X"EC",X"1E",X"ED",
		X"4F",X"35",X"50",X"39",X"BD",X"3F",X"B1",X"4C",X"EF",X"86",X"00",X"BD",X"48",X"02",X"84",X"F0",
		X"8A",X"0C",X"A7",X"0C",X"BD",X"76",X"35",X"BD",X"6C",X"67",X"EC",X"1E",X"DD",X"78",X"BD",X"46",
		X"BB",X"75",X"56",X"A1",X"97",X"39",X"8E",X"A1",X"74",X"CC",X"6B",X"68",X"7E",X"46",X"AA",X"34",
		X"76",X"AE",X"9F",X"50",X"35",X"0D",X"96",X"26",X"05",X"BD",X"6C",X"67",X"20",X"03",X"BD",X"6C",
		X"6A",X"35",X"76",X"39",X"34",X"06",X"FC",X"A1",X"A5",X"ED",X"88",X"14",X"4F",X"A7",X"88",X"13",
		X"A7",X"88",X"1C",X"CC",X"FF",X"FF",X"ED",X"88",X"18",X"CC",X"00",X"00",X"ED",X"88",X"16",X"86",
		X"00",X"A7",X"88",X"1D",X"86",X"00",X"BD",X"48",X"02",X"A7",X"0C",X"EC",X"1E",X"ED",X"88",X"11",
		X"FD",X"A1",X"A5",X"BD",X"46",X"DB",X"61",X"6B",X"08",X"A1",X"74",X"ED",X"04",X"EC",X"1E",X"AE",
		X"98",X"04",X"ED",X"0D",X"35",X"86",X"34",X"06",X"FC",X"A1",X"A7",X"ED",X"88",X"14",X"4F",X"A7",
		X"88",X"13",X"A7",X"88",X"1C",X"CC",X"FF",X"FF",X"ED",X"88",X"18",X"CC",X"00",X"00",X"ED",X"88",
		X"16",X"86",X"00",X"A7",X"88",X"1D",X"86",X"00",X"BD",X"48",X"02",X"34",X"20",X"31",X"84",X"BD",
		X"6A",X"3C",X"35",X"20",X"A7",X"0C",X"EC",X"1E",X"ED",X"88",X"11",X"FD",X"A1",X"A7",X"BD",X"46",
		X"DB",X"66",X"12",X"08",X"A1",X"74",X"ED",X"04",X"EC",X"1E",X"AE",X"98",X"04",X"ED",X"0D",X"35",
		X"06",X"39",X"34",X"46",X"CC",X"00",X"00",X"ED",X"88",X"13",X"ED",X"88",X"15",X"4F",X"5F",X"EE",
		X"04",X"11",X"83",X"4D",X"2D",X"26",X"05",X"0D",X"96",X"26",X"01",X"5C",X"ED",X"88",X"11",X"EC",
		X"1E",X"BD",X"46",X"DB",X"76",X"4F",X"08",X"A1",X"5F",X"ED",X"04",X"EC",X"1E",X"AE",X"98",X"04",
		X"ED",X"0D",X"35",X"46",X"39",X"34",X"56",X"EE",X"04",X"A6",X"49",X"A7",X"0C",X"A6",X"C8",X"21",
		X"33",X"86",X"4F",X"5F",X"ED",X"C1",X"ED",X"C1",X"ED",X"C1",X"A7",X"C4",X"35",X"56",X"39",X"7F",
		X"A1",X"BE",X"7A",X"A1",X"BE",X"7E",X"76",X"75",X"7F",X"A1",X"BE",X"CC",X"A1",X"38",X"10",X"A3",
		X"24",X"26",X"09",X"8E",X"A1",X"89",X"CC",X"76",X"75",X"7E",X"46",X"AA",X"8E",X"A1",X"97",X"CC",
		X"76",X"75",X"7E",X"46",X"AA",X"34",X"20",X"10",X"AE",X"B8",X"04",X"AE",X"24",X"A6",X"88",X"1D",
		X"97",X"00",X"86",X"00",X"97",X"01",X"9B",X"00",X"97",X"02",X"8E",X"7A",X"48",X"E6",X"86",X"96",
		X"01",X"30",X"A8",X"11",X"E1",X"86",X"22",X"0E",X"96",X"01",X"27",X"03",X"7E",X"77",X"C5",X"86",
		X"01",X"97",X"01",X"7E",X"76",X"86",X"E6",X"86",X"86",X"06",X"3D",X"D7",X"03",X"96",X"02",X"8E",
		X"7A",X"5C",X"E6",X"86",X"D0",X"03",X"D7",X"04",X"CB",X"40",X"D7",X"05",X"86",X"01",X"97",X"06",
		X"4F",X"5F",X"DD",X"07",X"96",X"01",X"48",X"8E",X"A1",X"A5",X"AE",X"86",X"7E",X"76",X"D2",X"AE",
		X"88",X"14",X"8C",X"00",X"00",X"27",X"66",X"AE",X"84",X"EC",X"88",X"11",X"10",X"A3",X"3E",X"27",
		X"EE",X"96",X"05",X"A1",X"88",X"13",X"23",X"E7",X"86",X"FF",X"A1",X"88",X"13",X"27",X"E0",X"A6",
		X"08",X"A1",X"28",X"2D",X"05",X"A0",X"28",X"7E",X"76",X"FE",X"A6",X"28",X"A0",X"08",X"E6",X"09",
		X"E1",X"29",X"2D",X"05",X"E0",X"29",X"7E",X"77",X"0D",X"E6",X"29",X"E0",X"09",X"DD",X"0B",X"BD",
		X"77",X"D4",X"97",X"09",X"9B",X"04",X"97",X"0A",X"EC",X"88",X"18",X"BD",X"77",X"D4",X"AB",X"88",
		X"13",X"97",X"0F",X"96",X"0A",X"91",X"0F",X"23",X"A6",X"91",X"06",X"23",X"A2",X"97",X"06",X"EC",
		X"1E",X"DD",X"07",X"DC",X"0B",X"DD",X"0D",X"96",X"09",X"81",X"F8",X"23",X"92",X"96",X"06",X"81",
		X"01",X"10",X"23",X"FF",X"53",X"AE",X"9F",X"98",X"07",X"EE",X"98",X"11",X"11",X"A3",X"98",X"FE",
		X"27",X"3C",X"96",X"01",X"8B",X"11",X"6A",X"C6",X"2A",X"01",X"3F",X"96",X"01",X"48",X"8B",X"13",
		X"EE",X"C6",X"11",X"A3",X"1E",X"26",X"0D",X"EE",X"98",X"11",X"33",X"C6",X"EC",X"88",X"16",X"ED",
		X"C4",X"7E",X"77",X"8E",X"EC",X"1E",X"EE",X"C4",X"10",X"A3",X"C8",X"16",X"27",X"0A",X"EE",X"D8",
		X"16",X"11",X"83",X"00",X"00",X"26",X"F1",X"3F",X"EC",X"88",X"16",X"ED",X"C8",X"16",X"96",X"01",
		X"8B",X"11",X"6C",X"A6",X"96",X"01",X"48",X"33",X"A8",X"13",X"33",X"C6",X"EC",X"C4",X"34",X"06",
		X"EC",X"1E",X"ED",X"C4",X"96",X"04",X"A7",X"88",X"13",X"EC",X"3E",X"ED",X"88",X"11",X"DC",X"0D",
		X"ED",X"88",X"18",X"35",X"06",X"ED",X"88",X"16",X"CE",X"7A",X"52",X"96",X"02",X"A6",X"C6",X"A7",
		X"88",X"1D",X"7E",X"76",X"98",X"35",X"20",X"B6",X"A1",X"BE",X"27",X"03",X"7E",X"76",X"58",X"EC",
		X"3E",X"DD",X"42",X"39",X"43",X"53",X"34",X"04",X"1F",X"89",X"3D",X"44",X"34",X"02",X"A6",X"61",
		X"E6",X"61",X"3D",X"44",X"AB",X"E4",X"32",X"62",X"C6",X"40",X"3D",X"39",X"6C",X"26",X"28",X"02",
		X"6A",X"26",X"A6",X"26",X"AE",X"B8",X"04",X"EE",X"0A",X"26",X"0A",X"81",X"10",X"25",X"0B",X"BD",
		X"6C",X"70",X"7E",X"78",X"2D",X"6F",X"26",X"7E",X"78",X"3D",X"A6",X"88",X"11",X"27",X"1E",X"96",
		X"2E",X"81",X"60",X"22",X"18",X"EE",X"98",X"13",X"86",X"0C",X"A1",X"C8",X"18",X"25",X"09",X"A1",
		X"C8",X"19",X"25",X"04",X"EC",X"4A",X"27",X"0A",X"EE",X"D8",X"16",X"26",X"EB",X"EC",X"3E",X"DD",
		X"42",X"39",X"BD",X"6C",X"70",X"1F",X"31",X"BD",X"6C",X"64",X"7E",X"78",X"2D",X"8E",X"A1",X"74",
		X"BD",X"46",X"A8",X"8D",X"41",X"96",X"2E",X"2B",X"05",X"EC",X"3E",X"DD",X"42",X"39",X"86",X"00",
		X"BD",X"48",X"08",X"8E",X"A1",X"5F",X"BD",X"46",X"A8",X"8D",X"2B",X"CC",X"26",X"B1",X"ED",X"C8",
		X"16",X"CC",X"43",X"B8",X"ED",X"C8",X"18",X"BD",X"38",X"91",X"4D",X"F7",X"CC",X"78",X"76",X"ED",
		X"22",X"EC",X"3E",X"DD",X"42",X"39",X"8D",X"0E",X"CC",X"26",X"A1",X"ED",X"C8",X"16",X"CC",X"43",
		X"B8",X"ED",X"C8",X"18",X"20",X"B7",X"AE",X"B8",X"04",X"EE",X"0A",X"27",X"01",X"39",X"32",X"62",
		X"8E",X"A1",X"89",X"CC",X"77",X"EC",X"7E",X"46",X"AA",X"AE",X"B8",X"04",X"EE",X"0A",X"26",X"3A",
		X"A6",X"88",X"11",X"27",X"35",X"A6",X"88",X"12",X"27",X"30",X"86",X"00",X"BD",X"48",X"02",X"81",
		X"B0",X"22",X"27",X"EE",X"98",X"15",X"86",X"20",X"A1",X"C8",X"18",X"25",X"1D",X"A1",X"C8",X"19",
		X"25",X"18",X"EE",X"98",X"13",X"86",X"20",X"A1",X"C8",X"18",X"25",X"09",X"A1",X"C8",X"19",X"25",
		X"04",X"EC",X"4A",X"27",X"0A",X"EE",X"D8",X"16",X"26",X"EB",X"EC",X"3E",X"DD",X"42",X"39",X"EC",
		X"48",X"1F",X"31",X"BD",X"6C",X"73",X"BD",X"74",X"95",X"7E",X"78",X"DA",X"34",X"20",X"10",X"8E",
		X"80",X"80",X"86",X"FF",X"97",X"7F",X"BD",X"79",X"00",X"35",X"20",X"EC",X"3E",X"DD",X"42",X"39",
		X"34",X"56",X"96",X"7F",X"27",X"25",X"4F",X"8E",X"A0",X"1B",X"E6",X"01",X"E0",X"84",X"23",X"07",
		X"34",X"04",X"AB",X"E0",X"24",X"01",X"3F",X"30",X"03",X"8C",X"A0",X"3C",X"25",X"EC",X"4D",X"27",
		X"41",X"44",X"44",X"44",X"27",X"05",X"8E",X"4E",X"28",X"A6",X"86",X"97",X"00",X"8E",X"7A",X"A8",
		X"CE",X"A0",X"1B",X"A6",X"41",X"A0",X"C4",X"23",X"20",X"D6",X"00",X"27",X"01",X"3D",X"4D",X"27",
		X"18",X"34",X"12",X"DC",X"73",X"10",X"83",X"06",X"00",X"2D",X"0C",X"AE",X"F8",X"01",X"1F",X"20",
		X"AD",X"98",X"05",X"6A",X"E4",X"26",X"EC",X"35",X"12",X"33",X"43",X"30",X"02",X"8C",X"7A",X"B6",
		X"26",X"D1",X"35",X"56",X"39",X"B6",X"A0",X"28",X"B1",X"00",X"20",X"2D",X"0B",X"86",X"02",X"B7",
		X"A0",X"28",X"B7",X"A0",X"25",X"7E",X"79",X"B6",X"86",X"00",X"BD",X"48",X"02",X"81",X"10",X"22",
		X"35",X"B6",X"00",X"20",X"B7",X"A0",X"28",X"B7",X"A0",X"25",X"86",X"20",X"BD",X"55",X"93",X"8E",
		X"7A",X"00",X"BD",X"55",X"83",X"C6",X"FF",X"86",X"60",X"BD",X"E2",X"0C",X"86",X"8D",X"BD",X"E2",
		X"0C",X"8E",X"76",X"00",X"BD",X"55",X"83",X"86",X"8E",X"BD",X"E2",X"0C",X"86",X"64",X"BD",X"E2",
		X"0C",X"BD",X"38",X"91",X"4D",X"E6",X"EC",X"3E",X"DD",X"42",X"39",X"34",X"06",X"FC",X"A0",X"16",
		X"10",X"83",X"4F",X"E2",X"27",X"16",X"0D",X"94",X"27",X"1E",X"86",X"02",X"BD",X"48",X"02",X"81",
		X"40",X"12",X"12",X"12",X"22",X"12",X"BD",X"5D",X"7B",X"7E",X"79",X"E8",X"86",X"02",X"BD",X"48",
		X"02",X"81",X"38",X"22",X"03",X"BD",X"6C",X"80",X"35",X"06",X"EC",X"3E",X"DD",X"42",X"39",X"34",
		X"02",X"86",X"00",X"BD",X"48",X"02",X"84",X"7F",X"BB",X"A1",X"BF",X"B7",X"A1",X"BF",X"81",X"28",
		X"22",X"07",X"BD",X"53",X"6C",X"03",X"7E",X"7A",X"39",X"81",X"50",X"22",X"07",X"BD",X"53",X"6C",
		X"04",X"7E",X"7A",X"39",X"81",X"78",X"22",X"07",X"BD",X"53",X"6C",X"05",X"7E",X"7A",X"39",X"81",
		X"A0",X"22",X"07",X"BD",X"53",X"6C",X"06",X"7E",X"7A",X"39",X"81",X"C8",X"22",X"07",X"BD",X"53",
		X"6C",X"07",X"7E",X"7A",X"39",X"BD",X"53",X"6C",X"08",X"35",X"02",X"39",X"86",X"01",X"BD",X"48",
		X"3E",X"A0",X"3F",X"EC",X"3E",X"DD",X"42",X"39",X"03",X"01",X"03",X"09",X"00",X"06",X"01",X"01",
		X"03",X"01",X"02",X"04",X"02",X"02",X"00",X"06",X"04",X"08",X"04",X"08",X"58",X"58",X"48",X"5B",
		X"00",X"54",X"70",X"70",X"68",X"5B",X"AE",X"B8",X"1C",X"CC",X"47",X"55",X"ED",X"02",X"30",X"A4",
		X"BD",X"43",X"86",X"7E",X"34",X"AA",X"BD",X"73",X"56",X"CC",X"47",X"4D",X"ED",X"22",X"39",X"43",
		X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"4C",X"B1",X"4C",X"D0",X"4B",X"E5",X"4C",X"07",
		X"4C",X"29",X"4C",X"4B",X"4C",X"6D",X"4C",X"8F",X"4D",X"2D",X"4C",X"EF",X"4B",X"C3",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"02",X"00",X"00",X"02",X"00",X"00",X"02",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"A0",
		X"19",X"06",X"59",X"A4",X"10",X"59",X"A7",X"F8",X"7B",X"AA",X"10",X"7B",X"AD",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"06",X"08",X"01",X"01",X"01",X"01",X"03",X"00",X"00",X"01",X"01",X"A0",
		X"19",X"06",X"59",X"A4",X"10",X"59",X"A7",X"FF",X"7B",X"AA",X"FF",X"7B",X"AD",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"10",X"03",X"0A",X"02",X"02",X"02",X"02",X"00",X"00",X"01",X"01",X"A0",
		X"19",X"0A",X"59",X"A4",X"10",X"59",X"A7",X"F8",X"7B",X"AA",X"10",X"7B",X"AD",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"04",X"0A",X"0A",X"02",X"02",X"02",X"02",X"00",X"00",X"01",X"01",X"A0",
		X"19",X"04",X"59",X"A4",X"10",X"59",X"A7",X"F8",X"7B",X"AA",X"10",X"7B",X"AD",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"06",X"08",X"10",X"02",X"10",X"02",X"05",X"00",X"00",X"01",X"01",X"A0",
		X"19",X"06",X"59",X"A4",X"0A",X"59",X"A7",X"10",X"7B",X"AA",X"10",X"7B",X"AD",X"03",X"59",X"AA",
		X"7F",X"59",X"AD",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"04",X"00",
		X"00",X"04",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"01",X"00",X"A0",X"19",X"06",X"59",X"A4",X"01",X"59",X"A7",X"01",X"7B",X"AA",
		X"01",X"7B",X"AD",X"03",X"59",X"AA",X"7F",X"59",X"AD",X"00",X"A0",X"22",X"00",X"A0",X"28",X"00",
		X"34",X"76",X"4F",X"5F",X"FD",X"A0",X"19",X"FD",X"A0",X"3C",X"0D",X"96",X"27",X"06",X"8E",X"7B",
		X"74",X"7E",X"7B",X"EB",X"B6",X"A0",X"3E",X"26",X"06",X"8E",X"7A",X"BE",X"7E",X"7B",X"EB",X"84",
		X"03",X"C6",X"20",X"3D",X"C3",X"7A",X"F4",X"1F",X"01",X"CE",X"A0",X"1B",X"A6",X"80",X"5F",X"ED",
		X"41",X"33",X"43",X"11",X"83",X"A0",X"3C",X"25",X"F3",X"20",X"0C",X"CE",X"A0",X"1B",X"CC",X"A0",
		X"3C",X"FD",X"A1",X"C0",X"BD",X"7C",X"4D",X"CE",X"A0",X"3F",X"CC",X"A0",X"54",X"FD",X"A1",X"C0",
		X"BD",X"7C",X"4D",X"F1",X"A0",X"3E",X"24",X"1D",X"D7",X"00",X"86",X"06",X"34",X"10",X"8E",X"CC",
		X"06",X"BD",X"4A",X"70",X"35",X"10",X"3D",X"1F",X"98",X"BD",X"48",X"3E",X"A0",X"3F",X"D6",X"00",
		X"CB",X"04",X"7E",X"7C",X"03",X"34",X"10",X"8E",X"CC",X"06",X"BD",X"4A",X"5F",X"35",X"10",X"BD",
		X"48",X"3E",X"A0",X"3F",X"B6",X"A0",X"3E",X"26",X"04",X"86",X"99",X"20",X"07",X"8E",X"50",X"DB",
		X"84",X"03",X"A6",X"86",X"B7",X"A0",X"18",X"BD",X"33",X"B4",X"35",X"76",X"39",X"E6",X"80",X"E7",
		X"C0",X"11",X"B3",X"A1",X"C0",X"25",X"F6",X"39",X"12",X"12",X"12",X"BD",X"46",X"DB",X"7C",X"64",
		X"08",X"A1",X"5F",X"39",X"7E",X"80",X"5E",X"7E",X"7E",X"29",X"7E",X"FF",X"90",X"34",X"76",X"86",
		X"07",X"97",X"1E",X"DC",X"73",X"10",X"83",X"01",X"F4",X"2D",X"5B",X"1F",X"13",X"BD",X"46",X"DB",
		X"7C",X"D8",X"F6",X"A1",X"66",X"6F",X"05",X"31",X"06",X"EC",X"45",X"34",X"06",X"86",X"3C",X"34",
		X"02",X"CC",X"02",X"0F",X"BD",X"47",X"FA",X"8B",X"F9",X"34",X"02",X"CC",X"00",X"07",X"BD",X"47",
		X"FA",X"8B",X"FD",X"35",X"04",X"ED",X"22",X"27",X"E8",X"CC",X"00",X"04",X"BD",X"47",X"FA",X"48",
		X"34",X"02",X"CC",X"02",X"04",X"BD",X"47",X"FA",X"35",X"04",X"E3",X"61",X"ED",X"A4",X"31",X"24",
		X"6A",X"E4",X"26",X"CD",X"32",X"63",X"DC",X"73",X"10",X"83",X"00",X"EA",X"2D",X"08",X"BD",X"46",
		X"DB",X"7D",X"85",X"71",X"A1",X"66",X"35",X"F6",X"A6",X"24",X"4C",X"84",X"03",X"A7",X"24",X"48",
		X"8E",X"7D",X"55",X"AE",X"86",X"BF",X"CA",X"02",X"CC",X"02",X"03",X"88",X"04",X"C8",X"04",X"FD",
		X"CA",X"06",X"E6",X"25",X"57",X"5C",X"C1",X"04",X"2F",X"02",X"C6",X"04",X"86",X"0F",X"3D",X"34",
		X"04",X"30",X"26",X"A6",X"E4",X"81",X"1E",X"26",X"0E",X"A6",X"25",X"84",X"04",X"44",X"12",X"CE",
		X"7D",X"75",X"EE",X"C6",X"FF",X"CA",X"02",X"EC",X"84",X"27",X"27",X"FD",X"CA",X"04",X"7F",X"CA",
		X"01",X"86",X"12",X"B7",X"CA",X"00",X"A6",X"84",X"E3",X"02",X"81",X"72",X"22",X"10",X"C1",X"F0",
		X"22",X"0C",X"ED",X"84",X"FD",X"CA",X"04",X"86",X"0E",X"B7",X"CA",X"00",X"20",X"04",X"6F",X"84",
		X"6F",X"01",X"30",X"04",X"6A",X"E4",X"26",X"BB",X"32",X"61",X"6C",X"25",X"10",X"2B",X"CA",X"05",
		X"EC",X"3E",X"DD",X"42",X"39",X"7D",X"5D",X"7D",X"63",X"7D",X"69",X"7D",X"6F",X"00",X"00",X"0C",
		X"00",X"00",X"00",X"C0",X"C0",X"0F",X"00",X"C0",X"C0",X"0F",X"00",X"F6",X"F0",X"0F",X"00",X"60",
		X"60",X"0B",X"00",X"60",X"60",X"7D",X"79",X"7D",X"7F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"8E",X"99",X"00",X"AE",X"05",X"30",X"89",X"01",X"02",X"86",X"03",
		X"34",X"12",X"30",X"25",X"86",X"02",X"4A",X"C6",X"06",X"C0",X"03",X"34",X"06",X"E3",X"63",X"ED",
		X"84",X"CC",X"00",X"08",X"BD",X"47",X"FA",X"47",X"24",X"01",X"40",X"A7",X"02",X"CC",X"02",X"0C",
		X"BD",X"47",X"FA",X"47",X"24",X"01",X"40",X"A7",X"03",X"30",X"04",X"35",X"06",X"5D",X"2A",X"D9",
		X"4D",X"2A",X"D3",X"6A",X"E4",X"26",X"CD",X"32",X"63",X"86",X"18",X"A7",X"24",X"CC",X"7D",X"D7",
		X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"6A",X"24",X"2A",X"06",X"BD",X"32",X"0F",X"7E",X"47",
		X"55",X"CC",X"05",X"05",X"FD",X"CA",X"06",X"CC",X"7E",X"1C",X"FD",X"CA",X"02",X"A6",X"24",X"47",
		X"CE",X"7E",X"1D",X"A6",X"C6",X"97",X"25",X"8E",X"00",X"1B",X"33",X"25",X"EC",X"C4",X"E3",X"42",
		X"4D",X"2B",X"0E",X"C1",X"F0",X"22",X"0A",X"ED",X"C4",X"FD",X"CA",X"04",X"86",X"0E",X"B7",X"CA",
		X"00",X"33",X"44",X"30",X"1F",X"26",X"E5",X"EC",X"3E",X"DD",X"42",X"39",X"70",X"00",X"48",X"91",
		X"CA",X"84",X"46",X"07",X"17",X"67",X"AF",X"FF",X"FF",X"34",X"76",X"DC",X"73",X"10",X"83",X"00",
		X"64",X"2D",X"63",X"1F",X"13",X"BD",X"46",X"DB",X"7E",X"98",X"2E",X"A1",X"66",X"6F",X"05",X"86",
		X"06",X"A7",X"04",X"31",X"06",X"DC",X"46",X"E3",X"4C",X"58",X"49",X"34",X"02",X"DC",X"44",X"E3",
		X"4E",X"58",X"49",X"34",X"02",X"EC",X"45",X"34",X"06",X"86",X"0A",X"34",X"02",X"CC",X"02",X"0F",
		X"BD",X"47",X"FA",X"8B",X"F9",X"34",X"02",X"CC",X"00",X"07",X"BD",X"47",X"FA",X"8B",X"FD",X"35",
		X"04",X"AB",X"63",X"EB",X"64",X"ED",X"22",X"27",X"E4",X"CC",X"00",X"04",X"BD",X"47",X"FA",X"48",
		X"34",X"02",X"CC",X"02",X"04",X"BD",X"47",X"FA",X"35",X"04",X"E3",X"61",X"ED",X"A4",X"31",X"24",
		X"6A",X"E4",X"26",X"C9",X"32",X"65",X"35",X"F6",X"A6",X"24",X"4A",X"48",X"8E",X"7F",X"03",X"AE",
		X"86",X"BF",X"CA",X"02",X"CC",X"03",X"05",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"6C",X"25",
		X"E6",X"25",X"57",X"25",X"02",X"6A",X"24",X"86",X"0A",X"34",X"02",X"30",X"26",X"EC",X"84",X"27",
		X"2F",X"FD",X"CA",X"04",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",X"6D",X"24",X"27",X"20",
		X"A6",X"84",X"E3",X"02",X"81",X"71",X"22",X"14",X"C1",X"10",X"25",X"10",X"C1",X"F0",X"22",X"0C",
		X"ED",X"84",X"FD",X"CA",X"04",X"86",X"0E",X"B7",X"CA",X"00",X"20",X"04",X"6F",X"84",X"6F",X"01",
		X"30",X"04",X"6A",X"E4",X"26",X"C7",X"32",X"61",X"6D",X"24",X"10",X"27",X"C8",X"57",X"EC",X"3E",
		X"DD",X"42",X"39",X"7F",X"3C",X"7F",X"2D",X"7F",X"1E",X"7F",X"0F",X"7F",X"0F",X"7F",X"0F",X"0A",
		X"0A",X"00",X"AA",X"AA",X"A0",X"0A",X"FA",X"00",X"AA",X"AA",X"A0",X"0A",X"0A",X"00",X"0A",X"0A",
		X"00",X"A1",X"D1",X"A0",X"0D",X"DD",X"00",X"A1",X"D1",X"A0",X"0A",X"0A",X"00",X"00",X"00",X"00",
		X"0C",X"CC",X"00",X"0C",X"0C",X"00",X"0C",X"CC",X"00",X"00",X"00",X"00",X"0D",X"0D",X"00",X"D0",
		X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"D0",X"0D",X"0D",X"00",X"34",X"76",X"BD",X"53",X"6C",
		X"09",X"12",X"12",X"12",X"12",X"12",X"12",X"BD",X"32",X"7E",X"BD",X"46",X"DB",X"7F",X"DE",X"05",
		X"A1",X"6D",X"CC",X"00",X"08",X"BD",X"47",X"FA",X"8B",X"00",X"10",X"8E",X"7F",X"D6",X"E6",X"A6",
		X"E7",X"04",X"BD",X"46",X"DB",X"7F",X"97",X"05",X"A1",X"5F",X"86",X"5A",X"A7",X"04",X"BD",X"46",
		X"DB",X"7F",X"B3",X"05",X"A1",X"66",X"86",X"0E",X"A7",X"04",X"7D",X"A1",X"BA",X"27",X"03",X"7C",
		X"A0",X"54",X"BD",X"59",X"B0",X"35",X"F6",X"7D",X"A1",X"BC",X"26",X"09",X"A6",X"24",X"4A",X"10",
		X"27",X"C7",X"B2",X"A7",X"24",X"C6",X"3F",X"47",X"24",X"02",X"C6",X"07",X"D7",X"1E",X"EC",X"3E",
		X"DD",X"42",X"39",X"AE",X"9F",X"98",X"78",X"AE",X"0A",X"27",X"16",X"EC",X"05",X"34",X"06",X"C3",
		X"0A",X"12",X"ED",X"05",X"BD",X"7C",X"67",X"35",X"06",X"ED",X"05",X"6A",X"24",X"10",X"27",X"C7",
		X"84",X"EC",X"3E",X"DD",X"42",X"39",X"00",X"FF",X"DE",X"EF",X"22",X"11",X"CD",X"BC",X"7D",X"A1",
		X"BC",X"26",X"18",X"CC",X"50",X"02",X"FD",X"A0",X"16",X"FD",X"A0",X"14",X"BD",X"46",X"DB",X"80",
		X"13",X"05",X"A1",X"5F",X"86",X"0E",X"A7",X"04",X"7E",X"47",X"55",X"CE",X"D8",X"70",X"8E",X"03",
		X"12",X"E6",X"C0",X"27",X"05",X"53",X"EB",X"24",X"E7",X"5F",X"30",X"1F",X"26",X"F3",X"EC",X"3E",
		X"DD",X"42",X"39",X"6A",X"24",X"27",X"08",X"BD",X"3C",X"D9",X"EC",X"3E",X"DD",X"42",X"39",X"CC",
		X"4F",X"B2",X"FD",X"A0",X"14",X"BD",X"32",X"0F",X"BD",X"32",X"7E",X"7E",X"47",X"55",X"43",X"4F",
		X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"BD",X"8B",X"58",X"7F",X"A1",X"BD",X"39",X"8E",X"CC",
		X"0A",X"BD",X"4A",X"5F",X"10",X"27",X"00",X"AA",X"7C",X"A1",X"BD",X"86",X"33",X"97",X"80",X"BD",
		X"32",X"45",X"B6",X"BF",X"FF",X"34",X"22",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"8E",
		X"82",X"2E",X"10",X"8E",X"CD",X"32",X"7C",X"A1",X"DB",X"BD",X"82",X"6C",X"31",X"28",X"8E",X"82",
		X"6A",X"BD",X"82",X"B1",X"8E",X"82",X"8A",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"8F",X"BD",X"E2",
		X"03",X"86",X"90",X"BD",X"E2",X"03",X"30",X"88",X"D6",X"B6",X"BF",X"FF",X"84",X"FB",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"86",X"27",X"BD",X"E2",X"00",X"8E",X"76",X"59",X"BD",X"2E",X"44",X"C6",
		X"DD",X"86",X"91",X"BD",X"E2",X"03",X"B6",X"BF",X"FF",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",
		X"00",X"8E",X"70",X"00",X"10",X"8E",X"CD",X"32",X"7F",X"A1",X"DB",X"BD",X"81",X"F2",X"8E",X"41",
		X"50",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"92",X"BD",X"E2",X"03",X"86",X"93",X"BD",X"E2",X"03",
		X"8E",X"3B",X"00",X"10",X"8E",X"DC",X"94",X"BD",X"81",X"F2",X"35",X"22",X"B7",X"BF",X"FF",X"B7",
		X"C9",X"00",X"BD",X"46",X"DB",X"81",X"DB",X"06",X"A1",X"5F",X"CC",X"01",X"2C",X"ED",X"04",X"BD",
		X"34",X"19",X"34",X"20",X"86",X"33",X"97",X"80",X"BD",X"32",X"45",X"BD",X"33",X"8E",X"8E",X"56",
		X"65",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"6C",X"BD",X"E2",X"03",X"8E",X"54",X"99",X"BD",X"2E",
		X"44",X"C6",X"DD",X"86",X"94",X"BD",X"E2",X"0C",X"C6",X"CC",X"8E",X"CE",X"D6",X"10",X"8E",X"34",
		X"25",X"BD",X"82",X"D7",X"C6",X"33",X"31",X"3F",X"BD",X"82",X"D7",X"C6",X"CC",X"8E",X"CF",X"0C",
		X"10",X"8E",X"2C",X"25",X"BD",X"82",X"D7",X"C6",X"22",X"31",X"3F",X"BD",X"82",X"D7",X"CC",X"01",
		X"C0",X"FD",X"A1",X"DC",X"35",X"20",X"8E",X"A1",X"5F",X"BD",X"46",X"A8",X"34",X"20",X"FC",X"A1",
		X"DC",X"83",X"00",X"01",X"FD",X"A1",X"DC",X"26",X"06",X"7F",X"A1",X"BD",X"7E",X"2E",X"D4",X"10",
		X"83",X"01",X"00",X"10",X"24",X"00",X"1D",X"86",X"00",X"BD",X"48",X"08",X"81",X"8E",X"22",X"F7",
		X"1F",X"01",X"CC",X"02",X"0C",X"BD",X"47",X"FA",X"8B",X"00",X"CE",X"81",X"CF",X"E6",X"C6",X"86",
		X"6C",X"BD",X"E2",X"03",X"8E",X"4A",X"2C",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"95",X"BD",X"E2",
		X"0C",X"86",X"96",X"BD",X"E2",X"0C",X"86",X"97",X"BD",X"E2",X"0C",X"86",X"98",X"BD",X"E2",X"0C",
		X"86",X"99",X"BD",X"E2",X"0C",X"BD",X"33",X"8E",X"35",X"20",X"EC",X"3E",X"DD",X"42",X"39",X"11",
		X"22",X"33",X"44",X"55",X"66",X"99",X"AA",X"BB",X"CC",X"DD",X"FF",X"EC",X"24",X"83",X"00",X"01",
		X"ED",X"24",X"10",X"27",X"C5",X"6F",X"BD",X"33",X"8E",X"86",X"48",X"97",X"1E",X"EC",X"3E",X"DD",
		X"42",X"39",X"4F",X"34",X"02",X"6C",X"E4",X"A6",X"E4",X"5F",X"34",X"04",X"1F",X"89",X"80",X"0A",
		X"2B",X"04",X"6C",X"E4",X"20",X"F6",X"35",X"02",X"4D",X"26",X"02",X"86",X"0A",X"34",X"06",X"30",
		X"88",X"18",X"C6",X"63",X"BD",X"E2",X"09",X"A6",X"61",X"BD",X"E2",X"09",X"86",X"2B",X"BD",X"E2",
		X"09",X"C6",X"FF",X"10",X"BC",X"A1",X"C3",X"27",X"12",X"10",X"BC",X"A1",X"C5",X"27",X"0C",X"10",
		X"BC",X"A1",X"C7",X"27",X"06",X"10",X"BC",X"A1",X"C9",X"26",X"06",X"C6",X"47",X"D7",X"2C",X"C6",
		X"EE",X"F7",X"A1",X"DE",X"30",X"03",X"31",X"28",X"BD",X"82",X"B1",X"30",X"88",X"10",X"31",X"38",
		X"BD",X"82",X"6C",X"31",X"2E",X"35",X"06",X"5D",X"27",X"06",X"30",X"89",X"FC",X"C9",X"20",X"95",
		X"81",X"03",X"27",X"06",X"30",X"89",X"1B",X"10",X"20",X"8B",X"35",X"82",X"34",X"36",X"C6",X"04",
		X"1E",X"12",X"BD",X"4A",X"5F",X"26",X"10",X"7D",X"A1",X"DB",X"26",X"04",X"31",X"28",X"20",X"02",
		X"31",X"2E",X"5A",X"26",X"ED",X"20",X"28",X"81",X"0F",X"22",X"02",X"8A",X"F0",X"34",X"04",X"1E",
		X"12",X"7D",X"A1",X"DB",X"26",X"08",X"F6",X"A1",X"DE",X"BD",X"E2",X"0F",X"20",X"05",X"C6",X"11",
		X"BD",X"E2",X"06",X"35",X"04",X"5A",X"27",X"07",X"1E",X"12",X"BD",X"4A",X"5F",X"20",X"DE",X"35",
		X"B6",X"34",X"36",X"C6",X"03",X"1E",X"12",X"BD",X"4A",X"5F",X"1E",X"12",X"34",X"04",X"7D",X"A1",
		X"DB",X"26",X"08",X"F6",X"A1",X"DE",X"BD",X"E2",X"09",X"20",X"05",X"C6",X"11",X"BD",X"E2",X"00",
		X"35",X"04",X"5A",X"26",X"E0",X"35",X"B6",X"34",X"36",X"86",X"1B",X"34",X"02",X"BD",X"4A",X"5F",
		X"1E",X"12",X"E6",X"62",X"BD",X"E2",X"00",X"1E",X"12",X"6A",X"E4",X"26",X"F0",X"32",X"61",X"35",
		X"B6",X"BD",X"8E",X"55",X"0D",X"96",X"27",X"10",X"BD",X"46",X"DB",X"83",X"09",X"05",X"A1",X"6D",
		X"BD",X"46",X"DB",X"84",X"8A",X"05",X"A1",X"6D",X"39",X"BD",X"84",X"72",X"86",X"96",X"A7",X"24",
		X"CC",X"83",X"1A",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"6A",X"24",X"27",X"55",X"34",X"36",
		X"8E",X"6D",X"4C",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"9A",X"BD",X"E2",X"0C",X"86",X"9B",X"BD",
		X"E2",X"0C",X"86",X"9C",X"BD",X"E2",X"0C",X"86",X"64",X"BD",X"E2",X"0C",X"8E",X"69",X"20",X"BD",
		X"2E",X"44",X"C6",X"FF",X"86",X"9D",X"BD",X"E2",X"0C",X"86",X"9E",X"BD",X"E2",X"0C",X"86",X"9B",
		X"BD",X"E2",X"0C",X"86",X"79",X"BD",X"E2",X"0C",X"86",X"9F",X"BD",X"E2",X"0C",X"86",X"A0",X"BD",
		X"E2",X"0C",X"86",X"A1",X"BD",X"E2",X"0C",X"86",X"A2",X"BD",X"E2",X"0C",X"35",X"36",X"EC",X"3E",
		X"DD",X"42",X"39",X"BD",X"84",X"72",X"86",X"96",X"A7",X"24",X"CC",X"83",X"84",X"ED",X"22",X"EC",
		X"3E",X"DD",X"42",X"39",X"6A",X"24",X"27",X"5C",X"34",X"36",X"8E",X"6D",X"2A",X"BD",X"2E",X"44",
		X"C6",X"FF",X"86",X"A3",X"BD",X"E2",X"0C",X"86",X"A4",X"BD",X"E2",X"0C",X"86",X"A5",X"BD",X"E2",
		X"0C",X"86",X"A6",X"BD",X"E2",X"0C",X"86",X"6B",X"BD",X"E2",X"0C",X"86",X"A7",X"BD",X"E2",X"0C",
		X"C6",X"DD",X"86",X"6C",X"BD",X"E2",X"0C",X"8E",X"69",X"32",X"BD",X"2E",X"44",X"C6",X"FF",X"86",
		X"A8",X"BD",X"E2",X"0C",X"86",X"A2",X"BD",X"E2",X"0C",X"86",X"A9",X"BD",X"E2",X"0C",X"86",X"A6",
		X"BD",X"E2",X"0C",X"86",X"AA",X"BD",X"E2",X"0C",X"86",X"AB",X"BD",X"E2",X"0C",X"35",X"36",X"EC",
		X"3E",X"DD",X"42",X"39",X"BD",X"84",X"72",X"86",X"C3",X"A7",X"24",X"CC",X"83",X"F5",X"ED",X"22",
		X"EC",X"3E",X"DD",X"42",X"39",X"6A",X"24",X"27",X"73",X"34",X"36",X"8E",X"6D",X"27",X"BD",X"2E",
		X"44",X"C6",X"FF",X"86",X"AC",X"BD",X"E2",X"0C",X"86",X"6B",X"BD",X"E2",X"0C",X"C6",X"DD",X"86",
		X"6C",X"BD",X"E2",X"0C",X"8E",X"6D",X"70",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"6E",X"BD",X"E2",
		X"0C",X"86",X"AD",X"BD",X"E2",X"0C",X"86",X"69",X"BD",X"E2",X"0C",X"86",X"AE",X"BD",X"E2",X"0C",
		X"86",X"AF",X"BD",X"E2",X"0C",X"86",X"B0",X"BD",X"E2",X"0C",X"8E",X"69",X"7C",X"BD",X"2E",X"44",
		X"C6",X"FF",X"86",X"B1",X"BD",X"E2",X"0C",X"8E",X"65",X"5C",X"BD",X"2E",X"44",X"C6",X"FF",X"86",
		X"69",X"BD",X"E2",X"0C",X"86",X"B2",X"BD",X"E2",X"0C",X"86",X"B3",X"BD",X"E2",X"0C",X"C6",X"DD",
		X"86",X"B4",X"BD",X"E2",X"0C",X"35",X"36",X"EC",X"3E",X"DD",X"42",X"39",X"BD",X"84",X"72",X"7E",
		X"47",X"55",X"34",X"06",X"CC",X"0F",X"FB",X"FD",X"CA",X"06",X"CC",X"65",X"00",X"FD",X"CA",X"04",
		X"7F",X"CA",X"01",X"86",X"11",X"B7",X"CA",X"00",X"35",X"86",X"6F",X"24",X"CC",X"84",X"96",X"ED",
		X"22",X"EC",X"3E",X"DD",X"42",X"39",X"34",X"20",X"B6",X"BF",X"1B",X"A1",X"24",X"27",X"16",X"A7",
		X"24",X"CC",X"00",X"FB",X"FD",X"CA",X"06",X"CC",X"17",X"00",X"FD",X"CA",X"04",X"7F",X"CA",X"01",
		X"86",X"11",X"B7",X"CA",X"00",X"8E",X"CC",X"0A",X"BD",X"4A",X"5F",X"27",X"2B",X"8E",X"1C",X"3E",
		X"BD",X"2E",X"44",X"C6",X"22",X"86",X"B5",X"BD",X"E2",X"0C",X"86",X"B6",X"BD",X"E2",X"0C",X"86",
		X"B7",X"BD",X"E2",X"0C",X"86",X"79",X"BD",X"E2",X"0C",X"86",X"B8",X"BD",X"E2",X"0C",X"86",X"B9",
		X"BD",X"E2",X"0C",X"86",X"BA",X"BD",X"E2",X"0C",X"B6",X"BF",X"1B",X"27",X"49",X"4A",X"27",X"28",
		X"8E",X"18",X"52",X"BD",X"2E",X"44",X"C6",X"22",X"86",X"B5",X"BD",X"E2",X"0C",X"86",X"52",X"BD",
		X"E2",X"0C",X"86",X"B1",X"BD",X"E2",X"0C",X"86",X"53",X"BD",X"E2",X"0C",X"86",X"51",X"BD",X"E2",
		X"0C",X"86",X"BB",X"BD",X"E2",X"0C",X"20",X"3A",X"8E",X"18",X"5C",X"BD",X"2E",X"44",X"C6",X"22",
		X"86",X"B5",X"BD",X"E2",X"0C",X"86",X"52",X"BD",X"E2",X"0C",X"86",X"51",X"BD",X"E2",X"0C",X"86",
		X"BB",X"BD",X"E2",X"0C",X"20",X"1C",X"8E",X"18",X"5E",X"BD",X"2E",X"44",X"C6",X"22",X"86",X"BC",
		X"BD",X"E2",X"0C",X"86",X"BD",X"BD",X"E2",X"0C",X"86",X"79",X"BD",X"E2",X"0C",X"86",X"BE",X"BD",
		X"E2",X"0C",X"35",X"20",X"EC",X"3E",X"DD",X"42",X"39",X"12",X"12",X"12",X"7F",X"A0",X"54",X"39",
		X"0D",X"96",X"26",X"1C",X"8D",X"3C",X"35",X"20",X"BD",X"34",X"19",X"7D",X"A0",X"54",X"27",X"0E",
		X"BD",X"46",X"DB",X"85",X"83",X"0A",X"A1",X"5F",X"7F",X"A0",X"54",X"BD",X"6C",X"7C",X"34",X"20",
		X"7E",X"2F",X"FC",X"BD",X"46",X"BB",X"5C",X"06",X"A1",X"6D",X"AE",X"1E",X"AF",X"28",X"CC",X"00",
		X"78",X"BD",X"34",X"19",X"AE",X"B8",X"08",X"CC",X"47",X"55",X"ED",X"02",X"BD",X"32",X"0F",X"7E",
		X"47",X"55",X"34",X"70",X"BD",X"38",X"91",X"4D",X"EB",X"BD",X"53",X"6C",X"0A",X"BD",X"32",X"7E",
		X"96",X"8A",X"4A",X"26",X"03",X"BD",X"32",X"0F",X"BD",X"33",X"B4",X"7D",X"A0",X"54",X"27",X"2C",
		X"8E",X"4E",X"4E",X"BD",X"2E",X"44",X"C6",X"11",X"86",X"68",X"BD",X"E2",X"03",X"8E",X"40",X"2B",
		X"BD",X"2E",X"44",X"C6",X"11",X"86",X"69",X"BD",X"E2",X"03",X"86",X"6A",X"BD",X"E2",X"03",X"86",
		X"6B",X"BD",X"E2",X"03",X"86",X"6C",X"BD",X"E2",X"03",X"7E",X"86",X"72",X"8E",X"58",X"53",X"BD",
		X"2E",X"44",X"C6",X"99",X"86",X"69",X"BD",X"E2",X"0C",X"86",X"BF",X"BD",X"E2",X"0C",X"34",X"06",
		X"B6",X"A0",X"13",X"BD",X"87",X"29",X"35",X"06",X"30",X"04",X"86",X"A2",X"BD",X"E2",X"0C",X"8E",
		X"52",X"52",X"BD",X"2E",X"44",X"C6",X"99",X"86",X"6C",X"BD",X"E2",X"0C",X"86",X"C0",X"BD",X"E2",
		X"0C",X"34",X"06",X"FC",X"A0",X"14",X"83",X"4F",X"B2",X"47",X"56",X"47",X"56",X"34",X"04",X"FC",
		X"A0",X"16",X"10",X"83",X"4F",X"E2",X"26",X"02",X"6C",X"E4",X"A6",X"E4",X"BD",X"87",X"29",X"EC",
		X"61",X"30",X"04",X"86",X"C1",X"BD",X"E2",X"0C",X"35",X"02",X"B1",X"A0",X"13",X"2F",X"21",X"8E",
		X"48",X"3C",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"78",X"BD",X"E2",X"0C",X"86",X"9B",X"BD",X"E2",
		X"0C",X"86",X"79",X"BD",X"E2",X"0C",X"86",X"7A",X"BD",X"E2",X"0C",X"86",X"A2",X"BD",X"E2",X"0C",
		X"32",X"62",X"BD",X"87",X"45",X"B6",X"A0",X"3E",X"27",X"33",X"8E",X"20",X"44",X"BD",X"2E",X"44",
		X"C6",X"55",X"86",X"69",X"BD",X"E2",X"0C",X"86",X"BF",X"BD",X"E2",X"0C",X"86",X"C2",X"BD",X"E2",
		X"0C",X"B6",X"A0",X"3E",X"BD",X"87",X"29",X"30",X"04",X"C6",X"55",X"86",X"6C",X"BD",X"E2",X"0C",
		X"B6",X"A0",X"3E",X"4A",X"27",X"07",X"30",X"1C",X"86",X"83",X"BD",X"E2",X"0C",X"B6",X"A0",X"3E",
		X"27",X"34",X"84",X"03",X"34",X"02",X"8E",X"1B",X"51",X"CE",X"87",X"21",X"E6",X"C6",X"30",X"85",
		X"CC",X"60",X"55",X"7D",X"A0",X"54",X"26",X"09",X"30",X"03",X"86",X"70",X"BD",X"E2",X"0C",X"86",
		X"71",X"BD",X"E2",X"0C",X"35",X"02",X"CE",X"87",X"25",X"A6",X"C6",X"C6",X"DD",X"BD",X"E2",X"0C",
		X"CC",X"65",X"55",X"BD",X"E2",X"0C",X"7D",X"A0",X"54",X"26",X"1E",X"FC",X"A0",X"16",X"10",X"83",
		X"4F",X"E2",X"26",X"1A",X"BD",X"53",X"6C",X"0B",X"BD",X"46",X"DB",X"87",X"37",X"05",X"A1",X"5F",
		X"86",X"B4",X"A7",X"04",X"CC",X"00",X"F0",X"20",X"08",X"CC",X"00",X"F0",X"20",X"11",X"CC",X"00",
		X"B4",X"34",X"06",X"BD",X"46",X"DB",X"87",X"65",X"06",X"A1",X"5F",X"35",X"06",X"ED",X"04",X"35",
		X"F0",X"0A",X"06",X"04",X"00",X"61",X"62",X"63",X"64",X"BD",X"4B",X"9E",X"85",X"F0",X"26",X"02",
		X"8A",X"F0",X"C6",X"DD",X"7E",X"E2",X"0F",X"6A",X"24",X"10",X"27",X"C0",X"18",X"BD",X"87",X"45",
		X"EC",X"3E",X"DD",X"42",X"39",X"34",X"06",X"86",X"1A",X"C6",X"31",X"88",X"04",X"C8",X"04",X"FD",
		X"CA",X"06",X"CC",X"2A",X"66",X"FD",X"CA",X"04",X"CC",X"D7",X"7C",X"FD",X"CA",X"02",X"86",X"0E",
		X"B7",X"CA",X"00",X"35",X"86",X"EC",X"24",X"83",X"00",X"01",X"ED",X"24",X"10",X"27",X"BF",X"E5",
		X"86",X"40",X"FE",X"A0",X"16",X"11",X"83",X"4F",X"E2",X"26",X"02",X"86",X"02",X"97",X"1E",X"EC",
		X"3E",X"DD",X"42",X"39",X"BD",X"8B",X"F4",X"8E",X"9F",X"FD",X"10",X"8E",X"A0",X"9A",X"B6",X"A0",
		X"0A",X"2A",X"02",X"1E",X"12",X"34",X"30",X"BD",X"31",X"49",X"BD",X"46",X"DB",X"87",X"B2",X"0E",
		X"A1",X"5F",X"35",X"60",X"10",X"AF",X"08",X"EF",X"0A",X"96",X"8A",X"A7",X"0D",X"0F",X"8A",X"7E",
		X"2E",X"DA",X"CC",X"00",X"3C",X"BD",X"34",X"19",X"8E",X"CC",X"0A",X"BD",X"4A",X"5F",X"27",X"59",
		X"1F",X"23",X"86",X"13",X"B7",X"A0",X"0A",X"10",X"AE",X"48",X"BD",X"88",X"22",X"A7",X"4C",X"1F",
		X"32",X"CC",X"87",X"DB",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"7D",X"A1",X"C2",X"26",X"05",
		X"EC",X"3E",X"DD",X"42",X"39",X"1F",X"23",X"A6",X"4D",X"4A",X"27",X"29",X"86",X"07",X"97",X"1E",
		X"86",X"B4",X"B7",X"A0",X"0A",X"10",X"AE",X"4A",X"BD",X"88",X"22",X"AA",X"4C",X"A7",X"4C",X"1F",
		X"32",X"CC",X"88",X"0B",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"7D",X"A1",X"C2",X"26",X"05",
		X"EC",X"3E",X"DD",X"42",X"39",X"6D",X"2C",X"26",X"06",X"CC",X"00",X"F0",X"BD",X"34",X"19",X"7E",
		X"2E",X"D4",X"34",X"74",X"7F",X"A1",X"C2",X"8E",X"CE",X"C8",X"BD",X"89",X"2A",X"25",X"0E",X"8E",
		X"DE",X"2A",X"BD",X"89",X"2A",X"25",X"06",X"4F",X"73",X"A1",X"C2",X"35",X"F4",X"34",X"30",X"BD",
		X"32",X"0F",X"BD",X"31",X"D8",X"8E",X"4D",X"4F",X"BD",X"2E",X"44",X"C6",X"99",X"86",X"68",X"BD",
		X"E2",X"03",X"8E",X"4E",X"4E",X"BD",X"2E",X"44",X"C6",X"FF",X"86",X"68",X"BD",X"E2",X"03",X"8E",
		X"46",X"49",X"BD",X"2E",X"44",X"C6",X"11",X"86",X"C3",X"BD",X"E2",X"03",X"86",X"BA",X"BD",X"E2",
		X"03",X"86",X"C4",X"BD",X"E2",X"03",X"8E",X"3E",X"49",X"BD",X"2E",X"44",X"C6",X"11",X"86",X"C5",
		X"BD",X"E2",X"03",X"86",X"6B",X"BD",X"E2",X"03",X"86",X"C6",X"BD",X"E2",X"03",X"86",X"C7",X"BD",
		X"E2",X"03",X"8E",X"36",X"53",X"BD",X"2E",X"44",X"C6",X"22",X"86",X"C8",X"BD",X"E2",X"03",X"86",
		X"C9",X"BD",X"E2",X"03",X"86",X"CA",X"BD",X"E2",X"03",X"BD",X"8A",X"88",X"BD",X"46",X"DB",X"8A",
		X"BA",X"32",X"A1",X"66",X"35",X"60",X"10",X"AF",X"0A",X"EF",X"0C",X"86",X"03",X"A7",X"88",X"2D",
		X"CC",X"88",X"D8",X"ED",X"88",X"2E",X"CC",X"1E",X"77",X"ED",X"88",X"30",X"86",X"0B",X"A7",X"09",
		X"CC",X"03",X"84",X"ED",X"0F",X"43",X"35",X"F4",X"AE",X"4A",X"8C",X"CE",X"C8",X"26",X"23",X"BD",
		X"89",X"4D",X"BE",X"A1",X"C3",X"26",X"06",X"10",X"BF",X"A1",X"C3",X"20",X"0F",X"10",X"BF",X"A1",
		X"C5",X"10",X"BC",X"A1",X"C3",X"22",X"05",X"30",X"0E",X"BF",X"A1",X"C3",X"BD",X"89",X"7B",X"8E",
		X"DE",X"2A",X"BD",X"89",X"4D",X"BE",X"A1",X"C7",X"26",X"06",X"10",X"BF",X"A1",X"C7",X"20",X"0F",
		X"10",X"BF",X"A1",X"C9",X"10",X"BC",X"A1",X"C7",X"22",X"05",X"30",X"0E",X"BF",X"A1",X"C7",X"BD",
		X"89",X"7B",X"73",X"A1",X"C2",X"1F",X"32",X"7E",X"47",X"55",X"34",X"36",X"C6",X"04",X"BD",X"4A",
		X"5F",X"A1",X"A0",X"25",X"05",X"22",X"07",X"5A",X"26",X"F4",X"1A",X"01",X"35",X"B6",X"1C",X"FE",
		X"35",X"B6",X"34",X"36",X"E6",X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"34",X"10",X"10",
		X"AE",X"4C",X"86",X"1E",X"34",X"02",X"6A",X"E4",X"27",X"09",X"30",X"12",X"BD",X"89",X"2A",X"25",
		X"F5",X"30",X"0E",X"34",X"10",X"AE",X"63",X"1F",X"12",X"86",X"0E",X"30",X"12",X"AC",X"E4",X"25",
		X"07",X"BD",X"89",X"42",X"31",X"32",X"20",X"F3",X"32",X"65",X"39",X"1F",X"21",X"10",X"AE",X"4C",
		X"C6",X"04",X"A6",X"A0",X"BD",X"4A",X"78",X"5A",X"26",X"F8",X"BD",X"8A",X"1A",X"39",X"EC",X"E4",
		X"FD",X"A1",X"DF",X"0F",X"80",X"BD",X"8E",X"3D",X"BD",X"46",X"DB",X"89",X"A3",X"32",X"A1",X"66",
		X"7E",X"2E",X"DA",X"7F",X"CA",X"01",X"BD",X"32",X"45",X"8E",X"4E",X"36",X"BD",X"2E",X"44",X"C6",
		X"11",X"86",X"CB",X"BD",X"E2",X"03",X"86",X"CC",X"BD",X"E2",X"03",X"86",X"CD",X"BD",X"E2",X"03",
		X"BD",X"8A",X"88",X"86",X"0A",X"C6",X"36",X"8E",X"CE",X"D6",X"BD",X"4A",X"78",X"5A",X"26",X"FA",
		X"A7",X"29",X"86",X"1B",X"A7",X"A8",X"2D",X"CC",X"89",X"F4",X"ED",X"A8",X"2E",X"CC",X"00",X"00",
		X"ED",X"2F",X"CC",X"38",X"18",X"ED",X"A8",X"30",X"BD",X"8A",X"70",X"CC",X"40",X"18",X"ED",X"A8",
		X"30",X"7E",X"8A",X"BA",X"8E",X"CE",X"D6",X"BD",X"8A",X"1A",X"CC",X"8A",X"09",X"ED",X"A8",X"2E",
		X"CC",X"38",X"18",X"ED",X"A8",X"30",X"7E",X"8A",X"BA",X"8E",X"CF",X"0C",X"BD",X"8A",X"1A",X"BD",
		X"31",X"49",X"10",X"CE",X"BF",X"00",X"6E",X"9F",X"A1",X"DF",X"34",X"26",X"31",X"C8",X"12",X"E6",
		X"C8",X"2D",X"A6",X"A0",X"BD",X"4A",X"78",X"5A",X"26",X"F8",X"35",X"A6",X"34",X"16",X"BD",X"8A",
		X"62",X"30",X"89",X"FE",X"00",X"86",X"33",X"BD",X"E2",X"00",X"35",X"96",X"34",X"76",X"BD",X"8A",
		X"62",X"A6",X"49",X"C6",X"FF",X"BD",X"E2",X"00",X"35",X"F6",X"34",X"16",X"BD",X"8A",X"62",X"BF",
		X"CA",X"04",X"8E",X"02",X"0C",X"BF",X"CA",X"06",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",
		X"35",X"96",X"34",X"06",X"A6",X"48",X"C6",X"08",X"3D",X"E3",X"C8",X"30",X"1F",X"01",X"35",X"86",
		X"34",X"46",X"1F",X"23",X"E6",X"A8",X"2D",X"E7",X"28",X"C6",X"99",X"6A",X"28",X"2B",X"05",X"BD",
		X"8A",X"2C",X"20",X"F7",X"6C",X"28",X"35",X"C6",X"34",X"36",X"8E",X"2E",X"50",X"BD",X"2E",X"44",
		X"C6",X"22",X"86",X"CE",X"BD",X"E2",X"03",X"86",X"CF",X"BD",X"E2",X"03",X"86",X"79",X"BD",X"E2",
		X"03",X"8E",X"26",X"46",X"BD",X"2E",X"44",X"C6",X"22",X"86",X"7A",X"BD",X"E2",X"03",X"86",X"D0",
		X"BD",X"E2",X"03",X"86",X"CD",X"BD",X"E2",X"03",X"35",X"B6",X"6F",X"28",X"86",X"0A",X"E6",X"A8",
		X"2D",X"33",X"A8",X"11",X"A7",X"C5",X"5A",X"26",X"FB",X"86",X"03",X"A7",X"2E",X"BD",X"8A",X"70",
		X"CC",X"8A",X"DA",X"ED",X"22",X"EC",X"3E",X"DD",X"42",X"39",X"1F",X"23",X"AE",X"4F",X"30",X"1F",
		X"26",X"03",X"6E",X"D8",X"2E",X"AF",X"4F",X"C6",X"11",X"BD",X"8A",X"2C",X"BD",X"8A",X"3C",X"6D",
		X"4E",X"27",X"04",X"6A",X"4E",X"20",X"5A",X"BD",X"48",X"F3",X"84",X"0F",X"27",X"53",X"C6",X"03",
		X"E7",X"4E",X"E6",X"49",X"81",X"01",X"27",X"37",X"81",X"02",X"27",X"3B",X"34",X"02",X"C6",X"12",
		X"E7",X"4E",X"C6",X"99",X"BD",X"8A",X"2C",X"E6",X"49",X"A6",X"48",X"8B",X"12",X"E7",X"C6",X"35",
		X"02",X"81",X"04",X"27",X"0B",X"A6",X"48",X"4C",X"A1",X"C8",X"2D",X"26",X"08",X"6E",X"D8",X"2E",
		X"A6",X"48",X"27",X"1D",X"4A",X"A7",X"48",X"8B",X"12",X"E6",X"C6",X"E7",X"49",X"20",X"12",X"5C",
		X"C1",X"2E",X"23",X"08",X"5F",X"20",X"05",X"5A",X"2A",X"02",X"C6",X"2E",X"E7",X"49",X"BD",X"8A",
		X"4A",X"1F",X"32",X"EC",X"3E",X"DD",X"42",X"39",X"BD",X"8E",X"5E",X"8E",X"DC",X"94",X"CC",X"00",
		X"01",X"7E",X"8B",X"9E",X"8E",X"CD",X"32",X"CC",X"00",X"03",X"BD",X"8B",X"9E",X"8E",X"DC",X"94",
		X"CC",X"00",X"01",X"BD",X"8B",X"9E",X"7F",X"CA",X"01",X"BD",X"32",X"45",X"8E",X"4D",X"30",X"BD",
		X"2E",X"44",X"C6",X"11",X"86",X"B9",X"BD",X"E2",X"03",X"86",X"BA",X"BD",X"E2",X"03",X"86",X"D1",
		X"BD",X"E2",X"03",X"86",X"D2",X"BD",X"E2",X"03",X"86",X"7F",X"BD",X"F0",X"09",X"39",X"34",X"76",
		X"CE",X"90",X"45",X"8E",X"CF",X"42",X"BD",X"4A",X"5F",X"4C",X"84",X"03",X"30",X"1E",X"BD",X"4A",
		X"78",X"48",X"10",X"8E",X"8C",X"03",X"10",X"AE",X"A6",X"AE",X"62",X"C6",X"1E",X"34",X"04",X"EC",
		X"61",X"BD",X"4A",X"84",X"1F",X"30",X"BD",X"4A",X"84",X"1E",X"89",X"8B",X"35",X"19",X"1E",X"89",
		X"8B",X"97",X"19",X"1F",X"03",X"C6",X"03",X"A6",X"A0",X"BD",X"4A",X"78",X"5A",X"26",X"F8",X"10",
		X"8C",X"8C",X"65",X"26",X"04",X"10",X"8E",X"8C",X"0B",X"6A",X"E4",X"26",X"D2",X"32",X"61",X"BD",
		X"8B",X"F4",X"35",X"F6",X"4F",X"5F",X"FD",X"A1",X"C3",X"FD",X"A1",X"C5",X"FD",X"A1",X"C7",X"FD",
		X"A1",X"C9",X"39",X"8C",X"14",X"8C",X"1A",X"8C",X"3B",X"8C",X"5C",X"11",X"19",X"0E",X"15",X"0B",
		X"23",X"12",X"0F",X"0D",X"1D",X"0B",X"17",X"15",X"20",X"0E",X"18",X"27",X"10",X"15",X"14",X"10",
		X"15",X"0B",X"11",X"10",X"1C",X"11",X"23",X"0B",X"15",X"14",X"14",X"15",X"15",X"10",X"16",X"1A",
		X"14",X"17",X"0E",X"19",X"0D",X"14",X"16",X"17",X"0F",X"27",X"24",X"26",X"17",X"26",X"1E",X"13",
		X"17",X"14",X"1C",X"18",X"1E",X"19",X"17",X"1A",X"10",X"24",X"1C",X"1E",X"1A",X"0C",X"10",X"0E",
		X"17",X"0C",X"1D",X"17",X"1C",X"1D",X"0F",X"14",X"1D",X"1D",X"1E",X"1F",X"21",X"13",X"1E",X"17",
		X"19",X"17",X"10",X"0B",X"0D",X"52",X"4F",X"42",X"45",X"52",X"54",X"20",X"4A",X"2E",X"20",X"4D",
		X"49",X"43",X"41",X"4C",X"86",X"00",X"BD",X"55",X"93",X"8E",X"7A",X"00",X"BD",X"55",X"83",X"C6",
		X"DD",X"86",X"4D",X"BD",X"E2",X"0C",X"86",X"4E",X"BD",X"E2",X"0C",X"39",X"EC",X"24",X"83",X"00",
		X"01",X"27",X"0E",X"ED",X"24",X"B6",X"A0",X"13",X"81",X"08",X"2C",X"05",X"EC",X"3E",X"DD",X"42",
		X"39",X"AE",X"9F",X"50",X"35",X"86",X"0A",X"A7",X"88",X"1D",X"DC",X"78",X"ED",X"88",X"11",X"86",
		X"FF",X"A7",X"88",X"13",X"0D",X"94",X"27",X"06",X"4F",X"5F",X"DD",X"81",X"DD",X"83",X"86",X"10",
		X"A7",X"24",X"8E",X"A1",X"74",X"BD",X"46",X"A8",X"BD",X"E1",X"D4",X"27",X"15",X"A6",X"24",X"27",
		X"0C",X"6A",X"24",X"84",X"03",X"CE",X"8C",X"EB",X"EC",X"C6",X"BD",X"74",X"95",X"EC",X"3E",X"DD",
		X"42",X"39",X"CC",X"00",X"1E",X"BD",X"34",X"19",X"7E",X"58",X"32",X"5F",X"5F",X"9F",X"9F",X"5F",
		X"BD",X"31",X"49",X"BD",X"46",X"DB",X"8D",X"0E",X"08",X"A1",X"5F",X"BD",X"46",X"DB",X"84",X"8A",
		X"05",X"A1",X"5F",X"BD",X"46",X"DB",X"52",X"8F",X"05",X"A1",X"5F",X"7E",X"2E",X"DA",X"34",X"20",
		X"86",X"33",X"97",X"80",X"BD",X"32",X"45",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",
		X"FF",X"B7",X"C9",X"00",X"8E",X"8E",X"11",X"10",X"8E",X"8E",X"1F",X"EE",X"81",X"27",X"1A",X"EC",
		X"C1",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",X"EC",X"C1",X"FD",X"CA",X"02",X"EC",X"A1",X"FD",
		X"CA",X"04",X"86",X"0E",X"B7",X"CA",X"00",X"20",X"E2",X"8E",X"80",X"60",X"BD",X"2E",X"44",X"C6",
		X"33",X"86",X"64",X"BD",X"E2",X"0C",X"C6",X"99",X"86",X"D3",X"BD",X"E2",X"0C",X"C6",X"55",X"86",
		X"D4",X"BD",X"E2",X"0C",X"8E",X"72",X"60",X"BD",X"2E",X"44",X"C6",X"33",X"86",X"62",X"BD",X"E2",
		X"0C",X"C6",X"99",X"86",X"D5",X"BD",X"E2",X"0C",X"C6",X"55",X"86",X"D4",X"BD",X"E2",X"0C",X"8E",
		X"64",X"60",X"BD",X"2E",X"44",X"C6",X"33",X"86",X"9B",X"BD",X"E2",X"0C",X"C6",X"99",X"86",X"D6",
		X"BD",X"E2",X"0C",X"C6",X"55",X"86",X"D4",X"BD",X"E2",X"0C",X"8E",X"56",X"60",X"BD",X"2E",X"44",
		X"C6",X"33",X"86",X"63",X"BD",X"E2",X"0C",X"C6",X"99",X"86",X"D7",X"BD",X"E2",X"0C",X"C6",X"55",
		X"86",X"D4",X"BD",X"E2",X"0C",X"8E",X"48",X"60",X"BD",X"2E",X"44",X"C6",X"33",X"86",X"6C",X"BD",
		X"E2",X"0C",X"86",X"C1",X"BD",X"E2",X"0C",X"C6",X"99",X"86",X"D7",X"BD",X"E2",X"0C",X"C6",X"55",
		X"86",X"D4",X"BD",X"E2",X"0C",X"8E",X"35",X"3E",X"BD",X"2E",X"44",X"C6",X"DD",X"86",X"AF",X"BD",
		X"E2",X"03",X"86",X"6B",X"BD",X"E2",X"03",X"86",X"6C",X"BD",X"E2",X"03",X"8E",X"2F",X"59",X"BD",
		X"2E",X"44",X"C6",X"99",X"86",X"D8",X"BD",X"E2",X"03",X"C6",X"55",X"86",X"D4",X"BD",X"E2",X"03",
		X"35",X"22",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"CC",X"01",X"A4",X"BD",X"34",X"19",X"7E",X"2E",
		X"D4",X"0C",X"CB",X"12",X"9D",X"E1",X"EB",X"19",X"E1",X"8E",X"2B",X"1E",X"13",X"00",X"00",X"7C",
		X"3A",X"71",X"40",X"65",X"44",X"54",X"3D",X"59",X"45",X"47",X"3E",X"02",X"01",X"8E",X"2F",X"42",
		X"20",X"BD",X"2F",X"1F",X"7E",X"2E",X"DA",X"5F",X"ED",X"06",X"7E",X"51",X"59",X"86",X"98",X"1F",
		X"8B",X"0F",X"8A",X"BD",X"2E",X"71",X"7E",X"31",X"49",X"F7",X"BF",X"1D",X"BD",X"2E",X"71",X"B6",
		X"C8",X"06",X"7E",X"2E",X"90",X"12",X"12",X"12",X"CC",X"00",X"7E",X"DD",X"51",X"39",X"12",X"12",
		X"12",X"7F",X"A1",X"B4",X"39",X"7D",X"A1",X"BA",X"10",X"27",X"CB",X"5C",X"BD",X"46",X"DB",X"8E",
		X"77",X"08",X"A1",X"5F",X"7E",X"59",X"D4",X"86",X"FF",X"B7",X"A1",X"BC",X"CC",X"00",X"87",X"BD",
		X"34",X"19",X"7F",X"A1",X"BC",X"7F",X"A1",X"B2",X"CC",X"4B",X"C3",X"FD",X"99",X"12",X"7E",X"47",
		X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"3E",X"BB",X"42",X"00",X"00",X"BB",X"45",X"13",X"1D",X"44",X"43",X"0E",X"52",X"11",X"86",
		X"4C",X"3E",X"22",X"45",X"00",X"00",X"22",X"47",X"39",X"2A",X"22",X"3D",X"2F",X"07",X"22",X"49",
		X"26",X"1F",X"22",X"CA",X"4C",X"26",X"99",X"C8",X"5F",X"23",X"33",X"25",X"00",X"00",X"33",X"CB",
		X"34",X"67",X"10",X"8E",X"E2",X"8F",X"20",X"06",X"34",X"67",X"10",X"8E",X"E2",X"25",X"1A",X"FF",
		X"F7",X"CA",X"01",X"8D",X"05",X"7F",X"CA",X"01",X"35",X"E7",X"BF",X"CA",X"04",X"48",X"81",X"6A",
		X"23",X"02",X"86",X"5C",X"10",X"AE",X"A6",X"EC",X"A1",X"88",X"04",X"C8",X"04",X"FD",X"CA",X"06",
		X"10",X"BF",X"CA",X"02",X"86",X"1A",X"B7",X"CA",X"00",X"C8",X"04",X"5C",X"4F",X"30",X"8B",X"39",
		X"34",X"67",X"10",X"8E",X"E2",X"8F",X"20",X"06",X"34",X"67",X"10",X"8E",X"E2",X"25",X"1A",X"FF",
		X"10",X"BF",X"BF",X"02",X"F7",X"CA",X"01",X"4D",X"2C",X"07",X"84",X"7F",X"CE",X"EB",X"7D",X"20",
		X"03",X"CE",X"EA",X"7D",X"33",X"C6",X"EE",X"C6",X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",
		X"BF",X"FF",X"B7",X"C9",X"00",X"A6",X"C4",X"10",X"BE",X"BF",X"02",X"BD",X"8E",X"EA",X"6D",X"C0",
		X"2A",X"F3",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"7F",X"CA",X"01",X"35",X"E7",X"34",
		X"67",X"10",X"8E",X"E2",X"8F",X"20",X"06",X"34",X"67",X"10",X"8E",X"E2",X"25",X"1A",X"FF",X"10",
		X"BF",X"BF",X"02",X"F7",X"CA",X"01",X"44",X"44",X"44",X"44",X"81",X"0A",X"2F",X"02",X"86",X"0A",
		X"10",X"BE",X"BF",X"02",X"BD",X"8E",X"EA",X"A6",X"61",X"84",X"0F",X"81",X"0A",X"2F",X"02",X"86",
		X"0A",X"10",X"BE",X"BF",X"02",X"BD",X"8E",X"EA",X"7F",X"CA",X"01",X"35",X"E7",X"7C",X"BF",X"1E",
		X"20",X"03",X"7F",X"BF",X"1E",X"CE",X"E2",X"0C",X"20",X"0B",X"7C",X"BF",X"1E",X"20",X"03",X"7F",
		X"BF",X"1E",X"CE",X"E2",X"03",X"10",X"8E",X"EF",X"8C",X"31",X"A6",X"10",X"AE",X"A6",X"34",X"02",
		X"B6",X"BF",X"FF",X"34",X"02",X"84",X"FB",X"B7",X"BF",X"FF",X"B7",X"C9",X"00",X"A6",X"61",X"EC",
		X"A1",X"27",X"02",X"1F",X"01",X"E6",X"A0",X"7D",X"BF",X"1E",X"27",X"01",X"5F",X"A6",X"A4",X"84",
		X"7F",X"AD",X"C4",X"6D",X"A0",X"2A",X"E8",X"A7",X"61",X"35",X"02",X"B7",X"BF",X"FF",X"B7",X"C9",
		X"00",X"35",X"02",X"39",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
