-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "F0FB9F0FF9C143EA14D4F4F5324BEB1495213340D89A2661875753315733751D";
    attribute INIT_01 of inst : label is "8AF6398AF5398563985539892E0536247149B5DF6820220AD5577B600CEAACF9";
    attribute INIT_02 of inst : label is "4B1E92011866CBFD621AEE4459DAB570485C001AE71B8E37319CAE5CA921695F";
    attribute INIT_03 of inst : label is "5324FEF7FBDF6BF716BF716BF400001C000086931C7468C6EB80AEB54C19C399";
    attribute INIT_04 of inst : label is "138ACB51594185E06150EFCDDEFFD77EB5E1615090A5132F905220200289A490";
    attribute INIT_05 of inst : label is "88C1B2E34AF349930E611440A5018AA96FDD24882835161A445D324A6494C902";
    attribute INIT_06 of inst : label is "DEA61E974D4DC814402958DFCDDC7576C24A94A653044A9E2A6A8558E76E3522";
    attribute INIT_07 of inst : label is "50245456B420A30204104280010815BDC000975AB02AB0822200002A49B4B57D";
    attribute INIT_08 of inst : label is "A2048105480AA40288AE0280410A00042056B3DE19028B01221A002AD6A24350";
    attribute INIT_09 of inst : label is "B6DD504ADD216D37640A346D56DBA02A84364C2922528B10110E905283A5A36A";
    attribute INIT_0A of inst : label is "DB2A2A2A2680DECBAC97F1A4C02CA68B14D08F46CA81290A0213A9BB2051B36A";
    attribute INIT_0B of inst : label is "250B531552A5EBE47EAF6F9DEA648FD5A3BC48241A7FC0F819209514A137AAC4";
    attribute INIT_0C of inst : label is "8855320C564182F4165714AD43CBCE15542456A523C5404A152D4B52D45DA84A";
    attribute INIT_0D of inst : label is "EADE6C002DCBCF20BD009100AA0677630A0A0C073102A13410243F02FF7E5E82";
    attribute INIT_0E of inst : label is "4C9AC571888621881C5A27EAAAAAAAADB6DB67FFFFF8DB6DB67FFFFF8DB6DB84";
    attribute INIT_0F of inst : label is "2D25A4B49692D25A4B49795AD62B2945CB162C58B162D58B5F00850264C99326";
    attribute INIT_10 of inst : label is "00A8881188055403100A2218010080FF7760F530E92D25A4B49692D25A4B4969";
    attribute INIT_11 of inst : label is "220110A0050020014443002A2018005110C00A88062014443002A2018005110C";
    attribute INIT_12 of inst : label is "70BC10008810028010028C228C08A8811000100C00A20400A004002888600500";
    attribute INIT_13 of inst : label is "E3055FF2A800AA05A2ED1768FB47DA3ED736A9B5EDAB6FAA69649253FE38A15B";
    attribute INIT_14 of inst : label is "943ACD64AC9592B2524A1B7EA7D4F29CA7A99A82A65B74073586C731CF438C38";
    attribute INIT_15 of inst : label is "6220853DB033B7B4EDE2CEB34928759AC94928759AC95929250EB3592B2564A4";
    attribute INIT_16 of inst : label is "2001AA148006908860001A812A1429000C9494A840B3DCD094A012044D554557";
    attribute INIT_17 of inst : label is "71D90761540485428FFC410C386652AA147FE208C3864051466802908D004546";
    attribute INIT_18 of inst : label is "222204645555462A00AA00D0C52DB2380AA314B7D591D4A095001005581E2C47";
    attribute INIT_19 of inst : label is "15F30808D1538E43F22AA9C54E3901100899911988811199955DD99DD5599840";
    attribute INIT_1A of inst : label is "528520409509BA00A0115044D34D31B99A00A0115044D26D3486F4014582AACD";
    attribute INIT_1B of inst : label is "55509AA954AA555DAAAA95554AAAA55555DAAAA95554AA55555DFBEAFFABFED4";
    attribute INIT_1C of inst : label is "A5558AAAA95554AAAA5508AAAA95554AAAA555508AA954AA5508AAAA95554AA5";
    attribute INIT_1D of inst : label is "8AAAA95554AAAA55555DAAAA954AAAA55555DAAAA95554AAAA55555DAA95554A";
    attribute INIT_1E of inst : label is "4AAAA5548AA954AA5508AA954AA5508AA95554AA555508AAAA95554AAAA55550";
    attribute INIT_1F of inst : label is "AA5555552AAAAAAAAAAAAA9555554DD838D1E799C2A95554AA55555DAAAA9555";
    attribute INIT_20 of inst : label is "555555552AAAAAAAAA95555555554AAAAAA9115555555554AAAAAAAAAAAAAAAA";
    attribute INIT_21 of inst : label is "22AAAAAAAAAAAA555555552AAAAA95555555554AAAABBAAAAAAAAAAAAAAAAA55";
    attribute INIT_22 of inst : label is "52AAE4555555555555552AAAAAAAAAAAAAAA95555555554AAAAAAAAAAAA55552";
    attribute INIT_23 of inst : label is "AAAAA555555555555152AAAAAAAAAAA955555554DDAAAAAAAA9555554AAAAAA5";
    attribute INIT_24 of inst : label is "AAAAA955555555555554AAAAAAAAAAB115555555555555555555554AAAAAAAAA";
    attribute INIT_25 of inst : label is "5554AAAAAAAAAAAAAAAAAA55555555276AAAAAAAAAA555555555555552AAAAAA";
    attribute INIT_26 of inst : label is "AAAAAA5555555555552AAAAAAAAAAC45555555555552AAAAAAAAAAAAA9555555";
    attribute INIT_27 of inst : label is "5555552AAAAAAAAAAA89DAAAAAAAAAAAAAAAAAA955555555555554AAAAAAAAAA";
    attribute INIT_28 of inst : label is "955555555555554AAAAAAAAAAAAB11555555555554AAAAAAAAAAAAAAAA555555";
    attribute INIT_29 of inst : label is "A55555555236AAAAAAAAAAAAAAAAAA5555555555555555552AAAAAAAAAAAAAAA";
    attribute INIT_2A of inst : label is "555555555555552AAAAAAAAAAAAAAAAA955555555555554AAAAAAAAAAAAAAAAA";
    attribute INIT_2B of inst : label is "555555554AAAAAAAAAAAAAAAAAAAA555555555555555555552AAAAAAA8EE5555";
    attribute INIT_2C of inst : label is "55555555555552AAAAAAAAAAAAAAA955555555C8AAAAAAAAAAAAAAAA95555555";
    attribute INIT_2D of inst : label is "AAAAAAAAA9555554AAAAAAAA1B95555555555555554AAAAAAAAAAAAAAAA55555";
    attribute INIT_2E of inst : label is "55555555555555772AAAAAAAAAAAAAAAAAA555555555555552AAAAAAAAAAAAAA";
    attribute INIT_2F of inst : label is "555555555555555552AAAAAAAAAAA955555555555555555554AAAAAAAAAAAAAA";
    attribute INIT_30 of inst : label is "AAAAAAAAA95555555555555554AAAAAAAA55555555555555552AAAAAAAAA8445";
    attribute INIT_31 of inst : label is "C6EE119BB91F33770F3B772BCCCBD77A9B7CE213DD9413CECB316182AAAAAAAA";
    attribute INIT_32 of inst : label is "DAA2862D0844FB7BD60D61C5AFCE2F63AD149C39323E34EA7BF7E117BF7EC1E1";
    attribute INIT_33 of inst : label is "26263C3115DACF849214572B0E000A07EBD1FF6D66DE3D005150465EAAEF064D";
    attribute INIT_34 of inst : label is "19090EBD81555BE8120650C0A51136CBE7EF87838D23319CCE13CE3BADEB436B";
    attribute INIT_35 of inst : label is "8ACDA82AA2A82DB6EAEAEAB22D214591694577A1006FD2C2B6E840464242E96A";
    attribute INIT_36 of inst : label is "9E4CE5362839B39CDEA683699529EAA166FABA9123DBAA4294550A420AA90A42";
    attribute INIT_37 of inst : label is "A4912881461D4A431BEE9873720AC92911028C1B7EEEEF534534CA94F450BA79";
    attribute INIT_38 of inst : label is "B5B63B66366487B7DE6366487DFDEEACDE7E36B69059E9A3D5475185CDC82AAA";
    attribute INIT_39 of inst : label is "F6BDEDB98E6398E63D694BDEF7DCC7318A639EF4A5296BE85218E6398B4AD2D7";
    attribute INIT_3A of inst : label is "42308CE52DCE6318E639EB4A5696BEC73988531CD4AD2F6BDF6318C5298E6A53";
    attribute INIT_3B of inst : label is "521EB5AD2F7B6E6398C531CF7A5294B5F731CC721CC38C63294E7B98E639CC61";
    attribute INIT_3C of inst : label is "9990A273998CC8403C88C5281C05901EFB42B98E6398E63D694BDEF7DCE7310B";
    attribute INIT_3D of inst : label is "8CA05038CC0201CCE6722144C623194826399CCA4131CCE50289CE6472890E73";
    attribute INIT_3E of inst : label is "45129CC4720904C73140A007399C884131CC8E44218E4728144E7339900A7311";
    attribute INIT_3F of inst : label is "738F33C4F9CE318CE33E3398E633C738CE38CA71C651C6719CEA18A975D7FCCC";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "DC400DC6C808B5C26C08056B02900F301C000BD4400B01E79D33117773577179";
    attribute INIT_01 of inst : label is "561640561340496410934118B02C256280192F75F7DFDFDFAAA3588D303FF580";
    attribute INIT_02 of inst : label is "180A9209150F50BD1802AECAB078D405803000170B2D5658806C1A3CA86822C2";
    attribute INIT_03 of inst : label is "235CBFE6FF9A79FFC71FF879FE00001C0000C20AA838B161A780D8DB109504A0";
    attribute INIT_04 of inst : label is "E7D75E22B8EFA7E9E8F232323101218B4A007FBF4F1A9EC0BAF64C926EE5325B";
    attribute INIT_05 of inst : label is "DC0420242DFBFC03D46A79AD09603915972618BE6F4AEAE95770E111C223844B";
    attribute INIT_06 of inst : label is "73CF7313E7A2592CBD95E9C4C7FE34C020835350681A23167EAB987DFFEA01B1";
    attribute INIT_07 of inst : label is "F275AF680B67BCA95BDB665294A73ECA5BD98C034BB503C22200000D00C11817";
    attribute INIT_08 of inst : label is "316032A3ED3FDBD6C5B4C6566D994A529CFB04A4C56E51D8B9696D950DE56EB9";
    attribute INIT_09 of inst : label is "100A6B2E05F2E3E115B94102E2014DB4F7817956B75BB473C9E2475BBD331817";
    attribute INIT_0A of inst : label is "2DD54CC459F9A410C906B7160340EA519D4B5C3003B2FDBDBF3A4F08ADCA0817";
    attribute INIT_0B of inst : label is "5509E7BADD0DBDAC81F9421570A9AAFAF55EAF16880009AD98564DA33F00F0E0";
    attribute INIT_0C of inst : label is "99E68379A87B3D06F79F21033DA6D37AAF56A8D7843EF7B5B846308C21705EBF";
    attribute INIT_0D of inst : label is "1F211268D5D8335DBA341E3D573808DEE3F737B80266DB037A53422500ED3698";
    attribute INIT_0E of inst : label is "30410A03D1AF7B5AAEAB590C4C4C4C5965965ACB2CB2B2CB2CE59659396596CB";
    attribute INIT_0F of inst : label is "584A08410C2584A08410CA210850126BD5BBF6EFDBBFCADF25B4EDF103040C10";
    attribute INIT_10 of inst : label is "B26916231624CBE62C9A5D31E4D57D0282829E7E82584A08410C2584A08410C2";
    attribute INIT_11 of inst : label is "C592F94792F9C7934BA63C9A5D3164D2F98F2697CC5934BA62C9A5D3164D2F98";
    attribute INIT_12 of inst : label is "5400A2C97CA2C97CA3D91845184BB74E2C912E98B25F28F65F38F26974C792E9";
    attribute INIT_13 of inst : label is "2C5CE002EB26E77ADD96ECB725B92DC968CB565A92D090D4823B6DB8006535E0";
    attribute INIT_14 of inst : label is "6EC0B05B0B616C2DADB7630118230C62188620FD56F25F280EA2539CA7ECB0C3";
    attribute INIT_15 of inst : label is "6F01B4AC46C0C68FA3EF002CB6DD8160B6B6DD8160B616D6DBB02C16C2D85B5B";
    attribute INIT_16 of inst : label is "D2C9954A4B276E668F2C99769BEA94964C4D6A459D3BFFEBF6E43ADCC1A49A4A";
    attribute INIT_17 of inst : label is "285D7765EE5A959BBFFE0B550A2EA044DDFFF05B50A2E4088CD52B4B42A563A0";
    attribute INIT_18 of inst : label is "775572BBBBAABB44CCC4CC998DEBA509934637AD2D2842484CB8CCC964D25404";
    attribute INIT_19 of inst : label is "7ED6693C47E73D2DB079F39F9CF0B4CDDDDDD555555CCAEEEEE662222AAEED37";
    attribute INIT_1A of inst : label is "1B13B1E65894257DF6CEB12960915800057DF6CEB129619155200AFBE98B9F59";
    attribute INIT_1B of inst : label is "66621B3198CC6675B33319998CCCC666675B33319998CC666675EEBFAAABFE90";
    attribute INIT_1C of inst : label is "C6620B33319998CCCC6620B33319998CCCC666620B3198CC6620B33319998CC6";
    attribute INIT_1D of inst : label is "5B33319998CCCC666620B333198CCCC666620B33319998CCCC666620B319998C";
    attribute INIT_1E of inst : label is "8CCCC6675B3198CC6675B3198CC6675B319998CC666675B33319998CCCC66667";
    attribute INIT_1F of inst : label is "CC6666663333333333333319999985F0C4B271A3B3319998CC666675B3331999";
    attribute INIT_20 of inst : label is "66666666333333333319999999998CCCCCC1419999999998CCCCCCCCCCCCCCCC";
    attribute INIT_21 of inst : label is "D6CCCCCCCCCCCC6666666633333319999999998CCCC142CCCCCCCCCCCCCCCC66";
    attribute INIT_22 of inst : label is "6333AF66666666666666333333333333333319999999998CCCCCCCCCCCC66667";
    attribute INIT_23 of inst : label is "CCCCC666666666666663333333333331999999985F333333331999998CCCCCC6";
    attribute INIT_24 of inst : label is "33333199999999999998CCCCCCCCCC1419999999999999999999998CCCCCCCCC";
    attribute INIT_25 of inst : label is "9998CCCCCCCCCCCCCCCCCC66666666782CCCCCCCCCC666666666666663333333";
    attribute INIT_26 of inst : label is "CCCCCC66666666666633333333333AF666666666666333333333333331999999";
    attribute INIT_27 of inst : label is "66666633333333333301F333333333333333333199999999999998CCCCCCCCCC";
    attribute INIT_28 of inst : label is "199999999999998CCCCCCCCCCCC141999999999998CCCCCCCCCCCCCCCC666666";
    attribute INIT_29 of inst : label is "C666666667C2CCCCCCCCCCCCCCCCCC6666666666666666663333333333333333";
    attribute INIT_2A of inst : label is "66666666666666333333333333333333199999999999998CCCCCCCCCCCCCCCCC";
    attribute INIT_2B of inst : label is "999999998CCCCCCCCCCCCCCCCCCCC66666666666666666666333333331AF6666";
    attribute INIT_2C of inst : label is "666666666666633333333333333331999999980A333333333333333319999999";
    attribute INIT_2D of inst : label is "3333333331999998CCCCCCCCB419999999999999998CCCCCCCCCCCCCCCC66666";
    attribute INIT_2E of inst : label is "666666666666667D6CCCCCCCCCCCCCCCCCC66666666666666333333333333333";
    attribute INIT_2F of inst : label is "66666666666666666333333333333199999999999999999998CCCCCCCCCCCCCC";
    attribute INIT_30 of inst : label is "33333333319999999999999998CCCCCCCC666666666666666633333333331056";
    attribute INIT_31 of inst : label is "9AA8BA280B890151790951564002D51BBE6426AAC7C89E407D78A83B33333333";
    attribute INIT_32 of inst : label is "DFCCE381694AAAD6B553AA9DE24389F3FDF9E9B4467CC06900040B801843F8A8";
    attribute INIT_33 of inst : label is "68DFA552305759324976015D44C0000102F508EBAF7E52BEFB2C8B854EA2289F";
    attribute INIT_34 of inst : label is "E3F3E4C81EB28497007C69BB7782A49E13082C9880B4341A0EA2AFF56B5A741D";
    attribute INIT_35 of inst : label is "7D327DF5FD7FF001DF5FDFD7E1EF3EBF06FE807ADB813F6F409FB7A9F5EF3FBF";
    attribute INIT_36 of inst : label is "F3D613C844AE404049557C96E9DAA326196DE7AB482679CEF7EB3BDEF5EF79CE";
    attribute INIT_37 of inst : label is "E805E425E4D1A9BC0089B9F57B57D40F484BC9A01A00A4AABA4B74ED509304B6";
    attribute INIT_38 of inst : label is "0817284FCA05288410BCA052878FFF75FE8DB6E81A0351B46ABCBBA3D5ED47CF";
    attribute INIT_39 of inst : label is "842148B98C7398A4398E6290855CC6398C4218C631CE522C7310842144210820";
    attribute INIT_3A of inst : label is "88431802058E631484298C6318E522E7398E6214E639884211731CC739486399";
    attribute INIT_3B of inst : label is "73084218C0002E631CC6210C6318E7291631CC731486318C42108B18C7318E51";
    attribute INIT_3C of inst : label is "0898C46201404E633440863918BF2EF04504B98C7398A4398E6290855CE731CF";
    attribute INIT_3D of inst : label is "40C462340F33118880503188C412818C6728100C6331008623118A2243118E42";
    attribute INIT_3E of inst : label is "062318A0439988E4298CC44620100C633904080639880439988C41281C8C7281";
    attribute INIT_3F of inst : label is "779F73DCFBCEF3BCEF3EF3B9EE77CF79DE7BCAF3DE57CEF3BCE21289D7DDD008";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "A4D09A4D14B033CD88EE659232F4802218008054424381041202240642246250";
    attribute INIT_01 of inst : label is "0ED7244ED72452725127251F0904107C48388088A0202A002A20214536555581";
    attribute INIT_02 of inst : label is "388A820914093994AAABAACCD1F0C3E57170000E8A5514A809B56050E12121DA";
    attribute INIT_03 of inst : label is "C99EBE22F88A31F1C31F1C39FC00001400008E7218B5E3C6AA0048C9582820B0";
    attribute INIT_04 of inst : label is "C4355A8CBB69A9EA7A3100110110180000009DA457309E50BA96104131B249A6";
    attribute INIT_05 of inst : label is "5727198938907C09E5385B696844EC4635628914EE4B3EE99627911FA33E445B";
    attribute INIT_06 of inst : label is "F94F2603F2B45C0A3B7870C114450711A10EBD9B8C230E08558C25DD73B8D741";
    attribute INIT_07 of inst : label is "D1172662B931389E63B6D338C63BDB64F676F35B88E7B32888AAAA9944CF6D77";
    attribute INIT_08 of inst : label is "31D3ECB34C9B9CCEE2EFBB99DB4CE318EF6DDE4F99DB168CE1D5DA46D3B992CC";
    attribute INIT_09 of inst : label is "A6D5CE82D9C385C6E76C4F6F34DABA06CCB67274E476C6D88DCDDC76C68D7B79";
    attribute INIT_0A of inst : label is "3EEEF66673A0DFFD2CB47C1D27CEFB17DF63B2F6FEECE9999E98AE373B627B79";
    attribute INIT_0B of inst : label is "1BE4A7825C7094AE64E77DE48EED051B376ACC1C893FC0C64C74166DBD4D7012";
    attribute INIT_0C of inst : label is "E9CCB1973F7BE7F6758F8D9B39E9DC7337A736E632B779D98BDAD6B5AD776733";
    attribute INIT_0D of inst : label is "5373BA70E05C74590B365C8C518F18929B9196338332C281331338010B2F4CC6";
    attribute INIT_0E of inst : label is "E5E9CBF3198E739CF8BB7BCE66EE66FDBFDBFFEDFEDBFB7FB7BFDBFDAFF6FFCF";
    attribute INIT_0F of inst : label is "D11A2364688991322444CB31AE5FBF6E5EDD3A76EDD30F4CB5E4E5E72E5EBD72";
    attribute INIT_10 of inst : label is "732C4629462773328CCB19946E00A8008A22CA7C88D11A2364688991322444C8";
    attribute INIT_11 of inst : label is "5198CC51B8CC519963328CCB19946658DCA372C6E519963729CCB1B946658CCA";
    attribute INIT_12 of inst : label is "7C6A68CC6629CC6668CC4C514C4EC6628CC18CCA731B9A331B8A332C6E51B8DC";
    attribute INIT_13 of inst : label is "0E76605BAE1DB39DE82E617A0B985E83F61F20FD87CC3CE1DAFD34DBFE34B1C1";
    attribute INIT_14 of inst : label is "B6C2211A22646889B4D376C6B2D752C8BA2CC38008A17F2D9ABB38C632AEB0E3";
    attribute INIT_15 of inst : label is "096E6690A2D9511745ED64889A6DC46226DA6D84423444DA4DB88C44C8D11369";
    attribute INIT_16 of inst : label is "998D46632635B3279998D46F0BCCC64C68E5B7260F2294B3DC30EBB6A2362362";
    attribute INIT_17 of inst : label is "0055D4527732C736CAAB23778B2B3931B655591B78B287262A998E639B31D9CD";
    attribute INIT_18 of inst : label is "E644C4515100400888800034B24E3791E652C939B9BCC702E0C264F1C8E38005";
    attribute INIT_19 of inst : label is "8A97CC79D8A7E531B25C53E29F95C3B99BB991111331115445544000011000E6";
    attribute INIT_1A of inst : label is "5C49E27074C0A6E4EC74E3C1E1F96CEC86E4EC74E3C1E1F9F5F3ADC9DC0BC55D";
    attribute INIT_1B of inst : label is "8787E3C1E0F07800BC3C1E1E0F0F078782A3C3C1E1E0F0787800FD77F5D60BC0";
    attribute INIT_1C of inst : label is "0787F3C3C1E1E0F0F07855BC3C1E1E0F0F078787F3C1E0F07855BC3C1E1E0F07";
    attribute INIT_1D of inst : label is "F3C3C1E1E0F0F0787855BC3C1E0F0F078787F3C3C1E1E0F0F0787855BC1E1E0F";
    attribute INIT_1E of inst : label is "0F0F0787F3C1E0F07855BC1E0F0787F3C1E1E0F0787855BC3C1E1E0F0F078787";
    attribute INIT_1F of inst : label is "F07878783C3C3C3C3C3C3C1E1E1E05FA67E05EE103C1E1E0F0787855BC3C1E1E";
    attribute INIT_20 of inst : label is "787878783C3C3C3C3C1E1E1E1E1E0F0F0F0155E1E1E1E1E0F0F0F0F0F0F0F0F0";
    attribute INIT_21 of inst : label is "A8F0F0F0F0F0F0787878783C3C3C1E1E1E1E1E0F0F0154F0F0F0F0F0F0F0F078";
    attribute INIT_22 of inst : label is "83C150787878787878783C3C3C3C3C3C3C3C1E1E1E1E1E0F0F0F0F0F0F078782";
    attribute INIT_23 of inst : label is "0F0F0787878787878783C3C3C3C3C3C1E1E1E1E1A03C3C3C3C1E1E1E0F0F0F07";
    attribute INIT_24 of inst : label is "C3C3C1E1E1E1E1E1E1E0F0F0F0F0F0EA9E1E1E1E1E1E1E1E1E1E1E0F0F0F0F0F";
    attribute INIT_25 of inst : label is "E1E0F0F0F0F0F0F0F0F0F078787878556F0F0F0F0F0787878787878783C3C3C3";
    attribute INIT_26 of inst : label is "F0F0F07878787878783C3C3C3C3C2AF7878787878783C3C3C3C3C3C3C1E1E1E1";
    attribute INIT_27 of inst : label is "7878783C3C3C3C3C3C01FBC3C3C3C3C3C3C3C3C1E1E1E1E1E1E1E0F0F0F0F0F0";
    attribute INIT_28 of inst : label is "1E1E1E1E1E1E1E0F0F0F0F0F0F0155E1E1E1E1E1E0F0F0F0F0F0F0F0F0787878";
    attribute INIT_29 of inst : label is "0787878782A8F0F0F0F0F0F0F0F0F07878787878787878783C3C3C3C3C3C3C3C";
    attribute INIT_2A of inst : label is "787878787878783C3C3C3C3C3C3C3C3C1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F";
    attribute INIT_2B of inst : label is "1E1E1E1E0F0F0F0F0F0F0F0F0F0F0787878787878787878783C3C3C3C3507878";
    attribute INIT_2C of inst : label is "87878787878783C3C3C3C3C3C3C3C1E1E1E1E1F53C3C3C3C3C3C3C3C1E1E1E1E";
    attribute INIT_2D of inst : label is "C3C3C3C3C1E1E1E0F0F0F0F0EA9E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0F078787";
    attribute INIT_2E of inst : label is "78787878787878556F0F0F0F0F0F0F0F0F0787878787878783C3C3C3C3C3C3C3";
    attribute INIT_2F of inst : label is "878787878787878783C3C3C3C3C3C1E1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F0";
    attribute INIT_30 of inst : label is "C3C3C3C3C1E1E1E1E1E1E1E1E0F0F0F0F078787878787878783C3C3C3C3C0057";
    attribute INIT_31 of inst : label is "F24DAEA91F829523729123FCA4199232080A76B90C8898A4557AA8EBC3C3C3C3";
    attribute INIT_32 of inst : label is "DF44F5B9CE725318C6E6AEF084A68E2A51A9EF24C67FB06E4207EB84A07C482E";
    attribute INIT_33 of inst : label is "6388C51CD5355DE9249814956780080446071F12AC7FBB7277388E8E4A463A9F";
    attribute INIT_34 of inst : label is "99C99ADFBCD0DB7E02F670B7A61896DC440FF89C24EE974FA7C142C58C6369D5";
    attribute INIT_35 of inst : label is "B9ED46C44C64E7BD3535B55781004ABC8372FD3D1D6C9C8CBE4E46377B74CE4C";
    attribute INIT_36 of inst : label is "CF5BA6FE4ED7F7544D677FDBBD7A63A61FBF9EB9FEBF42942588129431821084";
    attribute INIT_37 of inst : label is "4A4DF121A7332EDBEE2F3E050B65148FE2434E4177AAA6B3BFEDDEBD30D30FDF";
    attribute INIT_38 of inst : label is "6315210B6C65F2105EF6C65B20346255FE1525085E365545B6D963F8142F81CD";
    attribute INIT_39 of inst : label is "84210AA10A4294A5635AC6B58C5085214A429084214A42284290A4215AC6B18C";
    attribute INIT_3A of inst : label is "25294250850A5294A42B18C631AD62A42948421484210842154214A5210A5291";
    attribute INIT_3B of inst : label is "529085290842284290A521508421294214214A42948D6B18C6B18A10A4210A54";
    attribute INIT_3C of inst : label is "00108042090408403400852010ABAFBEAFEBA10A4294A5214A42948454852949";
    attribute INIT_3D of inst : label is "00A050300D120100A0512900850281080520144A402944840201082042094A42";
    attribute INIT_3E of inst : label is "24029480528144842904800420900840210048042948042810484028940A4201";
    attribute INIT_3F of inst : label is "BDCF9DF67CF7B9CF7B9F3DECF3BDE79EF73CF3B9E79DE73DEE6A3A0B7777D008";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "70B8970978E027D5486629921CE4E602700898104C06038E3C40600446620042";
    attribute INIT_01 of inst : label is "42441402431400415403155805044060287A008A82282A28A28BA15CBC519C09";
    attribute INIT_02 of inst : label is "7A80920910CDD15041020EC885B060E100A400062E065C0CA8008110A8282048";
    attribute INIT_03 of inst : label is "F8C701080424A0090A8094A81A0000100000A2E10D40A1450200CA795404A028";
    attribute INIT_04 of inst : label is "F021C6B8865819E6760200000000000000003DF65630EE63918078E31D9F6FBE";
    attribute INIT_05 of inst : label is "6E42399C36780D0837025D293C06D7E2C9121765776664E50B59F1936226C44F";
    attribute INIT_06 of inst : label is "8665510D0CD2450E33B050CBD2233AB591AD6B12CEF3AD5F870779A59C79C6C0";
    attribute INIT_07 of inst : label is "D11AE72E99315F8EF3B49B19CE31992CE6E69349F8C79BFDDDF5557144052D2A";
    attribute INIT_08 of inst : label is "91B8CC93659B98C564733BBDD26C6738C66496CFCEB312A8D5ADBA45B3B9DB8C";
    attribute INIT_09 of inst : label is "46638EA2CFFA8BC25ACC456668CC7A8458B2F75CDDACC598A8E49BACC5892B33";
    attribute INIT_0A of inst : label is "1323332333B0B6592DBCEE5B0BC75313EA633672CECCECB98E956F12D6622B33";
    attribute INIT_0B of inst : label is "1AAF32B25DDF67A2B6736DA48ACC65132662C5DB092A0096C01406677E461980";
    attribute INIT_0C of inst : label is "79F895A624FDC48F63A0A54ABE499E7F77BBF57AB7F779D389CE7394A56FE73B";
    attribute INIT_0D of inst : label is "7BB59B78FC2CB6F9877A4F9C7199297BD5F19F908EF4599133136E010B924F5A";
    attribute INIT_0E of inst : label is "F5C8EB2B55EF6BDABFBF7BEBA3B23A369A4D3D269B4F49A6D2D369A4B4DA69C7";
    attribute INIT_0F of inst : label is "911222644C8911222444D998C4595BEE4C99B264CD93266C1FEEFDF7AE5EB972";
    attribute INIT_10 of inst : label is "2B55C5B9C5EBBF338BD5799C5688888A80A2332EA8D91B2344688D91B2364688";
    attribute INIT_11 of inst : label is "717BDC715BDC717AAF738AD57B9C5EABCCE2B55E6717AAF338BD5799C5EABCCE";
    attribute INIT_12 of inst : label is "314E39BDE678BDE638ADCB71CB457E638BDDBCCE2F7B8E2B7B8E2F55EE715BDC";
    attribute INIT_13 of inst : label is "3EE670556519338BFC1FC0F607B83FC1F84FC27A93D49AF44E5DA4D9502CD6FB";
    attribute INIT_14 of inst : label is "374A311B2264488D3693B2D3782E05C1785E6B5555A9376F13881084229E7BCF";
    attribute INIT_15 of inst : label is "04902590AE71211545E4C68CD26ED44234D26ED44224469B4DD28C44C8911A6D";
    attribute INIT_16 of inst : label is "18ABDCE162AE4B47319BBDCE09B9C2CDDDEA0F67CE5B584B0B1E91F46722F22D";
    attribute INIT_17 of inst : label is "E75EB27763B272E4EFFF26B9931CA9BF277FF9359931C537CC738C720E719D0F";
    attribute INIT_18 of inst : label is "EECC44115544002AAAA22276F346139DFE7BCD18989C9F71ECF56AFCF2F5B3B9";
    attribute INIT_19 of inst : label is "F3D1E7BCBF32F8BF4555997CCBE6F1999BBBB333311110444555511110000066";
    attribute INIT_1A of inst : label is "35C97E576EDD8C74E4D86371F05E64C9AC74E4D86371F05C799338E9CA7559C6";
    attribute INIT_1B of inst : label is "0007D3FC00FF005D3FFFC01FEFFFF007FFFBFC0001FE00007FD77FF77FFDDF80";
    attribute INIT_1C of inst : label is "F00573FFFDFFFE00FF007FBFFFC01FEFF00007FD500000FF005D003FC01FEFF0";
    attribute INIT_1D of inst : label is "53FFFDFFFE0000007FFF3FFFC00FFFF007FF53FC01FFFEFF00007FFF001FFFEF";
    attribute INIT_1E of inst : label is "0FFFF007F001FE007FDD3FC00FF005D801FE00FF007FFDBFFFDFFFEFFFF00005";
    attribute INIT_1F of inst : label is "FF007F80003FC03FC03FC0001FE007D9F1D7222B2BFDFFFEFF0000573FFFC000";
    attribute INIT_20 of inst : label is "FF807FFF803FC03FC0001FE01FFFE00FF0051001FE01FE000000FF00FF00FF00";
    attribute INIT_21 of inst : label is "80FF00FF00FFFF007F807FBFC03FC0001FE01FEFF004400000FF00FF0000007F";
    attribute INIT_22 of inst : label is "FBFC44007F807F80007F803FC03FC03FC0000000001FE000000FF00FF007F802";
    attribute INIT_23 of inst : label is "000007F807F807F807F803FC03FFFC000001FFFE200000003FC0001FE0000007";
    attribute INIT_24 of inst : label is "0003FDFE01FFFE01FFFE00FF00FF0014401FFFE01FE01FE01FE01FEFFFF00FF0";
    attribute INIT_25 of inst : label is "FE0000FF0000FF00FF00FF7F80007F888FF00FF0000007F807F800000003FFFC";
    attribute INIT_26 of inst : label is "00FFFF7F807F807F803FC03FC0000517F807F80007FBFC0003FC03FFFDFE01FF";
    attribute INIT_27 of inst : label is "7FFF80003FC03FC0001E0003FC03FC03FFFC03FC01FE0001FFFE0000FF0000FF";
    attribute INIT_28 of inst : label is "DFFFFFFFFFFFE00FF00FF00FF00FE801FE01FFFE0000FF0000FF00FF00007F80";
    attribute INIT_29 of inst : label is "07FFFFF805DEFF0000FF00FF00FF00007F80007F80007F80003FFFC03FC03FFF";
    attribute INIT_2A of inst : label is "80007F8000007F803FC03FC0003FC000001FE0001FE000000FFFF00FF00FFFF0";
    attribute INIT_2B of inst : label is "1FE01FFFE00FF00FF00FF00FFFFFF7FFF80007F8000007F80000000003FF007F";
    attribute INIT_2C of inst : label is "07F807F807F803FC03FC03FC03FFFC01FFFE015FBFFFC0000000000000001FE0";
    attribute INIT_2D of inst : label is "FC03FFFFFDFFFFFEFFFF0000BE80001FFFFFE01FFFE00000000FFFFFFFF007F8";
    attribute INIT_2E of inst : label is "7F807F807FFF807F400FF00FFFFFFFF00FF007F80007FFF80003FC03FC0003FF";
    attribute INIT_2F of inst : label is "0007F800000007F8000003FC03FFFDFE01FFFE01FE01FFFE000000FFFFFFFF00";
    attribute INIT_30 of inst : label is "0003FFFFFDFFFE00000001FE0000FF00FF007FFF80007F807FBFC03FC03FD510";
    attribute INIT_31 of inst : label is "7CE43883918F14223F10229FC449622764BC56150E2ABFC46710E0F00003FFFC";
    attribute INIT_32 of inst : label is "E1F5FA12B53C518C6324E27A47C7449D17CC8783104BD41753021985A0213AE0";
    attribute INIT_33 of inst : label is "03E8CC4B9471CCF9A6D811C723C00002C4020410E05F4E3A73BBC5CA74E5A215";
    attribute INIT_34 of inst : label is "93D2A965FB9092DCBDEBA8E73A9B124C640460DE70D78241226D6100C631FD87";
    attribute INIT_35 of inst : label is "365BE4FE4FC4D96FA5A52671554A138AA367267ADADA3D2D6C1EB6E4F4AC9E95";
    attribute INIT_36 of inst : label is "4599282F11B1698D657952DB1A34CFF705968B3464D9E294A5FC5084BF021084";
    attribute INIT_37 of inst : label is "54BBF455BBF7278B4624850205B1297FA8AB77EFE4E632BCA96D8D1A66FB82CB";
    attribute INIT_38 of inst : label is "001433022E2993B04A32C39DB012511C41016B46A8A05AD56389203008149DB9";
    attribute INIT_39 of inst : label is "210800A10A5210846B18C6B1AD508529085200000000002A5214842900000420";
    attribute INIT_3A of inst : label is "10852948550A52148428020004200A84294852918D6B5AC6B14214A421480081";
    attribute INIT_3B of inst : label is "420020084000A842948429108421084214214A5290A94A5094250A9484214842";
    attribute INIT_3C of inst : label is "AA34A8D623051A413540856291FBBEFAEAFBA10A5210844A1084A12954A42109";
    attribute INIT_3D of inst : label is "418A44301C02011188D42151A412035A2C223118C16111AD52A358AA46AB0AC6";
    attribute INIT_3E of inst : label is "0546B582568B01856154A8046A350A5161510AA42908A46A9518D56A3008D601";
    attribute INIT_3F of inst : label is "38EF98E33C633CC671DF38CE7118F78CE79C671DE718F339C72038837F5DF51A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "A1F9BA1D3080A5CE28EC71DA30C8AE8C21190ED2A48C21AEB846464006464464";
    attribute INIT_01 of inst : label is "1403521400521B3521B0520734A9381CA541C0288A08A28A2080ABD73C455D23";
    attribute INIT_02 of inst : label is "4250004021EC6021B0A1012661881660B5800018006800D0A4451125434B4280";
    attribute INIT_03 of inst : label is "2D4381AA06AA900C8900C8900200000000000C8034A0508A0480100207B9940F";
    attribute INIT_04 of inst : label is "2555D66685D61615858A0000000000000000139B61CED92C0161469AC4440049";
    attribute INIT_05 of inst : label is "5434229425CEC58D11A269AD0A0893319D3A26554908AA8F97024A9495292A6B";
    attribute INIT_06 of inst : label is "816C500002D151ACA546AD32C6EE30A4D0C9425D284A095054E149314A494481";
    attribute INIT_07 of inst : label is "6A508F09224584295ACB6C73B5E53EDA09496C904295225D7D5FFFC581031A42";
    attribute INIT_08 of inst : label is "112312A8A36C52B4521464572DB1CED794FB6DA2542450A8912125B50CC5242B";
    attribute INIT_09 of inst : label is "2092297415C381C590914108A41245D43284727095091622A82B130915520845";
    attribute INIT_0A of inst : label is "2666666662CF240248219212B70A6050CC0A5814311294656B600E2C848A0845";
    attribute INIT_0B of inst : label is "5154B628992A962892180952B9EEF567CF68C312542AAD65E816C8E133820B20";
    attribute INIT_0C of inst : label is "1162A170AA7615677000614225B6F0589EE19C31A409ED2528C6318C636214A4";
    attribute INIT_0D of inst : label is "4742204C964042C5CE704229452E900431253CA3432E184A5AD243B54A2DB43C";
    attribute INIT_0E of inst : label is "95298B621B4AC234B5BB621766EFF66DBFFB6B6FF6DEDBFDB7B7FF6DADFFDBCC";
    attribute INIT_0F of inst : label is "620441A81506A0541A810BB18C5B9B6D5860C081020CAC32319CD994A950A142";
    attribute INIT_10 of inst : label is "A6C117A215B099A428B84D214DD77D7FD55DCB67106A0541A815062044188110";
    attribute INIT_11 of inst : label is "451669451669471609A428B04D21C582690A2C134851609A428B04D21C582690";
    attribute INIT_12 of inst : label is "6088A28B3CA29B3CA28B17C513E133CA28B92790A6CD28A2CD28E2C134851669";
    attribute INIT_13 of inst : label is "2AC8EA5841B2472C10E087043829C34E0E3071830C1864330632496A55538C2F";
    attribute INIT_14 of inst : label is "5B841A0D40A811020925D445C4B89F13CCF32A4009ED626F1BB99CE739A8A28A";
    attribute INIT_15 of inst : label is "CC6D9A59EBF109B96E14C50224B708140824B7081408810496E1068150220412";
    attribute INIT_16 of inst : label is "D2A8315ACAA1F2C68D2A8314D122B195425BF2C58D20D433C78E00D800A18A19";
    attribute INIT_17 of inst : label is "CE0075058ADA319B3AAA8FB70E02B4ECD9D5547D70E0369D88053B5BD0A776E0";
    attribute INIT_18 of inst : label is "66444555110000AAAAA2221B11CE7B1BA34C473BDBD8A2DE58B459D468D2A318";
    attribute INIT_19 of inst : label is "6BD5232D36B6992DB4535B5ADA60BBBBB99991111111155554444000000002EE";
    attribute INIT_1A of inst : label is "711314CC4C979149374FE52FB64C608F9149374BE53FB64C718222926E2935D4";
    attribute INIT_1B of inst : label is "F807580000007FDF000000000FF007FFFDD80001FFFEFF7F805DF7F55DDD7700";
    attribute INIT_1C of inst : label is "00077803FC01FE00000077003FDFE00FF007F80773FC00007FF5BFC0001FE007";
    attribute INIT_1D of inst : label is "7000000000FF0000005D803FC0000007F807D80001FE0000FF007FF700000000";
    attribute INIT_1E of inst : label is "E00007FDD00000FF7FF58000000005F3FDFFFE000000753FC0001FEFF0000007";
    attribute INIT_1F of inst : label is "FF00007F803FFFC0003FFFC0001FE7D428A882A90000000000007FF700001FFF";
    attribute INIT_20 of inst : label is "80007FFF803FFFC0001FFFFFE00000000001440001FE00000000FFFF0000FFFF";
    attribute INIT_21 of inst : label is "0800FF00FF00FF007FFF803FC03FC01FE01FFFE00000060000FFFF000000007F";
    attribute INIT_22 of inst : label is "03FD457F807F80000000003FFFC0003FFFFFC01FE0001FE0000FFFF00007F800";
    attribute INIT_23 of inst : label is "FFF0000007FFF80007FBFFFFFC03FC01FE0001FE08003FC03FC01FFFE00FFFF0";
    attribute INIT_24 of inst : label is "FFFC01FFFFFFFFFE0000FFFF00FF0051000000001FFFE0001FFFE00FF0000FFF";
    attribute INIT_25 of inst : label is "FE0000000000FFFFFF00FF007F807FAA0FFFF0000000000007FFFFFFF80003FF";
    attribute INIT_26 of inst : label is "0000007FFF80007FFFBFC0003FC00047F807F807FFFBFFFFFC03FFFFFDFE0001";
    attribute INIT_27 of inst : label is "FFFF8000003FC000000A280003FC0003FFFC03FC0001FFFFFFFE000000FFFF00";
    attribute INIT_28 of inst : label is "C0001FE01FFFE00FF0000FFFF001440000000001FE00000000FF00FFFF007FFF";
    attribute INIT_29 of inst : label is "07FFFFF8008AFF0000FFFF00FFFF000000007F8000007F8000003FFFC0003FFF";
    attribute INIT_2A of inst : label is "807F80007FFF803FFFC03FFFC03FFFFFDFE01FFFE0001FEFFFFFFFF0000FFFF0";
    attribute INIT_2B of inst : label is "E01FFFE0000FFFF0000FFFF00FFFF7F807F8000007F807F803FC03FC01457FFF";
    attribute INIT_2C of inst : label is "FFFFF807F80003FFFFFFFFFFFC0001FFFFFE00A03FC03FC0003FC03FC01FFFFF";
    attribute INIT_2D of inst : label is "FFFC03FC01FFFFFE00FF000054001FFFE01FFFE01FE00FF0000FFFF00FF007FF";
    attribute INIT_2E of inst : label is "0000007F80007FA20FF0000FF00FFFF00FF00007FFFFFFF80003FFFFFFFC0003";
    attribute INIT_2F of inst : label is "07F80007F807F80003FC03FC03FC01FFFE00000001FE00000000FFFF0000FF00";
    attribute INIT_30 of inst : label is "03FFFC03FDFE0000000001FFFE00FFFF00007F80007F80000000003FC03FFFE0";
    attribute INIT_31 of inst : label is "4B4F1AAFBD9615A73611A78D8400FA79B7D844155B8C9D843752E89003FFFC00";
    attribute INIT_32 of inst : label is "31BD64A023095FFEF706EC4FED856BD051EDC4A394C25C8149A4A094024BA06E";
    attribute INIT_33 of inst : label is "4A5D9D422905D892D96020177262A05091A46BA2EA0050A49BB30E9E474E2A94";
    attribute INIT_34 of inst : label is "39983A52122AE9B1A44A0D0A41D2D6E45088F018409CD06C342D7717FF7B7117";
    attribute INIT_35 of inst : label is "E1B60180180184D05454557452F7BBA2948AD1B313B6D9C9D26CE48E6609ECE1";
    attribute INIT_36 of inst : label is "8E183E275C11334CAC6CD24B9B70514764B79E3860A607BDEF00F7BDE01EF7BD";
    attribute INIT_37 of inst : label is "5B99CC9DA2C0A12E888801AD8115372E993B4584DA2656366925CDB829A3B25B";
    attribute INIT_38 of inst : label is "6B19472924718AF252126718AAD6B75D000540CB884688390A2CB862B6045925";
    attribute INIT_39 of inst : label is "200840CA5084212942128421286528421294B58D6358D630842529421AC6B18C";
    attribute INIT_3A of inst : label is "358C631AC650842129410A5214852B29421284A0010042008194A10842120001";
    attribute INIT_3B of inst : label is "8431AC631AD6329421094A4200802008194A1084250C6358D6358CA5294A1096";
    attribute INIT_3C of inst : label is "8230A042815018D07110842A10AABFAAFEFACA50842129631AC631AC61084253";
    attribute INIT_3D of inst : label is "10A050350D468140A04429408506A10A0C6A140A506140A502810A88D28108C2";
    attribute INIT_3E of inst : label is "050210A84223408D2B41A20428140A5063450A04230A052234085062150846A1";
    attribute INIT_3F of inst : label is "518702C438CE118CE30E30906012C308CA18C251C210C25084A0B8A3F7F7D40A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "D142AD16C9192BCCCAA94D22A6933D8080222950381805451004046200200674";
    attribute INIT_01 of inst : label is "400000400000400004000040002101000100088A082082A028A3525630AAA032";
    attribute INIT_02 of inst : label is "0010000005EC4000000000000180006400040000000040000004010000404000";
    attribute INIT_03 of inst : label is "6B64C07F01FBDE02FDE02FDE0000000400002000000000000000000003800407";
    attribute INIT_04 of inst : label is "67DA0366A5F2361D8DA20000000000000000179B7168BA0BA9244CB2EEEDB6DB";
    attribute INIT_05 of inst : label is "9CA4A0C6A4B9453B1D6169AD0B19933195AB044DDB08A2B9D6F250D4A1A943DB";
    attribute INIT_06 of inst : label is "06805C815D0D832DA544D9B01D54448686991259290A59D7FEB90B39EF6C6C92";
    attribute INIT_07 of inst : label is "72D48FC8226D6C294AC926529CEF6CDB1949E4124295225F75C00005D0610840";
    attribute INIT_08 of inst : label is "7D2732A4F92E529FCA94E65324994A73BDBA4DB2576EF08A9D29249504E52629";
    attribute INIT_09 of inst : label is "A490292693FBF1F43DBBE148B492049592A5F87091DBB6368B6833DBB4130A45";
    attribute INIT_0A of inst : label is "9554555444CBA492480593526B2BEEF0FDDE5814B1B29F252B303FA1EDDF0A45";
    attribute INIT_0B of inst : label is "5007402CD9206841C891094D4AA80A82055AB9D2265D09E5DB96DDE177020F60";
    attribute INIT_0C of inst : label is "9D62A560A2F0146E68C86102AD2402589EED9DB4AD0DED2528421084217014A6";
    attribute INIT_0D of inst : label is "874A654A95C94A47BAB0B229452E5206352530872FE79C225A52432536092190";
    attribute INIT_0E of inst : label is "08112A5E1D18D295A4AF448DDC54555B64925ED92493B64924EC92493B2492C8";
    attribute INIT_0F of inst : label is "0F01E01C0380700E01C02A2109525269523469D3A74E893A2595DB90C183060C";
    attribute INIT_10 of inst : label is "AE5B37E735AC89AE6A96CD7354A28A22088A7406D80F01E03C0780F01E03C078";
    attribute INIT_11 of inst : label is "4D526B4D726B4D72D9AE6B96CD735CB66B9AA5B35CD72D9AE6A96CD7354B66B9";
    attribute INIT_12 of inst : label is "5031A6A935A6A935A6A93FCD3BD9135A6B9566B9AA4D69AA4D69AA5B35CD526B";
    attribute INIT_13 of inst : label is "D95DA9BEDB36ED6A3611B08D846421201B00D806C03603108216DB2AE871A528";
    attribute INIT_14 of inst : label is "CAB60700E11C2784DB6D4A684B49692F43D0BE40008A42A8240494A52A1B6DB6";
    attribute INIT_15 of inst : label is "202490A52B421623881C09856D956C2E136D956C2E13C26DB2AD81C2384F09B6";
    attribute INIT_16 of inst : label is "528A11484A2802764528A1149922909450480654AC8C00035224264D98AD8ADB";
    attribute INIT_17 of inst : label is "11A3288CCA4A94899AAA4BF52A51B2644CD5525F52A51E4C9105294E10A53308";
    attribute INIT_18 of inst : label is "EECCCC5555444408888000098CEBA125914633AD0D097A4FCA954ACB2ACA4846";
    attribute INIT_19 of inst : label is "3421292C134093A5BD71A04D024E93BBBBBBB3333333315555555111111110EE";
    attribute INIT_1A of inst : label is "4B36B1AD4AB40149B5567D59A09741940149B5567D49A0975D06C2936D631A05";
    attribute INIT_1B of inst : label is "F8000BFC00FF7FA000001FFFEFF00007FA0803FDFFFE007FFFA088822A22AA80";
    attribute INIT_1C of inst : label is "07F8280000000000000002803FC0000FF0000000280000FF7F80BFC01FE00007";
    attribute INIT_1D of inst : label is "8000000000000000002080001FE0000007F8080001FE0000007FFF8280000000";
    attribute INIT_1E of inst : label is "E00007F8A80000007F80801FE00002000000000000002A3FC0001FEFF0000002";
    attribute INIT_1F of inst : label is "007F8000003FFFFFFFC0001FE01FF2257555777E5BFC0000FF0000028000001F";
    attribute INIT_20 of inst : label is "80007F80003FFFFFFFDFFFFFFFFFE00FF00AEC01FFFFFE00FF00FFFFFFFF0000";
    attribute INIT_21 of inst : label is "D400FFFF00000000007F803FFFC000001FE0000FFFFBB800FFFFFFFFFF00FF7F";
    attribute INIT_22 of inst : label is "03FFAF00007FFFFF807F803FFFFFFFC0003FC0001FE01FEFF00FFFFFFFF007FF";
    attribute INIT_23 of inst : label is "F00FF00007FFFFFFF803FFFFFFFFFFFDFE01FFFFFD803FC000001FFFEFFFFFF0";
    attribute INIT_24 of inst : label is "FFFFFDFFFE01FFFFFFFEFF0000FFFFAF801FE0001FFFFFFFE0001FEFF0000FFF";
    attribute INIT_25 of inst : label is "FFFE00FFFF000000FFFF00007F800057CFFFFFFFF00007F807FFF807F803FFFF";
    attribute INIT_26 of inst : label is "FF00FF007FFFFF800000003FC03FFFE00007FFFFF803FFFC0003FC03FDFFFE01";
    attribute INIT_27 of inst : label is "007FFF80003FFFC03FD5F803FFFFFFFC03FFFC0001FE01FE01FFFE00FF00FFFF";
    attribute INIT_28 of inst : label is "07E01FFFE01FFFE0000FF00FFFFBE801FE01FE01FE00FFFF00FF00FFFF000000";
    attribute INIT_29 of inst : label is "F7F807FFFDDCFFFF00FFFFFF00FFFF007FFFFFFFFF807FFF803FFFFFFFFFFFC0";
    attribute INIT_2A of inst : label is "007FFFFF807FFFBFC0003FFFFFC0003FDFFFE01FFFFFFFEFF00FFFFFFFF00FFF";
    attribute INIT_2B of inst : label is "FFE01FFFE00FF000000FFFF00FF007FFF80007FFF80007FFF80003FFFEAE7F80";
    attribute INIT_2C of inst : label is "07F80007FFFFFBFFFC0003FFFFFFFDFE01FFFF55BFFFC0003FC0003FC0001FFF";
    attribute INIT_2D of inst : label is "000003FFFDFE000000FFFFFFFAC01FFFFFE000001FE00FFFF00FFFFFF007F800";
    attribute INIT_2E of inst : label is "00007F8000007FF74FFFF00FFFF00FFFF00007F807F807FFF803FFFC000003FC";
    attribute INIT_2F of inst : label is "07F80007FFF807FFFBFC03FFFC0001FFFFFE0001FE0001FFFE00FF000000FFFF";
    attribute INIT_30 of inst : label is "FC03FFFC01FFFFFE01FE01FFFE00FFFFFF7F80007F8000007F80003FFFC02BE0";
    attribute INIT_31 of inst : label is "4AAA491829A92355B927550E4990D5500024A77A90EABA488809819003FC0003";
    attribute INIT_32 of inst : label is "253D6FAD6B4AA210840903488A488007AD90348A20C270192C912082D9100383";
    attribute INIT_33 of inst : label is "1E4A80A67C4A0292DB3275681A4200000AF5AAE502A0D0A4DB200A965EAAE452";
    attribute INIT_34 of inst : label is "39993B5B1232E931FD4BC98A6CB6AC849BA2E1190A9CB9D86F12AA2508426228";
    attribute INIT_35 of inst : label is "65A61991991996902A2A2A806884240344CAD9B39324D989D26CE48F6749CCC9";
    attribute INIT_36 of inst : label is "8A504348650A4A200945F48289143DF6092596A9433419CE732339CE646739CE";
    attribute INIT_37 of inst : label is "FA3DC417EA48A92EB9C083F5770AF46EC82FD4B4931004A2FA41448A1EFB0492";
    attribute INIT_38 of inst : label is "0858480D494D0C00841494D04FAD2AA020BD286A381B9A1ACA2E206FD5DC7962";
    attribute INIT_39 of inst : label is "294A52C210842108084210842161084210840421084210B08421084202108421";
    attribute INIT_3A of inst : label is "A5294A529610842108425294A5294B0842108421294A5294A5842108421094A5";
    attribute INIT_3B of inst : label is "8425294A5294B0842108421294A5294A5842108421094A5294A52C2108421084";
    attribute INIT_3C of inst : label is "8894A2528B454A513544A568944110140445C2108421084A5294A52961084211";
    attribute INIT_3D of inst : label is "44AA55344D568944AA556B44A552A94A2568955AD12B55A512894A2A528B5AD2";
    attribute INIT_3E of inst : label is "2D12B5A256A955A52B45A22528B44A5129445A252B5A252A945A512AB54AD289";
    attribute INIT_3F of inst : label is "538733C4784E308C611E1190E410C308CA184A11C650C6108CB5C57480A2144A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "A5D03A5D58E006D50044219010E4E48A0080984B60401218633111111311315B";
    attribute INIT_01 of inst : label is "9FFFFE9FFFFE9FFFE9FFFE9FFFDEFA7FFEFFD0A00A80A8002A032305B455D40B";
    attribute INIT_02 of inst : label is "FFE4FFFFE813BFEDFFFF4FFFEC7FFF8DFFEDFFFF4FFE9FFD3FE9FA7FDB9B9BFE";
    attribute INIT_03 of inst : label is "9982822A08AE80100801008004FFFFE9FFFF6FFFFFE9FFFF6FFFF4FEDC7FF9B8";
    attribute INIT_04 of inst : label is "D1654298263C780E0E3800000000000000004D7613380E0889CFB34911124924";
    attribute INIT_05 of inst : label is "67531D083A8843692326C718260E6CC6460C0C18C6270EED0A59F983F347E63F";
    attribute INIT_06 of inst : label is "A74595115E944486183A3C6934458B1D0D066D86C6318608070630D04A508361";
    attribute INIT_07 of inst : label is "8D0B7535BD901BC63136D9084258C16CF63616DDBC61BB357F4000384404236A";
    attribute INIT_08 of inst : label is "99D8EC1B26D18C6A7167998CDB642109630CB6CD9C912200E1C5DB609718D9C6";
    attribute INIT_09 of inst : label is "96CBC6D0D9C283D67244A46F12D97B406C367156E72441C800CC8D2440CC2378";
    attribute INIT_0A of inst : label is "02222222332616C96DB6FC1D83CE71224E258646CE6C64D8D4C64EB392252378";
    attribute INIT_0B of inst : label is "8107A2CB3EA2F4A241632DB486EC250B176AC61C6D3FE6764E0DB2043D270922";
    attribute INIT_0C of inst : label is "619C31870C70E18767A884083ADBD9677583706B50E358D8C108421084FBCA11";
    attribute INIT_0D of inst : label is "72A51060CC44A13088320984308129718190961092304399A18B1FD0FE76DC67";
    attribute INIT_0E of inst : label is "64C8CB32D96B5EF7B6B372722233222DB6DB736DB6DCDB6DB636DB6D8DB6DB86";
    attribute INIT_0F of inst : label is "911222444889112224449918C4590BEDCB870E1C3870C5C31B40E1C3264C9932";
    attribute INIT_10 of inst : label is "0306E21CE0036619C1C1B0CE0628A0280A083A28A89112224448891122244488";
    attribute INIT_11 of inst : label is "38198638398638383619C0C1B0CE0E0D8670706C338383619C1C1B0CE0E0D867";
    attribute INIT_12 of inst : label is "604F1C0CC31C0CC31C0CE438E006CC31C0C1D8670330C70330C70306C3383986";
    attribute INIT_13 of inst : label is "86221FF904891081ED8F687B63DA1ED9F2CF947CB3E51AECC84DB6C3FF1E5AD9";
    attribute INIT_14 of inst : label is "B06A351B23646C8DB6D833997B6F65EE7B1EC1BBB639602D1A88421084C61861";
    attribute INIT_15 of inst : label is "10DB6F9182D131334C1C468DDB60D46A36DB60D46A3646DB6C1A8D46C8D91B6D";
    attribute INIT_16 of inst : label is "8801CE2320064B07B8801CE345DC46400FE04F074F7B39CB2C5A71B0F7027025";
    attribute INIT_17 of inst : label is "2118C67B31B16B76655721DC990CA99BB32AB90FC990C5336CF886304F10CC27";
    attribute INIT_18 of inst : label is "664444111100000888800076734E3391EE39CD39999C8700E0EA64F4D0F58080";
    attribute INIT_19 of inst : label is "DA50D6B0CDA2613A505CD1368980E19999999111111110444444400000000066";
    attribute INIT_1A of inst : label is "4EECC33070C88E24407261C9E0D864E88E24407661D9E0D861933C48840DCD42";
    attribute INIT_1B of inst : label is "07F8080000007FAABFC0000000000000000BFC0000000000002A02808A28A000";
    attribute INIT_1C of inst : label is "07F8280001FFFE00007FA83FC00000000FF000002BFC00007FAA000000000000";
    attribute INIT_1D of inst : label is "000001FFFE00FF7F802A3FC01FEFF00000000BFFFDFE00FF000000283FDFE000";
    attribute INIT_1E of inst : label is "0FF007F8ABFC0000002A001FE007F8000001FEFF7F802A80001FE000000007F8";
    attribute INIT_1F of inst : label is "0000007F803FFFFFFFFFFFC0001FEA80088082AA2BFC01FE007F80283FC00000";
    attribute INIT_20 of inst : label is "00007FFF803FFFFFC0001FFFFFE00FF0000105FE01FFFFFE0000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "A000FFFFFFFF007F807FFF80003FDFE01FFFE0000FF416FF00FFFFFFFFFF0000";
    attribute INIT_22 of inst : label is "F8000500007FFFFFFF80003FFFFFFFFFFFC01FE01FFFE000000FFFFFFFF007F8";
    attribute INIT_23 of inst : label is "FFF0000007FFFFFFFFF803FFFFFC00000001FE0020BFFFFFC01FFFE0000FF007";
    attribute INIT_24 of inst : label is "FC0000000001FFFFFE00000000FFFF441FE000001FFFFFFFFFFFE00000000FFF";
    attribute INIT_25 of inst : label is "0000FF000000FFFF0000007F80007FA20FFFFFFFFFF7F80007FFFFF803FC03FF";
    attribute INIT_26 of inst : label is "FFFF00007FFFFFFFFF80003FFFC011000007FFF8000000000003FFFC01FFFFFE";
    attribute INIT_27 of inst : label is "7F80003FC03FFFFFC00883FC03FFFFFFFC000001FE0001FFFE0000FF0000FFFF";
    attribute INIT_28 of inst : label is "00001FFFFFE00000000FFFF0000051FE0001FFFE00FF000000FFFF00007F8000";
    attribute INIT_29 of inst : label is "07FFF80002AA000000FFFFFFFF00007F80007FFFFFFF80003FC03FFFFFFFC000";
    attribute INIT_2A of inst : label is "007FFFFFFF80000000003FFFFFFFFFC00000001FFFFFE000000FFFFFFFFFF000";
    attribute INIT_2B of inst : label is "FFFFE0000FF00000000FFFFFF0000000000007FFFFFFF800000003FFFC400000";
    attribute INIT_2C of inst : label is "07FFFFF800000000000003FFFFFC000001FFFE88800000003FFFFFC01FE01FFF";
    attribute INIT_2D of inst : label is "FFFFFC00000001FE00FFFF00451FE01FFFFFFFFFE00FF000000FF00000000000";
    attribute INIT_2E of inst : label is "7FFF8000007F80002000000FFFFFF0000007F80007FFF80003FC0000000003FF";
    attribute INIT_2F of inst : label is "F8000007FFFFF800000003FFFFFFFC0000000001FFFFFE0000FF000000FF0000";
    attribute INIT_30 of inst : label is "FFFC00000000000001FFFE0000FFFFFFFF0000007FFFFFFF8000003FFFFFD107";
    attribute INIT_31 of inst : label is "364E44C9380B19270B1D2702C7499272092C62F91C88DAC75508A06BFC000003";
    attribute INIT_32 of inst : label is "3706705AD4B65318C626A2348EC6AE2157A8833E52A9B146D8F7E02D877C44A0";
    attribute INIT_33 of inst : label is "01A8E4098465406D24CC11D51182804266A36FBAA0219F122000465C064E531A";
    attribute INIT_34 of inst : label is "C3E2C665DDC8365E80743671830996C270EFC4DE30E79249A46962018C63E9D5";
    attribute INIT_35 of inst : label is "BA4BE6EE6EE6EB6FF5F5F7519718CA8C33312EFCDC5B7E6E6DBF1770F8B61F16";
    attribute INIT_36 of inst : label is "6599B06E20B361844D6576DB9932C3060DB6493664DBE6B5ADDCD6B5BB9AD6B5";
    attribute INIT_37 of inst : label is "560FF015A5A716C1466CE4AB01352C1FE02B4B6B2DC226B2BB6DCC99618306DB";
    attribute INIT_38 of inst : label is "109319006C219B91DE46C219BAF462D4205407860820D9EBF1C30632AC04C56D";
    attribute INIT_39 of inst : label is "42108498C6318C6310842108424C6318C631884210842126318C6318C4210842";
    attribute INIT_3A of inst : label is "0842108424C6318C631884210842126318C6318C4210842109318C6318C62109";
    attribute INIT_3B of inst : label is "31884210842126318C6318C4210842109318C6318C6210842108498C6318C631";
    attribute INIT_3C of inst : label is "3319CC6711898CE27998C67138445105140498C6318C6310842108424C6318C7";
    attribute INIT_3D of inst : label is "98C4E2388E231188C4663198CE27119CCE31188C627188CE67319C4CE3338CE3";
    attribute INIT_3E of inst : label is "C66339C4E73388C67199CC4633198CE671988CCE338C4E33398C6673188C6711";
    attribute INIT_3F of inst : label is "1BCFA8E2BD6338C6B1AF3ACC751AE3BC671C6B78E378E758D6208A80A828998C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "2490124958C002D8004424901240E808004018002000031C713333333311314F";
    attribute INIT_01 of inst : label is "4000004000004000040000400000010000000A000AAA00002AA92105A4408089";
    attribute INIT_02 of inst : label is "0002000004000000000020000000000400040000200040000004010000000000";
    attribute INIT_03 of inst : label is "1806401100450200102001020000000000002000000000002000000040000080";
    attribute INIT_04 of inst : label is "10000A1020202008082400000000000000004140306010000804A00020200000";
    attribute INIT_05 of inst : label is "3050100022180008070004002400008441020C10482405060C7910222004402F";
    attribute INIT_06 of inst : label is "060215115C140804006058AB00000C3000007002000000085208000410A00000";
    attribute INIT_07 of inst : label is "140C454590202300000002010040136CC00096CE30019A2A80155560C0042328";
    attribute INIT_08 of inst : label is "21008000680200028186020000080401004D92CC0D020200810D0001B6200300";
    attribute INIT_09 of inst : label is "924B000249822392740824241249600080126346834081100104814081812120";
    attribute INIT_0A of inst : label is "133333332200B2CB6492E010020682025040024248800D0000166C93A0412120";
    attribute INIT_0B of inst : label is "0407010878AAE08441836D848244250912224810043FC2F44000040431250A00";
    attribute INIT_0C of inst : label is "811011040460808742280408224BC9444404408C41C440000108421084FB8002";
    attribute INIT_0D of inst : label is "628400408C0883A084601110201021E30100000002208110000A0F40FE725C87";
    attribute INIT_0E of inst : label is "448C99227339CE73939322F333222224924931249248492492124924C4924984";
    attribute INIT_0F of inst : label is "0300600C0180300600C0199CE4C919E5CB162C58B162E58B9F08C18224489122";
    attribute INIT_10 of inst : label is "0608829180C50403008220180C2A002AA00AB010380300600C0180300600C018";
    attribute INIT_11 of inst : label is "2031002011002010440301822018041100C0608806010440301822018041100C";
    attribute INIT_12 of inst : label is "302C10188010088010088DA0890A08010181100C022004022004060880601100";
    attribute INIT_13 of inst : label is "08041FFA08002003001800C026013001820C106093049A0048400001FE386319";
    attribute INIT_14 of inst : label is "000E0700600C01800000011B632C658C63188001423920251002421086C82082";
    attribute INIT_15 of inst : label is "18000190829131124418478100001C0E0000001C0E00C000000381C018030000";
    attribute INIT_16 of inst : label is "011088020442DA04201108800D10040887C0DE040851295A3062520444044047";
    attribute INIT_17 of inst : label is "0109022040018C40855404CA1405A002042AA026A140440044601000CC020166";
    attribute INIT_18 of inst : label is "EECCCC555544442AAAA22240C004161108230010B0B08600C080408110840084";
    attribute INIT_19 of inst : label is "100218A0C101012254408084040083BBBBBBB3333333315555555111111110EE";
    attribute INIT_1A of inst : label is "48808020408C88008056C15C804920AC88008052C14C80492482B001042E080B";
    attribute INIT_1B of inst : label is "F8000801FE00002ABFC01FE00FF007F802A3FC01FE00007F80000A8A28228200";
    attribute INIT_1C of inst : label is "F0002BFC01FE00FF00002ABFC01FE00FF007F8028001FEFF00003FC01FE00007";
    attribute INIT_1D of inst : label is "03FC01FE00FF007F802ABFC0000FF007F802A3FC000000FF007F8000001FE00F";
    attribute INIT_1E of inst : label is "0FF00000A8000000002ABFC0000002A801FE00FF7F80003FC01FE00FF007F800";
    attribute INIT_1F of inst : label is "007FFF803FC000000000001FFFE002A8AA22A8088801FE00FF7F80003FC01FE0";
    attribute INIT_20 of inst : label is "FFFF80003FC00000001FE00000000FFFFFF151FFFE000000FFFF000000000000";
    attribute INIT_21 of inst : label is "00FF00000000007FFF80003FFFC01FFFE000000FF00542FFFF0000000000007F";
    attribute INIT_22 of inst : label is "03FC057FFF80000000003FC00000000000001FFFE000000FFFF000000007F802";
    attribute INIT_23 of inst : label is "000007FFF80000000003FC0000000001FFFE00002A3FC000001FE0000FF00000";
    attribute INIT_24 of inst : label is "000001FFFFFE00000000FFFFFF0000055FFFFFFFE00000000000000FFFFFF000";
    attribute INIT_25 of inst : label is "0000FFFFFFFF00000000007FFFFF8002A00000000007FFFFF800000003FFFC00";
    attribute INIT_26 of inst : label is "0000007F80000000003FFFC000000157FFF800000003FFFFFFFC000000000000";
    attribute INIT_27 of inst : label is "8000003FFFC000000000ABFFFC00000000000001FFFFFE00000000FFFFFF0000";
    attribute INIT_28 of inst : label is "1FFFE0000000000FFFF00000000455FFFFFE000000FFFFFFFF000000007FFFFF";
    attribute INIT_29 of inst : label is "00000000020AFFFFFF0000000000007FFFFF8000000000003FFFC00000000000";
    attribute INIT_2A of inst : label is "FF8000000000003FFFFFC000000000001FFFFFE00000000FFFF0000000000000";
    attribute INIT_2B of inst : label is "000000000FFFFFFFFFF00000000007FFFFFFF8000000000003FFFC0000507FFF";
    attribute INIT_2C of inst : label is "F8000000000003FFFFFFFC00000001FFFE00000A3FFFFFFFC00000001FFFE000";
    attribute INIT_2D of inst : label is "0000000001FFFE00FF000000055FFFE000000000000FFFFFFFF000000007FFFF";
    attribute INIT_2E of inst : label is "7FFFFFFFFF8000282FFFFFF0000000000007FFFFF800000003FFFFFFFFFFFC00";
    attribute INIT_2F of inst : label is "FFFFFFF80000000003FFFC00000001FFFFFFFFFE0000000000FFFFFFFF000000";
    attribute INIT_30 of inst : label is "0000000001FFFFFFFE00000000FF0000007FFFFF80000000003FFFC000001407";
    attribute INIT_31 of inst : label is "864442A9100B15220B112202C549D220012C50E908089AC4002C0403FFFFFFFC";
    attribute INIT_32 of inst : label is "0404404318C651084204068406C4AE0307804838C114300858F7E005877C0286";
    attribute INIT_33 of inst : label is "382000D55C5009049250310024280002D0006F0005201C00410044490A444A92";
    attribute INIT_34 of inst : label is "03830E65D11036C8044042C02401924170EFC25000838140A22960008421E140";
    attribute INIT_35 of inst : label is "024B800800800B6E202022022400001120412E70505938286C9C1440E0C01C18";
    attribute INIT_36 of inst : label is "24C8B026203121C44521E2493060C3040492CB9722D980000010000002000000";
    attribute INIT_37 of inst : label is "161F801580141801206CBA0302102C3CC02B000B6CE22290F124983061820249";
    attribute INIT_38 of inst : label is "4210190024248B91DE424248B0700080A0D022061010108BC10303880C084540";
    attribute INIT_39 of inst : label is "2942108000000000425084A508400000000021094A1084220004000012942129";
    attribute INIT_3A of inst : label is "252842508400000400021294A109420000020085094A129421000001004084A1";
    attribute INIT_3B of inst : label is "10A12942128420000000001084A508421000000084284A1094A1080000000014";
    attribute INIT_3C of inst : label is "A890AA42215448553000A42A90EEEEAFEAFE8000000000425084A50840000043";
    attribute INIT_3D of inst : label is "448855310C42A910885123548442A90AA4221548D52110AC42A9088056214842";
    attribute INIT_3E of inst : label is "A4429088520154846B10AAA4221548D521110AA42908856015484428910A4221";
    attribute INIT_3F of inst : label is "308710C438C6118C230E10886030C7184238C230C611C231843D5D55FFD5710A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
