-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_3H is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_3H is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_3H_0 : RAMB16_S2
	generic map (
		INIT_00 => x"042054760AF14FFFFFFFFFFFFFFFD445E649FFFFFFFFFF7DFDEEFFDFF52FFFCF",
		INIT_01 => x"5937A59342555454554B7CE81450C17BE9E33C88DF35423D82C2F135D3413C81",
		INIT_02 => x"925235392948D7111176496150508DE8A416A1CC895751552DFCE8174A464276",
		INIT_03 => x"B445E69C65E69368919091A35D41C65F9A48DC6559279A7195649E698D04445D",
		INIT_04 => x"FF3FB7BB33B7359EC28E6D8FBE09D02F0FF64CCCFD108D82EE36B445D9242350",
		INIT_05 => x"1C45E70709D445B59249E79A48D48DD71979B76496F1951161CE8D649F47B773",
		INIT_06 => x"7F6358D63564DE1D54D6561BDD5F75937D6561BDF97559376495117E9D776707",
		INIT_07 => x"04755116DF9A7197E6DBF9A54BE94155CC8954763519095DE6564D445D925746",
		INIT_08 => x"64DF3F9B7CF64DF3F9B7CF64D445D925F8DCFD5607751CE3811555F1D1C9E772",
		INIT_09 => x"748D2715E1422492C492C492C41415055F7792561D4957B15154458D64DFB60F",
		INIT_0A => x"505E2370BFD9B5115D05C236D25C2370BD977195D05C236DA5C237E64D445741",
		INIT_0B => x"4400000000002021FFFFFFFFFFFF9292D9999F5F5073F25E69E79C15586D5C49",
		INIT_0C => x"F2F0200F200200F2F10020211000F1F10F0F210000F2F0200F2F8A8A8A8A8A88",
		INIT_0D => x"6DCF8ACCAAA75B38BAF428EA6684F200CDEE8EA0000F000000F000002F2F0000",
		INIT_0E => x"0DFFF074FC81EC4FC40DFFD07CF801EFAE4E48451451444361CC0440C30C3003",
		INIT_0F => x"C00CCFFF40EC043C003FE3771DB0C83F4F609090365CFA08080365CF2E5C5FCC",
		INIT_10 => x"2ECCFC00C3FC0F8FF43EC00DEC6C6C6C6C6C6B8C361CE1B1B1B1B1B1ACC0361C",
		INIT_11 => x"C3F0C1CFC20F3F0C3CD400FB51CC5C80EC624E31730BB78C5CC2EDC604C7F000",
		INIT_12 => x"AAC6C6C6C6C67939393936036D0DA86C6C6C6C6C64E4E4E4E4E603690DB69960",
		INIT_13 => x"2A4E75B7D00C79D6DF4031E75BDBD0C79C6DF431DD4144C68F5C41E68F5CC1ED",
		INIT_14 => x"33F00FB03BF303A9F774A0C719ED80F50200E7F508035E4A0C0FC01EC0FC40EE",
		INIT_15 => x"0C330C03E1E30C30C3003E1E0ACC003C103B01FF080C0CFC03EE4ACC17FC2030",
		INIT_16 => x"CF2C63104100E0321CC003212C31C2334480F3CB18C41040380C87333BDB1F0C",
		INIT_17 => x"50420321CC303723101034744C4E18F2C045141080C873000C84B0C708CD1203",
		INIT_18 => x"0000BC00C4C404C4BC8C68480000C0C80C8730C0DC8C4041D1D1313863CB0114",
		INIT_19 => x"0F434F03254A8F70B0F0F2F2F0C0C0C951A2CC2030307878F0F03254DF28501C",
		INIT_1A => x"080C8626BAC7100C861E892043218DF79D6138B3083012300C953E1C8283C7CB",
		INIT_1B => x"3A1E1E0020F0083C3C6AF8EBAE78EFAEF4E74C354CFFA961DA22130CB62EB9B7",
		INIT_1C => x"1E007140E3103D010B2048060F3383C3C07002CC02C0201A00E0088DC0CCE87B",
		INIT_1D => x"CCE0F1183C3CABFCFBEF7CFFEFF8F78C35408307818CC87C6009CC8828791A1E",
		INIT_1E => x"00E7007C001B7008C2CBC0B2F2F07CC3DC0EC4302B002008B1D0446CBD1B2F2F",
		INIT_1F => x"20F0F3E3C32CF1C30CF0F72F70C50313058188886C700A00842435190D0D0431",
		INIT_20 => x"3D042C8120183CCE0F0F01C00B300B008068038022370333A1ECE878780083C0",
		INIT_21 => x"E7D76D34D77D35D74D70D4020307818CC87C6009CC8828791A1E1E007140E310",
		INIT_22 => x"95C42130EDC0C8C3072108043410DDCC4320C007001C20400DE1D30D101DC300",
		INIT_23 => x"8BBBD62901125C122450641655AA882BEA9559219247472879B7D34D30C53DEE",
		INIT_24 => x"80000820082A81444989AF8EB8EB0C5082D36820A0BB6866002420A2282AEB58",
		INIT_25 => x"A06C198122450CE08CE0A0649498BA39E39E30C5082208820A8190601A066048",
		INIT_26 => x"E45B41224506016A22006C78425A990128DB3EF3FF30D84082209C71EC1906C1",
		INIT_27 => x"0CB0E0F3CF0D533DA674483A2208820A3AC981276D46840A28E9E386CB8E9E36",
		INIT_28 => x"E40A1759D19020E7CF9F3B00A4A279A82B2A0A0A886ACD561D561646763C4714",
		INIT_29 => x"2F5A0A05ECAA8297E6A9F9AA44AA8297E6A9F9AA4E1C5F11D31C71CF0D9400DC",
		INIT_2A => x"810800802A8A0AA885545AA166A8692A69354C576D74D34C3542524A94282819",
		INIT_2B => x"81825815902A9E0AA886A886A186AC2E82A69B58C576D76DB6C3254033382680",
		INIT_2C => x"30F790D54A20BDCE002390D47600BDCE002390D636D0BDCE592BAA9A00362926",
		INIT_2D => x"2368003DCFEF78EFEE683802F4A0D6392F7380086C35002C7380086C3500B1CE",
		INIT_2E => x"0500F73C8DF000F73CBC6F02003DCF2328003DCF200A3100F73CBC6F02003DCF",
		INIT_2F => x"3838C2378F0C9738CC84C4BCC404C414400C4C0440C404C000C8731C2F743CB2",
		INIT_30 => x"904437B3301C070D734DA344383A6CC9112C079C00C87380F42358D230325CE0",
		INIT_31 => x"E70607602715B4FE7060404C000D0340D73880823213DBB1F904D81F913DBB1F",
		INIT_32 => x"0701C35CE2C2CDCC836307E410A0B29836307E411C2300304C1035CE2C3F5B4F",
		INIT_33 => x"A281286417E3381361B4AA13227080C87396C9E2A5438808A04528A0510DECCC",
		INIT_34 => x"A5628A168BA9639A14321CAA8B466155844CBC2C814A116C83CA0EC321C5ACA4",
		INIT_35 => x"CD604C1C2D6826CAB2A0DB0E62ECEF3B4D80E626CEF3B4280E622B6D28E4CA4A",
		INIT_36 => x"CFFFF7EF70C872A3D439088601A3BCE01886011693D18C6018D3884631804325",
		INIT_37 => x"CC9C298D2C2AE3620A234A2332314B4F271605F509C698D2D3AE3670A63762FF",
		INIT_38 => x"5F4631846D20084631847FD4228061112088601844325C2A81880283C8C582DF",
		INIT_39 => x"C0325C38D284810F9706AC645208A262266E9950A0A2A989A266E990C97028C4",
		INIT_3A => x"1C6AE1B04321CDE55C7DA45816A8681AC691AC681E7B4E91AC6810C8702239CD",
		INIT_3B => x"16EC0F51EEC0F61E7FFC55D40C871A11A47433ACF40321C4A6619D8888236032",
		INIT_3C => x"9003BAEE4003D48ABA9B6A626503D48A39B86643D4E38A1807A975A18DC810C6",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8ABEBFB9A505664354886298",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_3H_1 : RAMB16_S2
	generic map (
		INIT_00 => x"00241E800980AFFFFFFFFFFFFFFFEDF73DFFFFFFFFFFFF9CFE13FFEBFA1DFFC4",
		INIT_01 => x"C30F433CC1ECDDE9EA8772FDB03640CDD0DCB84C67338390B9B9806C73E0A050",
		INIT_02 => x"7BD92E0707ACB3DD75E5DFA0B005CB00340C7880461EA7AA1D02FF83C9CDCDC1",
		INIT_03 => x"F5D7DFF5D75DF1D4F2727512E0C7DF7B7FC4B5D7A7BD77C71E5DF1CF4B479E7A",
		INIT_04 => x"84C40C44888C94CD6324D38AA584BAB48EE3EAAABD06CB4FD52CCDF7B7FC92E0",
		INIT_05 => x"02C94D028369E72D77E77D77ECB44B0C71C30F1CF337DD75E3B957DFFF4344C4",
		INIT_06 => x"D7B2ECB92ECF3E70E09E7A7000D9FB3CF0E7A7008B43B3CFDFF871DD0E1F8D02",
		INIT_07 => x"01E5975CB873C71FCF32C73E876F881E804471412E37378713ECF3DF7F7FE1C3",
		INIT_08 => x"4D3DB830F668E3DB934F664D3DF7F7FCC4B6EE000AA82AB8807560B30A036EA3",
		INIT_09 => x"26CB383B3EC3197301730173022C0B0035F1F5EF04D77440C0EDF74B8E3C9F26",
		INIT_0A => x"B22892D0554F9D75DF009B2D7BCA92D354F9C71DF02AB2D7BEA92D13E71C77C0",
		INIT_0B => x"0000000020321100FFFFFFFFFFFFE7A35C6D6FB288EEE5B5DF3E340B6CD7BE0F",
		INIT_0C => x"F0F0302F000001F0F01020200000F0F00F3F000102F0F0202F0F556677445560",
		INIT_0D => x"200DA64CFA8FA9B9571EC48BA84859B864764640000F100300F100003F0F0003",
		INIT_0E => x"0EFFE078FC01FC8FC40EFFE07CFC01FD544D0A0492492402200E0A0451451402",
		INIT_0F => x"EA84CFFF40FC043C003B6993201450B44D0747482240D0747482240D944CBFC4",
		INIT_10 => x"2FC8FF00C3FC030FF40FEEA4C80156A801568A9822C0C0055AA0055A889022C0",
		INIT_11 => x"C3F001CFC0033F000CFC103F400CFC00FE1B4D33F007C74CFC01F1E594CBF000",
		INIT_12 => x"80156A80156A95402A954002200EC00156A80156AA5500AA550002200E0828B0",
		INIT_13 => x"184D402A0B0A3644006C28D4022200A364400428E59628480FFC42F80FFC02FE",
		INIT_14 => x"B3F10BF03FFC03D2142A154681E0B0C12120831684820E694C0FC42FC0FC40FE",
		INIT_15 => x"141514022CC14514514022CEE84C023C103F01FF000C2CFC42FEAA4C27FC0030",
		INIT_16 => x"79CB4DECB2D3542200ECE605C45E7422AB339E72D37B2CB4D508803D6C92C80C",
		INIT_17 => x"9CB502200EDE1A0E61D72A957BB4D39CB779E72D408803B398171179D08AACCE",
		INIT_18 => x"E3432B73BB77777B2B3B43734373577508803B786839875DAA55EED34E72DDDB",
		INIT_19 => x"1995550A240E1997545454646545428903C449D1515151515554A240F4E3CC0E",
		INIT_1A => x"8708A0005855A708A0044A0642280F8C38D0011274989899288034551D119951",
		INIT_1B => x"E44444331514C54545F34F38F34F34F34F38F0A40C0D38F001205908900C595A",
		INIT_1C => x"44669E9E92A51A7A86069765516E545456A21449E1A147945E5579468BBB9112",
		INIT_1D => x"775192E46464E30E34E30E30E30E34E0A406227A7A665787879565725112E444",
		INIT_1E => x"5E5995955DA5A257A199AE666666565665E56967861E5078556B775999D66666",
		INIT_1F => x"15151743040043040040340342801AA579795217A7A784657A1999D666666A5E",
		INIT_20 => x"1A7A191A5D9545B951515A88512786851E517955E51A2EEE444B911110CC5453",
		INIT_21 => x"020420400430430000028018867A7A665787879565725112E44444669E9E92A5",
		INIT_22 => x"00418596965B30B96A0EE1B32AA6A68A9A07B96A215547B86A456EC56DEA4DE0",
		INIT_23 => x"B9956A26D21564A5D7575A245A0117096816A65E6A555544100100100080300C",
		INIT_24 => x"4C1DD75DD754797775B00010830808017E5D434D4E959AA9C2E840041B4855A2",
		INIT_25 => x"6E5796795DBA775D775D6D5B5B6B30000820808017E4D0B2C9355E5754C55E57",
		INIT_26 => x"5665495D757522468509559A5A9122094400430C30C088017E2CA79E5756E575",
		INIT_27 => x"518501C71C0903510604145922C8B2C856615929966A48912266491551244499",
		INIT_28 => x"65BA84044446EA111044446E92A05113A584E92117802155E155E56544701C80",
		INIT_29 => x"5055AA00116AA954029A0098416AA954029A0098547010871071C71C08901B96",
		INIT_2A => x"48A7AA66EAA5EA9979566A9E5AA7A6A6610462104104104024065254002AA804",
		INIT_2B => x"796A579556E551E5557AAA801E8044664844184521C71C6186022406E088567A",
		INIT_2C => x"D7695192521CA40CC7026192966CA40CC74261912A6CA40D9750410406EAAA51",
		INIT_2D => x"E2816C240D175541841C335D5541902A290331C15460FF281331C15460FCA04C",
		INIT_2E => x"55B0903F8AA0B0903F969A21EC240FE2016C240FE66195B0903F965A21EC240F",
		INIT_2F => x"E06785E97928A03B7B3777277B3777277377B74BB77B3B534288039244143F94",
		INIT_30 => x"6981995DD525490A03820A2C3B514A4529552965828803B7955E67A1E0A280ED",
		INIT_31 => x"9A491955D5665999A4900951DD164590A037474C2C556556669B555555565566",
		INIT_32 => x"49524280DD5D7A78155455555D11150155455555060233158560280DD5D66599",
		INIT_33 => x"0059C094A6569559855A04590558408A03B61A24A2C374740565440550665775",
		INIT_34 => x"5554455506535265342200A106B9AEA94A45665825815A9825846542280B184B",
		INIT_35 => x"0FDD79E3492C2CB12C43AD0A020B9AE6B5D0A028B56D574C0A024696C09A7054",
		INIT_36 => x"82492882808802C95462861595426A9856159594219A695854A97695A5614220",
		INIT_37 => x"7769167158459C50551C54CEED26B695D955DA55555957156655C5A459C64D24",
		INIT_38 => x"A5659569555596559569695548655959486159565422005475510D06B49A75A5",
		INIT_39 => x"B02280E356141D0BA03856555450055155555555001545555555555088034696",
		INIT_3A => x"80D185614A280FDC71D30F343C52545595655A549996A5695A549088034C2A86",
		INIT_3B => x"30CC28030CC28034AAABAAAB28A030AA6A86D96646CA280F1659917596645CA2",
		INIT_3C => x"57B565595ECA40D1645685915A0A40F19596564A40FCF34D0F15A945565452A0",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF16829515A0A544A00D19164",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_3H_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0A30C8478C064FFFFFFFFFFFFFFFC34DB249FFFFFFFFFF92FC99FFC9F114FFCC",
		INIT_01 => x"5D7508D343466C082A8A98FC83B2C2ED0EE0B140E42B3731E4380610C13BC8C0",
		INIT_02 => x"9A59040D0D24103DD76659245344C11D702516D8F1AE65AA2AA8FF60034B4B43",
		INIT_03 => x"F75DA6975D249368D0D0D330410F34D8924C134D4514924D35145249412FB6DA",
		INIT_04 => x"40CCC840C84028E2BF934DD4C02013318883733310E541232004834D8925805C",
		INIT_05 => x"7317DB0A36C34D211455549248128111D74D3565932DB5D7753004A6942B8C88",
		INIT_06 => x"432048120434D4D00234D0DED02370D3500D0DEE84800D352491D7502C371B0A",
		INIT_07 => x"08230D3488925D7534D05964450D45A4D8E298CB042D2D0D234B6D34D4924373",
		INIT_08 => x"34D490D352434D480D352075D34D49240C12CCC7BEA4D30BC204CCAB4432EAA7",
		INIT_09 => x"0AC1034EB397408008843880295C551493ECF31753CC900ACE434D41B6D6B768",
		INIT_0A => x"5061984F802D3CF3C0253B84F7609C4C83D3CF3C0342BC4FB50904234F3CF001",
		INIT_0B => x"0000203211000000FFFFFFFFFFFF688DDF33659E0D4CC05249366C2503CF5F4D",
		INIT_0C => x"F0F0100F000381F0F0100C000303F0F00F3F000100F0F0000F0F210321103210",
		INIT_0D => x"333C430C50146640545303013230430131303334203F040302F000201F0F0303",
		INIT_0E => x"23FFC00CFC403CCFF023FFC00CFC403C800CC8CA540FE883333CC8CA540FE883",
		INIT_0F => x"C800CFFD013C153C105F2043632A51F00CF0102C7333C70102C7333C810CDFF0",
		INIT_10 => x"03CCFF8233FE00CFF803CC10CC00000155554688F333C00000055555468CF333",
		INIT_11 => x"CBF0002FC000BF0002D4000F33385E013C430F317400CFCC5C0033C810CFF080",
		INIT_12 => x"32AAAABFFFFFFFFFEAAAA88B333C3000000155555555550000000B333C400000",
		INIT_13 => x"400CA215201CF288A88073CA211121CF288A8873C8100301CF5E0030CF5E003C",
		INIT_14 => x"3FF001F07FFC01F22A95144733CC00CCC873CF2232CF3CC20C0FC003C0FC013C",
		INIT_15 => x"AB95A8C333CEA540FE88333C810C273C009F00FF00044FFC007CC10C03FC0091",
		INIT_16 => x"CF0C0330C30000B333C10455155145440044000414004105112CCCF30820410C",
		INIT_17 => x"F0C00B333C00405045144000000000010000004112CCCF000C00000000CFF003",
		INIT_18 => x"08A89488444444449484A888A888A8822CCCF0C0FC0CC000FFFF333CF3C3333C",
		INIT_19 => x"0CC0000B3333C00000000000001012CCCCB11004040404040404B333C420C10C",
		INIT_1A => x"203CCCD31115103CCCD310544F333C0304005C89021212122CCCC3000000CCC0",
		INIT_1B => x"0111114444451111112CB3CB3C73C73CF1CB1CB33D400C206C45513CCCDB1115",
		INIT_1C => x"11C44040491C400010543044444011111C047110040710014005011010000444",
		INIT_1D => x"0004040101013CF0CF0CB0CB0C32CF2CB33C4401011470101011470444440111",
		INIT_1E => x"40451C000000043004000000000C003000000300004005010000000000000000",
		INIT_1F => x"00000037D74D76D77D75CF4CF2CCF0000101147000001147004000000000C040",
		INIT_20 => x"0F0C0003C00000CC000033C0C030030C00000300003F0333000CC00000000000",
		INIT_21 => x"76D74DF6D77DF6D36D32CCF0030000003000000003000000000000C00000040C",
		INIT_22 => x"41032A2844708A41C5A10B08951C556471A842C58B222002C555512551156109",
		INIT_23 => x"C0FFFF330300003C000000400054700FFC0000C0000000004DB4DB7DB3CCF618",
		INIT_24 => x"000330C330F303CCC304D37D76D73CCF0000000000000000100000000C0C0000",
		INIT_25 => x"E0F83E03C0CF08830883E0F838206DF6D35D33CCF00000C30FC3F0FC3F1FC0F0",
		INIT_26 => x"545151C0450445511C51444471544451516DF5DF4DF3CCCF0030FCF3F83E0F83",
		INIT_27 => x"5DB5CDB6D33CCF41451831548411041151451140000011144451515444462514",
		INIT_28 => x"47001551111C0044451111C0040555440011004470000000000000001B6CDF33",
		INIT_29 => x"C55555AA8B15555554355500CF157BBBAA79EA84D34CD736D36D34DB3CCCF014",
		INIT_2A => x"1100000C0000000300000000000000005D334CDB7DB4D34CF33C547155400151",
		INIT_2B => x"000000000C00000003000015401511001115DF34CD76D77DF7CF333C0511C000",
		INIT_2C => x"30FF33CC0000733C000333CC0000733C105403CC4000733DC51061060C0000C0",
		INIT_2D => x"041540F33DC51071441830C0FF33CC331CCF082A88F3001CCF041544F300733C",
		INIT_2E => x"5503CCF0255A03CCF03CCF0000F33C030000F33C00030303CCF000004400F33C",
		INIT_2F => x"00300000002CCCF00044444000444440044444500444845412CCCF6106143015",
		INIT_30 => x"144C00000000003CCF7147143018A461918A862A22CCCF003CC0F03000B333C0",
		INIT_31 => x"CF0C0FCC0F3F3CFCF0C0C000000C0303CCF02022915111511144511115111511",
		INIT_32 => x"33CCCF33C04045414445444511444454445444513C0300330CC0F33C0C3FF3CF",
		INIT_33 => x"551115010000000000000000000003CCCF41C51441C30202AA8AA2AAA3CFFCCF",
		INIT_34 => x"C8CA2C8CA1C8C91C8CF3334C500000000000300C00C003CC03C00CCF3337C110",
		INIT_35 => x"3D071441861C13000000F33CCDF0CC33CF33CCD70CC33CF33CCD71442A444AA2",
		INIT_36 => x"7D77D36D33CCCDF155441C4F131400313C4F13154400C0F131000C0F03C4CF33",
		INIT_37 => x"00007003C11C00C51C40F11000400000000030000003003C00C00C01C00DB4D7",
		INIT_38 => x"000303C0C0000C0F03C0C00000C0F03000C0F03C0CF333F10314505001000C00",
		INIT_39 => x"8CF3335CFCFFF33FCCD3C8CAAAAAA8B08C8B23AAAA8B2322C8C8B233CCCDBC0C",
		INIT_3A => x"336F13C4CB333DC71841871813C8F23C4F13C4F234514713C4F233CCCDF3E2BA",
		INIT_3B => x"DF332CCDB222CCD3114415102CCCDB11C44C11C44C0B3337C47113011C44C0B3",
		INIT_3C => x"30000C00C00F334F01301C04C04F336F030C0C0F33D0618407F00003C00032CC",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4F169513C5A544CF336C0701",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_3H_3 : RAMB16_S2
	generic map (
		INIT_00 => x"41041CD843D8CFFFFFFFFFFFFFFFF1C711C7FFFFFFFFFFFFFF11FFFFFC06FFC7",
		INIT_01 => x"C71F0071E0CFFD414001F3F5063090C7C8701CC07F2003E632F1D82C32F24000",
		INIT_02 => x"71C13F030304F3E471C1C7F330074F620D0C33C000FF05000703F633C0C0D0C0",
		INIT_03 => x"F1C71C71C71C71FC703030D3F3F91C7071F4F1C7071C71C71C1C71C78F091C70",
		INIT_04 => x"8844444400003CC30F81C7C33004F0342331CCCCFC8CCF03373CB1C7071C13D2",
		INIT_05 => x"F3D71E0307B1C73C71C71C71F4F04F3C71C71F1C73C71C71F0CC031C7F31C888",
		INIT_06 => x"DBE3FCFF3F1C7C33F00C3C3473F1FC71F3C3C347C3CFC71F1C7C71FC0F1FDE03",
		INIT_07 => x"017FC71CFC71C71F1C75C71F018700FFC003FC3F3F0343C731F1C71C7C71F1E1",
		INIT_08 => x"1C7C1C71F071C7C1C71F071C71C7C71CF8F07FFF27300CC2405FFFF000079F30",
		INIT_09 => x"F04F0F0711E00CF860F050F0530C0323F1C873CF41CFFC14D8F1C7CF1C7C1D07",
		INIT_0A => x"323C17D8EA971C71CB13C17C75FC13D8E871C71CB03C13C71FC13D31C71C72C0",
		INIT_0B => x"2032110000000000FFFFFFFFFFFF76676688AA88FC333031C71F7803F1C73D07",
		INIT_0C => x"F0F0080F080040F0F0080C000383F0F02F0F000080F0F0080F0F222111110000",
		INIT_0D => x"333C030C03212311303023003230222133223034282F040081F040180F0F0280",
		INIT_0E => x"03FFC00CFC003ECFF003FFC00CFC003C410E64E555500207333E64E555500207",
		INIT_0F => x"C000EFFF003E003C000F30C3939559F30CB8989C3333CB8989C3333C820EFFF0",
		INIT_10 => x"03ECFF0033FC00CFF003C410E1555555555565643333E5555555555565643333",
		INIT_11 => x"EFF0003FC000FF0003FC000F933CFF003CC20FB3FC00CFECFF0033C820EFF000",
		INIT_12 => x"795555555555555555555643333C39555555555555555555555643333C820400",
		INIT_13 => x"000E5995980CF966566033E5999990CF96656433CC30C202EFFF0032EFFF003C",
		INIT_14 => x"3FFC00F23FFC08F99555964333C410E66670CF9999C33C000E0FF003E0FF003C",
		INIT_15 => x"0055564733E555550020733CC30E033C000F84FF10100FFF003C820E03FC4000",
		INIT_16 => x"001050010414643333E12555155145555444514514445145190CCCF00C20400E",
		INIT_17 => x"010643333E12555155145555444514514445145190CCCF849154554515100110",
		INIT_18 => x"200000000000000000000000000000080CCCF809014114510000000000040000",
		INIT_19 => x"622666433332E65899999999999990CCCCB996266666666666643333C030820E",
		INIT_1A => x"980CCCC79995980CCCCB995643333C8104103E20888888880CCCCF9962662226",
		INIT_1B => x"1999994466651999992CB1C70CB1C70C33C33C333CC308200E20080CCCCB9995",
		INIT_1C => x"99E66262659E658999567866665199999E567996266798996265899558446665",
		INIT_1D => x"4466651999992CB2C71CB2C71C73C33C333E6589899678989899678666651999",
		INIT_1E => x"62659E666199567866665199999E567996266798996265899558446665199999",
		INIT_1F => x"666664F2CB2C72CB1C71CF1CF0CCF9998989967898989967866665199999E662",
		INIT_20 => x"60826558E199990266667819E648989E62658896264060009990266665119994",
		INIT_21 => x"F1C71C31C70C30C30C30CCF9988989967898989967866665199999E66262659E",
		INIT_22 => x"1083808222380008E0002380008E0002380008E023888888E000000000000020",
		INIT_23 => x"090000482456658E2458665555567850015559E1995555592CF3CB2CB0CCF008",
		INIT_24 => x"916008E008F883000881CB1C71C70CCF82515451925566561625555560915996",
		INIT_25 => x"C0F03C83E20080238023C0F030882CF3CF3CF0CCF82515041303C0F03C0F20F8",
		INIT_26 => x"020808E2008220088E08222238020008080C71C31C30CCCF82410000303C0F03",
		INIT_27 => x"1C71CC30C30CCF20800C38022000000008208800202080820208080222208082",
		INIT_28 => x"67899559999E2666659999E2665555649999266678956556255626664F0CC733",
		INIT_29 => x"E00000002380000000300020CF80000000300020CB3CC333C33CF3CB0CCCF896",
		INIT_2A => x"9958959E2556256789565562655899990C732CC71C71C71C333E023800000008",
		INIT_2B => x"899958959E25562567895655625599959992CB30CCF3CF2CB2C3333E2599E589",
		INIT_2C => x"080080CE5660333E185480CE5660333E185590CE5660333C820810400E2599E5",
		INIT_2D => x"255560333C410400000C38220080CD480CCF82002033880CCF8200203320333E",
		INIT_2E => x"0080CCF8800080CCF882206620333E245560333E26679380CCF896656620333E",
		INIT_2F => x"25889625890CCCF84444445444444454444444544444445490CCCF0003083880",
		INIT_30 => x"964D95511665990CCF100204388202080820208080CCCF8882220886243333E2",
		INIT_31 => x"20926022208082020924D95511625890CCF89891515999599964599995999599",
		INIT_32 => x"88220333E2624545666566659166665666566659325444489224333E22000820",
		INIT_33 => x"559915659565995955965959565990CCCF308204008388880020080003200000",
		INIT_34 => x"E0E08E0E08E0E08E0C33330E598662559655866165165821641962033332E598",
		INIT_35 => x"3C030C20010C0F866196080CCCB822082080CCCB822082080CCC782200220008",
		INIT_36 => x"3CF2CB2CB0CCCCF955559E4F939596793E4F93955559E4F939598E4F93E4C333",
		INIT_37 => x"44967983E59E60E59E60F91112594965259635555967983E59E60E59E60C70CF",
		INIT_38 => x"556793E4E5659E4F93E4D55559E4F93959E4F93E4C3333F98396525949658E55",
		INIT_39 => x"2033333E0200080FCCCBE0E0000002320E23830000238388E0E23830CCCC3E4E",
		INIT_3A => x"331F93E4C3333CC30C30810403E0F83E0F83E0F832082383E0F830CCCCF80800",
		INIT_3B => x"CF880CCCF880CCCF996495980CCCCB99E64E19E64E033331E67993899E64E033",
		INIT_3C => x"38899E64E203331F99399E64E643330F939E4E4333C8004103F95593D55930CC",
		INIT_3D => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2F800083E00020C3331E6799",
		INIT_3E => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
		INIT_3F => x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
