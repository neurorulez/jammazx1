-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity PROM4_DST is
port (
	ADDR : in  std_logic_vector(9 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of PROM4_DST is

	signal rom_addr : std_logic_vector(11 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(9 downto 0) <= ADDR;
	end process;

	p_rom : process(rom_addr)
	begin
			DATA <= (others => '0');
			case rom_addr is
				when x"000" => DATA <= x"00";
				when x"001" => DATA <= x"00";
				when x"002" => DATA <= x"00";
				when x"003" => DATA <= x"00";
				when x"004" => DATA <= x"00";
				when x"005" => DATA <= x"05";
				when x"006" => DATA <= x"03";
				when x"007" => DATA <= x"01";
				when x"008" => DATA <= x"00";
				when x"009" => DATA <= x"05";
				when x"00A" => DATA <= x"02";
				when x"00B" => DATA <= x"01";
				when x"00C" => DATA <= x"00";
				when x"00D" => DATA <= x"05";
				when x"00E" => DATA <= x"06";
				when x"00F" => DATA <= x"01";
				when x"010" => DATA <= x"00";
				when x"011" => DATA <= x"05";
				when x"012" => DATA <= x"07";
				when x"013" => DATA <= x"01";
				when x"014" => DATA <= x"00";
				when x"015" => DATA <= x"05";
				when x"016" => DATA <= x"0A";
				when x"017" => DATA <= x"01";
				when x"018" => DATA <= x"00";
				when x"019" => DATA <= x"05";
				when x"01A" => DATA <= x"0B";
				when x"01B" => DATA <= x"01";
				when x"01C" => DATA <= x"00";
				when x"01D" => DATA <= x"05";
				when x"01E" => DATA <= x"0C";
				when x"01F" => DATA <= x"01";
				when x"020" => DATA <= x"00";
				when x"021" => DATA <= x"05";
				when x"022" => DATA <= x"0D";
				when x"023" => DATA <= x"01";
				when x"024" => DATA <= x"00";
				when x"025" => DATA <= x"05";
				when x"026" => DATA <= x"04";
				when x"027" => DATA <= x"01";
				when x"028" => DATA <= x"00";
				when x"029" => DATA <= x"03";
				when x"02A" => DATA <= x"06";
				when x"02B" => DATA <= x"01";
				when x"02C" => DATA <= x"00";
				when x"02D" => DATA <= x"03";
				when x"02E" => DATA <= x"02";
				when x"02F" => DATA <= x"01";
				when x"030" => DATA <= x"00";
				when x"031" => DATA <= x"03";
				when x"032" => DATA <= x"07";
				when x"033" => DATA <= x"01";
				when x"034" => DATA <= x"00";
				when x"035" => DATA <= x"03";
				when x"036" => DATA <= x"05";
				when x"037" => DATA <= x"01";
				when x"038" => DATA <= x"00";
				when x"039" => DATA <= x"02";
				when x"03A" => DATA <= x"03";
				when x"03B" => DATA <= x"01";
				when x"03C" => DATA <= x"00";
				when x"03D" => DATA <= x"00";
				when x"03E" => DATA <= x"00";
				when x"03F" => DATA <= x"00";
				when x"040" => DATA <= x"00";
				when x"041" => DATA <= x"08";
				when x"042" => DATA <= x"03";
				when x"043" => DATA <= x"01";
				when x"044" => DATA <= x"00";
				when x"045" => DATA <= x"09";
				when x"046" => DATA <= x"02";
				when x"047" => DATA <= x"05";
				when x"048" => DATA <= x"00";
				when x"049" => DATA <= x"08";
				when x"04A" => DATA <= x"05";
				when x"04B" => DATA <= x"0D";
				when x"04C" => DATA <= x"04";
				when x"04D" => DATA <= x"04";
				when x"04E" => DATA <= x"04";
				when x"04F" => DATA <= x"04";
				when x"050" => DATA <= x"00";
				when x"051" => DATA <= x"00";
				when x"052" => DATA <= x"00";
				when x"053" => DATA <= x"00";
				when x"054" => DATA <= x"00";
				when x"055" => DATA <= x"00";
				when x"056" => DATA <= x"00";
				when x"057" => DATA <= x"00";
				when x"058" => DATA <= x"00";
				when x"059" => DATA <= x"02";
				when x"05A" => DATA <= x"02";
				when x"05B" => DATA <= x"02";
				when x"05C" => DATA <= x"00";
				when x"05D" => DATA <= x"03";
				when x"05E" => DATA <= x"03";
				when x"05F" => DATA <= x"03";
				when x"060" => DATA <= x"00";
				when x"061" => DATA <= x"06";
				when x"062" => DATA <= x"06";
				when x"063" => DATA <= x"06";
				when x"064" => DATA <= x"00";
				when x"065" => DATA <= x"07";
				when x"066" => DATA <= x"07";
				when x"067" => DATA <= x"07";
				when x"068" => DATA <= x"00";
				when x"069" => DATA <= x"0A";
				when x"06A" => DATA <= x"0A";
				when x"06B" => DATA <= x"0A";
				when x"06C" => DATA <= x"00";
				when x"06D" => DATA <= x"0B";
				when x"06E" => DATA <= x"0B";
				when x"06F" => DATA <= x"0B";
				when x"070" => DATA <= x"00";
				when x"071" => DATA <= x"01";
				when x"072" => DATA <= x"01";
				when x"073" => DATA <= x"01";
				when x"074" => DATA <= x"00";
				when x"075" => DATA <= x"05";
				when x"076" => DATA <= x"05";
				when x"077" => DATA <= x"05";
				when x"078" => DATA <= x"08";
				when x"079" => DATA <= x"09";
				when x"07A" => DATA <= x"0A";
				when x"07B" => DATA <= x"0B";
				when x"07C" => DATA <= x"0C";
				when x"07D" => DATA <= x"0D";
				when x"07E" => DATA <= x"0E";
				when x"07F" => DATA <= x"0F";
				when x"080" => DATA <= x"00";
				when x"081" => DATA <= x"00";
				when x"082" => DATA <= x"00";
				when x"083" => DATA <= x"00";
				when x"084" => DATA <= x"00";
				when x"085" => DATA <= x"03";
				when x"086" => DATA <= x"07";
				when x"087" => DATA <= x"0D";
				when x"088" => DATA <= x"00";
				when x"089" => DATA <= x"0C";
				when x"08A" => DATA <= x"0F";
				when x"08B" => DATA <= x"0B";
				when x"08C" => DATA <= x"00";
				when x"08D" => DATA <= x"0C";
				when x"08E" => DATA <= x"0E";
				when x"08F" => DATA <= x"0B";
				when x"090" => DATA <= x"00";
				when x"091" => DATA <= x"0C";
				when x"092" => DATA <= x"06";
				when x"093" => DATA <= x"0B";
				when x"094" => DATA <= x"00";
				when x"095" => DATA <= x"0C";
				when x"096" => DATA <= x"07";
				when x"097" => DATA <= x"0B";
				when x"098" => DATA <= x"00";
				when x"099" => DATA <= x"0C";
				when x"09A" => DATA <= x"03";
				when x"09B" => DATA <= x"0B";
				when x"09C" => DATA <= x"00";
				when x"09D" => DATA <= x"0C";
				when x"09E" => DATA <= x"08";
				when x"09F" => DATA <= x"0B";
				when x"0A0" => DATA <= x"00";
				when x"0A1" => DATA <= x"0C";
				when x"0A2" => DATA <= x"0D";
				when x"0A3" => DATA <= x"0B";
				when x"0A4" => DATA <= x"00";
				when x"0A5" => DATA <= x"0C";
				when x"0A6" => DATA <= x"04";
				when x"0A7" => DATA <= x"0B";
				when x"0A8" => DATA <= x"00";
				when x"0A9" => DATA <= x"0C";
				when x"0AA" => DATA <= x"09";
				when x"0AB" => DATA <= x"0B";
				when x"0AC" => DATA <= x"00";
				when x"0AD" => DATA <= x"0C";
				when x"0AE" => DATA <= x"05";
				when x"0AF" => DATA <= x"0B";
				when x"0B0" => DATA <= x"00";
				when x"0B1" => DATA <= x"0C";
				when x"0B2" => DATA <= x"02";
				when x"0B3" => DATA <= x"0B";
				when x"0B4" => DATA <= x"00";
				when x"0B5" => DATA <= x"0C";
				when x"0B6" => DATA <= x"0B";
				when x"0B7" => DATA <= x"02";
				when x"0B8" => DATA <= x"00";
				when x"0B9" => DATA <= x"08";
				when x"0BA" => DATA <= x"0C";
				when x"0BB" => DATA <= x"02";
				when x"0BC" => DATA <= x"00";
				when x"0BD" => DATA <= x"08";
				when x"0BE" => DATA <= x"0F";
				when x"0BF" => DATA <= x"02";
				when x"0C0" => DATA <= x"00";
				when x"0C1" => DATA <= x"03";
				when x"0C2" => DATA <= x"02";
				when x"0C3" => DATA <= x"01";
				when x"0C4" => DATA <= x"00";
				when x"0C5" => DATA <= x"02";
				when x"0C6" => DATA <= x"0F";
				when x"0C7" => DATA <= x"03";
				when x"0C8" => DATA <= x"00";
				when x"0C9" => DATA <= x"0F";
				when x"0CA" => DATA <= x"0E";
				when x"0CB" => DATA <= x"02";
				when x"0CC" => DATA <= x"00";
				when x"0CD" => DATA <= x"0E";
				when x"0CE" => DATA <= x"07";
				when x"0CF" => DATA <= x"0F";
				when x"0D0" => DATA <= x"00";
				when x"0D1" => DATA <= x"07";
				when x"0D2" => DATA <= x"06";
				when x"0D3" => DATA <= x"0E";
				when x"0D4" => DATA <= x"00";
				when x"0D5" => DATA <= x"06";
				when x"0D6" => DATA <= x"05";
				when x"0D7" => DATA <= x"07";
				when x"0D8" => DATA <= x"00";
				when x"0D9" => DATA <= x"05";
				when x"0DA" => DATA <= x"00";
				when x"0DB" => DATA <= x"06";
				when x"0DC" => DATA <= x"00";
				when x"0DD" => DATA <= x"00";
				when x"0DE" => DATA <= x"0B";
				when x"0DF" => DATA <= x"05";
				when x"0E0" => DATA <= x"00";
				when x"0E1" => DATA <= x"0B";
				when x"0E2" => DATA <= x"0C";
				when x"0E3" => DATA <= x"00";
				when x"0E4" => DATA <= x"00";
				when x"0E5" => DATA <= x"0C";
				when x"0E6" => DATA <= x"0D";
				when x"0E7" => DATA <= x"0B";
				when x"0E8" => DATA <= x"00";
				when x"0E9" => DATA <= x"0D";
				when x"0EA" => DATA <= x"08";
				when x"0EB" => DATA <= x"0C";
				when x"0EC" => DATA <= x"00";
				when x"0ED" => DATA <= x"08";
				when x"0EE" => DATA <= x"09";
				when x"0EF" => DATA <= x"0D";
				when x"0F0" => DATA <= x"00";
				when x"0F1" => DATA <= x"09";
				when x"0F2" => DATA <= x"0A";
				when x"0F3" => DATA <= x"08";
				when x"0F4" => DATA <= x"00";
				when x"0F5" => DATA <= x"0A";
				when x"0F6" => DATA <= x"01";
				when x"0F7" => DATA <= x"09";
				when x"0F8" => DATA <= x"00";
				when x"0F9" => DATA <= x"01";
				when x"0FA" => DATA <= x"04";
				when x"0FB" => DATA <= x"0A";
				when x"0FC" => DATA <= x"00";
				when x"0FD" => DATA <= x"04";
				when x"0FE" => DATA <= x"03";
				when x"0FF" => DATA <= x"01";
				when x"100" => DATA <= x"00";
				when x"101" => DATA <= x"00";
				when x"102" => DATA <= x"00";
				when x"103" => DATA <= x"00";
				when x"104" => DATA <= x"00";
				when x"105" => DATA <= x"03";
				when x"106" => DATA <= x"07";
				when x"107" => DATA <= x"0D";
				when x"108" => DATA <= x"00";
				when x"109" => DATA <= x"0C";
				when x"10A" => DATA <= x"0F";
				when x"10B" => DATA <= x"0B";
				when x"10C" => DATA <= x"00";
				when x"10D" => DATA <= x"0C";
				when x"10E" => DATA <= x"0E";
				when x"10F" => DATA <= x"0B";
				when x"110" => DATA <= x"00";
				when x"111" => DATA <= x"0C";
				when x"112" => DATA <= x"06";
				when x"113" => DATA <= x"0B";
				when x"114" => DATA <= x"00";
				when x"115" => DATA <= x"0C";
				when x"116" => DATA <= x"07";
				when x"117" => DATA <= x"0B";
				when x"118" => DATA <= x"00";
				when x"119" => DATA <= x"0C";
				when x"11A" => DATA <= x"03";
				when x"11B" => DATA <= x"0B";
				when x"11C" => DATA <= x"00";
				when x"11D" => DATA <= x"0C";
				when x"11E" => DATA <= x"08";
				when x"11F" => DATA <= x"0B";
				when x"120" => DATA <= x"00";
				when x"121" => DATA <= x"0C";
				when x"122" => DATA <= x"0D";
				when x"123" => DATA <= x"0B";
				when x"124" => DATA <= x"00";
				when x"125" => DATA <= x"0C";
				when x"126" => DATA <= x"04";
				when x"127" => DATA <= x"0B";
				when x"128" => DATA <= x"00";
				when x"129" => DATA <= x"0C";
				when x"12A" => DATA <= x"09";
				when x"12B" => DATA <= x"0B";
				when x"12C" => DATA <= x"00";
				when x"12D" => DATA <= x"0C";
				when x"12E" => DATA <= x"05";
				when x"12F" => DATA <= x"0B";
				when x"130" => DATA <= x"00";
				when x"131" => DATA <= x"0C";
				when x"132" => DATA <= x"02";
				when x"133" => DATA <= x"0B";
				when x"134" => DATA <= x"00";
				when x"135" => DATA <= x"0C";
				when x"136" => DATA <= x"0B";
				when x"137" => DATA <= x"02";
				when x"138" => DATA <= x"00";
				when x"139" => DATA <= x"08";
				when x"13A" => DATA <= x"0C";
				when x"13B" => DATA <= x"02";
				when x"13C" => DATA <= x"00";
				when x"13D" => DATA <= x"08";
				when x"13E" => DATA <= x"0F";
				when x"13F" => DATA <= x"02";
				when x"140" => DATA <= x"00";
				when x"141" => DATA <= x"03";
				when x"142" => DATA <= x"02";
				when x"143" => DATA <= x"01";
				when x"144" => DATA <= x"00";
				when x"145" => DATA <= x"02";
				when x"146" => DATA <= x"0F";
				when x"147" => DATA <= x"03";
				when x"148" => DATA <= x"00";
				when x"149" => DATA <= x"0F";
				when x"14A" => DATA <= x"0E";
				when x"14B" => DATA <= x"02";
				when x"14C" => DATA <= x"00";
				when x"14D" => DATA <= x"0E";
				when x"14E" => DATA <= x"07";
				when x"14F" => DATA <= x"0F";
				when x"150" => DATA <= x"00";
				when x"151" => DATA <= x"07";
				when x"152" => DATA <= x"06";
				when x"153" => DATA <= x"0E";
				when x"154" => DATA <= x"00";
				when x"155" => DATA <= x"06";
				when x"156" => DATA <= x"05";
				when x"157" => DATA <= x"07";
				when x"158" => DATA <= x"00";
				when x"159" => DATA <= x"05";
				when x"15A" => DATA <= x"00";
				when x"15B" => DATA <= x"06";
				when x"15C" => DATA <= x"00";
				when x"15D" => DATA <= x"00";
				when x"15E" => DATA <= x"0B";
				when x"15F" => DATA <= x"05";
				when x"160" => DATA <= x"00";
				when x"161" => DATA <= x"0B";
				when x"162" => DATA <= x"0C";
				when x"163" => DATA <= x"00";
				when x"164" => DATA <= x"00";
				when x"165" => DATA <= x"0C";
				when x"166" => DATA <= x"0D";
				when x"167" => DATA <= x"0B";
				when x"168" => DATA <= x"00";
				when x"169" => DATA <= x"0D";
				when x"16A" => DATA <= x"08";
				when x"16B" => DATA <= x"0C";
				when x"16C" => DATA <= x"00";
				when x"16D" => DATA <= x"08";
				when x"16E" => DATA <= x"09";
				when x"16F" => DATA <= x"0D";
				when x"170" => DATA <= x"00";
				when x"171" => DATA <= x"09";
				when x"172" => DATA <= x"0A";
				when x"173" => DATA <= x"08";
				when x"174" => DATA <= x"00";
				when x"175" => DATA <= x"0A";
				when x"176" => DATA <= x"01";
				when x"177" => DATA <= x"09";
				when x"178" => DATA <= x"00";
				when x"179" => DATA <= x"01";
				when x"17A" => DATA <= x"04";
				when x"17B" => DATA <= x"0A";
				when x"17C" => DATA <= x"00";
				when x"17D" => DATA <= x"04";
				when x"17E" => DATA <= x"03";
				when x"17F" => DATA <= x"01";
				when x"180" => DATA <= x"0F";
				when x"181" => DATA <= x"00";
				when x"182" => DATA <= x"0F";
				when x"183" => DATA <= x"00";
				when x"184" => DATA <= x"0F";
				when x"185" => DATA <= x"00";
				when x"186" => DATA <= x"0F";
				when x"187" => DATA <= x"00";
				when x"188" => DATA <= x"0F";
				when x"189" => DATA <= x"00";
				when x"18A" => DATA <= x"0F";
				when x"18B" => DATA <= x"00";
				when x"18C" => DATA <= x"0F";
				when x"18D" => DATA <= x"00";
				when x"18E" => DATA <= x"0F";
				when x"18F" => DATA <= x"00";
				when x"190" => DATA <= x"0F";
				when x"191" => DATA <= x"00";
				when x"192" => DATA <= x"0F";
				when x"193" => DATA <= x"00";
				when x"194" => DATA <= x"0F";
				when x"195" => DATA <= x"00";
				when x"196" => DATA <= x"0F";
				when x"197" => DATA <= x"00";
				when x"198" => DATA <= x"0F";
				when x"199" => DATA <= x"00";
				when x"19A" => DATA <= x"0F";
				when x"19B" => DATA <= x"00";
				when x"19C" => DATA <= x"0F";
				when x"19D" => DATA <= x"00";
				when x"19E" => DATA <= x"0F";
				when x"19F" => DATA <= x"00";
				when x"1A0" => DATA <= x"0F";
				when x"1A1" => DATA <= x"00";
				when x"1A2" => DATA <= x"0F";
				when x"1A3" => DATA <= x"00";
				when x"1A4" => DATA <= x"0F";
				when x"1A5" => DATA <= x"00";
				when x"1A6" => DATA <= x"0F";
				when x"1A7" => DATA <= x"00";
				when x"1A8" => DATA <= x"0F";
				when x"1A9" => DATA <= x"00";
				when x"1AA" => DATA <= x"0F";
				when x"1AB" => DATA <= x"00";
				when x"1AC" => DATA <= x"0F";
				when x"1AD" => DATA <= x"00";
				when x"1AE" => DATA <= x"0F";
				when x"1AF" => DATA <= x"00";
				when x"1B0" => DATA <= x"0F";
				when x"1B1" => DATA <= x"00";
				when x"1B2" => DATA <= x"0F";
				when x"1B3" => DATA <= x"00";
				when x"1B4" => DATA <= x"0F";
				when x"1B5" => DATA <= x"00";
				when x"1B6" => DATA <= x"0F";
				when x"1B7" => DATA <= x"00";
				when x"1B8" => DATA <= x"0F";
				when x"1B9" => DATA <= x"00";
				when x"1BA" => DATA <= x"0F";
				when x"1BB" => DATA <= x"00";
				when x"1BC" => DATA <= x"0F";
				when x"1BD" => DATA <= x"00";
				when x"1BE" => DATA <= x"0F";
				when x"1BF" => DATA <= x"00";
				when x"1C0" => DATA <= x"0F";
				when x"1C1" => DATA <= x"00";
				when x"1C2" => DATA <= x"0F";
				when x"1C3" => DATA <= x"00";
				when x"1C4" => DATA <= x"0F";
				when x"1C5" => DATA <= x"00";
				when x"1C6" => DATA <= x"0F";
				when x"1C7" => DATA <= x"00";
				when x"1C8" => DATA <= x"0F";
				when x"1C9" => DATA <= x"00";
				when x"1CA" => DATA <= x"0F";
				when x"1CB" => DATA <= x"00";
				when x"1CC" => DATA <= x"0F";
				when x"1CD" => DATA <= x"00";
				when x"1CE" => DATA <= x"0F";
				when x"1CF" => DATA <= x"00";
				when x"1D0" => DATA <= x"0F";
				when x"1D1" => DATA <= x"00";
				when x"1D2" => DATA <= x"0F";
				when x"1D3" => DATA <= x"00";
				when x"1D4" => DATA <= x"0F";
				when x"1D5" => DATA <= x"00";
				when x"1D6" => DATA <= x"0F";
				when x"1D7" => DATA <= x"00";
				when x"1D8" => DATA <= x"0F";
				when x"1D9" => DATA <= x"00";
				when x"1DA" => DATA <= x"0F";
				when x"1DB" => DATA <= x"00";
				when x"1DC" => DATA <= x"0F";
				when x"1DD" => DATA <= x"00";
				when x"1DE" => DATA <= x"0F";
				when x"1DF" => DATA <= x"00";
				when x"1E0" => DATA <= x"0F";
				when x"1E1" => DATA <= x"00";
				when x"1E2" => DATA <= x"0F";
				when x"1E3" => DATA <= x"00";
				when x"1E4" => DATA <= x"0F";
				when x"1E5" => DATA <= x"00";
				when x"1E6" => DATA <= x"0F";
				when x"1E7" => DATA <= x"00";
				when x"1E8" => DATA <= x"0F";
				when x"1E9" => DATA <= x"00";
				when x"1EA" => DATA <= x"0F";
				when x"1EB" => DATA <= x"00";
				when x"1EC" => DATA <= x"0F";
				when x"1ED" => DATA <= x"00";
				when x"1EE" => DATA <= x"0F";
				when x"1EF" => DATA <= x"00";
				when x"1F0" => DATA <= x"0F";
				when x"1F1" => DATA <= x"00";
				when x"1F2" => DATA <= x"0F";
				when x"1F3" => DATA <= x"00";
				when x"1F4" => DATA <= x"0F";
				when x"1F5" => DATA <= x"00";
				when x"1F6" => DATA <= x"0F";
				when x"1F7" => DATA <= x"00";
				when x"1F8" => DATA <= x"0F";
				when x"1F9" => DATA <= x"00";
				when x"1FA" => DATA <= x"0F";
				when x"1FB" => DATA <= x"00";
				when x"1FC" => DATA <= x"0F";
				when x"1FD" => DATA <= x"00";
				when x"1FE" => DATA <= x"0F";
				when x"1FF" => DATA <= x"00";
				when x"200" => DATA <= x"00";
				when x"201" => DATA <= x"0F";
				when x"202" => DATA <= x"00";
				when x"203" => DATA <= x"0F";
				when x"204" => DATA <= x"00";
				when x"205" => DATA <= x"0F";
				when x"206" => DATA <= x"00";
				when x"207" => DATA <= x"0F";
				when x"208" => DATA <= x"00";
				when x"209" => DATA <= x"0F";
				when x"20A" => DATA <= x"00";
				when x"20B" => DATA <= x"0F";
				when x"20C" => DATA <= x"00";
				when x"20D" => DATA <= x"0F";
				when x"20E" => DATA <= x"00";
				when x"20F" => DATA <= x"0F";
				when x"210" => DATA <= x"00";
				when x"211" => DATA <= x"0F";
				when x"212" => DATA <= x"00";
				when x"213" => DATA <= x"0F";
				when x"214" => DATA <= x"00";
				when x"215" => DATA <= x"0F";
				when x"216" => DATA <= x"00";
				when x"217" => DATA <= x"0F";
				when x"218" => DATA <= x"00";
				when x"219" => DATA <= x"0F";
				when x"21A" => DATA <= x"00";
				when x"21B" => DATA <= x"0F";
				when x"21C" => DATA <= x"00";
				when x"21D" => DATA <= x"0F";
				when x"21E" => DATA <= x"00";
				when x"21F" => DATA <= x"0F";
				when x"220" => DATA <= x"00";
				when x"221" => DATA <= x"0F";
				when x"222" => DATA <= x"00";
				when x"223" => DATA <= x"0F";
				when x"224" => DATA <= x"00";
				when x"225" => DATA <= x"0F";
				when x"226" => DATA <= x"00";
				when x"227" => DATA <= x"0F";
				when x"228" => DATA <= x"00";
				when x"229" => DATA <= x"0F";
				when x"22A" => DATA <= x"00";
				when x"22B" => DATA <= x"0F";
				when x"22C" => DATA <= x"00";
				when x"22D" => DATA <= x"0F";
				when x"22E" => DATA <= x"00";
				when x"22F" => DATA <= x"0F";
				when x"230" => DATA <= x"00";
				when x"231" => DATA <= x"0F";
				when x"232" => DATA <= x"00";
				when x"233" => DATA <= x"0F";
				when x"234" => DATA <= x"00";
				when x"235" => DATA <= x"0F";
				when x"236" => DATA <= x"00";
				when x"237" => DATA <= x"0F";
				when x"238" => DATA <= x"00";
				when x"239" => DATA <= x"0F";
				when x"23A" => DATA <= x"00";
				when x"23B" => DATA <= x"0F";
				when x"23C" => DATA <= x"00";
				when x"23D" => DATA <= x"0F";
				when x"23E" => DATA <= x"00";
				when x"23F" => DATA <= x"0F";
				when x"240" => DATA <= x"00";
				when x"241" => DATA <= x"0F";
				when x"242" => DATA <= x"00";
				when x"243" => DATA <= x"0F";
				when x"244" => DATA <= x"00";
				when x"245" => DATA <= x"0F";
				when x"246" => DATA <= x"00";
				when x"247" => DATA <= x"0F";
				when x"248" => DATA <= x"00";
				when x"249" => DATA <= x"0F";
				when x"24A" => DATA <= x"00";
				when x"24B" => DATA <= x"0F";
				when x"24C" => DATA <= x"00";
				when x"24D" => DATA <= x"0F";
				when x"24E" => DATA <= x"00";
				when x"24F" => DATA <= x"0F";
				when x"250" => DATA <= x"00";
				when x"251" => DATA <= x"0F";
				when x"252" => DATA <= x"00";
				when x"253" => DATA <= x"0F";
				when x"254" => DATA <= x"00";
				when x"255" => DATA <= x"0F";
				when x"256" => DATA <= x"00";
				when x"257" => DATA <= x"0F";
				when x"258" => DATA <= x"00";
				when x"259" => DATA <= x"0F";
				when x"25A" => DATA <= x"00";
				when x"25B" => DATA <= x"0F";
				when x"25C" => DATA <= x"00";
				when x"25D" => DATA <= x"0F";
				when x"25E" => DATA <= x"00";
				when x"25F" => DATA <= x"0F";
				when x"260" => DATA <= x"00";
				when x"261" => DATA <= x"0F";
				when x"262" => DATA <= x"00";
				when x"263" => DATA <= x"0F";
				when x"264" => DATA <= x"00";
				when x"265" => DATA <= x"0F";
				when x"266" => DATA <= x"00";
				when x"267" => DATA <= x"0F";
				when x"268" => DATA <= x"00";
				when x"269" => DATA <= x"0F";
				when x"26A" => DATA <= x"00";
				when x"26B" => DATA <= x"0F";
				when x"26C" => DATA <= x"00";
				when x"26D" => DATA <= x"0F";
				when x"26E" => DATA <= x"00";
				when x"26F" => DATA <= x"0F";
				when x"270" => DATA <= x"00";
				when x"271" => DATA <= x"0F";
				when x"272" => DATA <= x"00";
				when x"273" => DATA <= x"0F";
				when x"274" => DATA <= x"00";
				when x"275" => DATA <= x"0F";
				when x"276" => DATA <= x"00";
				when x"277" => DATA <= x"0F";
				when x"278" => DATA <= x"00";
				when x"279" => DATA <= x"0F";
				when x"27A" => DATA <= x"00";
				when x"27B" => DATA <= x"0F";
				when x"27C" => DATA <= x"00";
				when x"27D" => DATA <= x"0F";
				when x"27E" => DATA <= x"00";
				when x"27F" => DATA <= x"07";
				when x"280" => DATA <= x"0F";
				when x"281" => DATA <= x"00";
				when x"282" => DATA <= x"0F";
				when x"283" => DATA <= x"00";
				when x"284" => DATA <= x"0F";
				when x"285" => DATA <= x"00";
				when x"286" => DATA <= x"0F";
				when x"287" => DATA <= x"00";
				when x"288" => DATA <= x"0F";
				when x"289" => DATA <= x"00";
				when x"28A" => DATA <= x"0F";
				when x"28B" => DATA <= x"00";
				when x"28C" => DATA <= x"0F";
				when x"28D" => DATA <= x"00";
				when x"28E" => DATA <= x"0F";
				when x"28F" => DATA <= x"00";
				when x"290" => DATA <= x"0F";
				when x"291" => DATA <= x"00";
				when x"292" => DATA <= x"0F";
				when x"293" => DATA <= x"00";
				when x"294" => DATA <= x"0F";
				when x"295" => DATA <= x"00";
				when x"296" => DATA <= x"0F";
				when x"297" => DATA <= x"00";
				when x"298" => DATA <= x"0F";
				when x"299" => DATA <= x"00";
				when x"29A" => DATA <= x"0F";
				when x"29B" => DATA <= x"00";
				when x"29C" => DATA <= x"0F";
				when x"29D" => DATA <= x"00";
				when x"29E" => DATA <= x"0F";
				when x"29F" => DATA <= x"00";
				when x"2A0" => DATA <= x"0F";
				when x"2A1" => DATA <= x"00";
				when x"2A2" => DATA <= x"0F";
				when x"2A3" => DATA <= x"00";
				when x"2A4" => DATA <= x"0F";
				when x"2A5" => DATA <= x"00";
				when x"2A6" => DATA <= x"0F";
				when x"2A7" => DATA <= x"00";
				when x"2A8" => DATA <= x"0F";
				when x"2A9" => DATA <= x"00";
				when x"2AA" => DATA <= x"0F";
				when x"2AB" => DATA <= x"00";
				when x"2AC" => DATA <= x"0F";
				when x"2AD" => DATA <= x"00";
				when x"2AE" => DATA <= x"0F";
				when x"2AF" => DATA <= x"00";
				when x"2B0" => DATA <= x"0F";
				when x"2B1" => DATA <= x"00";
				when x"2B2" => DATA <= x"0F";
				when x"2B3" => DATA <= x"00";
				when x"2B4" => DATA <= x"0F";
				when x"2B5" => DATA <= x"00";
				when x"2B6" => DATA <= x"0F";
				when x"2B7" => DATA <= x"00";
				when x"2B8" => DATA <= x"0F";
				when x"2B9" => DATA <= x"00";
				when x"2BA" => DATA <= x"0F";
				when x"2BB" => DATA <= x"00";
				when x"2BC" => DATA <= x"0F";
				when x"2BD" => DATA <= x"00";
				when x"2BE" => DATA <= x"0F";
				when x"2BF" => DATA <= x"00";
				when x"2C0" => DATA <= x"0F";
				when x"2C1" => DATA <= x"00";
				when x"2C2" => DATA <= x"0F";
				when x"2C3" => DATA <= x"00";
				when x"2C4" => DATA <= x"0F";
				when x"2C5" => DATA <= x"00";
				when x"2C6" => DATA <= x"0F";
				when x"2C7" => DATA <= x"00";
				when x"2C8" => DATA <= x"0F";
				when x"2C9" => DATA <= x"00";
				when x"2CA" => DATA <= x"0F";
				when x"2CB" => DATA <= x"00";
				when x"2CC" => DATA <= x"0F";
				when x"2CD" => DATA <= x"00";
				when x"2CE" => DATA <= x"0F";
				when x"2CF" => DATA <= x"00";
				when x"2D0" => DATA <= x"0F";
				when x"2D1" => DATA <= x"00";
				when x"2D2" => DATA <= x"0F";
				when x"2D3" => DATA <= x"00";
				when x"2D4" => DATA <= x"0F";
				when x"2D5" => DATA <= x"00";
				when x"2D6" => DATA <= x"0F";
				when x"2D7" => DATA <= x"00";
				when x"2D8" => DATA <= x"0F";
				when x"2D9" => DATA <= x"00";
				when x"2DA" => DATA <= x"0F";
				when x"2DB" => DATA <= x"00";
				when x"2DC" => DATA <= x"0F";
				when x"2DD" => DATA <= x"00";
				when x"2DE" => DATA <= x"0F";
				when x"2DF" => DATA <= x"00";
				when x"2E0" => DATA <= x"0F";
				when x"2E1" => DATA <= x"00";
				when x"2E2" => DATA <= x"0F";
				when x"2E3" => DATA <= x"00";
				when x"2E4" => DATA <= x"0F";
				when x"2E5" => DATA <= x"00";
				when x"2E6" => DATA <= x"0F";
				when x"2E7" => DATA <= x"00";
				when x"2E8" => DATA <= x"0F";
				when x"2E9" => DATA <= x"00";
				when x"2EA" => DATA <= x"0F";
				when x"2EB" => DATA <= x"00";
				when x"2EC" => DATA <= x"0F";
				when x"2ED" => DATA <= x"00";
				when x"2EE" => DATA <= x"0F";
				when x"2EF" => DATA <= x"00";
				when x"2F0" => DATA <= x"0F";
				when x"2F1" => DATA <= x"00";
				when x"2F2" => DATA <= x"0F";
				when x"2F3" => DATA <= x"00";
				when x"2F4" => DATA <= x"0F";
				when x"2F5" => DATA <= x"00";
				when x"2F6" => DATA <= x"0F";
				when x"2F7" => DATA <= x"00";
				when x"2F8" => DATA <= x"0F";
				when x"2F9" => DATA <= x"00";
				when x"2FA" => DATA <= x"0F";
				when x"2FB" => DATA <= x"00";
				when x"2FC" => DATA <= x"0F";
				when x"2FD" => DATA <= x"00";
				when x"2FE" => DATA <= x"0F";
				when x"2FF" => DATA <= x"0D";
				when x"300" => DATA <= x"00";
				when x"301" => DATA <= x"0F";
				when x"302" => DATA <= x"00";
				when x"303" => DATA <= x"0F";
				when x"304" => DATA <= x"00";
				when x"305" => DATA <= x"0F";
				when x"306" => DATA <= x"00";
				when x"307" => DATA <= x"0F";
				when x"308" => DATA <= x"00";
				when x"309" => DATA <= x"0F";
				when x"30A" => DATA <= x"00";
				when x"30B" => DATA <= x"0F";
				when x"30C" => DATA <= x"00";
				when x"30D" => DATA <= x"0F";
				when x"30E" => DATA <= x"00";
				when x"30F" => DATA <= x"0F";
				when x"310" => DATA <= x"00";
				when x"311" => DATA <= x"0F";
				when x"312" => DATA <= x"00";
				when x"313" => DATA <= x"0F";
				when x"314" => DATA <= x"00";
				when x"315" => DATA <= x"0F";
				when x"316" => DATA <= x"00";
				when x"317" => DATA <= x"0F";
				when x"318" => DATA <= x"00";
				when x"319" => DATA <= x"0F";
				when x"31A" => DATA <= x"00";
				when x"31B" => DATA <= x"0F";
				when x"31C" => DATA <= x"00";
				when x"31D" => DATA <= x"0F";
				when x"31E" => DATA <= x"00";
				when x"31F" => DATA <= x"0F";
				when x"320" => DATA <= x"00";
				when x"321" => DATA <= x"0F";
				when x"322" => DATA <= x"00";
				when x"323" => DATA <= x"0F";
				when x"324" => DATA <= x"00";
				when x"325" => DATA <= x"0F";
				when x"326" => DATA <= x"00";
				when x"327" => DATA <= x"0F";
				when x"328" => DATA <= x"00";
				when x"329" => DATA <= x"0F";
				when x"32A" => DATA <= x"00";
				when x"32B" => DATA <= x"0F";
				when x"32C" => DATA <= x"00";
				when x"32D" => DATA <= x"0F";
				when x"32E" => DATA <= x"00";
				when x"32F" => DATA <= x"0F";
				when x"330" => DATA <= x"00";
				when x"331" => DATA <= x"0F";
				when x"332" => DATA <= x"00";
				when x"333" => DATA <= x"0F";
				when x"334" => DATA <= x"00";
				when x"335" => DATA <= x"0F";
				when x"336" => DATA <= x"00";
				when x"337" => DATA <= x"0F";
				when x"338" => DATA <= x"00";
				when x"339" => DATA <= x"0F";
				when x"33A" => DATA <= x"00";
				when x"33B" => DATA <= x"0F";
				when x"33C" => DATA <= x"00";
				when x"33D" => DATA <= x"0F";
				when x"33E" => DATA <= x"00";
				when x"33F" => DATA <= x"0F";
				when x"340" => DATA <= x"00";
				when x"341" => DATA <= x"0F";
				when x"342" => DATA <= x"00";
				when x"343" => DATA <= x"0F";
				when x"344" => DATA <= x"00";
				when x"345" => DATA <= x"0F";
				when x"346" => DATA <= x"00";
				when x"347" => DATA <= x"0F";
				when x"348" => DATA <= x"00";
				when x"349" => DATA <= x"0F";
				when x"34A" => DATA <= x"00";
				when x"34B" => DATA <= x"0F";
				when x"34C" => DATA <= x"00";
				when x"34D" => DATA <= x"0F";
				when x"34E" => DATA <= x"00";
				when x"34F" => DATA <= x"0F";
				when x"350" => DATA <= x"00";
				when x"351" => DATA <= x"0F";
				when x"352" => DATA <= x"00";
				when x"353" => DATA <= x"0F";
				when x"354" => DATA <= x"00";
				when x"355" => DATA <= x"0F";
				when x"356" => DATA <= x"00";
				when x"357" => DATA <= x"0F";
				when x"358" => DATA <= x"00";
				when x"359" => DATA <= x"0F";
				when x"35A" => DATA <= x"00";
				when x"35B" => DATA <= x"0F";
				when x"35C" => DATA <= x"00";
				when x"35D" => DATA <= x"0F";
				when x"35E" => DATA <= x"00";
				when x"35F" => DATA <= x"0F";
				when x"360" => DATA <= x"00";
				when x"361" => DATA <= x"0F";
				when x"362" => DATA <= x"00";
				when x"363" => DATA <= x"0F";
				when x"364" => DATA <= x"00";
				when x"365" => DATA <= x"0F";
				when x"366" => DATA <= x"00";
				when x"367" => DATA <= x"0F";
				when x"368" => DATA <= x"00";
				when x"369" => DATA <= x"0F";
				when x"36A" => DATA <= x"00";
				when x"36B" => DATA <= x"0F";
				when x"36C" => DATA <= x"00";
				when x"36D" => DATA <= x"0F";
				when x"36E" => DATA <= x"00";
				when x"36F" => DATA <= x"0F";
				when x"370" => DATA <= x"00";
				when x"371" => DATA <= x"0F";
				when x"372" => DATA <= x"00";
				when x"373" => DATA <= x"0F";
				when x"374" => DATA <= x"00";
				when x"375" => DATA <= x"0F";
				when x"376" => DATA <= x"00";
				when x"377" => DATA <= x"0F";
				when x"378" => DATA <= x"00";
				when x"379" => DATA <= x"0F";
				when x"37A" => DATA <= x"00";
				when x"37B" => DATA <= x"0F";
				when x"37C" => DATA <= x"00";
				when x"37D" => DATA <= x"0F";
				when x"37E" => DATA <= x"00";
				when x"37F" => DATA <= x"07";
				when x"380" => DATA <= x"0F";
				when x"381" => DATA <= x"00";
				when x"382" => DATA <= x"0F";
				when x"383" => DATA <= x"00";
				when x"384" => DATA <= x"0F";
				when x"385" => DATA <= x"00";
				when x"386" => DATA <= x"0F";
				when x"387" => DATA <= x"00";
				when x"388" => DATA <= x"0F";
				when x"389" => DATA <= x"00";
				when x"38A" => DATA <= x"0F";
				when x"38B" => DATA <= x"00";
				when x"38C" => DATA <= x"0F";
				when x"38D" => DATA <= x"00";
				when x"38E" => DATA <= x"0F";
				when x"38F" => DATA <= x"00";
				when x"390" => DATA <= x"0F";
				when x"391" => DATA <= x"00";
				when x"392" => DATA <= x"0F";
				when x"393" => DATA <= x"00";
				when x"394" => DATA <= x"0F";
				when x"395" => DATA <= x"00";
				when x"396" => DATA <= x"0F";
				when x"397" => DATA <= x"00";
				when x"398" => DATA <= x"0F";
				when x"399" => DATA <= x"00";
				when x"39A" => DATA <= x"0F";
				when x"39B" => DATA <= x"00";
				when x"39C" => DATA <= x"0F";
				when x"39D" => DATA <= x"00";
				when x"39E" => DATA <= x"0F";
				when x"39F" => DATA <= x"00";
				when x"3A0" => DATA <= x"0F";
				when x"3A1" => DATA <= x"00";
				when x"3A2" => DATA <= x"0F";
				when x"3A3" => DATA <= x"00";
				when x"3A4" => DATA <= x"0F";
				when x"3A5" => DATA <= x"00";
				when x"3A6" => DATA <= x"0F";
				when x"3A7" => DATA <= x"00";
				when x"3A8" => DATA <= x"0F";
				when x"3A9" => DATA <= x"00";
				when x"3AA" => DATA <= x"0F";
				when x"3AB" => DATA <= x"00";
				when x"3AC" => DATA <= x"0F";
				when x"3AD" => DATA <= x"00";
				when x"3AE" => DATA <= x"0F";
				when x"3AF" => DATA <= x"00";
				when x"3B0" => DATA <= x"0F";
				when x"3B1" => DATA <= x"00";
				when x"3B2" => DATA <= x"0F";
				when x"3B3" => DATA <= x"00";
				when x"3B4" => DATA <= x"0F";
				when x"3B5" => DATA <= x"00";
				when x"3B6" => DATA <= x"0F";
				when x"3B7" => DATA <= x"00";
				when x"3B8" => DATA <= x"0F";
				when x"3B9" => DATA <= x"00";
				when x"3BA" => DATA <= x"0F";
				when x"3BB" => DATA <= x"00";
				when x"3BC" => DATA <= x"0F";
				when x"3BD" => DATA <= x"00";
				when x"3BE" => DATA <= x"0F";
				when x"3BF" => DATA <= x"00";
				when x"3C0" => DATA <= x"0F";
				when x"3C1" => DATA <= x"00";
				when x"3C2" => DATA <= x"0F";
				when x"3C3" => DATA <= x"00";
				when x"3C4" => DATA <= x"0F";
				when x"3C5" => DATA <= x"00";
				when x"3C6" => DATA <= x"0F";
				when x"3C7" => DATA <= x"00";
				when x"3C8" => DATA <= x"0F";
				when x"3C9" => DATA <= x"00";
				when x"3CA" => DATA <= x"0F";
				when x"3CB" => DATA <= x"00";
				when x"3CC" => DATA <= x"0F";
				when x"3CD" => DATA <= x"00";
				when x"3CE" => DATA <= x"0F";
				when x"3CF" => DATA <= x"00";
				when x"3D0" => DATA <= x"0F";
				when x"3D1" => DATA <= x"00";
				when x"3D2" => DATA <= x"0F";
				when x"3D3" => DATA <= x"00";
				when x"3D4" => DATA <= x"0F";
				when x"3D5" => DATA <= x"00";
				when x"3D6" => DATA <= x"0F";
				when x"3D7" => DATA <= x"00";
				when x"3D8" => DATA <= x"0F";
				when x"3D9" => DATA <= x"00";
				when x"3DA" => DATA <= x"0F";
				when x"3DB" => DATA <= x"00";
				when x"3DC" => DATA <= x"0F";
				when x"3DD" => DATA <= x"00";
				when x"3DE" => DATA <= x"0F";
				when x"3DF" => DATA <= x"00";
				when x"3E0" => DATA <= x"0F";
				when x"3E1" => DATA <= x"00";
				when x"3E2" => DATA <= x"0F";
				when x"3E3" => DATA <= x"00";
				when x"3E4" => DATA <= x"0F";
				when x"3E5" => DATA <= x"00";
				when x"3E6" => DATA <= x"0F";
				when x"3E7" => DATA <= x"00";
				when x"3E8" => DATA <= x"0F";
				when x"3E9" => DATA <= x"00";
				when x"3EA" => DATA <= x"0F";
				when x"3EB" => DATA <= x"00";
				when x"3EC" => DATA <= x"0F";
				when x"3ED" => DATA <= x"00";
				when x"3EE" => DATA <= x"0F";
				when x"3EF" => DATA <= x"00";
				when x"3F0" => DATA <= x"0F";
				when x"3F1" => DATA <= x"00";
				when x"3F2" => DATA <= x"0F";
				when x"3F3" => DATA <= x"00";
				when x"3F4" => DATA <= x"0F";
				when x"3F5" => DATA <= x"00";
				when x"3F6" => DATA <= x"0F";
				when x"3F7" => DATA <= x"00";
				when x"3F8" => DATA <= x"0F";
				when x"3F9" => DATA <= x"00";
				when x"3FA" => DATA <= x"0F";
				when x"3FB" => DATA <= x"00";
				when x"3FC" => DATA <= x"0F";
				when x"3FD" => DATA <= x"00";
				when x"3FE" => DATA <= x"0F";
				when x"3FF" => DATA <= x"0D";
				when others => DATA <= (others => '0');
			end case;
	end process;
end RTL;
