-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "69AD0A038EAFFAA494D989FC43493C9349217FDC4999176122F3FCE50FAFF354";
    attribute INIT_01 of inst : label is "621A4B0F756E8DF9FFFCD8112C2901E7692495574C9724E9BC93CB3D74DA466E";
    attribute INIT_02 of inst : label is "58344EFC08D139F1A277E34842A98B338CB4F43090000DBBF1A41520F6127C83";
    attribute INIT_03 of inst : label is "333A333A333A333B3F7DF7D345900008689DF8D13BF02344EFC183C5E2F0783C";
    attribute INIT_04 of inst : label is "1E19419E76208F557B22F400E64CFF4620FF800036F03435F77761A6333A333A";
    attribute INIT_05 of inst : label is "0218E9ED555223382C80178B2005D03BE392ECA12AC2633502000001C19D04EA";
    attribute INIT_06 of inst : label is "0298251EB79FFF7DF9B9FE761D875DBF3607B65F65B651E35F967C9360100804";
    attribute INIT_07 of inst : label is "62193ABD41832EC196E5437C0CB7FFCF9A7FF4DFA59F592C5FF9334E9951D300";
    attribute INIT_08 of inst : label is "798F19E4F6E9377499FC603ACE1AD0D742658A9A9B0B5C7234CE649098A13108";
    attribute INIT_09 of inst : label is "B5684A0000000042B1298D216CF2568D13944E11A2728980344ED0A99A421556";
    attribute INIT_0A of inst : label is "ADA691B458AED52473446777B60CCCC99910CEC2D84162B3374C8526C5407F7F";
    attribute INIT_0B of inst : label is "BEE38E39F5C44C6431B3343091DE53366FB3646C9864C606490DA4993A491100";
    attribute INIT_0C of inst : label is "F4CF8270FEB0D0D4D563CBF0CAA862F0F173337B498B2498514A1FD78E6FBF6B";
    attribute INIT_0D of inst : label is "1EADDFD1EADB8D0A429036032BCF019FCDAA228BE3F1DBB7ACBC34D5563B379F";
    attribute INIT_0E of inst : label is "FFFE0000000000000000EE91D737DF1F7ED1D1FFFCDB668E8DC6C8CABDD5FBC7";
    attribute INIT_0F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "D896822A853189EA748A06B8C30BA1092DADAD1B7856FD4D90C38EB8C30BA109";
    attribute INIT_11 of inst : label is "0000000240001C18600000000082910960279BC2842C0280BD8EB0EA1AF42129";
    attribute INIT_12 of inst : label is "0625138B6052ABA8CB8000000067A00000001EC162C5498E8A002C000007D109";
    attribute INIT_13 of inst : label is "4C0602C0701C42008460180E0B84603C0500C12008120000D3384BA69045F101";
    attribute INIT_14 of inst : label is "C67054740788C2FC8D02C0500816100541681A1782116C8C07038EF011F71109";
    attribute INIT_15 of inst : label is "6F1382E1B80E1B81C5079479450BD0028200000000186165FDD5F5777755D109";
    attribute INIT_16 of inst : label is "1000645804458064300643A012419189A79450BD0505141E1C56DD4D3CF2A189";
    attribute INIT_17 of inst : label is "1AC0B1080A020838186061E1C40030471000645804458064300643A004003047";
    attribute INIT_18 of inst : label is "3C8E07946258962187945CC72DC107940715C47118560580200A08AA2AA20109";
    attribute INIT_19 of inst : label is "014514358143143396396030D63814338EDAE850CEDAEDAEDAE850CE9AE9210D";
    attribute INIT_1A of inst : label is "01451441259229229213B6396030D63814338E58E050CE58E58E58E050CE18E1";
    attribute INIT_1B of inst : label is "FFFF404125922922D32D32CC32C3210914338E58E050CE58E58E58E050CE18E1";
    attribute INIT_1C of inst : label is "500C370E060CE78E62E878CE7A0E3780EB7B6FAEABCAAAAEABAEBACEBAEB210D";
    attribute INIT_1D of inst : label is "FFFF4000000000000000FFFFFE2BF41FE7D1FE7D1F47F9FEF8C50BD00BB4E0D3";
    attribute INIT_1E of inst : label is "FFFF4000000000000000FFFFFFFFFFFFFFFF4000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "A9FE2800000000000000FFFFFFFFFFFFFFFF400000000000401EC0B082F04DE0";
    attribute INIT_20 of inst : label is "730469CC767B21096B2ED00828FFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "67AAF59A8C4426A856B3D57AED462215B67AA9EB351A880ED67A699EB3635205";
    attribute INIT_22 of inst : label is "BB0FC9BC9B5E64A59AB763D925926BDC94F756EF618A6E53327272C13988906D";
    attribute INIT_23 of inst : label is "F15D5BA054212002B18000003E4D649AD6B410F9293EADDE7E4D649AFF2537D5";
    attribute INIT_24 of inst : label is "BFB41804E7B44004FFB40004FFB4000FEDEF3E298E397E764D56191875499721";
    attribute INIT_25 of inst : label is "842652C23FFE6F2BE60000106C69208574E80A512848304170BF168B5A208AF4";
    attribute INIT_26 of inst : label is "32FCC00A2CC0023C701377B073F64F003875996C97734FCF6A30600364EE90F4";
    attribute INIT_27 of inst : label is "E0A983889E1E61A08869430E2923CC304D0B2182A60E227879868221A687188A";
    attribute INIT_28 of inst : label is "FDF4D31CB97FEA479BAB7BAF1C72E4D32BE27471123CC304D0C38A48F30C1342";
    attribute INIT_29 of inst : label is "D1DB9D98352DD9C6EE0F9CB1D43E83A554CCCE90350DE663A0A733880E46A0E6";
    attribute INIT_2A of inst : label is "30C5599BD2D8CEE90506E35BC89C131CC31E9B66A8FF9CEA64C350E6C294A74C";
    attribute INIT_2B of inst : label is "AC96400FFC94D5651D744777B0DB68D8C77F78144E9FCF3BFF36CC9CFD91A154";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000009C9BD81FEF379";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "51851501470E896823406861427FFFFFFFFF0000000000000000FFE35CEB3505";
    attribute INIT_31 of inst : label is "E5261693AC3D29932D4534826609A469228122A101EB8ACE608410286ADB2243";
    attribute INIT_32 of inst : label is "FC8AAB5E5635EFFF60CEE0D619D244D893A50AD2900F0952EEA9C7CDC8DD9ED2";
    attribute INIT_33 of inst : label is "45923950ACBCA333328CCCAACF083BD5FC3478A07C7A55418043F803487F1FF3";
    attribute INIT_34 of inst : label is "A28486A383CE5BFB7515B7FB32CC91254E53DBCD4F5325646CCDEA1414592391";
    attribute INIT_35 of inst : label is "E5089147315A20B1B8D4D5C5057EA1D197C6F138826500844EA000A2E6FD5144";
    attribute INIT_36 of inst : label is "A10C29966474F18B032186066AB063EC6668B8AFE19C04E863F001FE70008A79";
    attribute INIT_37 of inst : label is "CEB906A33F5C5A11E1212031566D65FA1FE5C8E7CB983E5BD2BE4C36A02D8D0A";
    attribute INIT_38 of inst : label is "00B852E14B802E14B802E00B852E00B852E00B852E14B802E00000BB23FF6C35";
    attribute INIT_39 of inst : label is "FFFF0102000301560000FF8100030333FFFF00010002001204004004010B802E";
    attribute INIT_3A of inst : label is "FF800002030101300001020201030131FF820002010301100000800301010377";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FF82000201030331";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000002000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "B1F7F299905001485D59D6487A0089460084C004A611A7EC86DE806DC4F07532";
    attribute INIT_01 of inst : label is "6651802248491AF6457F8281B64528C0DE71E7AEF7FDFF46BE43E43FD21D6A93";
    attribute INIT_02 of inst : label is "C5BE19B73EF864DDF0CD96FB1D60C50BD1D2154500000319A8E182FD47FB5B73";
    attribute INIT_03 of inst : label is "81BD81BD81BD81BC2596596CEF7000037C3366F864DCFBE19363108844231188";
    attribute INIT_04 of inst : label is "425C89AE036A46AB905FA1D80EC4AA85F7FFD0002A47681E22A2B8E181BD81BD";
    attribute INIT_05 of inst : label is "0E08B08808BA005E75D0169D70049A064058249237A780F80E000003009E0822";
    attribute INIT_06 of inst : label is "0051A7AFBDE002491111010CC336E4400C908C90CC8C9058EFB61105A030380C";
    attribute INIT_07 of inst : label is "19199B34AC996E5CE75F7CB644D3FC2A680011209B64928DDB6E88F0547CBC00";
    attribute INIT_08 of inst : label is "00E9D01364300413506E32078EC1AEC4AFAB22E3DBED60E1B0484A9B98C51C88";
    attribute INIT_09 of inst : label is "2FD7FE0000FEEEAFFF405BEC4A01C76F864EF87DF0C9DF0DBE19BB5737D8EB3D";
    attribute INIT_0A of inst : label is "59486870E1F8A1C35DBE952687C206A0466F8F93323387E0A02A7B38F9F2120A";
    attribute INIT_0B of inst : label is "AAC638E09B088AA9C56C1544255068202B152AB12D493534729148D1AB86F7AC";
    attribute INIT_0C of inst : label is "0B4050EF35C005010C7C7808C5F7FF6030E1116994246DE3AEBD716FFC592962";
    attribute INIT_0D of inst : label is "577B303556BEABFDEFFF93939C00F681DFDF77C5E70502ED576A513FFAA15AB8";
    attribute INIT_0E of inst : label is "FFFF0000000000000000D969FE4804E01366EE0002000915508A1131227E0B95";
    attribute INIT_0F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "1FED139D1E13402219B300AA0A2E3801D050D041C70C6E10828AA0AA0A2E3801";
    attribute INIT_11 of inst : label is "00000000800022220AA8A8A88A82A801A6B8420038B868020020A28A0280A801";
    attribute INIT_12 of inst : label is "010330EC11310310D08000010102E0000000421250A1D8508600120A80820805";
    attribute INIT_13 of inst : label is "0C03038431085A1285210805118010300500416058060082A3408A2800809801";
    attribute INIT_14 of inst : label is "C8B20CC82F0470540119C10110141081715C5C0B02F19C10000418E200862805";
    attribute INIT_15 of inst : label is "85340F02D8B6358D80282002003E030A82A22A2A2AA088880A02202000000805";
    attribute INIT_16 of inst : label is "220088420886A088200A8221AA82A801002003E0383820603899E11C71467805";
    attribute INIT_17 of inst : label is "124290082AAAAAA2E28A8A8ED882A1A8220088420886A088200A82219882A1A8";
    attribute INIT_18 of inst : label is "B00803850140500403856018120483855812048044490044298A802AA0A29801";
    attribute INIT_19 of inst : label is "00AEAA8620AAAA82A8AA882A0AA20A82A0E2086A00C20C20C2084A00E20EB801";
    attribute INIT_1A of inst : label is "00AEAAC0CF2CA2CA2C8228AA882A0AA20A82A2EA286A02CA2CA2CA284A02EA2E";
    attribute INIT_1B of inst : label is "FFFF0040CF2CA2CA4C12C1304B04B8010A82A2EA286A02CA2CA2CA284A02EA2E";
    attribute INIT_1C of inst : label is "4200862086A02EA2EA086A02E20286A008638C20A609A69A46186138E38CB801";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE2A00E0A8000A8000082A00800C064206058000";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "C6AB9000000000000000FFFFFFFFFFFFFFFF0000000000007DC1024F900FB21E";
    attribute INIT_20 of inst : label is "8721E40FDF67A7B7D492FCA1BF7FFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "A87D8EE056D2FBF5F1D43EC7702B697F8C07501D40AFA5BE3A07B681D425F66B";
    attribute INIT_22 of inst : label is "3020004004AF2CC849260600080095E5996924C0D7FFC0CF767661CC85F1D363";
    attribute INIT_23 of inst : label is "1CE3F2F4DC4298CB27098889400200253C6BC9EB321A4981000200257D665349";
    attribute INIT_24 of inst : label is "D9A081A0FE30A635418541853E153E1048085E962AAE816ED2A83B3AC77F2C88";
    attribute INIT_25 of inst : label is "C7A82125FFF3B037170002DF6F96FBEEEFDE9DB773F6BA6DABC3BF9F9F3E7700";
    attribute INIT_26 of inst : label is "AD8EC2DDDEC2D5DE8098551BF408A1B9C98B62916F848000DEAF4634A6A918F8";
    attribute INIT_27 of inst : label is "ED3D55D4544760AA908B55226A11EC1250534AB4F55751511D82AA422DA85071";
    attribute INIT_28 of inst : label is "820B2C5743C01C56543716039E4364240CB55233351EC12555489A847B049414";
    attribute INIT_29 of inst : label is "9E4A199F84A48DBE1F296CC55CFF7A7ADAAA8213A6291545D7D6A7BDAEF4FA90";
    attribute INIT_2A of inst : label is "FEFBFD0B4DB5AAFBF5E2DF3FDB410086FE6F55D8DA9FD73BDE8A6A94FB7F73AA";
    attribute INIT_2B of inst : label is "596C8C70166188629EFD88663A1B7E67FE4D472AB5AB545265D94CA102AA56FB";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000001F461DC04A492";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "BBD1B6F6AD19FED138221606B0FFFFFFFFFF0000000000000000FFE014020081";
    attribute INIT_31 of inst : label is "F42E3B28DBBF9E1399FB6F7376165A7EF675F2FFEA58092175F7BA761DC7DDAC";
    attribute INIT_32 of inst : label is "54DFF8A16B5A8FAAC571A67919CC635FACBF5339EEFFFE2155DA88D3854C9A42";
    attribute INIT_33 of inst : label is "1621203BC90EF59333D66EDFAF1FAB1A03FF7FAB047EFFECC8420DCCB4AA9543";
    attribute INIT_34 of inst : label is "A04E2DF3D4407EE9A26A07FCA85D8AC084AB4D4085A3BF228445A3E796112116";
    attribute INIT_35 of inst : label is "42D5A96AEBF5F36C7F6E0839F781DEAA6A2BCD8315C2B510BA56A2AF0901F025";
    attribute INIT_36 of inst : label is "A71FF753A81B3312185714B98D3A7C11DFB157781182AD1C945B9954C293654E";
    attribute INIT_37 of inst : label is "3A42A29C4121995304E5DA4112A28AE9DBFF7DBD7AF9ABD7B31354BA12BA1F31";
    attribute INIT_38 of inst : label is "400150040010005401500540100040015005401000400100041F82C200AAB51A";
    attribute INIT_39 of inst : label is "FFFF09C9490808320000FF89C9084835FFFF00098988C8151241451253001500";
    attribute INIT_3A of inst : label is "FFC949C948C888560049490948488877FF89C909C80848F60000C9894888C813";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFC9C94948C84857";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0800000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "0800000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "D902A4BD0C10B8705451C565D7400CA840007FFD41442068000A822D815F5580";
    attribute INIT_01 of inst : label is "223A020A514A0C9D674E3E81842608E1104904148765D96A28A28A2A555253FA";
    attribute INIT_02 of inst : label is "8AA55A5A2A95696D2AD2D59294156300BD00017D00002FD0EF6230A554957D21";
    attribute INIT_03 of inst : label is "BFD9A659A659BFD89EFBEFBE0D00002B4AB4B6956B78AA55ADB25128944A2512";
    attribute INIT_04 of inst : label is "02E184A034209F13DD2730898A817B8AB2AA800038D23274BB332F61A659BFD9";
    attribute INIT_05 of inst : label is "020828A1C1C2400B3990264E60099048449C2849F6F764668600000140850424";
    attribute INIT_06 of inst : label is "03EDB2FF39CFF36D9DDD835ED7A6ACFF1EBB9F91EC9F92F3EFA61506E0100804";
    attribute INIT_07 of inst : label is "D18809194810E80865D1347060D6AA26B0303DB7E1B6DB009FF01A87EC542100";
    attribute INIT_08 of inst : label is "7D756DB7BE781A32A8BFD204268F94144C8C29D212517A9904022C53140579C4";
    attribute INIT_09 of inst : label is "BA0B42000048200A5685564AF6FA84A95E90EA552BD2150AA57A42952C94A0A1";
    attribute INIT_0A of inst : label is "ADFC55E29542FFF7F6D6F31324AAEBDD5BD2A690575A550AFFF5A5BE9113F97E";
    attribute INIT_0B of inst : label is "D81DF7D8610CE4CF56D1816C26D6700004020EC561BFBB3A7FBDFC68DBE50911";
    attribute INIT_0C of inst : label is "30C320AC1D68D5150D49D9DA828D489397108032DAA84922804153AD27EDB9B2";
    attribute INIT_0D of inst : label is "6AD67BE6AD77365294A5071A160301863484CC4E14A68A7BF8C661006C90EA25";
    attribute INIT_0E of inst : label is "FFFE0000000000000000C4FD79224D4935BFBF124A492DDDDC0C4199B7AAF852";
    attribute INIT_0F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "12559B119407808C191002A0A8A8A1107FFFFF9EEA7495DF8AA80AA0A8A8A110";
    attribute INIT_11 of inst : label is "00000003C0002A28288882A2028A811080900A00128880080282AA2A2A8A9510";
    attribute INIT_12 of inst : label is "041110C840110B3C0900000000B4C00000202BD12C5858D2C800660AA800B110";
    attribute INIT_13 of inst : label is "30450004D0300C1300C1301A1CC03004060080A0280A01C321F0A2A200A22110";
    attribute INIT_14 of inst : label is "07A1B03A040320841C1404907C3010C32138571C07C0E002008302AA380AA110";
    attribute INIT_15 of inst : label is "311B44D1384E038002A2802802A0AA02A2808A82222828A8A282820A2A2AA110";
    attribute INIT_16 of inst : label is "AA2220EA228C0228802008A20A00011002802A0AA2B2A00A4B220A0002898110";
    attribute INIT_17 of inst : label is "15C1701408228A2A4A29282C5A888200AA2220EA228C0228802008A21A888200";
    attribute INIT_18 of inst : label is "440F0FF2B12C4B028FF2641916458FF2091244910C7300C4012808282AA22110";
    attribute INIT_19 of inst : label is "2384180CA38018081A81A880380A38081ACBA8C03ACBACBAEBA8E03AEBAEA110";
    attribute INIT_1A of inst : label is "23841843841819819808BA81A880380A3808184180C0384184186180E0386186";
    attribute INIT_1B of inst : label is "FFFF004384181981D84B84A02A02A1103808184180C0384184186180E0386186";
    attribute INIT_1C of inst : label is "883A8ABB8A0382182BA8A0382A380A03A8AA28BA9826186138E38CA28A2AA110";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE280AC00002000020A8000A81A8188A38882388";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "E37C9800000000000000FFFFFFFFFFFFFFFF00000000000063FEFFFF7FF1FFE3";
    attribute INIT_20 of inst : label is "4A0224C9444A242242A890A11D7FFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "6980353EAD54A5494530C01ABF56AA522818006A7D5AA940A6186186A7EB5452";
    attribute INIT_22 of inst : label is "8FD07E67E714CA5431B1FA0FCCFCE2894AE2363F4250BF91454542849D23920A";
    attribute INIT_23 of inst : label is "CA96020488E2B049A74CDCD943F33F38A4858D32950C6C7E83F33F38A652B18D";
    attribute INIT_24 of inst : label is "799079905F805F805E005E0078107810C92B429B26947D08D005E222826128E8";
    attribute INIT_25 of inst : label is "730752A40009FFB6650000184901048150291A032B003B6CEAA13A9D122A7CB0";
    attribute INIT_26 of inst : label is "9FC02089F02089E2D248002A961AE01979AE2BD5C8BFC7B66895362FC2474E0A";
    attribute INIT_27 of inst : label is "8A2197DDC848132A106B57264A160263545A2B28865F7721204CA841AC2FCB7A";
    attribute INIT_28 of inst : label is "8BFFB74A250228944F3238FC0000C07F26B732D23560263555C992858098D516";
    attribute INIT_29 of inst : label is "54B09112439800D4F1E6D274D8C1A9414E665E07D324D33F6A1494294A528252";
    attribute INIT_2A of inst : label is "A49054819648E4362D406A6C5B75AB89977DC82CAA51C9918A49B25292A84AE6";
    attribute INIT_2B of inst : label is "6FB7EC5BD4315844E28C6751A8D2481A9112122553E4924895FDE8B40D812546";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000AA405E4CBEDF";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "A109150C30610459B432D4C426FFFFFFFFFF0000000000000000FFE0A4561B44";
    attribute INIT_31 of inst : label is "44052DB565025080A8D048205448A049048CA0690079DA2761852414D0D48560";
    attribute INIT_32 of inst : label is "A82AA55FA188005565AA85535010041291B429A501AA5037323E62046D840CC0";
    attribute INIT_33 of inst : label is "E22A00928690001280006A75201C414D4141520EB90C8D52C0421D8CDCD582A0";
    attribute INIT_34 of inst : label is "049BA9505E1A2D1093DB655F91D15B0CC7B0C4CCC6B29406C200C9A57833811E";
    attribute INIT_35 of inst : label is "6422864511800238C7FCCCD4A50295B339575C9B16202110C604322D7FFD4240";
    attribute INIT_36 of inst : label is "261DECD56AEDBA19954492A22AA5402719F9CAAF950045C8EB5398AAA012289B";
    attribute INIT_37 of inst : label is "A5B221FC56DDAF6200201033FE9B6F7BDEBBF0F9F3EB9FBCE9BB54B8B23F9A11";
    attribute INIT_38 of inst : label is "D5BB06EC1BB06ED5BB56ED5BB56ED5BB06EC1BB06EC1BB06EC1F8B07AA01F55F";
    attribute INIT_39 of inst : label is "FFFF00048004005A0000FF84000400FDFFFF00048004807C0A080282003BB56E";
    attribute INIT_3A of inst : label is "FF840084008400DE000480040004807FFF840004008480FE000080040004807B";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FF8480848084005F";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "EDBA183A9410A8426840C32C1B600C826014540EFDFC102016104183C4108100";
    attribute INIT_01 of inst : label is "547A04A80900500500021A01BD06A0324A28A9D751F47D60740DC0F7416B0DED";
    attribute INIT_02 of inst : label is "AB97664A2E5D9B2CBB32502084072208420850880000380D4BF0B08C0E44AC0A";
    attribute INIT_03 of inst : label is "000019800000000232CB2CB15900003D2ECC965D9B28B9766CB2552A954AA552";
    attribute INIT_04 of inst : label is "5063EC200887589201A40AB5CE664832AAFF3000094ACB6200808BF019801980";
    attribute INIT_05 of inst : label is "020820802082519A3080020C20009050451E220036A60561060000010344004D";
    attribute INIT_06 of inst : label is "00DEFA314A250924CCCCC2769DF9AC68769936E77A37E8C4D79A0D04E0100804";
    attribute INIT_07 of inst : label is "777F92FD41B37C59AD871545468FFD0DB00827D520B2CB5F6DB812D09FC8B400";
    attribute INIT_08 of inst : label is "4F0F1DA5DEDC1E2AF8D2FB96A307D72D4AA10550E960773DCE39DF617CF2AABB";
    attribute INIT_09 of inst : label is "974B4A000049355852A70082FC9E72E5D9B58A5CBB36B14B9766569101042014";
    attribute INIT_0A of inst : label is "AC775F1AD5EA3A7CEF5726FFAAE979EF1D92EA29D1CB57AE7A6EA50E587149E5";
    attribute INIT_0B of inst : label is "4612CB2CA044466619F1109925C44082A472AD045B6EB6B71DE8765CB0C58065";
    attribute INIT_0C of inst : label is "2481A005487254D5B6650CA91AA52FB3A7D139FACAC22CA88049148793249C9A";
    attribute INIT_0D of inst : label is "D8866A7588612E1084A5ED71F7020103B2E44C5A01C59818E8863C00493F660F";
    attribute INIT_0E of inst : label is "FFFF0000000000000000E4A3A1324DC9371515924E4938888CC4D28896A89C27";
    attribute INIT_0F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "80414549538B40E6243B828222AA860CD9D9D9D2CE94D0598AA2228222AA860C";
    attribute INIT_11 of inst : label is "0000000280002A2820A0A0888A02260C24200A00822A0080200288A80A02240C";
    attribute INIT_12 of inst : label is "001000080003CB91078000060061E00000001F90000151DA8E000E000080A00C";
    attribute INIT_13 of inst : label is "60081240100404010000008000C0720C000000220802000831502A8000222008";
    attribute INIT_14 of inst : label is "02E0402E04C4215C00100401105000052018140E0100800A02858A880800840C";
    attribute INIT_15 of inst : label is "27118461084210850290000002AAAA0880A2220A0A0828A8A2A2808A8222240C";
    attribute INIT_16 of inst : label is "2800800A0A0020A8600886A02882240C00002AAAA2A2A0000228A2082AAA240C";
    attribute INIT_17 of inst : label is "004011042B0A28A888A222204A0220A82800800A0A0020A8600886A00A0220A8";
    attribute INIT_18 of inst : label is "4C4C1380010040101380340D034493800D0344D11C0711C4280AA022A022A408";
    attribute INIT_19 of inst : label is "8028A280A02EA28622E2286A00EA0286228A280A028A28A28A280A02AA2A860C";
    attribute INIT_1A of inst : label is "8028A2C008A0E20E2086A2E2286A00EA02862082080A0082082082080A00A20A";
    attribute INIT_1B of inst : label is "FFFF004008A0E20E402A02A02802866C02862082080A0082082082080A00A20A";
    attribute INIT_1C of inst : label is "0202008280A008208A2802008A008020280AAAA2E218E38CA28A2AAAAAAA860C";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE2A0A000828008280A0020A802002880280A000";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "DB04F000000000000000FFFFFFFFFFFFFFFF00000000000042203F00FD000201";
    attribute INIT_20 of inst : label is "4B3A566C8761D569460AD9D9457FFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "488211B2D9C6B4E96DA04548F96CE35A6E08A82365BB0D61B40849023657615D";
    attribute INIT_22 of inst : label is "5B14586586305D4415CB628B0CB0C61BA8E6B96C495848DABEEABBCCC99A6A9B";
    attribute INIT_23 of inst : label is "02531A876B59D76DCA999A8D22C32C31D424BBB7510D72D8A2C32C3186EA31AE";
    attribute INIT_24 of inst : label is "A1B5A1B580258025A7B5A7B5A035A0389461E0D92C31D218E84A35FFEBAD1C60";
    attribute INIT_25 of inst : label is "84A29CE20000C92C5300008925C0A68F10653062916430C2C4D11349DB455A85";
    attribute INIT_26 of inst : label is "B66D5E8D6D5E8D60A492F5A6BD16D375696D5B0D80A642492DB76FB65CE23081";
    attribute INIT_27 of inst : label is "8BCC869BDE3AEFA90FD9C63D79EF5DF2CC1EE3AD321A6F78EBBEA43F618D5D5C";
    attribute INIT_28 of inst : label is "0D4CB218FC398793199FE427716E9416322679FA32F5DF2CF18F5E7BD77CB307";
    attribute INIT_29 of inst : label is "E6F6CD8B5FF9CBD6AF0C91E192C0CBE944ECC449310C67632A9BB40D647632F6";
    attribute INIT_2A of inst : label is "97DD71EFDFEFCD002C7BEB600530B486D9349EFE34E09FC5A0F39EF6D8DD6A4E";
    attribute INIT_2B of inst : label is "66B35F5A688ED8CB818276A97DAFAF72DBDAFA3566ADA79EDA65853D4922A552";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF000000000000000B555433291ACD";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "843061A524C82514552AD2E5967FFFFFFFFF0000000000000000FFE21CC12009";
    attribute INIT_31 of inst : label is "B88BCD95652B5ADE001FBD2A2FC0822C1084B60D4045F82705398742C2802424";
    attribute INIT_32 of inst : label is "ACBB31280611E055758A815D2280D07B01A6B5F5A0A76A5A662AE68F7798FEC8";
    attribute INIT_33 of inst : label is "08880058F495AD737FBDC5714070842D6122FB848200059AC04D13EECAD51AA6";
    attribute INIT_34 of inst : label is "800981481020E035BD5FA80932AF8F554A7DE9954A73D7BBED67E8A9E7EAB200";
    attribute INIT_35 of inst : label is "25890C9B3552EA58C197754C39C291D51B44087F562021DEC6042BA44CA06000";
    attribute INIT_36 of inst : label is "D694DDE64125CB153B5DF682B3172E3E40CAD9AA7231584C2CA75AAB7CDADA91";
    attribute INIT_37 of inst : label is "6C98CD350248E3739232290667C92C3365E8D36AD5A1D6AD614ACA7739E3DE1D";
    attribute INIT_38 of inst : label is "14045011404501000400100040010004001000400100040010002C11A7FEDC93";
    attribute INIT_39 of inst : label is "FFFF0004848080800000FF8484808083FFFF0004848000A20828A20A2AA04501";
    attribute INIT_3A of inst : label is "FF8080848400008400000084840080A5FF8080048400002400008084848080A1";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFDFFFFFFFF0000000000000000FF80000484000085";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFD7FFFFFFF";
    attribute INIT_3D of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFDFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFDFFFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFDFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "493214BC1354A5409E11E4014EA8100AA81695568E9799C117302BB98855580A";
    attribute INIT_01 of inst : label is "A554C6B10A215A95444A1540976EA8C50000049D856559282882080205034A4A";
    attribute INIT_02 of inst : label is "CB0200962C0800481004B4B290A0100EC2335B0A10000110A2840A95044C801D";
    attribute INIT_03 of inst : label is "E67FE67FE67FE67D56DB6DB26C20000004012C080249B0200922190C86432190";
    attribute INIT_04 of inst : label is "60E1EEE10052028B549622900206AA15CFAA1000214A6A13A22AA287E67FE67F";
    attribute INIT_05 of inst : label is "3A28BEF8901313FC0C5F7FC313DFCA97E942FCD9CB4E89E88F80601DE0120F2D";
    attribute INIT_06 of inst : label is "018ED2346325536D9DDD9335EC606D6AF5F9F1871BF18C9690506312E0502874";
    attribute INIT_07 of inst : label is "3702A8D26932DA1973061091C02AAA743065289551B6DBC7692110018B8C0000";
    attribute INIT_08 of inst : label is "18244A012419102240A8A22435079F0068052AD2503F8A95C5200F79304B1B82";
    attribute INIT_09 of inst : label is "200D64000065A66B5AA032DA403034408806A2581100D45B02209ADC25948520";
    attribute INIT_0A of inst : label is "156048228542B5605249634A50408080101B34A41008100024E4368C88383648";
    attribute INIT_0B of inst : label is "DB210410402EF4CC94ADDB98E4C02B4A55060F16412C129258C1614A92E4A120";
    attribute INIT_0C of inst : label is "200100A4186ED5700045048D3334C4652AAAA8A4DAAA4002166DC185176DB3BB";
    attribute INIT_0D of inst : label is "49CE53449CE326318CE7E550570A00229017777400E4B939C1CE7CBFAA1A2407";
    attribute INIT_0E of inst : label is "FFFE0000000000000000CDB83B66DF1B7C373736D8DB6199980DC999B52ADC02";
    attribute INIT_0F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "014DD3011202E0AC1353020888AA04E46666E6DCB6EA959E0A888A0888AA14E4";
    attribute INIT_11 of inst : label is "00000000000020A8888A82A2028894E486804802A08082F0A00A0221C80084C4";
    attribute INIT_12 of inst : label is "003000300200080C5480000280122000002002D250A084005200500AA80284E0";
    attribute INIT_13 of inst : label is "4848008060181300C1701C9524080030040189D0741D20C3010080808280A4E4";
    attribute INIT_14 of inst : label is "010088150904410003194531446910C2C06009004070141906400A23D08224E0";
    attribute INIT_15 of inst : label is "101C4711D4751D44202000800AAA2A0222808A82A2222A088880A2220A0A14E0";
    attribute INIT_16 of inst : label is "03DC032BC0B29C2B01C2309C020094640800AAA2A2A2A080082082082AAAB460";
    attribute INIT_17 of inst : label is "1F87E0100020820A0A2828A8C0F08C0003DC032BC0B29C2B01C2309C00F08C00";
    attribute INIT_18 of inst : label is "9040100000C05014100040500C0510005004000160281604082820A8822A84E0";
    attribute INIT_19 of inst : label is "3C020042BC00004082882F01020BC0408A28A7210A08A08A28A7210A08A024E0";
    attribute INIT_1A of inst : label is "3C02005C02800800806082882F01020BC0408A28A7210A08A08A28A7210A08A0";
    attribute INIT_1B of inst : label is "FFFF005C02800800C028028022023484C0408A28A7210A08A08A28A7210A08A0";
    attribute INIT_1C of inst : label is "09C8C22AF210A28A2AA7290A29CA429CA428228A0A028A2AAAAAAA8A28A224E0";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE080080A0020A002008280A00882A83CAC0BC8C";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "C4AB5000000000000000FFFFFFFFFFFFFFFF0000000000005E3F7F10FDEE42FD";
    attribute INIT_20 of inst : label is "02288648C04201A00AA80DD9847FFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "08A21530C1A4B50B6800510AB860DA5A400A202A61836B69400A0802A6106A58";
    attribute INIT_22 of inst : label is "F0D0D26D06508068A11E1A1A4DA0CA000D7023C342420294C8585A8CC9188010";
    attribute INIT_23 of inst : label is "8A12E27D8A4D1E4D722AA9BB0693683280A6B9201A2847868693683284035508";
    attribute INIT_24 of inst : label is "064A064A27DA27DA27DA27DA205A2054D5E660C98614558081500204022C0118";
    attribute INIT_25 of inst : label is "0146843000044A08410000484089365864C9D242A169D8B18849E35191A6581A";
    attribute INIT_26 of inst : label is "9409928D71138D62802100A2A694D613714D5349A8B6C2B66C972276EA662100";
    attribute INIT_27 of inst : label is "8925C71C4C80803D2E0DE6A049F198034C9A1326979C71321300A43822CE0A58";
    attribute INIT_28 of inst : label is "484D93082C2042168B36146C20A100926747222B33110076F1A8337C4401DB06";
    attribute INIT_29 of inst : label is "428510414855068931C5BF40C0C189408C664F411BA4D2276650946D6232105E";
    attribute INIT_2A of inst : label is "620880C520160592983144A56B01E0A00BB5CA001A5108118A493042084842E6";
    attribute INIT_2B of inst : label is "6D3684DB5084AA9A60063048050007010E85A1332387024C2424A2340800359A";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF00000000000000140046100D34DA";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "82192494B0E014DD312210A480FFFFFFFFFF0000000000000000FFE280D239CC";
    attribute INIT_31 of inst : label is "CCC819B1D2180024A808001C40AA2505223C9404DD0232882C35A75081109440";
    attribute INIT_32 of inst : label is "AC111D4C0021105585820809A794B531540293000792303632B87CBA85D4694C";
    attribute INIT_33 of inst : label is "0000888C4DB8C62AEB1882D43091C618508451C80BA4A5D8C0CE509EDCD52AB0";
    attribute INIT_34 of inst : label is "9A70245C32382460938B6D5319F70B0CF63F448CF6B01202EAA2908580000888";
    attribute INIT_35 of inst : label is "6C88084C2201C678809CECC41592D1B331457801B644E73ECA9CA38444A969AE";
    attribute INIT_36 of inst : label is "661EE4B00264B3351D1CF2AA29020420084988B21A60CB8FCC413AAB949271B3";
    attribute INIT_37 of inst : label is "25B06C9332DCC92344848255101967682EA9D2E9D3A9CC9CE9DCAB4565019A91";
    attribute INIT_38 of inst : label is "1404501140450114045011404501140450114045011404501140300381545083";
    attribute INIT_39 of inst : label is "FFFF7581418181240000FFB141919125FFFF003161A1C1258FB0CB8D37C04501";
    attribute INIT_3A of inst : label is "FF95F50121A1C1000055951191A14101FFB5C5B10191F1200000F511E1A11105";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFA5C58131818101";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "0000000000000000FFFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "DA3296BC57536D6CBEE1EC414CD2791BC236FA509024567036E1A63395A97B0A";
    attribute INIT_01 of inst : label is "154617B80700D1F598FA5010B37FA985210414990D63589BC1B41B402DA348D8";
    attribute INIT_02 of inst : label is "91C22583E708960E112C1EFA52582359880E3520A000002220052ABD284DEC98";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFDAD92D9222CA00001844B0708940F9C22503EB2492C924B24";
    attribute INIT_04 of inst : label is "6B7AEDAE546290CA26144C95112C0C405BAA10000C6A4F5244C46007FFFFFFFF";
    attribute INIT_05 of inst : label is "360830C0A0A303CC001F030003C0C200E0006000020200200380601B8000083F";
    attribute INIT_06 of inst : label is "018ADAB6F7BE96C937550D84C16C1474849E85B45B85B906B07C20A2E030186C";
    attribute INIT_07 of inst : label is "1144CDA42B34C99A6A13B2705162AA282084C9BB4534D34A0928210D8B8A4300";
    attribute INIT_08 of inst : label is "18244A000019306A418806286E1F8EA22854A8CAD0200203AC852ADB935E08A4";
    attribute INIT_09 of inst : label is "4A2D6E000065A66B5AC81BF908301C708162A54E102C54B9C2058A54F7D292E2";
    attribute INIT_0A of inst : label is "1F6948078F47B16006CE618C98400010321BAEC0880C381000E5376D8F702691";
    attribute INIT_0B of inst : label is "FAE104104098A98824A6950034C000102B448018832D1212DA13684896D4A529";
    attribute INIT_0C of inst : label is "D6C712EC9C6B605804870D89B194C64C38ECCC48012B40124B25498D176DBBF0";
    attribute INIT_0D of inst : label is "CD29948CD28B677BDE738D1457456D8E948C4CC408C480AD5528404055062746";
    attribute INIT_0E of inst : label is "FFFE0000000000000000C90202449636C826626591964113360A0111287523A0";
    attribute INIT_0F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "414D1731D20AC53E5355800222A804004040C0E0560728108AA2200222A81400";
    attribute INIT_11 of inst : label is "FFFFFFFC3FFE22A282828A8A2A282400E6206002A2228A82A028088000022400";
    attribute INIT_12 of inst : label is "011110C411125D7BFEFFFFFAFE1FBFFFFFFF84607CFBD3BDFBFF81802880A400";
    attribute INIT_13 of inst : label is "80300C0300C0300C0300C0A0200B83C0380E0B02C0B00E0001002808A8220404";
    attribute INIT_14 of inst : label is "00000000000000002010060180401F0000802000000000300C00080800009400";
    attribute INIT_15 of inst : label is "400802008020080202802A82AAA02A0828A8A2A282828A880222808A82A22400";
    attribute INIT_16 of inst : label is "2800880A0A0220A822088200288A2400482AAA02A2A2AA8002200220AA2A8400";
    attribute INIT_17 of inst : label is "080000E022082080808202004A0220A82800880A0A0220A8220882000A0220A8";
    attribute INIT_18 of inst : label is "0070100201C0300C1002C0300C071002300C0700E0001E02202AAA8208020404";
    attribute INIT_19 of inst : label is "A02AA282A02AA28222A2282A00AA02822820802A0800800800800A0820828400";
    attribute INIT_1A of inst : label is "A02AA2C00AA0AA0AA08202A2282A00AA028228A2882A0882882882880A08A28A";
    attribute INIT_1B of inst : label is "FFFF00400AA0AA0AC022022088088400028228A2882A0882882882880A08A28A";
    attribute INIT_1C of inst : label is "000A008A80A088288A80020880088020800002082A0AAAAA8A28A22820808400";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE0A0A00082A0082A0A0020000A0AA080A0080A0";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "BAAAA800000000000000FFFFFFFFFFFFFFFF000000000000401E421090E042E0";
    attribute INIT_20 of inst : label is "32A496D0A59000B024A51AB554FFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "6319E2A9A08D981338B58CF174D046CED4B112C5D341193B16B165AC553823CA";
    attribute INIT_22 of inst : label is "E4CBB7CB752D1178457C9976B96AA5A22F68AF933AD6A6B4448486AADE1701B1";
    attribute INIT_23 of inst : label is "2B1C1086085F5D4E7608889915BA5BA902938A645E595F265DAEDAE9688BDA2B";
    attribute INIT_24 of inst : label is "279027902790279027902790201020134A00FDD24101A965848C04410AA48000";
    attribute INIT_25 of inst : label is "4B056B20FFFC94D9B90001BB40A4924C1224912A1524FA3B0A6DEB15A16D5C70";
    attribute INIT_26 of inst : label is "0D1897A56896A57C490500D66E683E555783E0F277C0053645020AA010152979";
    attribute INIT_27 of inst : label is "9B6D545705E44E5FF99635F1539D89CA9BD6DA6DB5D15C1791392F664EEA065E";
    attribute INIT_28 of inst : label is "14802480C5CBADB683768D4B6D8CD825455407B1A7D89CEB857C75E76273AED5";
    attribute INIT_29 of inst : label is "1763322136B6231E4EE1218C2FF96005CA000A0902C080054ED087852130B400";
    attribute INIT_2A of inst : label is "6209E0624D3102DFBB788F178984951C0B354699BE1F8737DE182E100AE086A0";
    attribute INIT_2B of inst : label is "5A653754958CA89A7C718CD46B3004410C4D637761023082654831A0358714CA";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF000000000000000000EDB3D4E994";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "E3132C94B22714D172BA8C14E47FFFFFFFFF0000000000000000FFE20080200E";
    attribute INIT_31 of inst : label is "C01C9006DA523144AC884898882F32859234B445DDC716DCCDB5A75C31BC9752";
    attribute INIT_32 of inst : label is "53331E7125292FAA850CDD89371625815E5636231698312500D018F3B5663201";
    attribute INIT_33 of inst : label is "0000000E4929CE762739F98AAF31D3B194D691A8ED76E08BE45A2AAC02AA6D4D";
    attribute INIT_34 of inst : label is "1B5806BBB29D37C602CA47FB05112A28B42A7028942CD6DA9331219580000000";
    attribute INIT_35 of inst : label is "4891084E1309CA4B3928A888958CD2A22089EECDD420E5588614FF4E805169B4";
    attribute INIT_36 of inst : label is "B75CE490614923DB580CF204694284C86E91013D1364CB0586555954C4B671A2";
    attribute INIT_37 of inst : label is "A5203ED00C96DD1B448482519A124B680ABD3C9D3A7529D6B515B9CE4F50DBD5";
    attribute INIT_38 of inst : label is "000400100040010A040010004001000400100040010004001000400AC55410EA";
    attribute INIT_39 of inst : label is "FFFF10B09090D0A00000FFD08090A0A1FFFF007090A080A08B2C2ACB80004001";
    attribute INIT_3A of inst : label is "FFC0A090A0D0B08000308090D0A09081FF808080E0B0A0800000809080F080A1";
    attribute INIT_3B of inst : label is "0000000080000000BFFFFFFF7FFFFFFF0000000080000000BFB0A0B0F0908081";
    attribute INIT_3C of inst : label is "0000000080000000BFFFFFFF7FFFFFFF0000000000000000BFFFFFFF7FFFFFFF";
    attribute INIT_3D of inst : label is "0000000080000000BFFFFFFF7FFFFFFF0000000000000000BFFFFFFF7FFFFFFF";
    attribute INIT_3E of inst : label is "0000000080000000BFFFFFFF7FFFFFFF0000000000000000BFFFFFFF7FFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000BFFFFFFF7FFFFFFF0000000080000000BFFFFFFF7FFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "D9CAC85BCF0FFC220E09A165B170C5C462923FCC4D9C10469224FE29875FD818";
    attribute INIT_01 of inst : label is "531B908C09814A9244491C41C92E84329EFBEA63F4D9364434434435821CA6DE";
    attribute INIT_02 of inst : label is "CEB8C2C97AE30935C616400189332E188C5AB23300001950E330B8488721FE4A";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF9FFF6DB386100019718592E30B24EB8C2C86793C964B2793";
    attribute INIT_04 of inst : label is "3EE0E49133085EA114422AC1CCE46AA31C55C000284320792A22A333FFFFFFFF";
    attribute INIT_05 of inst : label is "CFEFAEB8B0B2FC2BFFE0FAFFFC3EBDFF5FFFBFFFFBFFFFBFFA7F9FE77FFFF765";
    attribute INIT_06 of inst : label is "00D8E2BC633FFB6DD999FF1244C24E7F927F920D21920ED2B862A602FFFFFF9F";
    attribute INIT_07 of inst : label is "C03339C9D9830CC185D879DC0C6557E4B03FEDBF79B6DB30849C93F4D8E1FD00";
    attribute INIT_08 of inst : label is "4B2CDB24965C93230CB8C49FA4687601C70A51653F8005BB8108EE1719C76018";
    attribute INIT_09 of inst : label is "9FD09000009A088435830016649617AE30985275C6130A5EB8C2E102000C49BC";
    attribute INIT_0A of inst : label is "C0646322F5F8366C76F237613718D8DB1B246586F0CBD7E6364DC88EE494C964";
    attribute INIT_0B of inst : label is "9E218618624466649D99B2204DFFFF7425366E67196C9606198865DB30C61285";
    attribute INIT_0C of inst : label is "7987E02F597A40D0D873D7EB8C4270B8F19BBB92DE94FFC9249025AAC66DB720";
    attribute INIT_0D of inst : label is "59CECFE59CF32E94A52980031697932EE4A40046058DC839D9CE20402CB3602C";
    attribute INIT_0E of inst : label is "FFFE0000000000000000ED818376DFBFFE9DDDB7FCDFF6ECC9C44088BCABF016";
    attribute INIT_0F of inst : label is "FFFE0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "8C24018D190280E42D1B00288AA8140019199942091214590A8A88288AA80400";
    attribute INIT_11 of inst : label is "00000001C00020A28AAA282080000400E0A0000200AA0A0280A822820080B400";
    attribute INIT_12 of inst : label is "052000CC5301A2BD9F0000050187C000000063937EFDCDDEDC007E0A80029400";
    attribute INIT_13 of inst : label is "7C0F03C0F03C0F03C0F03C9F2FC8733CC721C8F23C8F21CBF3F8882A82809400";
    attribute INIT_14 of inst : label is "CBF2FCBF2FCFF2FC9F1FC5F17C7F10C3F07C1F0FC3F0FC8F23C3802218822400";
    attribute INIT_15 of inst : label is "BF27C9F27C9F27C9E022AAAAAAA02A0000020828AAA28A0A0828A8A2A2828400";
    attribute INIT_16 of inst : label is "020028080082802028020200002094004AAAAA02A2A2AA8A08220AA28AA80400";
    attribute INIT_17 of inst : label is "07C3F01C0220820202080888C080A0000200280800828020280202000080A000";
    attribute INIT_18 of inst : label is "FC4F0000F03C0F0380003C0F03C480004F13C0F01C3F11C42A0A28A28A2AB400";
    attribute INIT_19 of inst : label is "8002000280020002822820200228000288208020080080080080000800800400";
    attribute INIT_1A of inst : label is "8002004002802002800202282020022800028A28A0200A08A08A08A0000A08A0";
    attribute INIT_1B of inst : label is "FFFF004002802002C08808822022140000028A28A0200A08A08A08A0000A08A0";
    attribute INIT_1C of inst : label is "2208822A0200A28A2A80280A200A028080200208280A28A22820808000021400";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE0A0080A0280A0280082800008AA822080200A0";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "80000000000000000000FFFFFFFFFFFFFFFF00000000000063FE7F5F7DE1F2E3";
    attribute INIT_20 of inst : label is "CF83CFCE4E6F22079252E4B93E7FFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "C3C479B2DF57E7EDC4E1E23CF96FAB71243C40F365BEADCC9CBCD30F3E67D6F5";
    attribute INIT_22 of inst : label is "D937CAECA796CC64311B26F95D94F2C98CE22364C73BC9DE666663E1F9C1904D";
    attribute INIT_23 of inst : label is "E4E71088E94B106CE7BBBBAD3643643CD94801B3190C46C9BE47E47CB2633888";
    attribute INIT_24 of inst : label is "D865D865D865D865D865D865DFE5DFEF84A2205B2CB27F184E261330E2321F60";
    attribute INIT_25 of inst : label is "BDF339E30006DB1EE700020CFE724921B9720C8241920E68EB3F2E371C105FB5";
    attribute INIT_26 of inst : label is "B2FCC0197CC019627EDF5F8023F2C531712C4B0788F6C7C970B86666CCC2F787";
    attribute INIT_27 of inst : label is "4411B75DDCDA212B18CB572CCFB7442678596B10465D77736884FCE339ACD95B";
    attribute INIT_28 of inst : label is "39EDB6593E0672CBD91F776C30C78D3763977AF57F744225DDCB12EDD1089636";
    attribute INIT_29 of inst : label is "E9B1999CD38D9860F10DB2658DC09BFA06CEE601B92E6763330FB83ADC974AF2";
    attribute INIT_2A of inst : label is "39E61DDC96DCEE80C09730615BBC8009E33C9B6C4AF159C1A0CB12F7E5373A6E";
    attribute INIT_2B of inst : label is "7CF64CDFE8218DC7838CE273399FF29CE3B31CF896ED965D9A6DEC347F09E221";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF000000000000000BFFDC007873D9";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "984082420810C2401822C2E6167FFFFFFFFF0000000000000000FFE1FC3F0FC1";
    attribute INIT_31 of inst : label is "E40E0DBD64EDCE3E53E7FF4E6611C87241C2CFF26600810230CA1D02CC024088";
    attribute INIT_32 of inst : label is "A9EEC19EDEF7E055759B876570E9EA4C231C61DCE84F9E13772EE3C665DDC4C0";
    attribute INIT_33 of inst : label is "000000632DBC6303318C0C756082010F7E286C81B9202776C579F19CD8553AA6";
    attribute INIT_34 of inst : label is "082587580008E133B92B2551B0998BC446B199C466B31872EEEE4FCA00000000";
    attribute INIT_35 of inst : label is "6F66B1B3FCF6E3A6C5B66677CA7F0D911BF440B33FEB5899FF63573DEDFE8082";
    attribute INIT_36 of inst : label is "8616C9CCC02DCB991901861BB43C7BECC0D89EC7D71F30F87BA33CAB2B5B8E31";
    attribute INIT_37 of inst : label is "EDB024321EDCC303F2322930445B6CB64FD9B4D9B3610D9CE119F9EC671B1619";
    attribute INIT_38 of inst : label is "400100040010004A010004001000400100040010004001000400001B80AAF40B";
    attribute INIT_39 of inst : label is "FFFF0D7DBDADAD800000FFAD3DED2D01FFFF002D3D9DBD81BC7FD7BF7D601000";
    attribute INIT_3A of inst : label is "FFBD3D7D8D8DAD80000D7D7D0D2DAD81FFBD1DFD0D8D0D000000BD6D2DADAD01";
    attribute INIT_3B of inst : label is "0000000000000000FFFFFFFFFFFFFFFF00000000000000007F9D9DFD8D0DED81";
    attribute INIT_3C of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "00000000000000007FFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "0000000000000000FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "48AAA852860FE82010588325D1C005A2C0007FED4D9C102002007E09870F81B0";
    attribute INIT_01 of inst : label is "401E901A0B41080044001801E02400625AAAAD56D294A5021C21C21F410AD64E";
    attribute INIT_02 of inst : label is "8894C6D922531B64A636C00004932B180C42B03000001954E320B02842912522";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFF9249249341100019298DB2531974894C65D6F578BD5E2D56";
    attribute INIT_04 of inst : label is "1E4084003694DA9114222AA1C444E226925520002002A064AAAA2323FFFFFFFF";
    attribute INIT_05 of inst : label is "06182180A0AB00080000060000018000400020000206006006000001000000E8";
    attribute INIT_06 of inst : label is "00D88291085FF924C888FF1645C42E3F9657971171971092A0642D0260101804";
    attribute INIT_07 of inst : label is "4011194918C10C608194656C046D57E5903FE49F20924932049A57D4D910F500";
    attribute INIT_08 of inst : label is "CB2D9B6CB64852A28AB8C01EA208420506815396AD40053A8000664E18842008";
    attribute INIT_09 of inst : label is "BF484A000049044200032000659612A531B40AC4A636814894C6D081000024B4";
    attribute INIT_0A of inst : label is "A92C532A54E8972C72563721329858CB1912E20640C953A6366CA5A455505B6D";
    attribute INIT_0B of inst : label is "16018618604464441991B02009C0007424122454186596164B992DDBB2451345";
    attribute INIT_0C of inst : label is "74D7A009493A40D0D82BB3EC1AA16999933999924892B6A8904814AAA2249E00";
    attribute INIT_0D of inst : label is "1884CFC188410C42108480011207498EC02000020189C810888420404431200C";
    attribute INIT_0E of inst : label is "FFFE0000000000000000E48081324D2DB4155593684DA08AA8C640889D81F006";
    attribute INIT_0F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "1800020D110384E92D1B008228A024002D2DAD4A695E134D8A28208228A02400";
    attribute INIT_11 of inst : label is "00000000000020A28AAAAAAAAAAAA400008002000288880200A08A0802028400";
    attribute INIT_12 of inst : label is "043C008842C000000000000000000000000003D0000000000000000AA8802400";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000040100000000000000100A20A28A20400";
    attribute INIT_14 of inst : label is "0000000000040100400000000000000000000000000000000000008A0000A400";
    attribute INIT_15 of inst : label is "000000000000000002A2AAAAAAA02A0AAAAAAAAAAAA28A080000020828AAA400";
    attribute INIT_16 of inst : label is "2A00A8020A82208802088220228A24004AAAAA02A2A2AA8A022A2AA28A280400";
    attribute INIT_17 of inst : label is "00000000282AAAA2828A0A084A8280A82A00A8020A822088020882200A8280A8";
    attribute INIT_18 of inst : label is "0040100001004010100000000004100040100401004000000020820820800400";
    attribute INIT_19 of inst : label is "202AA282202AA2822082080A0082028020A2082A00A20A2082080A00A20A2400";
    attribute INIT_1A of inst : label is "202AA2C02AA2822A22822082080A0082028020A2082A00A20A2082080A00A20A";
    attribute INIT_1B of inst : label is "FFFF00402AA2822A4220220882882400028020A2082A00A20A2082080A00A20A";
    attribute INIT_1C of inst : label is "2A0280A080A00820880802008200802008028A20A00820808000020082082400";
    attribute INIT_1D of inst : label is "FFFF0000000000000000FFFFFE200A800802008020A80200802AA02A00020028";
    attribute INIT_1E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFC";
    attribute INIT_1F of inst : label is "FFFFF800000000000000FFFFFFFFFFFFFFFF0000000000005C0182A0121E0F1C";
    attribute INIT_20 of inst : label is "4D0345C51A2501054A4850A3317FFFFFFFFE0000000000000000FFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "63A27592C81783E50EB1D13AE9640B41643A20EB25902D0D963A698EBA6206C7";
    attribute INIT_22 of inst : label is "89074AA4A352C464313120E954946A588CE626240D2B495A22222340B8A100D9";
    attribute INIT_23 of inst : label is "E2D71080E942106994AAAABD3251251AF524009119044C483A55A55A92233889";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000F8CA240890C317F108D16311062291F60";
    attribute INIT_25 of inst : label is "95B339EA80064B10E2000112B569249354A9424221494E68CABC28140A284EB0";
    attribute INIT_26 of inst : label is "367CC2012CC2012048075F8207F657113165194EA07247C92835622246C25282";
    attribute INIT_27 of inst : label is "4A28F248D8DE630A1043136CC682CC6631492928A3492363798C78C11B249B49";
    attribute INIT_28 of inst : label is "39E49218B9066A4DD92967241042C41323536C516C2CC6214CDB10A0B3188472";
    attribute INIT_29 of inst : label is "F590888A118C8854E02C9061898093E966EEE520310E7763288BBC231447A0F2";
    attribute INIT_2A of inst : label is "B5554DCC965C6E0021532A4012BC80095194DB2CA0E0D9C122C390F756BD6A6E";
    attribute INIT_2B of inst : label is "34D2444FECA50E0D01046631198DAABAD1B73AE4564C861DBB24A4947D858150";
    attribute INIT_2C of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000019C1078D349";
    attribute INIT_2D of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFF0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "94A145210408A1002422C2C5167FFFFFFFFF0000000000000000FFE000000000";
    attribute INIT_31 of inst : label is "22420C912DA75A1A4A97BD262209A42928A2AB4911418086482D3002CA822084";
    attribute INIT_32 of inst : label is "A880215E4A52E055748204158265695A131001F5A42F5A9376A4E64CE4CC84A4";
    attribute INIT_33 of inst : label is "00000052A49CE731339CC4606091010C7D643A8039000000C479F88848D512A2";
    attribute INIT_34 of inst : label is "0125820810084111B9393009B8DD89466298CDC66291142246664D2D00000000";
    attribute INIT_35 of inst : label is "252253D355D2628080924656AD7E85911BD420B112A1481157214618E4FF4012";
    attribute INIT_36 of inst : label is "A41299CC6024DA991101860ABA142BE40048DAAFD83D104023B114AB2D7A8A11";
    attribute INIT_37 of inst : label is "EC9028621E4C8602E0000030CE4925B647D0A450A1418508410D318826111C11";
    attribute INIT_38 of inst : label is "000428100040010A042810004001000400100042810004281000001990AA4009";
    attribute INIT_39 of inst : label is "FFFF2000207010000000FF8020B05081FFFF000020709080C38A00C08A204001";
    attribute INIT_3A of inst : label is "FFA0808070B01000002000A030509001FFE0A080B0F01080000080A030905081";
    attribute INIT_3B of inst : label is "00000002800000007FFFFFFF7FFFFFFF0000000000000000FFE0208030701081";
    attribute INIT_3C of inst : label is "00000002800000007FFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "00000002800000007FFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "80000002800000007FFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "80000002800000007FFFFFFF7FFFFFFF0000000000000000FFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
