library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity eprom_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of eprom_4 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"06",X"0C",X"18",X"0C",X"06",X"03",X"80",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",
		X"00",X"00",X"80",X"C0",X"60",X"30",X"18",X"0C",X"C0",X"E0",X"B0",X"98",X"9C",X"9E",X"9F",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",
		X"FF",X"0F",X"38",X"E0",X"80",X"00",X"00",X"00",X"FF",X"F0",X"9C",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"40",
		X"00",X"03",X"0F",X"1E",X"3F",X"7F",X"5F",X"EE",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"81",X"81",X"81",X"81",X"81",X"81",
		X"BF",X"BF",X"FF",X"6E",X"7F",X"7F",X"7F",X"2E",X"FF",X"FF",X"FF",X"EE",X"FF",X"FF",X"FF",X"EE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"C0",X"40",X"40",X"40",X"60",X"20",X"30",
		X"BF",X"BF",X"9F",X"CE",X"4F",X"67",X"33",X"18",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"08",X"0C",X"06",X"03",X"01",X"00",
		X"0E",X"03",X"00",X"00",X"00",X"00",X"80",X"E0",X"7F",X"DF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",
		X"38",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"9C",X"F0",X"FF",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"01",X"03",X"06",X"0C",X"9F",X"9F",X"FF",X"DF",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"0C",
		X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"9F",X"9E",X"9C",X"98",X"B0",X"FF",X"9F",X"9F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"01",X"00",X"18",X"30",X"60",X"C0",X"80",X"FF",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"B0",X"98",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"3F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"9C",X"9E",X"9F",X"9F",X"9F",X"9F",X"9F",X"DF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",
		X"00",X"00",X"20",X"70",X"D8",X"8C",X"06",X"03",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"03",X"07",
		X"FC",X"F8",X"F0",X"F0",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"80",X"C0",X"60",X"30",X"18",X"8F",X"DF",X"FF",X"BF",X"9F",X"9F",X"9F",X"9F",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",
		X"0C",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"FF",X"01",X"03",X"06",X"0C",X"18",X"30",
		X"00",X"DF",X"8C",X"06",X"03",X"01",X"00",X"00",X"9F",X"FF",X"01",X"03",X"07",X"8F",X"DF",X"FF",
		X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FE",X"80",X"C0",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"C0",X"60",X"31",X"FB",X"80",
		X"00",X"00",X"20",X"70",X"D8",X"8C",X"FE",X"00",X"BF",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"9F",
		X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"FF",X"B0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"98",X"9C",X"9E",X"9F",X"9F",X"9F",X"9F",X"9F",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"F0",X"F8",X"F0",X"E0",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1C",X"1C",X"1C",X"1C",X"1C",X"1E",X"1C",X"1C",X"1C",X"1C",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"17",X"01",X"00",X"00",X"00",X"1E",X"1C",X"1F",X"1F",X"1F",X"1E",X"1E",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"01",X"17",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"10",X"00",
		X"1C",X"1C",X"1C",X"1C",X"1E",X"00",X"00",X"10",X"1C",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1C",
		X"00",X"00",X"00",X"1E",X"1C",X"1C",X"1C",X"1C",X"1E",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"03",
		X"1E",X"1E",X"1C",X"1C",X"1C",X"1C",X"1C",X"1E",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"1F",X"1F",
		X"FF",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"01",X"00",X"FD",X"EC",X"8C",X"0C",X"0C",X"8C",X"EC",X"FD",
		X"00",X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",
		X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"0F",X"E0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"1F",
		X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"7F",X"7F",X"00",X"7F",X"00",X"00",
		X"00",X"FE",X"FF",X"FF",X"00",X"00",X"FE",X"00",X"00",X"FF",X"AA",X"AA",X"55",X"55",X"FF",X"00",
		X"00",X"3F",X"7F",X"7F",X"00",X"40",X"3F",X"00",X"2C",X"2C",X"2F",X"27",X"20",X"1F",X"00",X"00",
		X"4E",X"4E",X"2C",X"00",X"2C",X"2C",X"2C",X"2C",X"72",X"4E",X"72",X"4E",X"4E",X"4E",X"4E",X"4E",
		X"4E",X"4E",X"4E",X"4E",X"72",X"4E",X"72",X"4E",X"2C",X"2C",X"2C",X"00",X"0C",X"4E",X"4E",X"4E",
		X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"2C",X"00",X"00",X"17",X"2F",X"2C",X"2C",X"2C",X"2C",
		X"00",X"80",X"FF",X"FF",X"80",X"FF",X"80",X"00",X"00",X"FE",X"FF",X"FF",X"00",X"00",X"FE",X"00",
		X"00",X"FF",X"FF",X"FF",X"55",X"55",X"FF",X"00",X"00",X"BF",X"FF",X"FF",X"80",X"C0",X"BF",X"00",
		X"00",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",X"80",X"DF",X"DF",X"00",X"1F",X"80",X"00",
		X"00",X"FF",X"BF",X"BF",X"40",X"40",X"FF",X"00",X"00",X"C1",X"80",X"80",X"41",X"41",X"C1",X"00",
		X"00",X"FF",X"FE",X"FE",X"01",X"01",X"FF",X"00",X"00",X"00",X"FD",X"FD",X"00",X"FD",X"00",X"00",
		X"00",X"E0",X"F7",X"F7",X"00",X"07",X"E0",X"00",X"00",X"7F",X"2F",X"2F",X"50",X"50",X"7F",X"00",
		X"00",X"FF",X"FA",X"FA",X"05",X"05",X"FF",X"00",X"00",X"03",X"F7",X"F7",X"00",X"F4",X"03",X"00",
		X"00",X"F8",X"FD",X"FD",X"00",X"01",X"F8",X"00",X"00",X"1F",X"0B",X"0B",X"14",X"14",X"1F",X"00",
		X"00",X"FC",X"E8",X"E8",X"14",X"14",X"FC",X"00",X"00",X"0F",X"DF",X"DF",X"00",X"D0",X"0F",X"00",
		X"00",X"FC",X"FE",X"FE",X"00",X"00",X"FC",X"00",X"00",X"1F",X"BF",X"BF",X"00",X"A0",X"1F",X"00",
		X"00",X"0F",X"D5",X"25",X"5A",X"8A",X"0F",X"00",X"00",X"00",X"D8",X"25",X"52",X"8D",X"00",X"00",
		X"00",X"F8",X"D0",X"D5",X"2A",X"2D",X"F8",X"00",X"00",X"0F",X"75",X"D5",X"8A",X"0A",X"0F",X"00",
		X"00",X"00",X"70",X"D8",X"8D",X"07",X"00",X"00",X"00",X"F8",X"D0",X"D0",X"2D",X"2F",X"F8",X"00",
		X"00",X"0F",X"85",X"55",X"2A",X"DA",X"0F",X"00",X"00",X"00",X"8D",X"52",X"25",X"D8",X"00",X"00",
		X"00",X"F8",X"D5",X"D2",X"2D",X"28",X"F8",X"00",X"00",X"0F",X"05",X"85",X"DA",X"7A",X"0F",X"00",
		X"00",X"00",X"07",X"8D",X"D8",X"70",X"00",X"00",X"00",X"F8",X"D7",X"D5",X"28",X"28",X"F8",X"00",
		X"46",X"46",X"24",X"00",X"2C",X"2C",X"2C",X"2C",X"62",X"46",X"62",X"46",X"46",X"46",X"46",X"46",
		X"46",X"46",X"46",X"46",X"62",X"46",X"62",X"46",X"2C",X"2C",X"2C",X"00",X"04",X"46",X"46",X"46",
		X"42",X"42",X"24",X"00",X"2C",X"2C",X"2C",X"2C",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",
		X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"2C",X"2C",X"2C",X"00",X"04",X"42",X"42",X"42",
		X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",
		X"81",X"81",X"42",X"00",X"2C",X"2C",X"2C",X"2C",X"00",X"81",X"00",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"00",X"81",X"00",X"81",X"2C",X"2C",X"2C",X"00",X"42",X"81",X"81",X"81",
		X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"2C",X"2C",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"02",X"00",X"FE",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"02",X"00",X"FE",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"02",X"00",X"FE",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"FE",X"7E",X"7E",X"7E",X"7E",X"FE",X"FE",
		X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"F2",X"00",X"FE",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"18",X"3C",X"00",X"7C",X"7C",X"7C",X"7C",X"00",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"00",X"7C",X"7C",X"7C",X"7C",X"7E",X"3C",X"18",
		X"F1",X"A0",X"F8",X"F8",X"F9",X"80",X"40",X"40",X"40",X"40",X"41",X"80",X"F8",X"F8",X"F9",X"AF",
		X"F1",X"A0",X"F8",X"F8",X"F9",X"80",X"40",X"40",X"40",X"40",X"41",X"80",X"F8",X"F8",X"F9",X"AF",
		X"00",X"20",X"F8",X"F8",X"F8",X"00",X"40",X"40",X"40",X"40",X"40",X"00",X"F8",X"F8",X"F8",X"20",
		X"FC",X"FC",X"F8",X"F8",X"FF",X"F7",X"E3",X"C3",X"3C",X"38",X"10",X"00",X"E0",X"E0",X"C0",X"C0",
		X"FC",X"FC",X"F8",X"F8",X"FF",X"F7",X"E3",X"C3",X"3C",X"38",X"10",X"00",X"E0",X"E0",X"C0",X"C0",
		X"81",X"E1",X"78",X"7E",X"3C",X"38",X"10",X"00",X"81",X"87",X"1E",X"7E",X"FC",X"FC",X"F8",X"F8",
		X"81",X"E1",X"78",X"7E",X"3C",X"38",X"10",X"00",X"81",X"87",X"1E",X"7E",X"FC",X"FC",X"F8",X"F8",
		X"E0",X"E0",X"C0",X"C0",X"81",X"87",X"1E",X"7E",X"FF",X"F7",X"E3",X"C3",X"81",X"E1",X"78",X"7E",
		X"E0",X"E0",X"C0",X"C0",X"81",X"87",X"1E",X"7E",X"FF",X"F7",X"E3",X"C3",X"81",X"E1",X"78",X"7E",
		X"78",X"6D",X"EF",X"F3",X"37",X"DE",X"DE",X"1E",X"E6",X"DE",X"BE",X"70",X"6F",X"DF",X"D8",X"F6",
		X"DD",X"19",X"C6",X"EE",X"6C",X"0D",X"6D",X"ED",X"C6",X"98",X"BB",X"33",X"BC",X"BF",X"BB",X"B4",
		X"36",X"F6",X"E3",X"5B",X"D9",X"B6",X"B7",X"83",X"F6",X"F7",X"7B",X"B8",X"C6",X"FF",X"39",X"06",
		X"EE",X"06",X"37",X"BB",X"B3",X"CD",X"CE",X"37",X"CE",X"EF",X"77",X"B8",X"DD",X"ED",X"61",X"06",
		X"1C",X"3E",X"37",X"A3",X"E3",X"E7",X"3C",X"19",X"6E",X"6D",X"23",X"3F",X"FE",X"E0",X"ED",X"CD",
		X"76",X"F0",X"EE",X"8F",X"6D",X"F1",X"C0",X"B3",X"F7",X"F3",X"2C",X"DE",X"EF",X"83",X"7C",X"7E",
		X"C1",X"D9",X"3D",X"FC",X"CB",X"33",X"76",X"7E",X"9F",X"B6",X"D6",X"C0",X"1F",X"7F",X"F1",X"E0",
		X"B7",X"DF",X"C9",X"B6",X"37",X"F3",X"EC",X"DD",X"9F",X"EF",X"F0",X"77",X"BF",X"0E",X"F6",X"F6",
		X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"00",X"FE",X"80",X"80",X"00",X"9F",X"90",X"90",
		X"04",X"C6",X"00",X"00",X"00",X"FF",X"00",X"0E",X"28",X"AD",X"00",X"00",X"00",X"EC",X"28",X"28",
		X"50",X"50",X"10",X"10",X"10",X"1B",X"40",X"7B",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"50",
		X"00",X"20",X"00",X"20",X"10",X"0A",X"00",X"00",X"08",X"A9",X"A8",X"A8",X"20",X"20",X"2F",X"88",
		X"00",X"7F",X"00",X"40",X"00",X"40",X"79",X"48",X"50",X"50",X"50",X"50",X"57",X"54",X"54",X"42",
		X"00",X"00",X"00",X"00",X"B2",X"A0",X"A6",X"00",X"28",X"80",X"28",X"28",X"A8",X"08",X"A8",X"28",
		X"48",X"05",X"00",X"00",X"01",X"50",X"50",X"00",X"50",X"5A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"C0",X"04",X"04",X"C4",X"04",X"04",X"04",X"28",X"28",X"28",X"28",X"28",X"28",X"28",X"28",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"22",X"15",X"11",X"17",X"14",X"F7",X"00",X"C0",X"41",
		X"00",X"00",X"DF",X"51",X"DF",X"00",X"1F",X"C4",X"10",X"10",X"50",X"50",X"5F",X"00",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"E2",X"00",X"40",X"40",X"41",X"41",X"40",X"40",X"41",X"04",X"00",X"08",
		X"33",X"88",X"64",X"12",X"8A",X"29",X"05",X"15",X"F0",X"10",X"F0",X"40",X"70",X"10",X"77",X"45",
		X"40",X"40",X"FC",X"05",X"04",X"05",X"04",X"05",X"08",X"08",X"00",X"C4",X"81",X"C0",X"00",X"41",
		X"17",X"10",X"05",X"29",X"8A",X"12",X"64",X"88",X"7D",X"05",X"F7",X"00",X"00",X"00",X"00",X"00",
		X"FD",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"C1",X"05",X"F5",X"11",X"15",X"15",X"11",X"15",
		X"30",X"20",X"3F",X"00",X"00",X"00",X"00",X"00",X"07",X"05",X"F5",X"15",X"17",X"10",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"24",X"12",X"01",X"01",X"19",X"A1",X"00",X"73",X"21",X"01",X"82",X"80",X"00",X"02",X"00",
		X"00",X"63",X"21",X"25",X"C4",X"00",X"01",X"03",X"00",X"80",X"80",X"A0",X"A4",X"78",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"05",X"1F",X"A1",X"00",X"7F",X"25",X"25",X"A2",X"80",X"00",X"23",X"21",
		X"25",X"67",X"25",X"25",X"FC",X"24",X"21",X"03",X"00",X"A0",X"A7",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"A5",X"7F",X"A5",X"00",X"FF",X"A5",X"25",X"FF",X"81",X"81",X"FB",X"A1",
		X"25",X"F7",X"25",X"A5",X"FD",X"A4",X"21",X"67",X"00",X"A5",X"EF",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"A5",X"FF",X"A5",X"00",X"FF",X"A5",X"A5",X"FF",X"A5",X"A5",X"FF",X"A5",
		X"A5",X"FF",X"A5",X"A5",X"FF",X"A5",X"A5",X"FF",X"00",X"A5",X"FF",X"A5",X"A5",X"7E",X"24",X"18",
		X"18",X"3C",X"7E",X"FD",X"FD",X"FF",X"FD",X"00",X"FF",X"A7",X"A7",X"FF",X"A7",X"A7",X"FF",X"A7",
		X"A7",X"FF",X"A7",X"A7",X"FF",X"A7",X"A7",X"FF",X"00",X"FD",X"FF",X"FD",X"FD",X"7E",X"3C",X"18",
		X"18",X"3C",X"00",X"7C",X"7C",X"7C",X"7C",X"00",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"00",X"7C",X"7C",X"7C",X"7C",X"7E",X"3C",X"18",
		X"00",X"00",X"00",X"18",X"3C",X"00",X"7C",X"7C",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"7C",X"7C",X"7E",X"3C",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"00",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"7E",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"A6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"2E",X"0E",X"00",X"A6",X"A6",X"A6",X"A6",X"A0",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A0",X"A6",X"A6",X"A6",X"A6",X"4E",X"0E",X"2E",X"14",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1C",X"2E",X"0E",X"4E",X"4E",X"00",X"A6",X"A6",X"A6",X"A6",X"A0",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"A0",X"A6",X"A6",X"A6",X"A6",X"4E",X"4E",X"4E",X"0E",X"2E",X"14",X"00",X"00",
		X"00",X"04",X"0E",X"0E",X"4E",X"4E",X"4E",X"00",X"AE",X"AE",X"AE",X"AE",X"AE",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"AE",X"AE",X"AE",X"AE",X"AE",X"4E",X"4E",X"4E",X"4E",X"0E",X"2E",X"14",X"00",
		X"0C",X"16",X"20",X"47",X"47",X"47",X"47",X"7E",X"AE",X"AE",X"AE",X"AE",X"AE",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"AE",X"AE",X"AE",X"AE",X"AE",X"7E",X"47",X"47",X"47",X"47",X"20",X"16",X"08",
		X"0C",X"1E",X"20",X"61",X"C3",X"C3",X"C3",X"00",X"AE",X"AE",X"AE",X"AE",X"AE",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"AE",X"AE",X"AE",X"AE",X"AE",X"00",X"C3",X"C3",X"C3",X"21",X"10",X"0A",X"04",
		X"0C",X"1E",X"22",X"67",X"CF",X"CB",X"CB",X"00",X"AE",X"AE",X"AE",X"AE",X"AE",X"A6",X"A6",X"A6",
		X"A6",X"A6",X"A6",X"AE",X"AE",X"AE",X"AE",X"AE",X"00",X"CB",X"CB",X"CF",X"27",X"12",X"0A",X"04",
		X"18",X"3C",X"00",X"5C",X"3C",X"7C",X"7C",X"00",X"86",X"A6",X"A6",X"A6",X"A2",X"A0",X"A6",X"A6",
		X"A6",X"A6",X"86",X"26",X"86",X"A6",X"A4",X"A2",X"00",X"78",X"78",X"5C",X"3C",X"7E",X"3C",X"18",
		X"18",X"3C",X"24",X"7C",X"7E",X"7D",X"7C",X"7E",X"A6",X"E6",X"E6",X"BE",X"E6",X"A6",X"AF",X"B6",
		X"B6",X"BF",X"A6",X"E7",X"A6",X"B7",X"AE",X"A6",X"7E",X"7C",X"7C",X"7E",X"7D",X"7E",X"3C",X"18",
		X"00",X"00",X"80",X"C0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"10",X"08",X"88",X"C0",X"80",X"00",X"06",X"06",X"80",X"C0",X"E2",X"42",
		X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"03",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"80",X"C0",X"80",X"00",X"80",X"80",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"80",X"80",
		X"01",X"83",X"11",X"20",X"03",X"01",X"00",X"00",X"00",X"19",X"3C",X"3C",X"18",X"03",X"07",X"01",
		X"00",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"10",X"02",X"04",X"00",X"00",X"00",X"00",X"81",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"30",X"00",
		X"00",X"18",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"10",X"00",X"80",X"40",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1C",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"30",X"10",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"04",X"08",X"00",X"00",X"00",X"00",X"01",X"70",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"70",X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"00",X"30",X"10",X"00",X"00",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"10",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"03",X"00",X"00",X"00",X"01",X"03",X"03",X"02",X"02",X"01",X"00",X"00",
		X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"E0",X"00",
		X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"F0",X"70",X"70",X"F8",X"FC",X"FC",X"7C",X"3C",X"F8",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"0B",X"09",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"7C",X"3C",X"F8",X"F0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1F",X"1F",X"17",X"13",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"BE",X"9E",X"FC",X"F8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"1F",X"17",X"13",X"0F",X"07",X"00",
		X"00",X"00",X"00",X"00",X"38",X"7C",X"FE",X"FE",X"BE",X"DE",X"FC",X"F8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1F",X"3F",X"3F",X"2F",X"27",X"1F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"7C",X"BC",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"1F",X"3F",X"3F",X"2F",X"27",X"1F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"70",X"F8",X"FC",X"FC",X"7C",X"BC",X"F8",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"03",X"1F",X"3E",X"7F",X"7F",X"5F",X"4F",X"3E",X"1C",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"78",X"F0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"60",X"20",X"00",X"00",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"18",X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"18",X"08",X"00",X"00",X"00",X"80",X"80",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"0C",X"04",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"02",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"20",X"00",X"10",X"00",X"00",X"10",X"00",X"02",
		X"40",X"00",X"08",X"00",X"00",X"08",X"00",X"04",X"00",X"00",X"08",X"00",X"00",X"88",X"00",X"40",
		X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"08",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"08",X"00",X"00",
		X"00",X"06",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"78",X"78",X"3C",X"3C",X"1E",X"1E",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"70",X"78",X"7C",X"7C",X"3C",X"1C",X"0C",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"7C",X"FE",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"07",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",X"07",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"08",X"0C",X"1E",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"7F",X"3F",X"1E",X"0E",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"1E",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1E",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"1C",X"3E",X"3E",X"7F",X"7F",X"7F",X"3E",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"7E",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3E",X"3F",X"3F",X"1F",X"1F",X"06",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"07",X"1C",X"33",X"E3",X"38",X"0E",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"A0",X"F0",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0F",X"3B",X"63",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",
		X"00",X"00",X"00",X"00",X"30",X"F0",X"30",X"20",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"30",X"12",X"18",X"08",X"0C",X"04",X"07",X"03",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"18",X"30",X"20",X"60",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"38",X"2E",X"33",X"13",X"13",X"18",X"08",X"08",X"0D",X"07",X"06",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"E0",X"38",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"02",X"06",X"07",X"05",X"0D",X"08",X"0B",X"1B",X"10",X"10",X"30",X"2F",X"38",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"60",X"20",X"10",X"F8",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"06",X"1C",X"33",X"E3",X"30",X"1C",X"06",X"03",X"00",X"00",X"00",
		X"00",X"00",X"60",X"E0",X"A0",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"A0",X"E0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0E",X"38",X"E0",X"32",X"1C",X"07",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"F0",X"A0",X"20",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"06",X"0C",X"18",X"30",X"63",X"3B",X"0F",X"01",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"20",X"30",X"F0",X"30",X"00",X"00",X"00",X"00",
		X"02",X"03",X"07",X"04",X"0C",X"08",X"18",X"13",X"33",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"C0",X"60",X"20",X"30",X"18",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"06",X"07",X"0D",X"08",X"08",X"18",X"13",X"13",X"33",X"2E",X"38",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"38",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"38",X"2F",X"30",X"10",X"10",X"18",X"0A",X"08",X"0D",X"05",X"07",X"06",X"02",X"00",
		X"00",X"00",X"00",X"80",X"F8",X"10",X"20",X"60",X"40",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"7F",X"7F",X"1F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"E0",X"FE",X"FE",X"FE",X"FE",X"FC",X"7C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"1F",X"7F",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"EC",X"FE",X"FE",X"FE",X"FE",X"FE",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"0E",X"1F",X"3F",X"7C",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3C",X"3C",X"3C",X"1E",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"1E",X"7E",X"FE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"10",X"38",X"38",X"3C",X"3C",X"3C",X"3E",X"3E",X"FE",X"FE",X"FE",X"7E",X"3C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"06",X"7F",X"7F",X"1F",X"07",X"00",X"00",X"00",X"00",
		X"00",X"00",X"18",X"3C",X"3C",X"7E",X"7E",X"7E",X"FE",X"FE",X"FE",X"FE",X"FC",X"7C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E3",X"7F",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"0E",X"0E",X"1E",X"1E",X"1E",X"FE",X"FC",X"FC",X"FC",X"F8",X"78",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"60",X"70",X"3C",X"3E",X"1C",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"78",X"78",X"F0",X"F0",X"F0",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"7C",X"3F",X"1F",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"70",X"F0",X"F0",X"F0",X"E0",X"F0",X"FC",X"FC",X"FC",X"F8",X"78",X"30",X"00",
		X"00",X"00",X"40",X"40",X"40",X"48",X"5C",X"5C",X"74",X"74",X"64",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"52",X"56",X"56",X"5C",X"5C",X"48",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"44",X"44",X"44",X"46",X"46",X"42",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"42",X"42",X"42",X"42",X"42",X"40",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"00",X"80",X"80",X"80",X"80",X"C0",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"00",X"80",X"C0",X"C0",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"60",X"70",X"70",X"D0",X"D0",X"D0",X"40",X"40",X"40",X"40",X"20",
		X"7C",X"FE",X"FE",X"FE",X"EA",X"E8",X"FC",X"DC",X"C4",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FA",X"FA",X"FE",X"F6",X"F0",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"7E",X"3E",X"BE",X"BE",X"BE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"BE",X"9E",X"DE",X"DE",X"5E",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"AE",X"A6",X"F6",X"76",X"16",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"00",X"00",X"40",X"40",X"40",X"44",X"44",X"44",X"44",X"7C",X"7C",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"5E",X"5E",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"46",X"46",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"42",X"42",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"C0",X"C0",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"50",X"50",X"50",X"10",X"F0",X"F0",X"40",X"40",X"40",X"40",X"20",
		X"7C",X"FE",X"FE",X"FE",X"DC",X"D4",X"D4",X"D4",X"D4",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"F6",X"F4",X"F4",X"F4",X"F4",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"BE",X"BE",X"BE",X"BE",X"BE",X"BE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"DE",X"DE",X"DE",X"DE",X"5E",X"DE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"76",X"56",X"56",X"56",X"56",X"F6",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"00",X"00",X"40",X"40",X"40",X"78",X"7C",X"44",X"44",X"7C",X"7C",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"4E",X"5E",X"50",X"50",X"5E",X"5E",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"42",X"46",X"44",X"44",X"46",X"46",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"42",X"42",X"42",X"42",X"42",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"40",X"00",X"80",X"80",X"80",X"80",X"C0",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"00",X"80",X"C0",X"40",X"40",X"C0",X"C0",X"40",X"40",X"40",X"40",X"20",
		X"00",X"00",X"40",X"40",X"00",X"E0",X"F0",X"50",X"10",X"F0",X"F0",X"40",X"40",X"40",X"40",X"20",
		X"7C",X"FE",X"FE",X"FE",X"EA",X"E8",X"FC",X"D4",X"D4",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FA",X"FA",X"FE",X"F4",X"F4",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"7E",X"3E",X"BE",X"BE",X"BE",X"BE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"BE",X"9E",X"DE",X"5E",X"5E",X"DE",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"7C",X"FE",X"FE",X"FE",X"AE",X"A6",X"F6",X"56",X"56",X"F6",X"FE",X"FE",X"FE",X"FE",X"FE",X"7C",
		X"00",X"18",X"7C",X"7C",X"64",X"70",X"78",X"78",X"78",X"7C",X"7C",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"78",X"7C",X"7E",X"76",X"72",X"7E",X"7E",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"7C",X"7E",X"7E",X"7C",X"7C",X"7E",X"7E",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"3C",X"BC",X"FC",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"7C",X"3C",X"BC",X"BC",X"9C",X"DC",X"FC",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"18",X"7C",X"7C",X"1C",X"CC",X"EC",X"6C",X"24",X"F4",X"FC",X"7C",X"7C",X"7C",X"58",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"80",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"80",X"20",
		X"00",X"80",X"20",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"80",X"00",
		X"54",X"AA",X"54",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"54",X"AA",X"54",
		X"00",X"00",X"00",X"0C",X"08",X"07",X"17",X"07",X"0B",X"1F",X"1F",X"00",X"0D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"40",X"80",X"90",X"B0",X"B0",X"20",X"40",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"05",X"07",X"0F",X"0B",X"01",X"07",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"40",X"A0",X"E0",X"F0",X"B0",X"A0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"1B",X"0C",X"0D",X"0F",X"1F",X"0B",X"0B",X"0D",X"0F",X"09",X"10",X"00",X"00",
		X"00",X"00",X"08",X"90",X"F0",X"B0",X"F0",X"D0",X"D8",X"F0",X"B0",X"F0",X"D8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"27",X"4C",X"41",X"17",X"13",X"03",X"07",X"09",X"0C",X"07",X"10",X"08",X"00",
		X"00",X"00",X"20",X"18",X"C8",X"50",X"E8",X"E8",X"E0",X"88",X"48",X"10",X"10",X"00",X"60",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"03",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"80",X"A0",X"C0",X"C0",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"00",X"00",X"00",X"00",X"01",X"00",X"F9",X"08",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"CB",X"4A",X"4A",X"4A",X"4A",X"7B",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"00",X"00",
		X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"7D",X"45",X"45",X"7D",X"01",X"7D",X"45",X"00",X"E0",X"20",X"20",X"00",X"03",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"45",X"7D",X"01",X"5D",X"15",X"15",X"5D",X"01",X"03",X"03",X"03",X"03",X"00",X"03",X"00",X"20",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"DD",X"55",X"DD",X"00",X"01",X"00",X"F9",X"08",X"20",X"60",X"E0",X"00",X"80",X"00",X"80",X"00",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"CB",X"4A",X"4A",X"4A",X"4A",X"7B",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"00",X"00",
		X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"01",X"01",X"00",X"04",X"07",X"04",X"A7",X"A4",
		X"22",X"22",X"06",X"90",X"F7",X"91",X"F1",X"90",X"20",X"00",X"00",X"20",X"20",X"00",X"EA",X"20",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A4",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"90",X"90",X"97",X"90",X"97",X"91",X"91",X"97",X"2E",X"2A",X"EE",X"00",X"7E",X"42",X"4E",X"48",
		X"00",X"00",X"00",X"00",X"01",X"00",X"F9",X"08",X"01",X"01",X"01",X"01",X"81",X"00",X"80",X"00",
		X"20",X"20",X"20",X"20",X"97",X"95",X"95",X"92",X"48",X"78",X"00",X"78",X"08",X"C8",X"60",X"F0",
		X"CB",X"4A",X"4A",X"4A",X"4A",X"7B",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"00",X"00",
		X"CB",X"49",X"48",X"48",X"48",X"00",X"00",X"00",X"38",X"48",X"9C",X"64",X"4E",X"32",X"2E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"00",X"AF",X"A5",
		X"29",X"65",X"53",X"CB",X"BE",X"E5",X"55",X"55",X"78",X"E3",X"8A",X"26",X"9C",X"58",X"72",X"E2",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",X"05",X"05",X"0F",X"00",X"06",X"09",X"04",
		X"57",X"5E",X"F0",X"17",X"91",X"71",X"21",X"EB",X"8A",X"0E",X"00",X"70",X"50",X"70",X"00",X"A8",
		X"00",X"00",X"00",X"00",X"01",X"00",X"F9",X"08",X"02",X"09",X"07",X"0E",X"88",X"00",X"80",X"00",
		X"C8",X"8B",X"0A",X"4A",X"4A",X"4B",X"48",X"4B",X"00",X"F8",X"08",X"08",X"18",X"F8",X"00",X"78",
		X"CB",X"4A",X"4A",X"4A",X"4A",X"7B",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"01",X"01",
		X"49",X"4B",X"C8",X"93",X"91",X"97",X"90",X"26",X"48",X"78",X"00",X"70",X"50",X"70",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"00",X"00",X"00",X"00",X"01",X"00",X"F9",X"08",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"03",
		X"CB",X"4A",X"4A",X"4A",X"4A",X"7B",X"00",X"00",X"C0",X"40",X"40",X"40",X"40",X"C0",X"00",X"00",
		X"18",X"18",X"18",X"00",X"01",X"06",X"0A",X"12",X"02",X"03",X"0E",X"3A",X"EA",X"AA",X"95",X"4F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"00",X"40",X"96",X"CC",X"28",X"98",X"51",X"36",X"00",X"00",X"08",X"18",X"24",X"53",X"AB",X"A6",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"30",X"1C",X"17",X"25",X"69",X"3A",
		X"BA",X"CA",X"A9",X"A5",X"97",X"7C",X"E0",X"80",X"9C",X"58",X"70",X"C0",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"E3",X"7F",X"AA",X"00",X"00",X"08",X"18",X"74",X"EB",X"56",X"AC",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"30",X"1C",X"17",X"25",X"69",X"3A",
		X"AA",X"AA",X"7F",X"00",X"00",X"00",X"00",X"00",X"B9",X"E1",X"05",X"77",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"00",X"06",X"00",X"00",X"00",X"0E",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"82",
		X"00",X"00",X"00",X"00",X"00",X"E3",X"7F",X"AA",X"00",X"00",X"08",X"18",X"74",X"EB",X"56",X"AC",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"02",X"0E",X"00",X"35",X"15",X"10",X"17",X"15",
		X"AA",X"AA",X"7F",X"00",X"00",X"00",X"00",X"00",X"B9",X"E1",X"05",X"77",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"00",X"06",X"00",X"00",X"00",X"77",X"00",X"07",X"05",X"BD",X"21",X"BF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EB",X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"03",X"03",X"03",X"00",X"03",X"00",X"00",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"00",X"00",X"19",X"17",X"19",X"17",X"19",X"17",X"00",X"00",X"C4",X"DC",X"E4",X"DC",X"E4",X"DC",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"19",X"17",X"19",X"17",X"19",X"0B",X"0C",X"0B",X"E4",X"DC",X"E4",X"CE",X"F2",X"EC",X"F0",X"EC",
		X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"6B",X"4C",X"4B",X"44",X"77",X"04",X"77",X"F0",X"EC",X"F0",X"FC",X"00",X"83",X"00",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"44",X"47",X"42",X"7B",X"02",X"4B",X"02",X"01",X"03",X"83",X"03",X"83",X"00",X"83",X"00",X"80",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"6D",X"29",X"6D",X"00",X"0E",X"08",X"08",X"0E",X"70",X"88",X"78",X"8E",X"BF",X"C7",X"5F",X"67",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"01",X"0B",X"03",X"07",X"0F",X"07",X"07",X"0F",X"5F",X"63",X"2F",X"B3",X"AF",X"B0",X"AC",X"90",
		X"18",X"18",X"18",X"00",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"00",X"02",X"00",X"02",X"00",X"DC",X"D0",X"DC",X"10",X"00",X"83",X"80",X"83",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"60",
		X"01",X"05",X"04",X"06",X"00",X"00",X"01",X"01",X"83",X"83",X"83",X"83",X"80",X"03",X"00",X"40",
		X"77",X"77",X"77",X"77",X"00",X"FF",X"00",X"88",X"60",X"60",X"60",X"60",X"00",X"E0",X"00",X"80",
		X"01",X"00",X"06",X"06",X"0E",X"0E",X"0B",X"09",X"40",X"08",X"E8",X"EE",X"E8",X"CE",X"11",X"1C",
		X"49",X"49",X"2A",X"00",X"3C",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"0F",X"00",X"6F",X"28",X"28",X"20",X"00",X"00",X"13",X"1D",X"93",X"A9",X"B5",X"00",X"00",X"00",
		X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"DF",X"3F",X"C7",X"47",X"FF",X"89",
		X"5D",X"79",X"51",X"77",X"6B",X"F3",X"A7",X"A7",X"10",X"10",X"FD",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"EF",X"B7",X"A7",X"E7",X"A7",X"BF",X"E7",X"A7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A7",X"E7",X"BF",X"A7",X"E7",X"A7",X"B7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A7",X"A7",X"F3",X"6B",X"77",X"51",X"79",X"5D",X"FB",X"E1",X"E1",X"E1",X"E3",X"FD",X"10",X"10",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"89",X"FF",X"47",X"C7",X"3F",X"DF",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",
		X"07",X"3F",X"D1",X"3F",X"C4",X"44",X"FE",X"89",X"FF",X"CB",X"2F",X"1F",X"BF",X"7F",X"7F",X"FF",
		X"5D",X"79",X"51",X"76",X"6A",X"F2",X"A4",X"A5",X"10",X"10",X"FD",X"23",X"21",X"21",X"21",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"B4",X"A4",X"E4",X"A7",X"BC",X"E4",X"A4",
		X"47",X"43",X"43",X"43",X"F3",X"4F",X"43",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",
		X"A4",X"E4",X"BC",X"A7",X"E4",X"A4",X"B4",X"EE",X"43",X"43",X"4F",X"F3",X"43",X"43",X"43",X"47",
		X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"A5",X"A4",X"F2",X"6A",X"76",X"51",X"79",X"5D",
		X"FB",X"21",X"21",X"21",X"23",X"FD",X"10",X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"89",X"FE",X"44",X"C4",X"3F",X"D1",X"3F",X"07",
		X"FF",X"7F",X"7F",X"BF",X"1F",X"2F",X"CB",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"0B",X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"D5",
		X"07",X"3F",X"D1",X"3F",X"C4",X"44",X"FE",X"89",X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",
		X"FC",X"37",X"2D",X"59",X"6F",X"5A",X"72",X"54",X"FF",X"A4",X"24",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"10",X"10",X"FD",X"23",X"21",X"21",X"21",X"FB",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A7",X"BD",X"E9",X"A9",X"A9",X"FF",X"A9",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F1",X"F1",
		X"46",X"42",X"42",X"42",X"F2",X"4E",X"42",X"42",X"00",X"00",X"00",X"07",X"0F",X"12",X"1F",X"14",
		X"A9",X"9F",X"F7",X"78",X"88",X"9F",X"F1",X"91",X"EB",X"47",X"8F",X"9F",X"BF",X"FF",X"FF",X"FF",
		X"42",X"42",X"4E",X"F2",X"42",X"42",X"42",X"46",X"14",X"1F",X"12",X"0F",X"07",X"00",X"00",X"00",
		X"91",X"F1",X"9F",X"88",X"78",X"F7",X"9F",X"A9",X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"47",X"EB",
		X"FB",X"21",X"21",X"21",X"23",X"FD",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"E9",X"A9",X"FF",X"A9",X"A9",X"E9",X"BD",X"A7",X"F1",X"F1",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"89",X"FE",X"44",X"C4",X"3F",X"D1",X"3F",X"07",X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",
		X"54",X"72",X"5A",X"6F",X"59",X"2D",X"37",X"FC",X"FF",X"FF",X"FF",X"FF",X"3F",X"24",X"A4",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",X"D5",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"D5",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"7F",
		X"FF",X"A4",X"24",X"3F",X"C8",X"88",X"88",X"9F",X"BF",X"FF",X"9F",X"9F",X"FF",X"9F",X"8B",X"89",
		X"F0",X"10",X"10",X"11",X"FE",X"1A",X"11",X"11",X"F9",X"FF",X"F9",X"F9",X"7D",X"FE",X"FE",X"FF",
		X"EB",X"47",X"8F",X"97",X"A7",X"47",X"27",X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"17",X"27",X"47",X"A7",X"97",X"8F",X"47",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"1A",X"FE",X"11",X"10",X"10",X"F0",X"FF",X"FE",X"FE",X"7D",X"F9",X"F9",X"FF",X"F9",
		X"9F",X"88",X"88",X"C8",X"3F",X"24",X"A4",X"FF",X"89",X"8B",X"9F",X"FF",X"9F",X"9F",X"FF",X"BF",
		X"D5",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"D5",X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"56",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",X"A4",X"24",X"3F",X"C8",X"88",X"88",X"9F",
		X"A9",X"FC",X"96",X"95",X"F2",X"9E",X"8B",X"89",X"7F",X"FF",X"5F",X"C4",X"7F",X"22",X"A2",X"7F",
		X"F0",X"10",X"10",X"11",X"FE",X"1A",X"11",X"11",X"F9",X"8F",X"89",X"F9",X"65",X"82",X"02",X"03",
		X"21",X"20",X"D0",X"7B",X"5F",X"BF",X"BB",X"39",X"EA",X"46",X"8C",X"94",X"A4",X"44",X"24",X"14",
		X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"79",X"77",X"F3",X"F3",X"F3",X"FB",X"FF",X"FE",
		X"14",X"24",X"44",X"A4",X"94",X"8C",X"46",X"EA",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",
		X"FE",X"FF",X"FB",X"F3",X"F3",X"F3",X"77",X"79",X"11",X"11",X"1A",X"FE",X"11",X"10",X"10",X"F0",
		X"03",X"02",X"82",X"65",X"F9",X"89",X"8F",X"F9",X"39",X"BB",X"BF",X"5F",X"7B",X"D0",X"20",X"21",
		X"9F",X"88",X"88",X"C8",X"3F",X"24",X"A4",X"FF",X"89",X"8B",X"9E",X"F2",X"95",X"96",X"FC",X"A9",
		X"7F",X"A2",X"22",X"7F",X"C4",X"5F",X"FF",X"7F",X"D5",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"56",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"56",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",X"A9",X"FC",X"96",X"95",X"F2",X"9E",X"8B",X"89",
		X"5F",X"E7",X"5F",X"C4",X"7F",X"22",X"A2",X"7F",X"FF",X"FF",X"C4",X"7F",X"C4",X"22",X"2F",X"FF",
		X"F9",X"8F",X"89",X"F9",X"65",X"82",X"02",X"03",X"21",X"20",X"D0",X"6B",X"55",X"AD",X"AB",X"29",
		X"0F",X"8F",X"87",X"FF",X"3F",X"1F",X"9F",X"9F",X"03",X"03",X"02",X"04",X"04",X"05",X"06",X"04",
		X"49",X"56",X"D3",X"52",X"D2",X"5A",X"57",X"52",X"6F",X"4F",X"47",X"A7",X"7F",X"A7",X"27",X"27",
		X"04",X"06",X"05",X"04",X"04",X"02",X"03",X"03",X"52",X"57",X"5A",X"D2",X"52",X"D3",X"56",X"49",
		X"27",X"27",X"A7",X"7F",X"A7",X"47",X"4F",X"6F",X"03",X"02",X"82",X"65",X"F9",X"89",X"8F",X"F9",
		X"29",X"AB",X"AD",X"55",X"6B",X"D0",X"20",X"21",X"9F",X"9F",X"1F",X"3F",X"FF",X"87",X"8F",X"0F",
		X"89",X"8B",X"9E",X"F2",X"95",X"96",X"FC",X"A9",X"7F",X"A2",X"22",X"7F",X"C4",X"5F",X"E7",X"5F",
		X"FF",X"2F",X"22",X"C4",X"7F",X"C4",X"FF",X"FF",X"56",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"5F",X"E4",X"5F",X"C4",X"7F",X"22",X"A2",X"7F",
		X"CF",X"7F",X"C4",X"7F",X"C4",X"22",X"2F",X"F1",X"FF",X"8F",X"3D",X"C4",X"03",X"0E",X"FE",X"FE",
		X"21",X"20",X"D0",X"6B",X"55",X"AD",X"AB",X"29",X"08",X"88",X"87",X"FE",X"22",X"11",X"91",X"9F",
		X"FF",X"7F",X"FF",X"3F",X"1F",X"1F",X"3F",X"CF",X"49",X"56",X"D3",X"52",X"D2",X"5A",X"57",X"52",
		X"68",X"48",X"44",X"A4",X"7F",X"A4",X"24",X"24",X"8F",X"8F",X"8F",X"9F",X"E7",X"47",X"47",X"47",
		X"52",X"57",X"5A",X"D2",X"52",X"D3",X"56",X"49",X"24",X"24",X"A4",X"7F",X"A4",X"44",X"48",X"68",
		X"47",X"47",X"47",X"E7",X"9F",X"8F",X"8F",X"8F",X"29",X"AB",X"AD",X"55",X"6B",X"D0",X"20",X"21",
		X"9F",X"91",X"11",X"22",X"FE",X"87",X"88",X"08",X"CF",X"3F",X"1F",X"1F",X"3F",X"FF",X"7F",X"FF",
		X"7F",X"A2",X"22",X"7F",X"C4",X"5F",X"E4",X"5F",X"F1",X"2F",X"22",X"C4",X"7F",X"C4",X"7F",X"CF",
		X"FE",X"FE",X"0E",X"03",X"C4",X"3D",X"8F",X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",X"00",X"00",X"00",X"00",X"00",X"0F",X"F7",X"17",
		X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",X"C8",X"7F",X"C4",X"7F",X"C4",X"22",X"2F",X"F1",
		X"79",X"8B",X"3D",X"C4",X"03",X"0E",X"F2",X"02",X"EF",X"FF",X"FF",X"FF",X"FE",X"BF",X"BF",X"9F",
		X"08",X"88",X"87",X"FE",X"22",X"11",X"91",X"9F",X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",
		X"FC",X"5C",X"5C",X"4D",X"4E",X"EA",X"3A",X"2E",X"68",X"48",X"44",X"A4",X"7F",X"A4",X"24",X"24",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",
		X"24",X"24",X"A4",X"7F",X"A4",X"44",X"48",X"68",X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",
		X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",X"9F",X"91",X"11",X"22",X"FE",X"87",X"88",X"08",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"2E",X"3A",X"EA",X"4E",X"4D",X"5C",X"5C",X"FC",
		X"F1",X"2F",X"22",X"C4",X"7F",X"C4",X"7F",X"C8",X"02",X"F2",X"0E",X"03",X"C4",X"3D",X"8B",X"79",
		X"9F",X"BF",X"BF",X"FE",X"FF",X"FF",X"FF",X"EF",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"17",X"F7",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"79",X"8B",X"3D",X"C4",X"03",X"0E",X"F2",X"02",X"6F",X"FF",X"7F",X"BF",X"FE",X"BF",X"AF",X"9F",
		X"83",X"4E",X"F1",X"21",X"11",X"11",X"3F",X"C9",X"F4",X"5C",X"54",X"4D",X"4E",X"EA",X"3A",X"2E",
		X"88",X"88",X"88",X"9F",X"E4",X"44",X"44",X"44",X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",
		X"44",X"44",X"44",X"E4",X"9F",X"88",X"88",X"88",X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",
		X"C9",X"3F",X"11",X"11",X"21",X"F1",X"4E",X"83",X"2E",X"3A",X"EA",X"4E",X"4D",X"54",X"5C",X"F4",
		X"02",X"F2",X"0E",X"03",X"C4",X"3D",X"8B",X"79",X"9F",X"AF",X"BF",X"FE",X"BF",X"7F",X"FF",X"6F",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",X"00",X"00",X"07",X"1F",X"7F",X"FC",X"E8",X"C7",
		X"6B",X"F4",X"7C",X"B3",X"F6",X"B9",X"A9",X"9B",X"0E",X"B2",X"C1",X"23",X"3F",X"7F",X"9F",X"1F",
		X"F4",X"5C",X"54",X"4D",X"4E",X"EA",X"3A",X"2E",X"8F",X"BF",X"CF",X"87",X"47",X"47",X"7F",X"C7",
		X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",X"47",X"47",X"47",X"47",X"7F",X"C7",X"47",X"47",
		X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",X"47",X"47",X"C7",X"7F",X"47",X"47",X"47",X"47",
		X"2E",X"3A",X"EA",X"4E",X"4D",X"54",X"5C",X"F4",X"C7",X"7F",X"47",X"47",X"87",X"CF",X"BF",X"8F",
		X"9B",X"A9",X"B9",X"F6",X"B3",X"7C",X"F4",X"6B",X"1F",X"9F",X"7F",X"3F",X"23",X"C1",X"B2",X"0E",
		X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",X"C7",X"E8",X"FC",X"7F",X"1F",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",X"00",X"00",X"07",X"18",X"73",X"9C",X"28",X"C7",
		X"00",X"C0",X"40",X"60",X"A0",X"10",X"70",X"88",X"6B",X"F4",X"7C",X"B3",X"F6",X"B9",X"A9",X"9B",
		X"0E",X"B2",X"C1",X"23",X"3D",X"70",X"90",X"10",X"08",X"08",X"78",X"84",X"04",X"84",X"8E",X"F2",
		X"F4",X"5C",X"54",X"4D",X"4E",X"EA",X"3A",X"2E",X"8F",X"B8",X"C8",X"84",X"44",X"47",X"7C",X"C4",
		X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",X"AB",X"AA",X"AA",X"FA",X"AE",X"AB",X"AA",X"AA",
		X"44",X"44",X"44",X"45",X"7E",X"C4",X"44",X"44",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"AA",X"AA",X"AB",X"AE",X"FA",X"AA",X"AA",X"AB",X"44",X"44",X"C4",X"7E",X"45",X"44",X"44",X"44",
		X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"2E",X"3A",X"EA",X"4E",X"4D",X"54",X"5C",X"F4",
		X"C4",X"7C",X"47",X"44",X"84",X"C8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"9B",X"A9",X"B9",X"F6",X"B3",X"7C",X"F4",X"6B",X"10",X"90",X"70",X"3D",X"23",X"C1",X"B2",X"0E",
		X"F2",X"8E",X"84",X"04",X"84",X"78",X"08",X"08",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"28",X"9C",X"73",X"18",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"60",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"43",X"2C",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"3E",X"7F",X"7F",X"3E",X"1C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"3C",X"3E",X"3E",X"1E",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"3C",X"1C",X"1E",X"0E",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"04",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"10",X"10",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"10",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"3E",X"7F",X"3E",X"1C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",X"7E",X"7F",X"3C",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"FF",X"78",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"D5",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FC",X"E8",X"C7",X"00",X"C0",X"C0",X"E0",X"A0",X"10",X"70",X"88",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"C7",X"C7",X"FF",X"89",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F9",X"EF",X"DB",X"F3",X"D7",
		X"FF",X"A4",X"24",X"3F",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"9F",X"9F",X"FF",X"9F",X"8B",X"89",
		X"FF",X"FF",X"DF",X"C4",X"FF",X"E2",X"E2",X"7F",X"FF",X"FF",X"C4",X"7F",X"C4",X"22",X"2F",X"FF",
		X"FF",X"8F",X"3D",X"C4",X"03",X"0E",X"FE",X"FE",X"EF",X"FF",X"FF",X"FF",X"FE",X"BF",X"BF",X"9F",
		X"0E",X"B2",X"C1",X"23",X"3F",X"7F",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"7D",X"79",X"71",X"77",X"6B",X"F3",X"E7",X"E7",X"10",X"10",X"FD",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A7",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F1",X"F1",X"F9",X"FF",X"F9",X"F9",X"FD",X"FE",X"FE",X"FF",
		X"21",X"20",X"D0",X"7B",X"5F",X"BF",X"BB",X"39",X"0F",X"8F",X"87",X"FF",X"3F",X"1F",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"DC",X"DC",X"CD",X"CE",X"EA",X"FA",X"EE",
		X"8F",X"BF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"BF",X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"88",X"9F",X"FF",X"FF",
		X"EB",X"C7",X"8F",X"9F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"79",X"77",X"F3",X"F3",X"F3",X"FB",X"FF",X"FE",X"EF",X"CF",X"C7",X"E7",X"FF",X"A7",X"27",X"27",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"EA",X"EA",X"FA",X"EE",X"EB",X"EA",X"EA",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"BF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"88",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"C7",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FB",X"F3",X"F3",X"F3",X"77",X"79",X"27",X"27",X"A7",X"FF",X"E7",X"C7",X"CF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"EA",X"EB",X"EE",X"FA",X"EA",X"EA",X"EB",
		X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E7",X"E7",X"F3",X"6B",X"77",X"71",X"79",X"7D",X"FB",X"E1",X"E1",X"E1",X"E3",X"FD",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"A7",
		X"F1",X"F1",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FD",X"F9",X"F9",X"FF",X"F9",
		X"39",X"BB",X"BF",X"5F",X"7B",X"D0",X"20",X"21",X"9F",X"9F",X"1F",X"3F",X"FF",X"87",X"8F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FA",X"EA",X"CE",X"CD",X"DC",X"DC",X"FC",
		X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"BF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"89",X"FF",X"C7",X"C7",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"F3",X"DB",X"EF",X"F9",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"24",X"A4",X"FF",X"89",X"8B",X"9F",X"FF",X"9F",X"9F",X"FF",X"BF",
		X"7F",X"E2",X"E2",X"FF",X"C4",X"DF",X"FF",X"FF",X"FF",X"2F",X"22",X"C4",X"7F",X"C4",X"FF",X"FF",
		X"FE",X"FE",X"0E",X"03",X"C4",X"3D",X"8F",X"FF",X"9F",X"BF",X"BF",X"FE",X"FF",X"FF",X"FF",X"EF",
		X"1F",X"9F",X"7F",X"3F",X"23",X"C1",X"B2",X"0E",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"D5",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E8",X"FC",X"7F",X"1F",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F5",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FC",X"E8",X"C7",X"00",X"C0",X"C0",X"E0",X"A0",X"10",X"70",X"88",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"C7",X"C7",X"FF",X"89",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F9",X"EF",X"DB",X"F3",X"D7",
		X"FF",X"A8",X"28",X"7F",X"FF",X"FF",X"FF",X"FF",X"EF",X"BF",X"97",X"F7",X"FB",X"FF",X"F9",X"F9",
		X"FF",X"FF",X"DF",X"C4",X"FF",X"E2",X"E1",X"7F",X"FF",X"FF",X"C4",X"7F",X"C4",X"22",X"2F",X"FF",
		X"FF",X"8F",X"3D",X"C4",X"03",X"0E",X"FE",X"FE",X"EF",X"FF",X"FF",X"FF",X"FE",X"BF",X"BF",X"9F",
		X"0E",X"B2",X"C1",X"23",X"3F",X"7F",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"7D",X"79",X"71",X"77",X"6B",X"F3",X"E7",X"E7",X"10",X"10",X"FD",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A7",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F1",X"F3",X"FC",X"FF",X"FD",X"FC",X"FC",X"FF",X"FF",X"FF",
		X"A0",X"A0",X"F8",X"B7",X"FB",X"BD",X"3E",X"7F",X"8F",X"8F",X"47",X"FF",X"1F",X"0F",X"8F",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"DC",X"DC",X"CD",X"CE",X"EA",X"FA",X"EE",
		X"8F",X"BF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"BF",X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"88",X"9F",X"FF",X"FF",
		X"EB",X"C7",X"8F",X"9F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FD",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"EF",X"E7",X"E3",X"F3",X"FF",X"D3",X"D3",X"93",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"EA",X"EA",X"FA",X"EE",X"EB",X"EA",X"EA",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"BF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"88",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"9F",X"8F",X"C7",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FD",X"7F",X"93",X"D3",X"D3",X"FF",X"F3",X"E3",X"E7",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"EA",X"EB",X"EE",X"FA",X"EA",X"EA",X"EB",
		X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E7",X"E7",X"F3",X"6B",X"77",X"71",X"79",X"7D",X"FB",X"E1",X"E1",X"E1",X"E3",X"FD",X"10",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"A7",
		X"F3",X"F1",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FD",X"FF",X"FC",
		X"7F",X"3E",X"BD",X"FB",X"B7",X"F8",X"A0",X"A0",X"DF",X"8F",X"0F",X"1F",X"FF",X"47",X"8F",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FA",X"EA",X"CE",X"CD",X"DC",X"DC",X"FC",
		X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"BF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"89",X"FF",X"C7",X"C7",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"F3",X"DB",X"EF",X"F9",X"FD",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"28",X"A8",X"FF",X"F9",X"F9",X"FF",X"FB",X"F7",X"97",X"BF",X"EF",
		X"7F",X"E1",X"E2",X"FF",X"C4",X"DF",X"FF",X"FF",X"FF",X"2F",X"22",X"C4",X"7F",X"C4",X"FF",X"FF",
		X"FE",X"FE",X"0E",X"03",X"C4",X"3D",X"8F",X"FF",X"9F",X"BF",X"BF",X"FE",X"FF",X"FF",X"FF",X"EF",
		X"1F",X"9F",X"7F",X"3F",X"23",X"C1",X"B2",X"0E",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F5",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"5F",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E8",X"FC",X"7F",X"1F",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F2",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FC",X"E8",X"C7",X"00",X"C0",X"C0",X"E0",X"A0",X"10",X"70",X"88",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"C7",X"CF",X"FF",X"91",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"CF",X"F3",X"D7",X"A7",X"AF",
		X"FF",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"5F",X"DF",X"FF",X"EB",X"E9",X"FF",X"FD",
		X"FF",X"FF",X"DF",X"C4",X"FF",X"E2",X"61",X"BF",X"FF",X"FF",X"C4",X"7F",X"C2",X"21",X"1F",X"FF",
		X"FF",X"8F",X"3D",X"C4",X"03",X"0E",X"FE",X"FE",X"EF",X"FF",X"FF",X"FF",X"FE",X"BF",X"BF",X"9F",
		X"0E",X"B2",X"C1",X"23",X"3F",X"7F",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"7D",X"7A",X"73",X"77",X"6F",X"F7",X"EF",X"EF",X"10",X"20",X"FD",X"E3",X"C1",X"C3",X"C3",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"D3",X"CF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"E0",X"A0",X"B8",X"B7",X"FB",X"BC",X"3E",X"7F",X"8F",X"87",X"47",X"FF",X"BF",X"1F",X"0F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"DC",X"DC",X"CD",X"CE",X"EA",X"FA",X"EE",
		X"8F",X"BF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"BF",X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"7F",X"FF",X"F9",X"93",X"FF",X"FF",X"FF",
		X"87",X"8F",X"1F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"C7",X"C3",X"E3",X"73",X"FF",X"29",X"29",X"29",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"EA",X"EA",X"FA",X"EE",X"EB",X"EA",X"EA",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"BF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"93",X"F9",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"1F",X"8F",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"7F",X"29",X"29",X"29",X"FF",X"73",X"E3",X"C3",X"C7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"EA",X"EB",X"EE",X"FA",X"EA",X"EA",X"EB",
		X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"F7",X"6F",X"77",X"73",X"7A",X"7D",X"FB",X"C3",X"C3",X"C1",X"E3",X"FD",X"20",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"BF",
		X"CF",X"D3",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"7F",X"3E",X"BC",X"FB",X"B7",X"B8",X"A0",X"E0",X"3F",X"0F",X"1F",X"BF",X"FF",X"47",X"87",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FA",X"EA",X"CE",X"CD",X"DC",X"DC",X"FC",
		X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"BF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"91",X"FF",X"CF",X"C7",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"A7",X"D7",X"F3",X"CF",X"F9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"FF",X"FD",X"FF",X"E9",X"EB",X"FF",X"DF",X"5F",X"F7",
		X"BF",X"61",X"E2",X"FF",X"C4",X"DF",X"FF",X"FF",X"FF",X"1F",X"21",X"C2",X"7F",X"C4",X"FF",X"FF",
		X"FE",X"FE",X"0E",X"03",X"C4",X"3D",X"8F",X"FF",X"9F",X"BF",X"BF",X"FE",X"FF",X"FF",X"FF",X"EF",
		X"1F",X"9F",X"7F",X"3F",X"23",X"C1",X"B2",X"0E",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"AF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E8",X"FC",X"7F",X"1F",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F2",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"AF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",
		X"00",X"00",X"07",X"1F",X"7F",X"FC",X"E8",X"C7",X"00",X"C0",X"C0",X"E0",X"A0",X"10",X"70",X"88",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"FF",X"FF",X"C7",X"CF",X"FF",X"91",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"CF",X"F3",X"D7",X"A7",X"AF",
		X"FF",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"5F",X"DF",X"FF",X"EB",X"E9",X"FF",X"FD",
		X"FF",X"FF",X"DF",X"C4",X"FF",X"E2",X"61",X"BF",X"FF",X"FF",X"C4",X"7F",X"C2",X"21",X"1F",X"FF",
		X"FF",X"8F",X"3D",X"C4",X"03",X"0E",X"FE",X"FE",X"EF",X"FF",X"FF",X"FF",X"FE",X"BF",X"BF",X"9F",
		X"0E",X"B2",X"C1",X"23",X"3F",X"7F",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"7D",X"7A",X"73",X"77",X"6F",X"F7",X"EF",X"EF",X"10",X"20",X"FD",X"E3",X"C1",X"C3",X"C3",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"D3",X"CF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"E0",X"A0",X"B8",X"B7",X"FB",X"B8",X"3E",X"7F",X"8F",X"87",X"47",X"FF",X"9F",X"EF",X"5F",X"2F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"DC",X"DC",X"CD",X"CE",X"EA",X"FA",X"EE",
		X"8F",X"BF",X"FF",X"FF",X"7F",X"7F",X"7F",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"BF",X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"7F",X"FF",X"F9",X"93",X"FF",X"FF",X"FF",
		X"87",X"8F",X"1F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FB",X"FD",X"FD",X"FA",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"EA",X"EA",X"FA",X"EE",X"EB",X"EA",X"EA",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"BF",X"BF",X"FF",X"BF",X"BF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"F2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"93",X"F9",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"1F",X"8F",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FE",X"FE",X"FE",X"FA",X"FD",X"FD",X"FB",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EA",X"EA",X"EB",X"EE",X"FA",X"EA",X"EA",X"EB",
		X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"F7",X"6F",X"77",X"73",X"7A",X"7D",X"FB",X"C3",X"C3",X"C1",X"E3",X"FD",X"20",X"10",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"FF",X"BF",
		X"CF",X"D3",X"F3",X"FB",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FE",X"FC",X"FC",
		X"7F",X"3E",X"B8",X"FB",X"B7",X"B8",X"A0",X"E0",X"2F",X"5F",X"EF",X"9F",X"FF",X"47",X"87",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FA",X"EA",X"CE",X"CD",X"DC",X"DC",X"FC",
		X"FF",X"7F",X"7F",X"7F",X"FF",X"FF",X"BF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"91",X"FF",X"CF",X"C7",X"FF",X"FF",X"3F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"A7",X"D7",X"F3",X"CF",X"F9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"FF",X"FD",X"FF",X"E9",X"EB",X"FF",X"DF",X"5F",X"F7",
		X"BF",X"61",X"E2",X"FF",X"C4",X"DF",X"FF",X"FF",X"FF",X"1F",X"21",X"C2",X"7F",X"C4",X"FF",X"FF",
		X"FE",X"FE",X"0E",X"03",X"C4",X"3D",X"8F",X"FF",X"9F",X"BF",X"BF",X"FE",X"FF",X"FF",X"FF",X"EF",
		X"1F",X"9F",X"7F",X"3F",X"23",X"C1",X"B2",X"0E",X"FE",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F2",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"AF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"C7",X"E8",X"FC",X"7F",X"1F",X"07",X"00",X"00",X"88",X"70",X"10",X"A0",X"E0",X"C0",X"C0",X"00",
		X"FF",X"FF",X"07",X"47",X"47",X"FF",X"4F",X"4F",X"4F",X"4F",X"4F",X"FF",X"47",X"47",X"47",X"FF",
		X"39",X"83",X"C3",X"C3",X"81",X"E1",X"78",X"7E",X"01",X"81",X"00",X"7E",X"60",X"60",X"68",X"78",
		X"0C",X"00",X"00",X"00",X"C0",X"80",X"00",X"40",X"6D",X"01",X"01",X"C3",X"01",X"01",X"08",X"46",
		X"81",X"87",X"1E",X"7E",X"7C",X"6C",X"68",X"68",X"3C",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"C0",
		X"E3",X"07",X"03",X"C3",X"81",X"01",X"78",X"7C",X"01",X"01",X"00",X"7E",X"0C",X"04",X"E0",X"F0",
		X"34",X"00",X"00",X"00",X"60",X"60",X"40",X"40",X"FF",X"F7",X"E3",X"C3",X"81",X"01",X"60",X"72",
		X"08",X"83",X"47",X"B8",X"DD",X"ED",X"61",X"06",X"06",X"80",X"81",X"33",X"20",X"21",X"29",X"34",
		X"8F",X"01",X"00",X"77",X"81",X"00",X"36",X"76",X"65",X"01",X"00",X"DE",X"01",X"01",X"0C",X"46",
		X"CE",X"EF",X"77",X"B8",X"5D",X"6D",X"61",X"04",X"44",X"00",X"83",X"33",X"BC",X"BF",X"BB",X"B4",
		X"83",X"07",X"00",X"77",X"83",X"00",X"74",X"74",X"65",X"01",X"00",X"DE",X"0F",X"03",X"60",X"70",
		X"46",X"01",X"01",X"B8",X"5D",X"6D",X"61",X"04",X"C6",X"98",X"BB",X"33",X"8C",X"09",X"21",X"30",
		X"08",X"81",X"80",X"A8",X"20",X"20",X"2F",X"88",X"20",X"81",X"00",X"00",X"00",X"60",X"28",X"28",
		X"08",X"00",X"00",X"28",X"00",X"00",X"20",X"20",X"28",X"00",X"00",X"28",X"00",X"00",X"88",X"00",
		X"08",X"A9",X"A8",X"A8",X"20",X"20",X"2D",X"08",X"28",X"01",X"00",X"00",X"00",X"EC",X"28",X"28",
		X"20",X"00",X"08",X"28",X"00",X"00",X"28",X"28",X"28",X"00",X"00",X"28",X"08",X"00",X"A0",X"20",
		X"00",X"01",X"00",X"A8",X"20",X"20",X"2D",X"08",X"28",X"AD",X"00",X"00",X"00",X"08",X"20",X"20",
		X"30",X"00",X"C0",X"40",X"70",X"10",X"77",X"45",X"10",X"00",X"40",X"50",X"41",X"00",X"6D",X"00",
		X"07",X"01",X"01",X"15",X"01",X"00",X"10",X"10",X"6D",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"10",X"F0",X"40",X"70",X"00",X"65",X"45",X"10",X"00",X"00",X"50",X"5F",X"00",X"FF",X"00",
		X"03",X"05",X"05",X"15",X"03",X"00",X"10",X"10",X"6D",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"70",X"00",X"00",X"40",X"70",X"00",X"65",X"45",X"10",X"10",X"50",X"50",X"0D",X"00",X"61",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FA",X"6E",X"00",X"00",X"00",X"FC",X"E7",X"00",X"C0",X"00",X"01",X"02",X"05",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",
		X"F9",X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"00",X"00",X"00",X"0C",X"10",X"01",
		X"00",X"00",X"0F",X"18",X"07",X"0F",X"07",X"C0",X"0B",X"1F",X"DF",X"7F",X"FF",X"FF",X"BF",X"37",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FF",X"F7",X"FF",X"F8",X"CF",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"DF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FC",X"FC",X"F8",X"F8",X"78",X"C8",X"0E",X"03",
		X"00",X"30",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"1C",X"00",X"00",X"00",X"08",X"00",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"23",X"13",X"01",X"08",X"00",X"08",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A8",X"F8",X"FB",X"05",X"08",X"F9",X"E9",X"E8",X"01",X"00",X"00",X"C0",X"00",X"80",X"01",X"07",
		X"80",X"C1",X"48",X"4A",X"40",X"00",X"02",X"34",X"00",X"90",X"34",X"18",X"C6",X"20",X"F8",X"DE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"04",X"00",X"00",X"00",X"00",X"20",X"10",X"08",X"00",
		X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"C2",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"0C",X"38",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"08",X"06",X"00",X"12",X"18",X"23",X"68",X"D7",X"2E",X"1B",X"44",X"FA",X"0E",X"B8",X"E0",X"CC",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"05",X"09",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"20",X"00",X"80",X"E1",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"01",X"DF",X"7F",X"80",X"E0",
		X"BF",X"3F",X"1F",X"0E",X"03",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"37",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"E0",X"FE",X"FF",X"FF",X"FF",X"03",X"03",X"01",X"00",X"00",X"C0",X"E1",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"F8",X"C6",X"30",X"10",X"FF",X"FF",X"FF",X"7F",X"FF",X"00",X"20",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",
		X"02",X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",X"00",X"00",X"20",X"07",X"38",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F8",X"E3",X"E0",X"CB",X"91",X"00",X"00",X"11",X"01",
		X"F8",X"2D",X"EF",X"FF",X"3D",X"79",X"E7",X"E0",X"FF",X"03",X"0C",X"00",X"06",X"1F",X"FF",X"40",
		X"FF",X"FF",X"FF",X"BE",X"4E",X"94",X"E9",X"67",X"00",X"00",X"02",X"0D",X"00",X"20",X"E6",X"CC",
		X"00",X"00",X"84",X"20",X"46",X"82",X"20",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F8",X"F8",X"FE",X"FF",X"FF",X"FF",X"23",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"80",X"EF",X"FB",X"EA",X"1F",X"FC",X"7F",X"00",X"28",X"00",X"83",X"81",X"00",X"00",X"41",
		X"03",X"02",X"83",X"84",X"0C",X"18",X"F0",X"E1",X"FB",X"FF",X"7F",X"7F",X"39",X"23",X"7F",X"C0",
		X"1A",X"63",X"FE",X"FF",X"FF",X"FB",X"E1",X"FF",X"00",X"80",X"38",X"C3",X"DF",X"FE",X"DF",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"BF",X"8F",X"C6",X"F0",X"FD",X"FF",
		X"BF",X"FF",X"FF",X"F8",X"43",X"1F",X"FF",X"FF",X"FF",X"79",X"CB",X"8F",X"3F",X"FF",X"FF",X"FF",
		X"9F",X"FF",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"80",X"40",X"00",X"20",X"00",X"00",X"30",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"07",X"A3",X"9F",X"97",X"CF",X"EF",X"E7",
		X"00",X"84",X"80",X"FF",X"57",X"BF",X"E0",X"F8",X"00",X"00",X"80",X"E8",X"40",X"80",X"00",X"7C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BB",X"04",X"80",X"FC",X"FF",X"FF",X"FF",X"FF",X"A0",X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"24",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"C7",X"B2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"C0",X"80",X"C0",X"00",X"80",
		X"41",X"30",X"03",X"00",X"08",X"00",X"00",X"00",X"FF",X"3F",X"C3",X"7C",X"0F",X"8F",X"0F",X"00",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"E0",X"0A",X"10",X"E0",X"8F",X"3F",X"7F",X"FF",X"E1",
		X"3F",X"0F",X"07",X"FF",X"E3",X"70",X"B0",X"A0",X"FF",X"FF",X"FF",X"DF",X"E7",X"08",X"07",X"67",
		X"FF",X"FE",X"FE",X"F7",X"EC",X"FF",X"FE",X"C0",X"00",X"00",X"20",X"98",X"08",X"04",X"12",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E1",X"C1",X"E9",X"E0",X"E0",X"E0",X"F0",X"F0",X"C1",X"C0",X"C0",X"60",X"30",X"1F",X"FF",X"3D",
		X"81",X"1F",X"00",X"01",X"87",X"A0",X"A0",X"E0",X"F7",X"BA",X"00",X"00",X"B0",X"30",X"01",X"0F",
		X"E0",X"F0",X"40",X"C0",X"C0",X"F0",X"E0",X"80",X"0C",X"0E",X"01",X"0F",X"18",X"00",X"00",X"00",
		X"80",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"1B",X"FF",X"4C",X"00",X"E3",X"FF",X"FF",
		X"E0",X"C3",X"FF",X"0C",X"3F",X"FF",X"FF",X"FF",X"1B",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"F8",X"E1",X"F4",X"F8",X"FC",X"FC",X"FE",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"C0",X"63",X"21",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"BF",X"70",X"FC",X"FF",X"FF",X"FF",X"FF",X"07",X"C0",X"00",X"7F",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"C0",X"E0",X"C0",X"F0",X"F8",X"F8",X"F6",X"00",X"01",X"03",X"03",X"03",X"03",X"03",X"01",
		X"00",X"80",X"C0",X"80",X"E0",X"F0",X"F0",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",
		X"01",X"01",X"01",X"81",X"80",X"C0",X"C0",X"E0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"7C",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"40",X"40",X"C1",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",
		X"00",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"80",X"83",X"83",X"87",X"87",X"8F",X"57",X"6B",
		X"E0",X"70",X"30",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"10",X"10",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"0B",X"1B",X"3B",X"37",X"37",X"07",X"0F",X"EF",X"DF",X"DE",X"DE",X"BE",X"BE",
		X"6B",X"6D",X"6D",X"3C",X"BC",X"DE",X"DE",X"DE",X"80",X"00",X"00",X"00",X"00",X"00",X"81",X"81",
		X"3E",X"3E",X"3F",X"5F",X"DF",X"EF",X"AF",X"B7",X"04",X"04",X"00",X"22",X"A1",X"91",X"D0",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"37",X"2F",X"2F",X"2F",X"1F",X"1E",X"1E",
		X"7E",X"7E",X"7F",X"7F",X"7D",X"6D",X"EE",X"F6",X"D6",X"F7",X"7B",X"7B",X"7D",X"BD",X"BE",X"BE",
		X"A3",X"D3",X"DB",X"D3",X"D5",X"F9",X"FA",X"FA",X"D7",X"DB",X"EB",X"ED",X"DD",X"DA",X"BA",X"BD",
		X"E8",X"E4",X"B4",X"70",X"D8",X"B0",X"E0",X"68",X"40",X"40",X"20",X"20",X"00",X"00",X"20",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"0E",X"06",X"02",X"01",X"01",X"01",X"01",X"D7",X"DF",X"EF",X"EF",X"FF",X"BE",X"BE",X"D6",
		X"5E",X"5E",X"5E",X"5E",X"3D",X"BD",X"AD",X"AD",X"F8",X"F4",X"B5",X"B5",X"DD",X"DD",X"EB",X"6B",
		X"7D",X"7B",X"3B",X"3F",X"9F",X"9F",X"CF",X"CF",X"5C",X"BC",X"FE",X"FE",X"BF",X"FF",X"FF",X"FF",
		X"10",X"18",X"08",X"0C",X"04",X"06",X"82",X"83",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"D6",X"DB",X"DB",X"DD",X"BD",X"BD",X"BD",X"BD",X"B7",X"B7",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"6B",X"AB",X"AB",X"DB",X"D7",X"D7",X"C7",X"87",X"E7",X"E7",X"F3",X"F3",X"FB",X"FB",X"FB",X"FB",
		X"FF",X"FF",X"FE",X"FC",X"F9",X"FA",X"FC",X"FD",X"C1",X"C1",X"E0",X"E0",X"70",X"70",X"B0",X"20",
		X"40",X"A0",X"A0",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",
		X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FE",X"7C",X"7C",X"BC",X"BC",
		X"40",X"80",X"00",X"00",X"28",X"28",X"34",X"34",X"00",X"00",X"00",X"00",X"60",X"60",X"30",X"30",
		X"00",X"00",X"00",X"00",X"86",X"86",X"43",X"43",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"BD",X"BF",X"7F",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DC",X"DC",X"E8",X"E8",X"F0",X"F0",X"F8",X"F8",X"39",X"38",X"7C",X"7C",X"7E",X"7E",X"7F",X"7F",
		X"FC",X"48",X"EC",X"EC",X"76",X"76",X"24",X"00",X"1F",X"04",X"0E",X"0E",X"07",X"07",X"02",X"00",
		X"C0",X"80",X"C0",X"C0",X"60",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"1E",X"1E",X"1E",X"1C",X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",X"FC",X"7C",X"3E",X"1E",X"0E",X"06",X"00",X"00",
		X"3F",X"3F",X"1F",X"1F",X"0E",X"0E",X"06",X"06",X"00",X"00",X"10",X"36",X"2E",X"3F",X"3F",X"3F",
		X"00",X"00",X"01",X"03",X"02",X"03",X"03",X"C3",X"00",X"00",X"00",X"60",X"E0",X"F0",X"F0",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"0D",X"0D",X"0D",X"0D",X"0D",X"03",X"02",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"1C",X"1C",X"08",X"08",X"04",X"04",X"02",X"23",X"11",X"11",X"08",X"08",X"10",X"10",X"20",
		X"E2",X"C1",X"C1",X"80",X"80",X"41",X"41",X"22",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"02",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",
		X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",
		X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",X"80",X"80",X"C0",X"40",X"20",X"20",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"40",X"80",X"09",X"09",X"0C",X"0C",X"1E",X"1E",X"00",X"00",X"00",X"00",X"80",X"A0",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"0F",X"1F",X"1F",X"5F",X"5F",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"1F",X"1F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"40",X"20",X"80",X"80",X"80",X"80",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"F7",X"F7",X"FB",X"FB",X"F9",X"F9",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"88",X"88",X"08",X"10",X"10",X"10",X"10",X"00",
		X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"7E",X"7E",X"BE",X"BE",X"DE",X"DE",X"EE",X"EF",
		X"00",X"00",X"00",X"00",X"30",X"70",X"F8",X"88",X"7E",X"7E",X"3E",X"3E",X"1E",X"1E",X"0C",X"0C",
		X"00",X"00",X"00",X"20",X"20",X"20",X"70",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F7",X"F7",X"FB",X"FB",X"7D",X"7D",X"3E",X"3E",X"04",X"04",X"04",X"04",X"88",X"F8",X"F8",X"F8",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"74",X"28",X"28",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"3F",X"6F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"78",X"78",X"B0",X"B0",X"D0",X"D0",X"E0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"7F",X"7F",X"B0",X"30",X"58",X"98",X"2C",X"48",X"90",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"C0",X"80",X"0A",X"0A",X"0D",X"0D",X"0E",X"0E",X"00",X"00",X"18",X"18",X"0C",X"0C",X"7F",X"12",
		X"00",X"00",X"21",X"21",X"10",X"10",X"07",X"01",X"00",X"00",X"80",X"80",X"C0",X"C0",X"F0",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",
		X"3B",X"3B",X"9D",X"9D",X"C9",X"C0",X"C0",X"C0",X"03",X"03",X"81",X"81",X"00",X"00",X"00",X"00",
		X"B0",X"B0",X"D8",X"D8",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"C4",X"CD",X"8B",X"8F",X"8F",X"8F",X"8F",X"87",
		X"00",X"80",X"80",X"C0",X"C0",X"F0",X"88",X"04",X"40",X"D8",X"B8",X"FC",X"FC",X"FF",X"F8",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"04",X"02",X"02",X"04",X"04",X"88",X"70",X"00",
		X"70",X"20",X"20",X"10",X"10",X"08",X"07",X"00",X"40",X"20",X"20",X"40",X"40",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"B9",X"BB",X"7F",
		X"0F",X"0F",X"07",X"37",X"7B",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"7F",X"33",X"4F",X"5F",X"6F",X"77",X"77",X"77",
		X"DD",X"EE",X"EE",X"F0",X"FA",X"FA",X"C3",X"D3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"77",X"7B",X"3F",X"2F",X"2D",X"2E",X"4F",X"DF",
		X"D3",X"C3",X"FF",X"FF",X"FF",X"EF",X"2F",X"CF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"EE",X"F6",X"EE",X"1D",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"00",X"B8",X"B9",X"BB",X"7B",
		X"0F",X"0F",X"07",X"37",X"7B",X"BB",X"BD",X"BD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"7B",X"31",X"4E",X"5F",X"6F",X"67",X"57",X"36",
		X"DD",X"EE",X"EE",X"70",X"7A",X"7A",X"03",X"D3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"75",X"7B",X"35",X"2D",X"2D",X"2E",X"4E",X"DE",
		X"D3",X"C3",X"EF",X"EF",X"EF",X"EF",X"2F",X"CF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DE",X"ED",X"E3",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"EE",X"F6",X"EE",X"1D",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"DC",X"CE",X"E6",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"DE",X"D0",X"78",X"78",X"F9",X"F3",X"E3",X"83",
		X"0F",X"0F",X"07",X"17",X"1B",X"9B",X"9D",X"CD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"81",X"C0",X"D8",X"FC",X"DE",X"4E",X"8E",X"CE",
		X"E5",X"E6",X"F2",X"72",X"38",X"08",X"19",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"EE",X"E8",X"60",X"41",X"4C",X"0C",X"5E",X"DE",
		X"01",X"63",X"E3",X"F3",X"F3",X"F3",X"73",X"27",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"FE",X"FE",X"FD",X"E1",X"E3",X"D9",X"D8",X"D8",
		X"06",X"86",X"C6",X"E6",X"E5",X"F1",X"ED",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8F",X"83",X"66",X"65",X"73",X"53",X"9C",X"92",X"11",X"60",X"E0",X"E2",X"63",X"41",
		X"0F",X"0F",X"07",X"97",X"9B",X"5B",X"59",X"8C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D1",X"C0",X"C0",X"80",X"80",X"80",X"C0",X"C0",X"C0",
		X"C4",X"66",X"3E",X"0E",X"04",X"04",X"05",X"09",X"7F",X"7F",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6C",X"6C",X"2D",X"2D",X"1F",X"1F",X"0F",X"0E",X"E0",X"60",X"40",X"40",X"40",X"00",X"40",X"C0",
		X"09",X"0B",X"13",X"19",X"1C",X"3C",X"3D",X"1B",X"7E",X"7C",X"7C",X"3C",X"18",X"18",X"18",X"58",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DC",X"D8",X"D8",X"E6",X"E1",X"D8",X"D8",X"DF",
		X"16",X"06",X"0E",X"1E",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"57",X"77",X"36",X"37",X"0F",X"0F",X"8F",X"CF",
		X"87",X"CF",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"E6",X"F9",X"FD",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"60",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"DC",X"8D",X"81",X"63",X"63",X"73",X"53",X"5C",X"D2",X"51",X"60",X"E0",X"E0",X"E0",X"C0",
		X"0F",X"CF",X"C5",X"C4",X"E2",X"62",X"71",X"71",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",
		X"35",X"06",X"1E",X"0E",X"04",X"04",X"05",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"6B",X"6B",X"7B",X"1F",X"0F",X"0E",X"F0",X"F0",X"40",X"40",X"40",X"40",X"60",X"E0",
		X"09",X"0B",X"13",X"17",X"17",X"13",X"15",X"09",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"58",
		X"06",X"06",X"08",X"19",X"1E",X"6E",X"EC",X"FC",X"FC",X"F8",X"F8",X"E6",X"81",X"18",X"18",X"D8",
		X"10",X"10",X"10",X"12",X"F5",X"FD",X"7D",X"1B",X"D9",X"DB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7B",X"7B",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"75",X"30",X"38",X"1C",X"09",X"8F",X"CF",
		X"07",X"8F",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EF",X"EF",X"EE",X"F6",X"F6",X"F4",X"B0",X"30",X"10",X"40",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"DC",X"D2",X"51",X"60",X"E0",X"E0",X"E0",X"C0",
		X"0D",X"0C",X"06",X"96",X"9B",X"5B",X"5D",X"4D",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"3F",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",
		X"25",X"16",X"1E",X"0E",X"04",X"04",X"05",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6C",X"29",X"29",X"1D",X"1F",X"0F",X"0E",X"F0",X"F0",X"40",X"40",X"40",X"40",X"60",X"E0",
		X"09",X"0B",X"13",X"17",X"17",X"17",X"17",X"17",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1A",X"1F",X"6D",X"EE",X"F6",X"FC",X"F8",X"F8",X"A6",X"01",X"98",X"D8",X"D8",
		X"16",X"16",X"0F",X"1F",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"B7",X"B4",X"98",X"98",X"98",X"98",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0C",X"8E",X"CE",
		X"07",X"8F",X"FF",X"FF",X"FF",X"7F",X"7F",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"74",X"30",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"DC",X"D2",X"51",X"60",X"E0",X"E0",X"E0",X"C0",
		X"0F",X"0F",X"07",X"97",X"9B",X"5B",X"5D",X"4D",X"DF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",
		X"25",X"16",X"1E",X"0E",X"04",X"04",X"05",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"37",X"37",X"1F",X"1F",X"0F",X"0E",X"F0",X"F0",X"40",X"40",X"40",X"40",X"60",X"E0",
		X"09",X"0B",X"13",X"17",X"17",X"17",X"17",X"17",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"FC",X"F8",X"F8",X"E6",X"E1",X"D8",X"D8",X"98",
		X"16",X"16",X"0E",X"1E",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"C8",X"C8",X"C8",X"C8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"C6",X"77",X"37",X"37",X"0F",X"0F",X"8C",X"CE",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"DC",X"D2",X"51",X"60",X"E0",X"E0",X"E0",X"C0",
		X"0F",X"0F",X"07",X"97",X"9B",X"5B",X"5D",X"4D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"C0",X"E0",
		X"25",X"16",X"1E",X"0E",X"04",X"04",X"05",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"F0",X"F0",X"40",X"40",X"40",X"40",X"60",X"E0",
		X"09",X"0B",X"13",X"17",X"17",X"17",X"17",X"17",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"FC",X"F8",X"F8",X"E6",X"E1",X"D8",X"D8",X"D8",
		X"16",X"16",X"0E",X"1E",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"BD",X"BF",X"7F",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"BD",X"BF",X"7F",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"7F",X"7F",X"7F",X"7F",X"7F",X"77",X"77",X"77",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"BD",X"BF",X"7F",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"7F",X"7F",X"77",X"67",X"63",X"63",X"63",X"63",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"63",X"63",X"33",X"37",X"3F",X"3F",X"5F",X"DF",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"BD",X"BF",X"77",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"67",X"63",X"63",X"63",X"63",X"61",X"61",X"61",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"61",X"71",X"31",X"31",X"31",X"39",X"5B",X"DF",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"DF",X"EF",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"FA",X"FA",X"FA",X"FA",X"EE",X"EE",X"ED",X"ED",X"F6",X"F6",X"F4",X"B0",X"B0",X"D0",X"C0",X"E0",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FD",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"DD",X"8D",X"81",X"63",X"63",X"73",X"53",X"C0",X"C0",X"40",X"18",X"BC",X"A5",X"A7",X"43",
		X"0F",X"0F",X"07",X"37",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5B",X"6B",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"43",X"41",X"41",X"41",X"41",X"41",X"40",X"40",
		X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",X"C3",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",X"7E",
		X"6E",X"6E",X"2F",X"2F",X"1F",X"1F",X"0F",X"0E",X"40",X"40",X"20",X"20",X"20",X"20",X"50",X"D1",
		X"DB",X"C3",X"FF",X"FF",X"FF",X"FF",X"BF",X"DF",X"7E",X"7C",X"7C",X"7C",X"78",X"78",X"78",X"78",
		X"06",X"06",X"0A",X"1B",X"1D",X"6D",X"EE",X"F6",X"D1",X"E9",X"E7",X"E1",X"E0",X"D8",X"D8",X"D8",
		X"EE",X"FE",X"FE",X"FE",X"FD",X"FD",X"7D",X"1B",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"7F",X"7E",X"5C",X"58",X"40",X"40",X"56",X"77",X"37",X"37",X"0F",X"0F",X"8F",X"CF",
		X"07",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E3",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"1A",X"2D",X"16",X"0A",X"05",X"05",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"28",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"1A",X"2D",X"17",X"0B",X"05",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"28",
		X"34",X"98",X"50",X"48",X"24",X"14",X"08",X"00",X"00",X"00",X"80",X"40",X"20",X"90",X"C8",X"64",
		X"04",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"36",X"9D",X"54",X"4A",X"25",X"14",X"0A",X"05",
		X"00",X"00",X"80",X"40",X"20",X"90",X"C8",X"64",X"90",X"40",X"40",X"20",X"90",X"48",X"28",X"10",
		X"00",X"00",X"80",X"40",X"20",X"90",X"48",X"28",X"09",X"04",X"02",X"01",X"01",X"00",X"00",X"00",
		X"9B",X"48",X"44",X"23",X"90",X"48",X"2C",X"1A",X"00",X"00",X"80",X"40",X"20",X"90",X"48",X"2C",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"20",X"90",X"48",X"28",
		X"00",X"80",X"40",X"20",X"90",X"48",X"28",X"10",X"10",X"02",X"05",X"04",X"02",X"01",X"01",X"00",
		X"05",X"84",X"42",X"41",X"20",X"90",X"48",X"28",X"00",X"80",X"40",X"20",X"90",X"48",X"28",X"12",
		X"48",X"24",X"12",X"12",X"0A",X"04",X"00",X"00",X"0A",X"04",X"00",X"80",X"40",X"20",X"20",X"90",
		X"00",X"80",X"40",X"20",X"90",X"48",X"24",X"12",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"24",X"12",X"12",X"0A",X"04",X"01",X"01",X"0A",X"05",X"01",X"81",X"40",X"20",X"20",X"90",
		X"00",X"80",X"40",X"20",X"90",X"48",X"24",X"12",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"10",X"90",X"48",X"24",X"22",X"11",X"09",X"04",X"08",X"04",X"02",X"01",X"00",X"80",X"40",X"20",
		X"80",X"40",X"20",X"10",X"88",X"44",X"22",X"11",X"40",X"40",X"40",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"40",X"80",X"00",X"00",X"00",
		X"08",X"04",X"02",X"02",X"01",X"00",X"00",X"00",X"40",X"40",X"50",X"A8",X"28",X"24",X"22",X"11",
		X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"50",X"AC",X"22",X"21",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"01",X"01",X"00",X"00",X"00",X"00",X"02",X"05",X"04",X"02",X"01",X"00",X"02",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"04",X"02",X"01",X"01",X"00",X"00",X"00",
		X"0B",X"08",X"04",X"03",X"00",X"00",X"04",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"02",X"05",X"04",X"02",X"01",X"01",X"00",X"05",X"04",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"10",X"28",X"28",X"24",X"22",X"11",X"08",X"04",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"2C",X"22",X"21",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"70",X"F8",X"88",X"3E",X"1C",X"1C",X"08",X"08",X"04",X"04",X"02",
		X"23",X"11",X"11",X"08",X"08",X"10",X"10",X"20",X"E2",X"C1",X"C1",X"80",X"80",X"41",X"41",X"22",
		X"04",X"04",X"04",X"04",X"88",X"F8",X"F8",X"F8",X"F9",X"FB",X"F7",X"F4",X"F8",X"F8",X"F8",X"F8",
		X"80",X"80",X"C0",X"40",X"20",X"20",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C4",X"CD",X"8B",X"8F",X"8F",X"8F",X"8F",X"87",X"00",X"80",X"80",X"C0",X"C0",X"F0",X"88",X"04",
		X"40",X"D8",X"B8",X"FC",X"FC",X"FF",X"F8",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"07",X"02",X"02",X"01",X"01",X"00",X"00",X"00",X"04",X"02",X"02",X"04",X"04",X"88",X"70",X"00",
		X"70",X"20",X"20",X"10",X"10",X"08",X"07",X"00",X"40",X"20",X"20",X"40",X"40",X"80",X"00",X"00",
		X"09",X"08",X"08",X"04",X"04",X"04",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"81",X"41",X"26",X"28",X"00",X"00",X"C1",X"6E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"10",X"20",X"20",X"60",X"00",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"06",X"04",X"04",X"08",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"83",X"00",X"00",X"14",X"64",X"82",X"81",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"20",X"20",X"20",X"10",X"10",X"90",
		X"12",X"12",X"11",X"01",X"18",X"08",X"08",X"04",X"06",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"80",X"83",X"6A",X"08",X"00",X"00",X"C2",X"6E",X"00",X"00",X"00",X"00",
		X"00",X"48",X"08",X"80",X"98",X"10",X"30",X"00",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"00",X"0C",X"08",X"19",X"01",X"10",X"12",X"00",
		X"00",X"00",X"00",X"00",X"76",X"43",X"00",X"00",X"10",X"56",X"C1",X"01",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"60",X"20",X"10",X"10",X"18",X"80",X"88",X"48",X"48",
		X"44",X"44",X"60",X"22",X"22",X"31",X"11",X"10",X"08",X"0C",X"04",X"03",X"01",X"00",X"00",X"00",
		X"80",X"40",X"02",X"04",X"00",X"00",X"01",X"41",X"6C",X"08",X"00",X"00",X"C3",X"7E",X"00",X"00",
		X"02",X"22",X"06",X"44",X"C4",X"0C",X"88",X"18",X"10",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"06",X"0C",X"08",X"18",X"11",X"30",X"23",X"22",X"60",X"44",X"40",
		X"00",X"00",X"7E",X"C3",X"00",X"00",X"10",X"36",X"82",X"80",X"00",X"00",X"20",X"40",X"02",X"01",
		X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"08",X"88",X"8C",X"44",X"44",X"06",X"22",X"22",
		X"89",X"89",X"88",X"CC",X"44",X"46",X"62",X"23",X"31",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"81",X"81",X"C3",X"66",X"3C",X"00",X"00",X"81",X"E7",X"3C",X"00",X"00",X"81",X"FF",X"1C",
		X"91",X"91",X"11",X"33",X"22",X"62",X"46",X"C4",X"8C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"31",X"23",X"62",X"46",X"44",X"CC",X"88",X"89",X"89",
		X"1C",X"FF",X"81",X"00",X"00",X"3C",X"E7",X"81",X"00",X"00",X"3C",X"66",X"C3",X"81",X"81",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"8C",X"C4",X"46",X"62",X"22",X"33",X"11",X"91",X"91",
		X"22",X"32",X"13",X"11",X"19",X"08",X"0C",X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"81",X"C3",X"7E",X"18",X"00",X"00",X"C3",X"7E",X"00",X"00",X"00",X"00",
		X"44",X"4C",X"C8",X"88",X"98",X"10",X"30",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"04",X"0C",X"08",X"19",X"11",X"13",X"32",X"22",
		X"00",X"00",X"00",X"00",X"7E",X"C3",X"00",X"00",X"18",X"7E",X"C3",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",X"30",X"10",X"98",X"88",X"C8",X"4C",X"44",
		X"88",X"88",X"88",X"CC",X"44",X"46",X"62",X"23",X"31",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"E7",X"3C",X"00",X"00",X"81",X"FF",X"1C",
		X"11",X"11",X"11",X"33",X"22",X"62",X"46",X"C4",X"8C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"31",X"23",X"62",X"46",X"44",X"CC",X"88",X"88",X"88",
		X"1C",X"FF",X"81",X"00",X"00",X"3C",X"E7",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"8C",X"C4",X"46",X"62",X"22",X"33",X"11",X"11",X"11",
		X"20",X"30",X"10",X"10",X"18",X"08",X"0C",X"04",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"7E",X"00",X"00",X"00",X"00",
		X"04",X"0C",X"08",X"08",X"18",X"10",X"30",X"20",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"06",X"04",X"0C",X"08",X"18",X"10",X"10",X"30",X"20",
		X"00",X"00",X"00",X"00",X"7E",X"C3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"20",X"30",X"10",X"18",X"08",X"08",X"0C",X"04",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"24",X"24",X"22",X"42",X"42",X"41",X"41",X"41",X"41",X"41",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"20",X"20",X"20",X"20",X"10",X"11",X"11",X"09",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"24",X"24",X"22",X"42",X"42",X"41",X"41",X"41",X"41",X"41",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"20",X"20",X"20",X"20",X"10",X"11",X"11",X"09",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"38",X"6C",X"6C",X"66",X"C6",X"C6",X"C3",X"C3",X"C3",X"C3",X"C3",X"C1",X"C1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C1",X"C1",X"61",X"61",X"61",X"61",X"31",X"33",X"33",X"1B",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"78",X"B4",X"B4",X"AA",X"4A",X"4A",X"45",X"45",X"45",X"45",X"45",X"42",X"42",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"42",X"42",X"A2",X"A2",X"A2",X"A2",X"52",X"55",X"55",X"2D",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"D8",X"24",X"24",X"32",X"52",X"52",X"49",X"49",X"49",X"49",X"49",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"02",X"02",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"44",X"24",X"24",X"24",X"24",X"94",X"99",X"99",X"49",X"36",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"03",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"D8",X"64",X"64",X"32",X"72",X"72",X"59",X"59",X"59",X"59",X"59",X"4C",X"4C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"06",X"06",X"03",X"03",X"03",X"03",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4C",X"4C",X"2C",X"2C",X"2C",X"2C",X"9C",X"99",X"99",X"D9",X"76",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"05",X"05",X"05",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",
		X"00",X"00",X"00",X"D8",X"A4",X"A4",X"72",X"52",X"52",X"69",X"69",X"69",X"69",X"69",X"54",X"54",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"0A",X"0A",X"05",X"05",X"05",X"05",X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"54",X"54",X"34",X"34",X"34",X"34",X"94",X"B9",X"B9",X"69",X"F6",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"09",X"09",X"09",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"00",X"00",X"00",X"D8",X"24",X"24",X"B2",X"D2",X"D2",X"49",X"49",X"49",X"49",X"49",X"64",X"64",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"12",X"12",X"09",X"09",X"09",X"09",X"04",X"04",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"64",X"64",X"24",X"24",X"24",X"24",X"B4",X"D9",X"D9",X"49",X"B6",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"0C",X"0C",X"06",X"06",X"06",X"03",X"03",X"03",X"03",X"03",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"03",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"14",X"14",X"0A",X"0A",X"0A",X"05",X"05",X"05",X"05",X"05",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"05",X"05",X"0D",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D8",X"24",X"24",X"12",X"12",X"12",X"09",X"09",X"09",X"09",X"09",X"04",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"09",X"09",X"09",X"36",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D8",X"64",X"64",X"32",X"32",X"32",X"19",X"19",X"19",X"19",X"19",X"0C",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"1C",X"19",X"19",X"19",X"76",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D8",X"A4",X"A4",X"52",X"52",X"52",X"29",X"29",X"29",X"29",X"29",X"14",X"14",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"29",X"29",X"29",X"F6",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"D8",X"24",X"24",X"92",X"92",X"92",X"49",X"49",X"49",X"49",X"49",X"24",X"24",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"49",X"49",X"49",X"B6",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"80",X"80",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"40",
		X"00",X"00",X"00",X"00",X"08",X"06",X"00",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",
		X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"40",X"C0",X"E0",X"F0",X"C0",X"C0",X"80",X"80",X"C0",
		X"00",X"00",X"10",X"08",X"04",X"06",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"2F",X"16",X"08",X"04",
		X"00",X"00",X"00",X"01",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"08",X"0C",X"0C",X"1E",X"1F",X"3F",X"5F",X"5F",X"2F",X"2C",X"10",X"10",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"80",X"80",X"80",X"80",X"C0",X"40",X"20",X"00",X"00",
		X"00",X"00",X"20",X"10",X"08",X"04",X"0C",X"0C",X"1D",X"3F",X"3F",X"3F",X"1F",X"1D",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",
		X"00",X"20",X"10",X"08",X"04",X"0C",X"1C",X"1E",X"1F",X"1E",X"0E",X"0F",X"11",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"08",X"04",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"18",X"18",X"1C",X"1E",X"1E",X"0C",X"16",X"02",X"02",X"02",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"0C",X"0C",X"0C",X"1E",X"1E",X"1D",X"05",X"05",X"05",X"08",X"08",X"00",
		X"00",X"00",X"00",X"40",X"60",X"70",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"01",X"03",X"07",X"03",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"60",X"60",X"C0",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"02",X"04",X"04",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"40",X"20",X"10",X"88",X"44",X"24",X"14",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"20",X"10",X"08",X"C4",X"24",X"14",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"40",X"20",X"10",X"88",X"44",X"24",X"14",X"08",X"00",X"01",X"01",X"01",X"01",X"00",
		X"40",X"20",X"10",X"08",X"C4",X"24",X"14",X"08",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"44",X"42",X"22",X"11",X"08",X"04",X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"20",X"20",X"10",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"30",X"08",X"84",X"42",X"21",X"10",X"08",
		X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"10",X"08",X"84",X"48",X"28",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"06",X"06",X"06",X"06",X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"00",X"40",X"E0",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"09",X"0D",X"0C",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"00",X"40",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"12",X"11",X"18",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"C0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"0C",X"09",X"00",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",
		X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"80",X"B0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"02",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"80",X"E0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"0E",X"06",X"01",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"40",X"C0",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"06",X"00",X"03",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"80",X"80",X"80",
		X"03",X"03",X"03",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"40",X"80",X"80",X"80",
		X"03",X"03",X"01",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",
		X"02",X"04",X"0C",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"80",
		X"07",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0F",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"00",X"02",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"80",X"00",X"00",
		X"01",X"00",X"04",X"02",X"00",X"04",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"04",X"02",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"00",X"80",X"40",X"80",
		X"01",X"02",X"04",X"03",X"00",X"04",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"40",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"05",X"02",X"05",X"02",X"01",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"80",X"40",X"80",X"40",X"80",
		X"05",X"06",X"05",X"03",X"02",X"04",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"40",X"80",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"07",X"07",X"02",X"07",X"07",X"07",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"80",X"C0",X"80",X"C0",X"80",
		X"07",X"07",X"07",X"07",X"02",X"07",X"07",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"80",X"C0",X"80",X"C0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"06",X"06",X"06",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",
		X"06",X"06",X"06",X"06",X"00",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"00",X"FF",X"FF",X"FF",X"C7",X"F8",X"FF",X"FF",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F0",X"E3",X"C0",X"E0",X"C3",X"58",X"00",X"00",
		X"FF",X"FF",X"00",X"04",X"82",X"FB",X"78",X"3F",X"FF",X"FF",X"00",X"00",X"7C",X"0B",X"F7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"FF",X"FF",X"FE",X"E0",X"87",X"00",X"00",X"00",
		X"FF",X"FF",X"0F",X"00",X"E0",X"00",X"12",X"B3",X"FF",X"FF",X"FF",X"FF",X"1F",X"CF",X"77",X"47",
		X"FF",X"F0",X"F0",X"F0",X"E0",X"F8",X"BF",X"FC",X"FC",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"F3",X"0F",X"F0",X"1A",X"03",X"10",X"02",X"00",
		X"F0",X"ED",X"C7",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"80",X"E0",X"61",X"7F",X"3C",X"1D",X"3A",
		X"0D",X"FF",X"80",X"E0",X"40",X"00",X"00",X"80",X"FF",X"F0",X"18",X"0C",X"06",X"02",X"03",X"01",
		X"D2",X"01",X"02",X"01",X"00",X"01",X"01",X"00",X"00",X"88",X"C0",X"C0",X"80",X"C0",X"E0",X"34",
		X"00",X"00",X"03",X"00",X"00",X"07",X"01",X"00",X"0C",X"02",X"80",X"00",X"3F",X"00",X"FF",X"03",
		X"C0",X"E0",X"E2",X"E7",X"F3",X"F3",X"F9",X"FC",X"3E",X"3A",X"F1",X"E0",X"81",X"C2",X"F2",X"07",
		X"80",X"00",X"80",X"00",X"00",X"00",X"C0",X"C0",X"41",X"40",X"E0",X"E1",X"E0",X"03",X"1F",X"FF",
		X"01",X"80",X"87",X"FF",X"98",X"40",X"40",X"80",X"80",X"03",X"1E",X"80",X"40",X"40",X"03",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"01",X"7F",X"22",X"0F",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"91",X"C4",X"E0",X"E6",X"E0",X"E8",X"F0",X"FC",X"C0",X"00",X"17",X"00",X"00",X"38",X"00",X"00",
		X"00",X"03",X"FF",X"00",X"7F",X"00",X"10",X"02",X"3B",X"B3",X"00",X"00",X"80",X"38",X"7F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"BF",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"00",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F1",X"E7",
		X"FF",X"FF",X"FC",X"81",X"3F",X"FF",X"FB",X"FB",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CF",X"D7",X"BE",X"FF",X"68",X"7E",X"70",X"E8",
		X"FF",X"89",X"A8",X"27",X"00",X"2F",X"04",X"00",X"7F",X"FD",X"9F",X"77",X"8B",X"F7",X"17",X"02",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"FF",X"E0",X"83",X"30",X"39",X"1D",X"03",X"0F",
		X"FF",X"00",X"C0",X"FF",X"C9",X"F0",X"A0",X"80",X"FF",X"FF",X"7F",X"DF",X"F7",X"0C",X"03",X"01",
		X"FE",X"FD",X"F9",X"F0",X"E4",X"FF",X"C0",X"C0",X"E4",X"A0",X"A0",X"00",X"20",X"09",X"80",X"00",
		X"01",X"08",X"00",X"00",X"00",X"02",X"00",X"00",X"FF",X"03",X"1F",X"0F",X"1F",X"1F",X"85",X"03",
		X"F8",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"F8",X"38",X"3C",X"0C",X"04",X"2E",X"1D",X"70",X"B3",
		X"A0",X"0F",X"38",X"00",X"1F",X"00",X"62",X"60",X"10",X"98",X"10",X"18",X"98",X"10",X"00",X"01",
		X"E0",X"E0",X"60",X"60",X"40",X"C0",X"C0",X"81",X"28",X"10",X"18",X"44",X"78",X"20",X"90",X"28",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"08",X"3F",X"01",X"0F",X"0F",X"1B",X"1F",X"03",X"2F",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"55",X"07",X"41",X"F0",X"FE",X"FE",X"FF",X"FF",
		X"A0",X"C0",X"CF",X"10",X"02",X"1F",X"FF",X"FF",X"07",X"3B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F6",X"E0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FF",X"73",X"90",X"E8",X"76",X"FE",X"7F",X"7F",X"7A",
		X"03",X"00",X"82",X"04",X"A2",X"FF",X"6D",X"EF",X"5F",X"BF",X"FF",X"7F",X"BF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"BF",X"9F",X"DF",X"CF",X"E7",X"F3",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"E6",X"EE",X"C8",X"95",X"EA",X"94",X"9A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"03",X"F0",X"FF",X"FF",X"FF",X"FF",X"C4",X"A4",X"E5",X"79",X"2F",X"C1",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"80",X"11",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"60",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"E1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"F0",X"E2",X"C0",X"C0",X"C0",X"E0",X"F0",X"E0",X"80",X"1F",X"0E",X"0F",X"1D",X"E6",X"73",X"18",
		X"77",X"FC",X"01",X"00",X"06",X"79",X"E8",X"9B",X"FF",X"7E",X"9F",X"45",X"3B",X"25",X"91",X"33",
		X"7F",X"FF",X"FF",X"FF",X"DF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"FE",X"FF",X"0F",X"0E",X"03",X"23",X"07",X"00",X"00",X"C3",
		X"F6",X"00",X"83",X"9F",X"F7",X"0F",X"7F",X"FF",X"63",X"C7",X"FF",X"CF",X"F7",X"FF",X"FB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"EB",X"FF",X"FF",X"FF",X"FF",X"98",X"CC",X"08",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FD",X"FB",X"FF",X"F7",X"EF",X"EF",X"01",X"0E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"3F",X"02",X"E0",X"FC",X"1E",X"83",X"E0",X"0F",X"E1",X"DE",X"67",X"FB",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"FB",X"FE",X"FF",X"FF",X"FF",X"C1",X"00",X"FF",X"87",X"3F",X"F3",
		X"FF",X"FF",X"FF",X"07",X"FB",X"5D",X"ED",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BE",X"2D",
		X"DF",X"BF",X"FF",X"FF",X"FF",X"FF",X"2F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"E0",X"F8",X"FC",X"FF",X"FF",X"FF",X"E0",
		X"F7",X"CF",X"9E",X"BE",X"FE",X"DE",X"FE",X"FF",X"C7",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"88",X"80",X"80",X"1A",X"04",X"00",X"08",X"00",X"0C",X"04",X"82",X"02",X"48",X"40",X"00",X"80",
		X"FF",X"7F",X"39",X"16",X"8F",X"1F",X"0F",X"75",X"FF",X"FC",X"83",X"7F",X"FF",X"FF",X"1F",X"FC",
		X"F8",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"0E",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"07",
		X"DE",X"CF",X"E7",X"F7",X"FB",X"FC",X"FE",X"FF",X"82",X"42",X"A3",X"F1",X"FD",X"FF",X"00",X"E3",
		X"88",X"80",X"40",X"01",X"F1",X"C7",X"1F",X"FF",X"08",X"98",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F2",X"E2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"E8",X"E7",X"FE",X"FE",X"FF",X"88",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"DE",X"FF",X"FE",X"DF",X"FF",X"FF",X"07",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FF",X"FF",X"FE",
		X"E7",X"FF",X"49",X"1F",X"FF",X"F8",X"80",X"1F",X"BF",X"FF",X"FF",X"FF",X"FE",X"0F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"E7",X"DF",X"3F",X"46",X"FE",X"7B",X"8F",X"FF",
		X"1F",X"FE",X"FF",X"CF",X"DC",X"F8",X"D8",X"D0",X"E3",X"3C",X"CB",X"FC",X"07",X"00",X"00",X"00",
		X"FF",X"FF",X"1F",X"C3",X"FF",X"F8",X"60",X"30",X"FF",X"FF",X"4F",X"F6",X"FF",X"1A",X"03",X"00",
		X"E0",X"98",X"E0",X"FF",X"87",X"40",X"01",X"47",X"FF",X"E7",X"07",X"03",X"C8",X"E0",X"F9",X"1F",
		X"F9",X"FA",X"FF",X"F7",X"FF",X"FF",X"FF",X"FB",X"F8",X"F8",X"EC",X"F2",X"F0",X"E0",X"F1",X"F1",
		X"C0",X"47",X"08",X"00",X"05",X"80",X"B0",X"B0",X"08",X"88",X"00",X"10",X"00",X"08",X"00",X"00",
		X"38",X"18",X"08",X"08",X"08",X"08",X"10",X"70",X"02",X"09",X"00",X"01",X"03",X"14",X"07",X"03",
		X"A2",X"B6",X"F8",X"88",X"61",X"C3",X"E0",X"C0",X"E7",X"7E",X"00",X"06",X"F0",X"F0",X"3C",X"0F",
		X"FB",X"FF",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"E9",X"F6",X"F9",X"FF",X"3F",X"80",X"FC",X"FF",
		X"90",X"F0",X"F8",X"FF",X"FF",X"7F",X"00",X"C9",X"00",X"01",X"07",X"F8",X"F9",X"47",X"1F",X"FF",
		X"E0",X"C0",X"E7",X"0F",X"FF",X"FF",X"FF",X"FF",X"0B",X"1F",X"EE",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"00",X"0D",X"FE",X"FF",X"80",X"F8",X"7C",X"97",X"23",X"FD",X"01",X"FB",X"0F",X"61",X"00",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F9",X"FF",X"FC",X"FE",X"FE",X"FF",
		X"FF",X"7F",X"00",X"87",X"3F",X"FC",X"F0",X"00",X"FF",X"FF",X"1F",X"8F",X"FF",X"7F",X"1F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"FE",X"03",X"87",X"F8",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"7F",X"78",X"FF",X"FF",X"F3",X"D3",X"67",X"FF",X"FF",X"2D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"83",X"F3",X"DA",X"8E",X"73",X"81",X"FF",
		X"47",X"87",X"EC",X"7F",X"39",X"8F",X"FE",X"FF",X"F8",X"7F",X"E7",X"BD",X"FF",X"3F",X"3F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F9",X"F2",X"FF",X"FF",X"FF",X"80",X"1F",X"60",X"83",X"7F",
		X"FF",X"FF",X"FF",X"17",X"00",X"FF",X"F7",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"06",
		X"FF",X"FD",X"FC",X"FF",X"FE",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"00",X"F7",X"FC",X"A4",
		X"FF",X"F1",X"80",X"FF",X"00",X"C0",X"73",X"73",X"E7",X"40",X"3F",X"C0",X"40",X"27",X"B8",X"C8",
		X"E8",X"CB",X"D4",X"D2",X"C5",X"C0",X"E3",X"F9",X"BF",X"BE",X"76",X"EC",X"50",X"70",X"E0",X"C2",
		X"D0",X"90",X"40",X"07",X"08",X"00",X"4F",X"C0",X"03",X"11",X"B8",X"DC",X"00",X"00",X"90",X"18",
		X"DF",X"C3",X"61",X"30",X"20",X"20",X"20",X"70",X"F2",X"81",X"FF",X"7F",X"7F",X"02",X"70",X"80",
		X"8C",X"20",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"19",X"17",X"FE",X"FF",X"7F",X"82",X"00",X"00",
		X"F8",X"F7",X"E5",X"FF",X"C9",X"FC",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"E0",X"00",X"0F",X"FF",
		X"30",X"B0",X"F0",X"F7",X"8B",X"19",X"FF",X"FF",X"00",X"07",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C1",X"87",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"F4",X"FC",X"12",X"90",X"C8",X"FF",X"FF",
		X"9E",X"71",X"71",X"CC",X"00",X"20",X"FF",X"FF",X"69",X"C7",X"45",X"A8",X"02",X"0F",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"EF",X"08",X"80",X"BB",X"EE",X"C2",X"B0",
		X"03",X"E0",X"FF",X"00",X"0B",X"38",X"28",X"40",X"00",X"1F",X"C0",X"00",X"3C",X"E3",X"27",X"1C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"B7",X"FF",X"F1",X"F6",X"FF",X"FF",X"FF",
		X"90",X"FF",X"FF",X"80",X"7F",X"9F",X"FF",X"FF",X"0B",X"FD",X"1F",X"FD",X"C7",X"FF",X"FB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F3",X"E0",X"F8",X"FF",X"FF",X"FF",X"1F",X"FF",X"7F",X"0F",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F9",X"FA",X"FF",X"FF",X"FC",X"E1",X"1F",X"7C",X"E7",X"3F",
		X"FF",X"FF",X"03",X"F9",X"7E",X"FC",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"7F",X"0E",X"C7",X"7F",
		X"C0",X"80",X"86",X"00",X"00",X"00",X"80",X"E0",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"07",X"03",X"06",X"82",X"03",X"14",
		X"F7",X"F3",X"FC",X"FF",X"FB",X"FF",X"FF",X"FF",X"F6",X"FA",X"86",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"9E",X"F2",X"E0",X"FA",X"1C",X"00",X"3C",X"46",X"73",X"1E",X"1E",X"22",X"03",X"0C",
		X"30",X"18",X"10",X"08",X"8C",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"FC",X"07",X"00",X"00",X"06",X"7F",
		X"FF",X"FB",X"FD",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"8F",X"E0",X"FF",
		X"C4",X"F8",X"FB",X"F8",X"F3",X"8F",X"1F",X"FF",X"3C",X"7F",X"BD",X"7F",X"FE",X"FF",X"FF",X"FF",
		X"00",X"C0",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"1F",X"03",X"03",X"02",X"02",X"02",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"E8",X"F4",X"FF",X"FC",X"FF",X"FF",X"03",X"01",X"13",X"08",X"00",X"90",X"7F",X"FF",
		X"F0",X"FF",X"7F",X"7F",X"FF",X"FB",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"70",X"00",X"F0",X"EE",X"18",X"34",X"30",X"29",X"24",X"50",
		X"F8",X"00",X"00",X"07",X"70",X"80",X"00",X"00",X"3F",X"1E",X"7C",X"A0",X"00",X"00",X"83",X"06",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"C0",X"00",X"50",X"90",X"A8",X"AF",X"FD",
		X"00",X"01",X"06",X"09",X"14",X"E0",X"80",X"F0",X"84",X"00",X"80",X"00",X"00",X"02",X"0C",X"03",
		X"00",X"0C",X"00",X"00",X"00",X"10",X"00",X"50",X"8B",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FC",X"F0",X"C0",X"80",X"00",X"00",X"80",
		X"FF",X"00",X"1C",X"02",X"01",X"00",X"00",X"00",X"FF",X"1B",X"9F",X"87",X"23",X"BC",X"3F",X"70",
		X"00",X"00",X"02",X"00",X"FF",X"7F",X"EF",X"7F",X"04",X"01",X"A0",X"00",X"00",X"C0",X"C0",X"E0",
		X"80",X"00",X"00",X"02",X"09",X"18",X"08",X"00",X"00",X"00",X"00",X"01",X"81",X"BC",X"2C",X"04",
		X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F8",X"F8",X"00",X"20",X"10",X"00",X"01",X"01",X"01",X"00",
		X"0E",X"0E",X"31",X"09",X"AA",X"23",X"04",X"03",X"00",X"00",X"00",X"80",X"08",X"08",X"80",X"80",
		X"1F",X"0D",X"07",X"03",X"03",X"87",X"86",X"CE",X"E0",X"60",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"08",X"00",X"03",X"0D",X"05",X"00",X"00",X"00",X"03",X"4F",X"C3",X"00",X"44",X"B7",X"FF",X"E0",
		X"F0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"C2",
		X"06",X"0B",X"0A",X"13",X"FF",X"76",X"FF",X"C0",X"02",X"23",X"E3",X"FC",X"C7",X"EC",X"71",X"D7",
		X"DC",X"FA",X"60",X"F0",X"70",X"F0",X"F8",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"C0",X"F8",X"FC",X"FC",X"FF",
		X"00",X"00",X"00",X"14",X"00",X"06",X"00",X"80",X"00",X"00",X"00",X"0C",X"03",X"1C",X"20",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
