library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity eprom_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of eprom_2 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"15",X"FF",X"1A",X"1A",X"1A",X"00",X"00",X"00",X"1A",X"1A",X"1A",X"FF",X"15",X"00",X"15",X"FF",
		X"1A",X"1A",X"1A",X"00",X"1A",X"1A",X"1A",X"FF",X"15",X"00",X"00",X"00",X"15",X"FF",X"1A",X"1A",
		X"19",X"1A",X"1A",X"FF",X"15",X"00",X"00",X"00",X"00",X"00",X"16",X"FF",X"1A",X"19",X"1A",X"FF",
		X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"FF",X"19",X"FF",X"15",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"1A",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"CD",X"17",X"21",X"CD",X"D0",X"21",X"21",X"7D",X"C4",X"11",X"7E",X"C4",X"01",X"40",
		X"00",X"36",X"00",X"ED",X"B0",X"3E",X"00",X"32",X"D5",X"C4",X"3A",X"11",X"EC",X"A7",X"20",X"10",
		X"2A",X"88",X"ED",X"E5",X"D1",X"13",X"01",X"EA",X"00",X"3E",X"01",X"77",X"ED",X"B0",X"18",X"0F",
		X"21",X"12",X"EC",X"ED",X"5B",X"88",X"ED",X"06",X"EA",X"7E",X"12",X"23",X"13",X"10",X"FA",X"E7",
		X"FD",X"21",X"0A",X"EC",X"FD",X"36",X"00",X"00",X"06",X"EA",X"AF",X"F5",X"C5",X"CD",X"40",X"84",
		X"C1",X"F1",X"3C",X"10",X"F6",X"21",X"02",X"E6",X"11",X"4D",X"86",X"AF",X"CD",X"F1",X"21",X"21",
		X"2A",X"E7",X"11",X"61",X"86",X"AF",X"CD",X"F1",X"21",X"21",X"2E",X"E7",X"11",X"79",X"86",X"AF",
		X"CD",X"F1",X"21",X"21",X"32",X"E7",X"11",X"8F",X"86",X"AF",X"CD",X"F1",X"21",X"21",X"36",X"E7",
		X"11",X"A5",X"86",X"AF",X"CD",X"F1",X"21",X"21",X"3A",X"E7",X"11",X"C0",X"86",X"AF",X"CD",X"F1",
		X"21",X"21",X"3E",X"E7",X"11",X"D6",X"86",X"AF",X"CD",X"F1",X"21",X"3A",X"7B",X"C4",X"CB",X"97",
		X"32",X"08",X"D0",X"3A",X"7C",X"C4",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"07",
		X"EC",X"3E",X"00",X"32",X"09",X"EC",X"32",X"0D",X"EC",X"3E",X"01",X"32",X"0C",X"EC",X"E7",X"3A",
		X"0C",X"D0",X"CB",X"57",X"20",X"1A",X"CD",X"17",X"21",X"21",X"12",X"EC",X"ED",X"5B",X"88",X"ED",
		X"06",X"EA",X"1A",X"77",X"13",X"23",X"10",X"FA",X"3E",X"FF",X"32",X"11",X"EC",X"3E",X"00",X"D7",
		X"CD",X"ED",X"82",X"3A",X"07",X"EC",X"47",X"4F",X"3A",X"7C",X"C4",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"B8",X"CA",X"0C",X"82",X"32",X"07",X"EC",X"30",X"48",X"F5",X"C5",X"CD",X"78",
		X"83",X"C1",X"F1",X"90",X"2F",X"3C",X"E6",X"0F",X"CB",X"5F",X"20",X"30",X"47",X"3A",X"09",X"EC",
		X"3D",X"FE",X"FF",X"20",X"02",X"3E",X"EA",X"32",X"09",X"EC",X"C5",X"CD",X"3F",X"83",X"C1",X"3E",
		X"01",X"DF",X"3A",X"09",X"EC",X"FE",X"EA",X"28",X"07",X"C5",X"CD",X"40",X"84",X"C1",X"18",X"05",
		X"C5",X"CD",X"A9",X"83",X"C1",X"10",X"D9",X"CD",X"BE",X"83",X"18",X"50",X"3A",X"07",X"EC",X"91",
		X"E6",X"0F",X"18",X"0E",X"F5",X"C5",X"CD",X"78",X"83",X"C1",X"F1",X"90",X"E6",X"0F",X"CB",X"5F",
		X"20",X"30",X"47",X"3A",X"09",X"EC",X"3C",X"FE",X"EB",X"20",X"02",X"3E",X"00",X"32",X"09",X"EC",
		X"C5",X"CD",X"3F",X"83",X"C1",X"3E",X"01",X"DF",X"3A",X"09",X"EC",X"FE",X"EA",X"28",X"07",X"C5",
		X"CD",X"40",X"84",X"C1",X"18",X"05",X"C5",X"CD",X"A9",X"83",X"C1",X"10",X"D6",X"CD",X"BE",X"83",
		X"18",X"0A",X"3A",X"07",X"EC",X"91",X"2F",X"3C",X"E6",X"0F",X"18",X"80",X"3A",X"0C",X"D0",X"CB",
		X"47",X"20",X"3C",X"3A",X"0D",X"EC",X"CB",X"47",X"20",X"3D",X"CB",X"C7",X"32",X"0D",X"EC",X"3A",
		X"09",X"EC",X"FE",X"EA",X"28",X"17",X"3A",X"0C",X"EC",X"3C",X"32",X"0C",X"EC",X"FE",X"14",X"20",
		X"05",X"3E",X"00",X"32",X"0C",X"EC",X"21",X"24",X"86",X"CD",X"A8",X"3D",X"E9",X"3A",X"72",X"ED",
		X"3C",X"FE",X"21",X"20",X"02",X"3E",X"00",X"32",X"72",X"ED",X"CD",X"A9",X"83",X"18",X"08",X"3A",
		X"0D",X"EC",X"E6",X"FE",X"32",X"0D",X"EC",X"3A",X"0C",X"D0",X"CB",X"4F",X"20",X"3C",X"3A",X"0D",
		X"EC",X"CB",X"4F",X"20",X"3D",X"CB",X"CF",X"32",X"0D",X"EC",X"3A",X"09",X"EC",X"FE",X"EA",X"28",
		X"17",X"3A",X"0C",X"EC",X"3D",X"32",X"0C",X"EC",X"FE",X"FF",X"20",X"05",X"3E",X"13",X"32",X"0C",
		X"EC",X"21",X"24",X"86",X"CD",X"A8",X"3D",X"E9",X"3A",X"72",X"ED",X"3D",X"FE",X"FF",X"20",X"02",
		X"3E",X"20",X"32",X"72",X"ED",X"CD",X"A9",X"83",X"18",X"08",X"3A",X"0D",X"EC",X"E6",X"FD",X"32",
		X"0D",X"EC",X"3A",X"10",X"D0",X"CB",X"47",X"C2",X"E2",X"82",X"3A",X"0D",X"EC",X"CB",X"57",X"C2",
		X"3E",X"81",X"CB",X"D7",X"32",X"0D",X"EC",X"CD",X"78",X"83",X"CD",X"D2",X"84",X"46",X"3A",X"09",
		X"EC",X"3C",X"FE",X"EA",X"28",X"16",X"FE",X"EB",X"20",X"02",X"3E",X"00",X"F5",X"C5",X"CD",X"BE",
		X"83",X"C1",X"F1",X"F5",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"70",X"F1",X"32",X"09",X"EC",X"C3",
		X"3E",X"81",X"3A",X"0D",X"EC",X"E6",X"FB",X"32",X"0D",X"EC",X"C3",X"3E",X"81",X"3A",X"08",X"EC",
		X"3C",X"32",X"08",X"EC",X"E6",X"0F",X"C0",X"3A",X"08",X"EC",X"CB",X"7F",X"28",X"41",X"AF",X"32",
		X"08",X"EC",X"3A",X"09",X"EC",X"FE",X"EA",X"CA",X"A9",X"83",X"FD",X"21",X"0A",X"EC",X"3A",X"09",
		X"EC",X"CD",X"40",X"84",X"CD",X"BE",X"83",X"C9",X"11",X"10",X"86",X"21",X"F0",X"0A",X"CD",X"D1",
		X"20",X"1A",X"85",X"6F",X"30",X"01",X"24",X"13",X"1A",X"B4",X"67",X"EB",X"3A",X"09",X"EC",X"D5",
		X"CD",X"CA",X"5A",X"D1",X"72",X"23",X"73",X"13",X"CD",X"03",X"21",X"72",X"23",X"73",X"C9",X"AF",
		X"CB",X"FF",X"32",X"08",X"EC",X"3A",X"09",X"EC",X"FE",X"EA",X"28",X"22",X"CD",X"D2",X"84",X"7E",
		X"A7",X"20",X"05",X"CD",X"18",X"83",X"18",X"0C",X"3A",X"09",X"EC",X"CD",X"CA",X"5A",X"11",X"4C",
		X"86",X"CD",X"1C",X"22",X"11",X"E8",X"86",X"21",X"7A",X"E3",X"CD",X"1C",X"22",X"C9",X"21",X"7E",
		X"E3",X"11",X"4C",X"86",X"CD",X"1C",X"22",X"C9",X"3A",X"09",X"EC",X"FE",X"EA",X"28",X"2A",X"2A",
		X"88",X"ED",X"CD",X"50",X"20",X"7E",X"A7",X"28",X"0F",X"FD",X"21",X"0A",X"EC",X"3A",X"09",X"EC",
		X"CD",X"40",X"84",X"AF",X"32",X"08",X"EC",X"C9",X"3A",X"09",X"EC",X"CD",X"CA",X"5A",X"11",X"4C",
		X"86",X"CD",X"1C",X"22",X"AF",X"32",X"08",X"EC",X"C9",X"3A",X"72",X"ED",X"3C",X"11",X"0E",X"EC",
		X"CD",X"A2",X"84",X"21",X"7E",X"E3",X"11",X"0E",X"EC",X"AF",X"CD",X"F1",X"21",X"C9",X"CD",X"D2",
		X"84",X"7E",X"E6",X"E3",X"21",X"2E",X"84",X"11",X"34",X"84",X"BE",X"28",X"05",X"23",X"13",X"13",
		X"18",X"F8",X"EB",X"5E",X"23",X"56",X"EB",X"E9",X"11",X"E8",X"86",X"CD",X"DC",X"84",X"AF",X"32",
		X"0C",X"EC",X"C9",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"CD",X"D2",X"84",X"7E",X"CB",X"3F",X"CB",
		X"3F",X"3C",X"32",X"0C",X"EC",X"C9",X"11",X"FA",X"86",X"CD",X"DC",X"84",X"CD",X"D2",X"84",X"7E",
		X"CB",X"3F",X"CB",X"3F",X"C6",X"09",X"32",X"0C",X"EC",X"C9",X"11",X"0C",X"87",X"CD",X"DC",X"84",
		X"3E",X"12",X"32",X"0C",X"EC",X"C9",X"11",X"03",X"87",X"CD",X"DC",X"84",X"3E",X"11",X"32",X"0C",
		X"EC",X"C9",X"11",X"15",X"87",X"CD",X"DC",X"84",X"3E",X"13",X"32",X"0C",X"EC",X"C9",X"00",X"01",
		X"02",X"03",X"E3",X"E2",X"D8",X"83",X"E3",X"83",X"F6",X"83",X"0A",X"84",X"16",X"84",X"22",X"84",
		X"F5",X"ED",X"5B",X"88",X"ED",X"CD",X"4A",X"20",X"1A",X"A7",X"28",X"4B",X"FE",X"FF",X"28",X"03",
		X"FD",X"34",X"00",X"E6",X"03",X"28",X"3E",X"FE",X"03",X"20",X"0D",X"1A",X"11",X"20",X"86",X"FE",
		X"FF",X"20",X"10",X"11",X"22",X"86",X"18",X"0B",X"1A",X"CB",X"3F",X"E6",X"0E",X"11",X"10",X"86",
		X"CD",X"4A",X"20",X"21",X"F0",X"0A",X"CD",X"D1",X"20",X"1A",X"85",X"6F",X"30",X"01",X"24",X"13",
		X"1A",X"B4",X"67",X"EB",X"F1",X"F5",X"D5",X"CD",X"CA",X"5A",X"D1",X"72",X"23",X"73",X"13",X"CD",
		X"03",X"21",X"72",X"23",X"73",X"F1",X"C9",X"F1",X"CD",X"CA",X"5A",X"11",X"4C",X"86",X"CD",X"1C",
		X"22",X"C9",X"06",X"00",X"FE",X"0A",X"38",X"05",X"04",X"D6",X"0A",X"18",X"F7",X"CB",X"20",X"CB",
		X"20",X"CB",X"20",X"CB",X"20",X"80",X"F5",X"3E",X"02",X"12",X"F1",X"F5",X"E6",X"F0",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"30",X"13",X"12",X"F1",X"E6",X"0F",X"C6",X"30",X"13",
		X"12",X"C9",X"3A",X"09",X"EC",X"2A",X"88",X"ED",X"CD",X"50",X"20",X"C9",X"21",X"7A",X"E3",X"AF",
		X"CD",X"F1",X"21",X"C9",X"CD",X"D2",X"84",X"3E",X"00",X"77",X"11",X"E8",X"86",X"CD",X"DC",X"84",
		X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"01",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",
		X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"05",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",
		X"82",X"CD",X"D2",X"84",X"3E",X"09",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",
		X"CD",X"D2",X"84",X"3E",X"0D",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",
		X"D2",X"84",X"3E",X"11",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",
		X"84",X"3E",X"15",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",
		X"3E",X"19",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",
		X"1D",X"77",X"11",X"F1",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"02",
		X"77",X"11",X"FA",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"06",X"77",
		X"11",X"FA",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"0A",X"77",X"11",
		X"FA",X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"0E",X"77",X"11",X"FA",
		X"86",X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"12",X"77",X"11",X"FA",X"86",
		X"CD",X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"16",X"77",X"11",X"FA",X"86",X"CD",
		X"DC",X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"1A",X"77",X"11",X"FA",X"86",X"CD",X"DC",
		X"84",X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"1E",X"77",X"11",X"FA",X"86",X"CD",X"DC",X"84",
		X"C3",X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"FF",X"77",X"11",X"03",X"87",X"CD",X"DC",X"84",X"C3",
		X"A2",X"82",X"CD",X"D2",X"84",X"3E",X"03",X"77",X"11",X"0C",X"87",X"CD",X"DC",X"84",X"C3",X"A2",
		X"82",X"CD",X"D2",X"84",X"3E",X"E2",X"77",X"11",X"15",X"87",X"CD",X"DC",X"84",X"C3",X"A2",X"82",
		X"00",X"C0",X"02",X"C0",X"04",X"C0",X"06",X"C0",X"08",X"C0",X"0A",X"C0",X"0C",X"C8",X"0E",X"C8",
		X"10",X"C8",X"10",X"D8",X"E4",X"84",X"F3",X"84",X"02",X"85",X"11",X"85",X"20",X"85",X"2F",X"85",
		X"3E",X"85",X"4D",X"85",X"5C",X"85",X"6B",X"85",X"7A",X"85",X"89",X"85",X"98",X"85",X"A7",X"85",
		X"B6",X"85",X"C5",X"85",X"D4",X"85",X"E3",X"85",X"F2",X"85",X"01",X"86",X"02",X"13",X"43",X"41",
		X"4E",X"20",X"59",X"4F",X"55",X"20",X"44",X"4F",X"20",X"42",X"45",X"54",X"54",X"45",X"52",X"20",
		X"3F",X"17",X"43",X"4F",X"4E",X"54",X"52",X"4F",X"4C",X"4C",X"45",X"52",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"50",X"4F",X"53",X"49",X"54",X"49",X"4F",X"4E",X"15",X"31",X"50",X"2D",X"32",X"50",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"2E",X"2E",X"2E",X"43",X"48",X"4F",X"49",X"43",X"45",X"15",
		X"53",X"48",X"4F",X"54",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"2E",X"2E",X"2E",X"2E",X"52",
		X"45",X"47",X"49",X"53",X"54",X"1A",X"53",X"45",X"52",X"56",X"49",X"43",X"45",X"20",X"53",X"57",
		X"2E",X"2E",X"2E",X"2E",X"2E",X"45",X"4E",X"44",X"20",X"4F",X"46",X"20",X"45",X"44",X"49",X"54",
		X"15",X"42",X"4C",X"4F",X"43",X"4B",X"20",X"4B",X"49",X"4E",X"44",X"2E",X"2E",X"2E",X"2E",X"2E",
		X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"11",X"52",X"4F",X"55",X"4E",X"44",X"2E",X"2E",X"2E",X"2E",
		X"2E",X"2E",X"2E",X"2E",X"2E",X"2E",X"30",X"31",X"08",X"42",X"4C",X"41",X"4E",X"4B",X"20",X"20",
		X"20",X"08",X"4E",X"4F",X"52",X"4D",X"41",X"4C",X"20",X"20",X"08",X"49",X"54",X"45",X"4D",X"20",
		X"20",X"20",X"20",X"08",X"49",X"4D",X"4F",X"54",X"41",X"52",X"54",X"59",X"08",X"48",X"41",X"52",
		X"44",X"20",X"20",X"20",X"20",X"08",X"4B",X"45",X"59",X"20",X"20",X"20",X"20",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1D",X"1D",X"1D",X"1D",X"1D",X"FF",X"00",X"FF",X"1D",X"1D",X"1D",X"1D",X"1D",X"19",
		X"19",X"19",X"19",X"19",X"FF",X"00",X"FF",X"19",X"19",X"19",X"19",X"19",X"FF",X"FF",X"02",X"FF",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"02",X"FF",X"FF",X"15",X"15",X"15",X"15",X"15",X"FF",X"00",
		X"FF",X"15",X"15",X"15",X"15",X"15",X"11",X"11",X"11",X"11",X"11",X"FF",X"00",X"FF",X"11",X"11",
		X"11",X"11",X"11",X"0D",X"0D",X"0D",X"0D",X"0D",X"FF",X"00",X"FF",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"03",X"03",X"02",X"03",X"03",X"FF",X"00",X"FF",X"03",X"03",X"02",X"03",X"03",X"09",X"09",X"09",
		X"09",X"09",X"FF",X"00",X"FF",X"09",X"09",X"09",X"09",X"09",X"05",X"05",X"05",X"05",X"05",X"FF",
		X"00",X"FF",X"05",X"05",X"05",X"05",X"05",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"FF",X"01",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"89",X"3E",X"06",X"CF",X"3E",X"0C",X"CD",X"AE",
		X"67",X"3A",X"7B",X"C4",X"CB",X"F7",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"2A",X"88",X"ED",X"E5",
		X"D1",X"13",X"01",X"EA",X"00",X"36",X"00",X"ED",X"B0",X"3E",X"FF",X"32",X"83",X"ED",X"AF",X"32",
		X"FE",X"EC",X"21",X"91",X"8E",X"06",X"00",X"3A",X"FE",X"EC",X"CB",X"27",X"CB",X"27",X"4F",X"09",
		X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"C5",X"E1",X"CD",X"D1",X"20",X"3E",X"88",X"06",X"04",
		X"0E",X"04",X"CD",X"55",X"22",X"3A",X"FE",X"EC",X"3C",X"32",X"FE",X"EC",X"FE",X"24",X"20",X"D2",
		X"11",X"C6",X"E0",X"06",X"07",X"21",X"10",X"1E",X"CD",X"D1",X"20",X"C5",X"06",X"00",X"0E",X"0C",
		X"09",X"06",X"04",X"0E",X"01",X"3E",X"88",X"CD",X"55",X"22",X"01",X"38",X"00",X"ED",X"42",X"EB",
		X"C1",X"10",X"E2",X"11",X"06",X"E7",X"06",X"07",X"21",X"10",X"1E",X"CD",X"D1",X"20",X"C5",X"06",
		X"04",X"0E",X"01",X"3E",X"88",X"CD",X"55",X"22",X"01",X"38",X"00",X"ED",X"42",X"EB",X"C1",X"10",
		X"E7",X"AF",X"32",X"FF",X"EC",X"11",X"FE",X"E0",X"06",X"1A",X"21",X"10",X"1E",X"CD",X"D1",X"20",
		X"C5",X"D5",X"11",X"21",X"8F",X"3A",X"FF",X"EC",X"83",X"30",X"01",X"14",X"5F",X"1A",X"4F",X"06",
		X"00",X"09",X"06",X"01",X"0E",X"01",X"3E",X"88",X"D1",X"CD",X"55",X"22",X"EB",X"3A",X"FF",X"EC",
		X"3C",X"FE",X"04",X"20",X"01",X"AF",X"32",X"FF",X"EC",X"C1",X"10",X"CE",X"CD",X"70",X"22",X"21",
		X"D0",X"2B",X"3E",X"80",X"CD",X"58",X"8B",X"21",X"0B",X"ED",X"11",X"0C",X"ED",X"01",X"5A",X"00",
		X"36",X"00",X"ED",X"B0",X"21",X"0B",X"ED",X"11",X"0B",X"00",X"19",X"11",X"0D",X"00",X"AF",X"06",
		X"07",X"77",X"3C",X"19",X"10",X"FB",X"3E",X"00",X"32",X"05",X"ED",X"32",X"07",X"ED",X"32",X"04",
		X"ED",X"32",X"6B",X"ED",X"3E",X"02",X"32",X"00",X"ED",X"3E",X"FF",X"32",X"01",X"ED",X"3E",X"80",
		X"32",X"06",X"ED",X"3E",X"FF",X"32",X"FD",X"EC",X"2A",X"44",X"C4",X"22",X"69",X"ED",X"E7",X"3A",
		X"FD",X"EC",X"A7",X"CA",X"3A",X"8A",X"CD",X"54",X"8D",X"CD",X"99",X"8D",X"CD",X"0A",X"8C",X"3A",
		X"05",X"ED",X"CB",X"6F",X"C4",X"BB",X"8B",X"CB",X"67",X"C4",X"D3",X"8B",X"CB",X"7F",X"20",X"2F",
		X"3A",X"00",X"ED",X"3D",X"32",X"00",X"ED",X"A7",X"20",X"CE",X"3E",X"FF",X"32",X"66",X"ED",X"32",
		X"67",X"ED",X"3A",X"05",X"ED",X"CB",X"FF",X"32",X"05",X"ED",X"3E",X"01",X"32",X"02",X"ED",X"3E",
		X"05",X"32",X"03",X"ED",X"21",X"D0",X"2E",X"3A",X"06",X"ED",X"CD",X"58",X"8B",X"18",X"A9",X"3A",
		X"66",X"ED",X"FE",X"FF",X"C2",X"E6",X"89",X"3A",X"03",X"ED",X"3D",X"32",X"03",X"ED",X"A7",X"20",
		X"97",X"3A",X"02",X"ED",X"3C",X"FE",X"06",X"28",X"76",X"32",X"02",X"ED",X"3A",X"04",X"ED",X"A7",
		X"20",X"03",X"CD",X"45",X"8B",X"3A",X"02",X"ED",X"FE",X"03",X"28",X"08",X"3E",X"05",X"32",X"03",
		X"ED",X"C3",X"28",X"89",X"3A",X"01",X"ED",X"FE",X"C0",X"38",X"1E",X"E6",X"38",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"A7",X"28",X"01",X"3D",X"21",X"97",X"8F",X"CD",X"50",X"20",X"7E",X"FE",X"06",
		X"30",X"02",X"3E",X"05",X"32",X"66",X"ED",X"18",X"05",X"3E",X"07",X"32",X"66",X"ED",X"3E",X"03",
		X"32",X"03",X"ED",X"C3",X"28",X"89",X"3A",X"03",X"ED",X"3D",X"32",X"03",X"ED",X"A7",X"C2",X"28",
		X"89",X"3E",X"18",X"32",X"03",X"ED",X"3A",X"66",X"ED",X"3D",X"32",X"66",X"ED",X"FE",X"FF",X"28",
		X"06",X"CD",X"1C",X"8E",X"C3",X"28",X"89",X"3E",X"12",X"32",X"03",X"ED",X"C3",X"28",X"89",X"3A",
		X"01",X"ED",X"D6",X"02",X"FE",X"0D",X"20",X"02",X"3E",X"10",X"32",X"01",X"ED",X"3E",X"3C",X"32",
		X"00",X"ED",X"3A",X"05",X"ED",X"CB",X"BF",X"32",X"05",X"ED",X"AF",X"32",X"02",X"ED",X"21",X"D0",
		X"2B",X"3A",X"06",X"ED",X"CD",X"58",X"8B",X"C3",X"28",X"89",X"3E",X"04",X"CF",X"3E",X"1C",X"CD",
		X"AE",X"67",X"21",X"85",X"C4",X"06",X"0A",X"23",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"10",
		X"F6",X"E7",X"3A",X"08",X"ED",X"A7",X"28",X"05",X"CD",X"D3",X"8B",X"18",X"F4",X"3A",X"02",X"ED",
		X"A7",X"28",X"10",X"3C",X"32",X"02",X"ED",X"FE",X"06",X"28",X"08",X"CD",X"45",X"8B",X"3E",X"05",
		X"DF",X"18",X"EA",X"21",X"D0",X"2B",X"3E",X"38",X"CD",X"58",X"8B",X"3E",X"28",X"32",X"03",X"ED",
		X"3E",X"FF",X"32",X"02",X"ED",X"E7",X"3A",X"03",X"ED",X"3D",X"32",X"03",X"ED",X"A7",X"20",X"F5",
		X"3A",X"02",X"ED",X"3C",X"32",X"02",X"ED",X"FE",X"0B",X"28",X"39",X"CB",X"27",X"F5",X"11",X"67",
		X"8F",X"CD",X"4A",X"20",X"1A",X"47",X"0E",X"08",X"13",X"1A",X"32",X"03",X"ED",X"F1",X"11",X"51",
		X"8F",X"CD",X"4A",X"20",X"1A",X"6F",X"13",X"1A",X"67",X"CD",X"D1",X"20",X"E5",X"21",X"3B",X"8F",
		X"3A",X"02",X"ED",X"CB",X"27",X"CD",X"50",X"20",X"5E",X"23",X"56",X"E1",X"3E",X"38",X"CD",X"55",
		X"22",X"C3",X"85",X"8A",X"3E",X"05",X"32",X"03",X"ED",X"AF",X"32",X"02",X"ED",X"21",X"7D",X"8F",
		X"7E",X"CD",X"80",X"8B",X"E7",X"3A",X"03",X"ED",X"3D",X"32",X"03",X"ED",X"20",X"F6",X"3E",X"05",
		X"32",X"03",X"ED",X"3A",X"02",X"ED",X"3C",X"FE",X"05",X"28",X"0F",X"32",X"02",X"ED",X"21",X"7D",
		X"8F",X"CD",X"50",X"20",X"7E",X"CD",X"80",X"8B",X"18",X"DA",X"21",X"20",X"00",X"11",X"0E",X"E3",
		X"06",X"0C",X"0E",X"08",X"3E",X"48",X"CD",X"66",X"8B",X"3E",X"DC",X"DF",X"3E",X"0F",X"CD",X"AE",
		X"67",X"3E",X"F0",X"DF",X"3E",X"00",X"32",X"C4",X"C4",X"3A",X"7B",X"C4",X"CB",X"EF",X"32",X"7B",
		X"C4",X"32",X"08",X"D0",X"CD",X"A6",X"A5",X"3E",X"01",X"32",X"62",X"EF",X"32",X"71",X"ED",X"3E",
		X"00",X"D7",X"AF",X"DF",X"E7",X"3A",X"02",X"ED",X"CB",X"27",X"11",X"2F",X"8F",X"CD",X"4A",X"20",
		X"1A",X"6F",X"13",X"1A",X"67",X"3A",X"06",X"ED",X"CD",X"D1",X"20",X"11",X"0E",X"E3",X"06",X"0C",
		X"0E",X"08",X"CD",X"55",X"22",X"C9",X"EB",X"C5",X"E5",X"CD",X"76",X"8B",X"E1",X"01",X"40",X"00",
		X"09",X"C1",X"0D",X"20",X"F2",X"C9",X"F5",X"B2",X"77",X"F1",X"23",X"73",X"23",X"10",X"F7",X"C9",
		X"21",X"0E",X"E3",X"06",X"0C",X"0E",X"08",X"C5",X"E5",X"CD",X"96",X"8B",X"E1",X"01",X"40",X"00",
		X"09",X"C1",X"0D",X"20",X"F2",X"C9",X"F5",X"7E",X"E6",X"07",X"57",X"F1",X"F5",X"B2",X"77",X"F1",
		X"23",X"23",X"10",X"F2",X"C9",X"21",X"D0",X"34",X"3E",X"F8",X"CD",X"58",X"8B",X"3E",X"02",X"32",
		X"0A",X"ED",X"3A",X"05",X"ED",X"CB",X"EF",X"32",X"05",X"ED",X"C9",X"F5",X"3A",X"0A",X"ED",X"3D",
		X"32",X"0A",X"ED",X"A7",X"20",X"0B",X"CD",X"45",X"8B",X"3A",X"05",X"ED",X"CB",X"AF",X"32",X"05",
		X"ED",X"F1",X"C9",X"F5",X"3A",X"07",X"ED",X"3D",X"32",X"07",X"ED",X"A7",X"20",X"25",X"3E",X"05",
		X"32",X"07",X"ED",X"3A",X"08",X"ED",X"3C",X"FE",X"0A",X"20",X"01",X"AF",X"32",X"08",X"ED",X"11",
		X"25",X"8F",X"CD",X"4A",X"20",X"1A",X"32",X"06",X"ED",X"CD",X"45",X"8B",X"3E",X"FF",X"32",X"04",
		X"ED",X"F1",X"C9",X"3E",X"00",X"32",X"04",X"ED",X"F1",X"C9",X"F5",X"3A",X"6B",X"C4",X"A7",X"CA",
		X"B5",X"8C",X"2A",X"44",X"C4",X"CD",X"B7",X"8C",X"30",X"22",X"3A",X"09",X"ED",X"CB",X"47",X"20",
		X"23",X"CB",X"C7",X"32",X"09",X"ED",X"3A",X"40",X"C4",X"CD",X"CE",X"8C",X"32",X"40",X"C4",X"3A",
		X"43",X"C4",X"CB",X"BF",X"32",X"43",X"C4",X"CD",X"15",X"8D",X"18",X"08",X"3A",X"09",X"ED",X"CB",
		X"87",X"32",X"09",X"ED",X"3A",X"6B",X"C4",X"3D",X"A7",X"28",X"6A",X"2A",X"50",X"C4",X"CD",X"B7",
		X"8C",X"30",X"22",X"3A",X"09",X"ED",X"CB",X"4F",X"20",X"23",X"CB",X"CF",X"32",X"09",X"ED",X"3A",
		X"4C",X"C4",X"CD",X"CE",X"8C",X"32",X"4C",X"C4",X"3A",X"4F",X"C4",X"CB",X"BF",X"32",X"4F",X"C4",
		X"CD",X"15",X"8D",X"18",X"08",X"3A",X"09",X"ED",X"CB",X"8F",X"32",X"09",X"ED",X"3A",X"6B",X"C4",
		X"D6",X"02",X"A7",X"28",X"30",X"2A",X"5C",X"C4",X"CD",X"B7",X"8C",X"30",X"20",X"3A",X"09",X"ED",
		X"CB",X"57",X"20",X"21",X"CB",X"D7",X"32",X"09",X"ED",X"3A",X"58",X"C4",X"CD",X"CE",X"8C",X"32",
		X"58",X"C4",X"3A",X"5B",X"C4",X"CB",X"BF",X"32",X"5B",X"C4",X"CD",X"15",X"8D",X"3A",X"09",X"ED",
		X"CB",X"97",X"32",X"09",X"ED",X"F1",X"C9",X"7D",X"FE",X"36",X"38",X"10",X"FE",X"96",X"30",X"0C",
		X"7C",X"FE",X"60",X"38",X"07",X"FE",X"9A",X"30",X"03",X"A7",X"37",X"C9",X"A7",X"C9",X"F5",X"7D",
		X"FE",X"8F",X"30",X"06",X"FE",X"3D",X"38",X"02",X"18",X"17",X"2A",X"69",X"ED",X"7D",X"FE",X"96",
		X"30",X"06",X"FE",X"36",X"38",X"02",X"18",X"22",X"F1",X"21",X"9E",X"8F",X"CD",X"50",X"20",X"7E",
		X"C9",X"7C",X"FE",X"93",X"30",X"06",X"FE",X"67",X"38",X"02",X"18",X"DE",X"2A",X"69",X"ED",X"7C",
		X"FE",X"9A",X"30",X"06",X"FE",X"60",X"38",X"02",X"18",X"DE",X"F1",X"21",X"9E",X"8F",X"CD",X"50",
		X"20",X"7E",X"EE",X"10",X"C9",X"3E",X"1B",X"CD",X"AE",X"67",X"3A",X"FD",X"EC",X"A7",X"28",X"2E",
		X"3A",X"6B",X"ED",X"3C",X"32",X"6B",X"ED",X"CB",X"67",X"20",X"23",X"3C",X"CB",X"67",X"28",X"10",
		X"3D",X"CB",X"E7",X"32",X"05",X"ED",X"3E",X"05",X"32",X"07",X"ED",X"3E",X"FF",X"32",X"08",X"ED",
		X"CD",X"A5",X"8B",X"3A",X"6B",X"ED",X"16",X"01",X"1E",X"00",X"CD",X"23",X"27",X"C9",X"3E",X"00",
		X"32",X"FD",X"EC",X"C9",X"DD",X"21",X"0B",X"ED",X"06",X"07",X"DD",X"CB",X"0B",X"7E",X"28",X"0B",
		X"CD",X"73",X"8D",X"30",X"06",X"3E",X"01",X"32",X"62",X"EF",X"C9",X"11",X"0D",X"00",X"DD",X"19",
		X"10",X"E8",X"C9",X"DD",X"7E",X"07",X"D6",X"E8",X"30",X"02",X"2F",X"3C",X"FE",X"08",X"30",X"17",
		X"3A",X"3A",X"C4",X"47",X"DD",X"7E",X"08",X"90",X"38",X"07",X"FE",X"10",X"30",X"09",X"A7",X"37",
		X"C9",X"2F",X"3C",X"FE",X"18",X"38",X"F7",X"A7",X"C9",X"06",X"07",X"DD",X"21",X"0B",X"ED",X"DD",
		X"E5",X"C5",X"DD",X"CB",X"0B",X"7E",X"28",X"2F",X"DD",X"7E",X"0B",X"E6",X"07",X"CD",X"E2",X"8D",
		X"DD",X"35",X"0C",X"DD",X"7E",X"0C",X"E6",X"0F",X"CC",X"EC",X"8D",X"FD",X"E5",X"E1",X"CD",X"4A",
		X"11",X"E5",X"FD",X"E1",X"FD",X"7E",X"00",X"FE",X"F0",X"38",X"0C",X"DD",X"CB",X"0B",X"BE",X"FD",
		X"36",X"00",X"00",X"FD",X"36",X"01",X"00",X"C1",X"DD",X"E1",X"11",X"0D",X"00",X"DD",X"19",X"10",
		X"BE",X"C9",X"21",X"82",X"8F",X"CD",X"A8",X"3D",X"E5",X"FD",X"E1",X"C9",X"DD",X"7E",X"0C",X"F6",
		X"05",X"C6",X"10",X"DD",X"77",X"0C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"0C",
		X"20",X"06",X"3E",X"05",X"DD",X"77",X"0C",X"AF",X"21",X"10",X"2B",X"CD",X"BA",X"20",X"5F",X"16",
		X"00",X"19",X"FD",X"75",X"03",X"3E",X"78",X"B4",X"FD",X"77",X"02",X"C9",X"DD",X"21",X"0B",X"ED",
		X"0E",X"07",X"DD",X"CB",X"0B",X"7E",X"20",X"0B",X"DD",X"CB",X"0B",X"FE",X"CD",X"3C",X"8E",X"CD",
		X"7C",X"8E",X"C9",X"0D",X"C8",X"11",X"0D",X"00",X"DD",X"19",X"18",X"E6",X"18",X"11",X"3A",X"01",
		X"ED",X"2F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"A7",X"20",X"02",X"3E",X"01",X"E6",X"07",X"3E",
		X"03",X"DD",X"77",X"02",X"3E",X"F5",X"DD",X"77",X"0C",X"3E",X"01",X"DD",X"77",X"04",X"3A",X"3B",
		X"C4",X"C6",X"20",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"A7",X"28",X"01",
		X"3D",X"21",X"90",X"8F",X"CD",X"50",X"20",X"7E",X"DD",X"77",X"03",X"C9",X"DD",X"7E",X"0B",X"E6",
		X"07",X"CD",X"E2",X"8D",X"FD",X"36",X"01",X"7E",X"FD",X"36",X"00",X"6A",X"AF",X"CD",X"08",X"8E",
		X"C9",X"06",X"E1",X"10",X"1E",X"0E",X"E1",X"10",X"1E",X"16",X"E1",X"10",X"1E",X"1E",X"E1",X"10",
		X"1E",X"26",X"E1",X"10",X"1E",X"2E",X"E1",X"10",X"1E",X"36",X"E1",X"10",X"1E",X"06",X"E2",X"10",
		X"20",X"0E",X"E2",X"90",X"20",X"16",X"E2",X"10",X"21",X"1E",X"E2",X"90",X"21",X"26",X"E2",X"10",
		X"22",X"2E",X"E2",X"10",X"1E",X"36",X"E2",X"10",X"1E",X"06",X"E3",X"90",X"1F",X"26",X"E3",X"90",
		X"22",X"2E",X"E3",X"10",X"1E",X"36",X"E3",X"10",X"1E",X"06",X"E4",X"10",X"1F",X"26",X"E4",X"10",
		X"23",X"2E",X"E4",X"10",X"1E",X"36",X"E4",X"10",X"1E",X"06",X"E5",X"10",X"1E",X"0E",X"E5",X"90",
		X"1E",X"16",X"E5",X"90",X"1E",X"1E",X"E5",X"90",X"1E",X"26",X"E5",X"10",X"1E",X"2E",X"E5",X"10",
		X"1E",X"36",X"E5",X"10",X"1E",X"06",X"E6",X"10",X"1E",X"0E",X"E6",X"10",X"1E",X"16",X"E6",X"10",
		X"1E",X"1E",X"E6",X"10",X"1E",X"26",X"E6",X"10",X"1E",X"2E",X"E6",X"10",X"1E",X"36",X"E6",X"10",
		X"1E",X"0C",X"00",X"04",X"08",X"80",X"10",X"18",X"20",X"28",X"30",X"28",X"20",X"18",X"10",X"D0",
		X"2B",X"D0",X"2E",X"D0",X"31",X"D0",X"34",X"D0",X"31",X"D0",X"2E",X"0E",X"E3",X"0E",X"E3",X"10",
		X"E3",X"16",X"E3",X"16",X"E3",X"18",X"E3",X"1A",X"E3",X"1C",X"E3",X"1E",X"E3",X"20",X"E3",X"20",
		X"E3",X"90",X"23",X"10",X"24",X"D0",X"24",X"D0",X"25",X"50",X"26",X"10",X"27",X"D0",X"27",X"90",
		X"28",X"50",X"29",X"D0",X"29",X"50",X"2A",X"02",X"05",X"03",X"05",X"04",X"05",X"02",X"05",X"03",
		X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"02",X"05",X"02",X"05",X"03",X"28",X"38",X"C0",X"C8",
		X"D0",X"D8",X"85",X"C4",X"89",X"C4",X"8D",X"C4",X"91",X"C4",X"95",X"C4",X"99",X"C4",X"9D",X"C4",
		X"13",X"12",X"11",X"10",X"0F",X"0E",X"0D",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"10",X"0F",
		X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"18",X"07",X"06",X"05",X"04",X"03",X"02",X"01",X"00",X"1F",
		X"1E",X"1D",X"1C",X"1B",X"1A",X"19",X"08",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"1A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",
		X"1A",X"16",X"12",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1A",X"16",X"12",
		X"0E",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1A",X"16",X"12",X"0E",X"0A",X"06",
		X"02",X"00",X"00",X"00",X"00",X"00",X"1E",X"1A",X"16",X"12",X"0E",X"0A",X"06",X"02",X"1E",X"1A",
		X"00",X"00",X"00",X"03",X"1A",X"16",X"12",X"0E",X"0A",X"06",X"02",X"1E",X"1A",X"16",X"12",X"00",
		X"00",X"FF",X"03",X"12",X"0E",X"0A",X"06",X"02",X"1E",X"1A",X"16",X"12",X"0E",X"00",X"00",X"00",
		X"FF",X"03",X"0A",X"06",X"02",X"1E",X"1A",X"16",X"12",X"0E",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"03",X"02",X"1E",X"1A",X"16",X"12",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",
		X"1A",X"16",X"12",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"12",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"12",X"00",
		X"16",X"00",X"1A",X"00",X"1E",X"00",X"02",X"00",X"06",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"16",X"00",X"12",X"00",X"0E",X"00",X"0A",X"00",X"06",
		X"00",X"02",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"0A",X"00",X"0E",X"00",X"12",X"00",X"16",X"00",X"1A",X"00",X"1E",X"00",X"02",X"03",X"00",X"03",
		X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"1A",X"00",X"16",X"00",X"12",
		X"00",X"0E",X"00",X"0A",X"00",X"06",X"00",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"06",X"00",X"0A",X"00",X"0E",X"00",X"12",X"00",X"16",X"00",X"1A",X"00",
		X"1E",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"1E",
		X"00",X"1A",X"00",X"16",X"00",X"12",X"00",X"0E",X"00",X"0A",X"00",X"00",X"03",X"00",X"03",X"00",
		X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"02",X"00",X"06",X"00",X"0A",X"00",X"0E",X"00",
		X"12",X"00",X"16",X"00",X"1A",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",X"03",
		X"00",X"03",X"AF",X"32",X"78",X"EF",X"21",X"00",X"90",X"01",X"00",X"10",X"3A",X"78",X"EF",X"86",
		X"32",X"78",X"EF",X"23",X"0B",X"78",X"B1",X"20",X"F3",X"3A",X"78",X"EF",X"21",X"73",X"A5",X"BE",
		X"28",X"0C",X"32",X"8A",X"ED",X"3D",X"32",X"61",X"EF",X"C6",X"16",X"32",X"34",X"C4",X"AF",X"32",
		X"C4",X"C4",X"CD",X"BF",X"95",X"E7",X"CD",X"17",X"21",X"3A",X"C1",X"C4",X"CB",X"57",X"CA",X"66",
		X"2A",X"3A",X"FF",X"BF",X"FE",X"76",X"C2",X"FE",X"91",X"3E",X"07",X"F7",X"E7",X"3E",X"87",X"32",
		X"00",X"EC",X"E7",X"3A",X"00",X"EC",X"A7",X"20",X"F9",X"3E",X"3C",X"DF",X"3E",X"88",X"32",X"00",
		X"EC",X"E7",X"3A",X"00",X"EC",X"A7",X"20",X"F9",X"3E",X"FF",X"DF",X"3E",X"07",X"CF",X"E7",X"CD",
		X"17",X"21",X"E7",X"18",X"2E",X"21",X"0D",X"D0",X"2B",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",
		X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"3E",X"72",X"86",X"E1",X"32",
		X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"72",X"ED",X"CB",X"27",X"57",X"3A",X"80",X"ED",X"82",
		X"32",X"18",X"D0",X"E5",X"D5",X"C5",X"21",X"2A",X"94",X"11",X"05",X"92",X"01",X"2E",X"00",X"1A",
		X"ED",X"A1",X"20",X"07",X"13",X"78",X"B1",X"20",X"F6",X"18",X"0C",X"ED",X"46",X"ED",X"5F",X"32",
		X"71",X"ED",X"32",X"86",X"ED",X"ED",X"47",X"C1",X"D1",X"E1",X"CD",X"BF",X"95",X"3E",X"01",X"32",
		X"D0",X"C4",X"3E",X"01",X"32",X"66",X"EF",X"3A",X"6C",X"ED",X"A7",X"28",X"22",X"3E",X"E9",X"ED",
		X"47",X"E7",X"3E",X"EA",X"ED",X"47",X"E7",X"3E",X"EB",X"ED",X"47",X"E7",X"3E",X"EC",X"ED",X"47",
		X"E7",X"3E",X"ED",X"ED",X"47",X"E7",X"3E",X"EE",X"ED",X"47",X"E7",X"3E",X"EF",X"ED",X"47",X"3E",
		X"01",X"F7",X"AF",X"DF",X"E7",X"3E",X"04",X"CF",X"3E",X"03",X"CF",X"3E",X"06",X"CF",X"3E",X"01",
		X"CF",X"3E",X"07",X"CF",X"E7",X"3A",X"32",X"C4",X"A7",X"28",X"BC",X"3A",X"80",X"ED",X"32",X"C4",
		X"C4",X"21",X"05",X"92",X"11",X"CB",X"92",X"06",X"1D",X"1A",X"BE",X"20",X"06",X"23",X"13",X"10",
		X"F8",X"18",X"25",X"AF",X"32",X"08",X"D0",X"39",X"E5",X"18",X"1D",X"21",X"0D",X"D0",X"2B",X"CB",
		X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",
		X"20",X"3E",X"72",X"86",X"E1",X"32",X"18",X"D0",X"3A",X"80",X"ED",X"32",X"66",X"EF",X"21",X"5C",
		X"E4",X"11",X"2B",X"9A",X"AF",X"CD",X"F1",X"21",X"21",X"11",X"93",X"E5",X"3A",X"32",X"C4",X"FE",
		X"01",X"11",X"46",X"9A",X"20",X"03",X"11",X"30",X"9A",X"21",X"62",X"E6",X"AF",X"CD",X"F1",X"21",
		X"C9",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",
		X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"E7",X"3A",X"6C",X"ED",
		X"A7",X"20",X"5F",X"CD",X"FC",X"92",X"3A",X"0C",X"D0",X"E6",X"03",X"28",X"D4",X"2F",X"E6",X"03",
		X"28",X"CF",X"47",X"3A",X"32",X"C4",X"90",X"38",X"C8",X"32",X"32",X"C4",X"78",X"CB",X"3F",X"CB",
		X"D7",X"32",X"6F",X"ED",X"3E",X"10",X"32",X"D0",X"C4",X"3A",X"C1",X"C4",X"E6",X"20",X"07",X"07",
		X"07",X"21",X"28",X"9A",X"CD",X"50",X"20",X"7E",X"32",X"76",X"ED",X"32",X"7B",X"ED",X"3E",X"EF",
		X"CD",X"AE",X"67",X"CD",X"15",X"27",X"3A",X"86",X"ED",X"A7",X"28",X"05",X"ED",X"5F",X"32",X"32",
		X"C4",X"3E",X"01",X"CD",X"C4",X"99",X"AF",X"32",X"75",X"EF",X"32",X"76",X"EF",X"21",X"77",X"ED",
		X"06",X"04",X"77",X"23",X"10",X"FC",X"21",X"7C",X"ED",X"06",X"04",X"77",X"23",X"10",X"FC",X"32",
		X"85",X"ED",X"32",X"87",X"ED",X"32",X"83",X"ED",X"32",X"62",X"EF",X"32",X"68",X"EF",X"32",X"69",
		X"EF",X"32",X"6A",X"EF",X"32",X"6B",X"EF",X"32",X"6C",X"EF",X"32",X"6E",X"EF",X"3E",X"20",X"32",
		X"6D",X"EF",X"32",X"6F",X"EF",X"CD",X"D0",X"21",X"CD",X"17",X"21",X"3A",X"6F",X"ED",X"CB",X"47",
		X"CA",X"89",X"94",X"CB",X"4F",X"CA",X"89",X"94",X"CD",X"BF",X"95",X"3A",X"FF",X"BF",X"FE",X"76",
		X"20",X"12",X"3A",X"C1",X"C4",X"CB",X"7F",X"28",X"0B",X"CD",X"45",X"96",X"3A",X"7B",X"C4",X"CB",
		X"D7",X"32",X"7B",X"C4",X"3E",X"01",X"32",X"D5",X"C4",X"3A",X"76",X"EF",X"A7",X"CC",X"74",X"A5",
		X"3E",X"FF",X"32",X"76",X"EF",X"3E",X"01",X"32",X"D5",X"C4",X"21",X"7B",X"ED",X"11",X"71",X"ED",
		X"01",X"05",X"00",X"ED",X"B0",X"21",X"76",X"EE",X"22",X"88",X"ED",X"3A",X"87",X"ED",X"32",X"83",
		X"ED",X"21",X"70",X"94",X"E5",X"A7",X"CA",X"5B",X"96",X"E1",X"21",X"0D",X"D0",X"2B",X"CB",X"76",
		X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",
		X"3E",X"72",X"86",X"E1",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"72",X"ED",X"CB",X"27",
		X"57",X"3A",X"80",X"ED",X"82",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"88",X"ED",X"32",
		X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"89",X"ED",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",
		X"3A",X"FF",X"BF",X"FE",X"76",X"20",X"0F",X"3A",X"C1",X"C4",X"CB",X"7F",X"20",X"08",X"3A",X"7B",
		X"C4",X"CB",X"97",X"32",X"7B",X"C4",X"C3",X"1A",X"95",X"3A",X"7B",X"C4",X"CB",X"97",X"32",X"7B",
		X"C4",X"CD",X"BF",X"95",X"3E",X"01",X"32",X"D5",X"C4",X"3A",X"75",X"EF",X"A7",X"CC",X"74",X"A5",
		X"3E",X"FF",X"32",X"75",X"EF",X"3E",X"01",X"32",X"D5",X"C4",X"E7",X"21",X"76",X"ED",X"11",X"71",
		X"ED",X"01",X"05",X"00",X"ED",X"B0",X"21",X"8B",X"ED",X"22",X"88",X"ED",X"3A",X"85",X"ED",X"32",
		X"83",X"ED",X"21",X"1A",X"95",X"E5",X"A7",X"CA",X"5B",X"96",X"3A",X"0C",X"D0",X"CB",X"77",X"28",
		X"F9",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"3E",
		X"72",X"86",X"E1",X"32",X"18",X"D0",X"3A",X"0C",X"D0",X"CB",X"77",X"28",X"F9",X"3A",X"84",X"ED",
		X"CB",X"27",X"CB",X"27",X"67",X"3A",X"72",X"ED",X"CB",X"27",X"84",X"32",X"18",X"D0",X"21",X"0C",
		X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"88",X"ED",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",
		X"89",X"ED",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"E1",X"3A",X"84",X"ED",X"32",X"CE",X"C4",
		X"E7",X"3E",X"04",X"F7",X"E7",X"AF",X"DF",X"E7",X"3E",X"04",X"CF",X"3E",X"00",X"32",X"C4",X"C4",
		X"CD",X"D0",X"21",X"3E",X"16",X"DF",X"3A",X"72",X"ED",X"FE",X"20",X"28",X"08",X"3A",X"7B",X"C4",
		X"CB",X"B7",X"32",X"7B",X"C4",X"3A",X"62",X"EF",X"A7",X"20",X"17",X"3A",X"72",X"ED",X"3C",X"67",
		X"3A",X"86",X"ED",X"84",X"32",X"72",X"ED",X"21",X"00",X"00",X"22",X"74",X"ED",X"CD",X"5B",X"96",
		X"18",X"B8",X"3A",X"8A",X"ED",X"32",X"62",X"EF",X"32",X"CE",X"C4",X"CD",X"D0",X"21",X"3A",X"71",
		X"ED",X"3D",X"32",X"71",X"ED",X"CC",X"74",X"97",X"3A",X"6F",X"ED",X"CB",X"47",X"28",X"0D",X"CB",
		X"4F",X"20",X"1C",X"CB",X"67",X"20",X"05",X"CB",X"CF",X"32",X"6F",X"ED",X"21",X"71",X"ED",X"11",
		X"76",X"ED",X"01",X"05",X"00",X"ED",X"B0",X"3A",X"83",X"ED",X"32",X"85",X"ED",X"18",X"1A",X"CB",
		X"5F",X"20",X"05",X"CB",X"8F",X"32",X"6F",X"ED",X"21",X"71",X"ED",X"11",X"7B",X"ED",X"01",X"05",
		X"00",X"ED",X"B0",X"3A",X"83",X"ED",X"32",X"87",X"ED",X"C3",X"CB",X"93",X"C3",X"5A",X"92",X"3A",
		X"7B",X"C4",X"E6",X"FC",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"3A",X"C1",X"C4",X"CB",X"4F",X"20",
		X"0B",X"3A",X"7B",X"C4",X"F6",X"03",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"E5",X"D5",X"C5",X"21",
		X"CA",X"94",X"11",X"0E",X"96",X"01",X"37",X"00",X"1A",X"ED",X"A1",X"20",X"07",X"13",X"78",X"B1",
		X"20",X"F6",X"18",X"0C",X"ED",X"5E",X"ED",X"5F",X"77",X"32",X"6E",X"ED",X"ED",X"47",X"18",X"FD",
		X"C1",X"D1",X"E1",X"C9",X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",X"38",X"39",X"3A",X"0C",
		X"D0",X"CB",X"77",X"28",X"F9",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",
		X"CD",X"50",X"20",X"3E",X"72",X"86",X"E1",X"32",X"18",X"D0",X"3A",X"0C",X"D0",X"CB",X"77",X"28",
		X"F9",X"3A",X"84",X"ED",X"CB",X"27",X"CB",X"27",X"67",X"3A",X"72",X"ED",X"CB",X"27",X"84",X"32",
		X"18",X"D0",X"21",X"0C",X"D0",X"3A",X"7B",X"C4",X"E6",X"03",X"2F",X"E6",X"03",X"47",X"3A",X"7B",
		X"C4",X"E6",X"FC",X"B0",X"32",X"7B",X"C4",X"32",X"08",X"D0",X"C9",X"21",X"0C",X"D0",X"CB",X"76",
		X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",
		X"3E",X"22",X"86",X"E1",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"72",X"ED",X"CB",X"27",
		X"57",X"3A",X"6C",X"ED",X"82",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"6C",X"ED",X"32",
		X"18",X"D0",X"CB",X"76",X"28",X"FC",X"3A",X"88",X"ED",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",
		X"3A",X"89",X"ED",X"32",X"18",X"D0",X"CB",X"76",X"28",X"FC",X"CB",X"7E",X"20",X"FC",X"ED",X"5F",
		X"28",X"F8",X"18",X"00",X"11",X"5C",X"9A",X"CD",X"4A",X"20",X"7E",X"22",X"81",X"ED",X"CB",X"7F",
		X"C2",X"00",X"00",X"3A",X"18",X"D0",X"5F",X"CB",X"7E",X"20",X"FC",X"ED",X"5F",X"28",X"F8",X"D5",
		X"01",X"6F",X"9A",X"7E",X"CB",X"7F",X"C2",X"00",X"00",X"CD",X"4A",X"20",X"22",X"81",X"ED",X"D1",
		X"3A",X"18",X"D0",X"57",X"CB",X"7E",X"20",X"FC",X"ED",X"5F",X"28",X"F8",X"D5",X"01",X"5C",X"9A",
		X"7E",X"CB",X"7F",X"C2",X"00",X"00",X"CD",X"4A",X"20",X"22",X"81",X"ED",X"D1",X"3A",X"18",X"D0",
		X"CD",X"4A",X"20",X"3A",X"6E",X"ED",X"CD",X"4A",X"20",X"CB",X"76",X"28",X"FC",X"3A",X"C1",X"C4",
		X"32",X"18",X"D0",X"EB",X"E7",X"ED",X"5B",X"88",X"ED",X"01",X"EA",X"00",X"ED",X"A0",X"1B",X"1A",
		X"FE",X"03",X"20",X"0A",X"3A",X"72",X"ED",X"CB",X"3F",X"C6",X"04",X"F6",X"03",X"12",X"3A",X"86",
		X"ED",X"A7",X"20",X"FD",X"13",X"78",X"B1",X"20",X"E3",X"3A",X"72",X"ED",X"FE",X"20",X"20",X"0F",
		X"3A",X"75",X"EE",X"2A",X"88",X"ED",X"06",X"EA",X"77",X"10",X"FD",X"3D",X"32",X"83",X"ED",X"3A",
		X"C1",X"C4",X"CB",X"5F",X"3E",X"03",X"20",X"0D",X"32",X"64",X"EF",X"AF",X"32",X"65",X"EF",X"26",
		X"D0",X"2E",X"18",X"7E",X"C9",X"21",X"17",X"D0",X"23",X"7E",X"32",X"64",X"EF",X"3A",X"6A",X"C6",
		X"32",X"65",X"EF",X"C9",X"3A",X"72",X"ED",X"FE",X"20",X"20",X"10",X"CD",X"17",X"21",X"3E",X"01",
		X"32",X"D5",X"C4",X"3A",X"7B",X"C4",X"CB",X"B7",X"32",X"7B",X"C4",X"3A",X"6F",X"ED",X"CB",X"47",
		X"CA",X"35",X"98",X"CB",X"4F",X"28",X"04",X"CB",X"E7",X"18",X"02",X"CB",X"DF",X"32",X"6F",X"ED",
		X"CD",X"D4",X"A0",X"CD",X"C9",X"28",X"3A",X"AE",X"EF",X"FE",X"00",X"20",X"05",X"3E",X"0E",X"CD",
		X"AE",X"67",X"E7",X"21",X"00",X"20",X"01",X"00",X"10",X"AF",X"32",X"60",X"EF",X"3A",X"60",X"EF",
		X"86",X"23",X"32",X"60",X"EF",X"0B",X"78",X"B1",X"20",X"F3",X"3A",X"60",X"EF",X"21",X"46",X"35",
		X"BE",X"28",X"0A",X"32",X"86",X"ED",X"32",X"75",X"EE",X"3E",X"EC",X"ED",X"47",X"06",X"B4",X"26",
		X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",
		X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"E7",X"10",X"E6",X"CD",X"D0",X"21",
		X"E7",X"CD",X"55",X"9B",X"3A",X"6F",X"ED",X"E6",X"18",X"FE",X"18",X"28",X"6D",X"21",X"00",X"40",
		X"01",X"00",X"10",X"AF",X"32",X"60",X"EF",X"3A",X"60",X"EF",X"86",X"23",X"32",X"60",X"EF",X"0B",
		X"78",X"B1",X"20",X"F3",X"3A",X"60",X"EF",X"21",X"74",X"55",X"BE",X"28",X"07",X"3E",X"EC",X"ED",
		X"47",X"32",X"6F",X"ED",X"C9",X"3E",X"02",X"CD",X"C4",X"99",X"AF",X"32",X"70",X"EF",X"3E",X"20",
		X"CD",X"C4",X"99",X"21",X"D7",X"C4",X"7E",X"CD",X"AB",X"99",X"23",X"7E",X"CD",X"AB",X"99",X"23",
		X"7E",X"CD",X"AB",X"99",X"23",X"3E",X"30",X"CD",X"C4",X"99",X"3E",X"03",X"CD",X"C4",X"99",X"3A",
		X"77",X"ED",X"3C",X"CD",X"92",X"99",X"CD",X"D4",X"A0",X"CD",X"55",X"9B",X"3A",X"AE",X"EF",X"FE",
		X"00",X"20",X"6F",X"3E",X"0E",X"CD",X"AE",X"67",X"18",X"68",X"3E",X"02",X"CD",X"C4",X"99",X"3E",
		X"20",X"CD",X"C4",X"99",X"AF",X"32",X"70",X"EF",X"21",X"D7",X"C4",X"7E",X"CD",X"AB",X"99",X"23",
		X"7E",X"CD",X"AB",X"99",X"23",X"7E",X"CD",X"AB",X"99",X"23",X"3E",X"30",X"CD",X"C4",X"99",X"3E",
		X"03",X"CD",X"C4",X"99",X"3A",X"77",X"ED",X"3C",X"CD",X"92",X"99",X"3E",X"04",X"CD",X"C4",X"99",
		X"AF",X"32",X"70",X"EF",X"3E",X"20",X"CD",X"C4",X"99",X"21",X"DB",X"C4",X"7E",X"CD",X"AB",X"99",
		X"23",X"7E",X"CD",X"AB",X"99",X"23",X"7E",X"CD",X"AB",X"99",X"23",X"3E",X"30",X"CD",X"C4",X"99",
		X"3E",X"05",X"CD",X"C4",X"99",X"3A",X"7C",X"ED",X"3C",X"CD",X"92",X"99",X"3E",X"01",X"32",X"D5",
		X"C4",X"E7",X"CD",X"17",X"21",X"3E",X"01",X"32",X"D5",X"C4",X"F5",X"CD",X"0A",X"29",X"F1",X"CD",
		X"BF",X"95",X"3E",X"0F",X"32",X"FF",X"C7",X"E7",X"AF",X"32",X"78",X"EF",X"21",X"00",X"80",X"01",
		X"00",X"10",X"3A",X"78",X"EF",X"86",X"32",X"78",X"EF",X"23",X"0B",X"78",X"B1",X"20",X"F3",X"3A",
		X"78",X"EF",X"21",X"DE",X"9D",X"BE",X"28",X"05",X"32",X"86",X"ED",X"ED",X"5E",X"06",X"F0",X"26",
		X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",
		X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"E7",X"10",X"E6",X"CD",X"D0",X"21",
		X"AF",X"32",X"6F",X"ED",X"3E",X"10",X"32",X"D5",X"C4",X"E7",X"3E",X"00",X"CD",X"AE",X"67",X"E7",
		X"CD",X"17",X"21",X"3E",X"EE",X"CD",X"AE",X"67",X"21",X"00",X"60",X"01",X"00",X"10",X"AF",X"32",
		X"60",X"EF",X"3A",X"60",X"EF",X"86",X"23",X"32",X"60",X"EF",X"0B",X"78",X"B1",X"20",X"F3",X"3A",
		X"60",X"EF",X"21",X"D7",X"75",X"BE",X"28",X"16",X"3E",X"07",X"F7",X"E7",X"3E",X"40",X"32",X"00",
		X"EC",X"E7",X"3A",X"00",X"EC",X"A7",X"18",X"F9",X"3E",X"0A",X"DF",X"ED",X"5E",X"E1",X"E1",X"C3",
		X"5A",X"92",X"E5",X"D5",X"C5",X"11",X"70",X"EF",X"CD",X"A2",X"84",X"21",X"71",X"EF",X"7E",X"CD",
		X"C4",X"99",X"23",X"7E",X"CD",X"C4",X"99",X"C1",X"D1",X"E1",X"C9",X"E5",X"D5",X"C5",X"11",X"70",
		X"EF",X"CD",X"F7",X"99",X"21",X"71",X"EF",X"7E",X"CD",X"C4",X"99",X"23",X"7E",X"CD",X"C4",X"99",
		X"C1",X"D1",X"E1",X"C9",X"C5",X"F5",X"3A",X"FF",X"C7",X"47",X"F1",X"32",X"FF",X"C7",X"0E",X"02",
		X"E7",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",
		X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"0D",X"28",X"06",X"3A",
		X"FF",X"C7",X"B8",X"28",X"DB",X"C1",X"C9",X"47",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"20",X"0A",X"1A",X"A7",X"3E",X"20",X"28",X"07",X"3E",X"30",X"18",X"03",X"C6",X"30",X"12",X"13",
		X"12",X"1B",X"78",X"E6",X"0F",X"20",X"0A",X"1A",X"A7",X"3E",X"20",X"28",X"07",X"3E",X"30",X"18",
		X"03",X"C6",X"30",X"12",X"13",X"13",X"12",X"C9",X"05",X"03",X"06",X"04",X"50",X"55",X"53",X"48",
		X"15",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"42",
		X"55",X"54",X"54",X"4F",X"4E",X"20",X"15",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"12",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"31",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"12",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"32",X"20",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",
		X"45",X"52",X"09",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"0E",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"31",X"20",X"52",X"45",X"41",X"44",X"59",X"0E",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"32",X"20",X"52",X"45",X"41",X"44",X"59",X"05",X"52",X"45",X"41",X"44",X"59",
		X"10",X"54",X"4F",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",X"55",X"45",X"20",X"47",X"41",X"4D",
		X"45",X"1A",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"41",X"44",X"44",X"49",X"54",X"49",X"4F",
		X"4E",X"41",X"4C",X"20",X"43",X"4F",X"49",X"4E",X"28",X"53",X"29",X"2C",X"19",X"48",X"4F",X"4C",
		X"44",X"20",X"46",X"49",X"52",X"45",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"20",X"41",X"4E",
		X"44",X"20",X"50",X"55",X"53",X"48",X"14",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"0D",X"4F",X"4E",X"4C",X"59",
		X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"06",X"42",X"45",X"46",X"4F",X"52",X"45",
		X"12",X"54",X"49",X"4D",X"45",X"52",X"20",X"52",X"45",X"41",X"43",X"48",X"45",X"53",X"20",X"22",
		X"30",X"22",X"2E",X"07",X"54",X"49",X"4D",X"45",X"20",X"20",X"39",X"3B",X"CB",X"76",X"28",X"FC",
		X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"3E",X"72",
		X"86",X"E1",X"32",X"18",X"D0",X"21",X"2E",X"94",X"11",X"3C",X"9B",X"01",X"19",X"00",X"1A",X"ED",
		X"A1",X"20",X"07",X"13",X"78",X"B1",X"20",X"F6",X"18",X"0A",X"ED",X"5F",X"32",X"6C",X"ED",X"32",
		X"32",X"C4",X"ED",X"47",X"3A",X"C1",X"C4",X"CB",X"47",X"C0",X"CD",X"17",X"21",X"CD",X"D0",X"21",
		X"3E",X"01",X"32",X"D5",X"C4",X"32",X"D0",X"C4",X"3A",X"72",X"ED",X"FE",X"20",X"C8",X"21",X"CA",
		X"E5",X"11",X"B0",X"9A",X"3E",X"01",X"CD",X"F1",X"21",X"3A",X"32",X"C4",X"A7",X"20",X"0A",X"21",
		X"D2",X"E6",X"11",X"C1",X"9A",X"AF",X"CD",X"F1",X"21",X"21",X"D6",X"E6",X"11",X"DC",X"9A",X"AF",
		X"CD",X"F1",X"21",X"21",X"DA",X"E6",X"11",X"F6",X"9A",X"AF",X"CD",X"F1",X"21",X"21",X"62",X"E6",
		X"11",X"19",X"9B",X"AF",X"CD",X"F1",X"21",X"21",X"66",X"E6",X"11",X"20",X"9B",X"AF",X"CD",X"F1",
		X"21",X"21",X"6C",X"E5",X"11",X"33",X"9B",X"3E",X"02",X"CD",X"F1",X"21",X"06",X"09",X"21",X"3C",
		X"00",X"22",X"73",X"EF",X"3A",X"0C",X"D0",X"E6",X"03",X"FE",X"03",X"20",X"47",X"3A",X"32",X"C4",
		X"A7",X"28",X"0C",X"21",X"D2",X"E6",X"11",X"C1",X"9A",X"AF",X"C5",X"CD",X"1C",X"22",X"C1",X"E7",
		X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",
		X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",X"32",X"18",X"D0",X"2A",X"73",X"EF",X"2B",X"22",
		X"73",X"EF",X"7C",X"B5",X"20",X"BE",X"78",X"C6",X"2F",X"32",X"ED",X"E3",X"10",X"B0",X"3E",X"10",
		X"32",X"D0",X"C4",X"C9",X"3A",X"6F",X"ED",X"CB",X"47",X"28",X"1A",X"CB",X"4F",X"28",X"16",X"3A",
		X"FF",X"BF",X"FE",X"76",X"20",X"0F",X"3A",X"C1",X"C4",X"CB",X"7F",X"28",X"08",X"3A",X"10",X"D0",
		X"CB",X"57",X"28",X"07",X"C9",X"3A",X"10",X"D0",X"CB",X"47",X"C0",X"3A",X"32",X"C4",X"A7",X"28",
		X"9E",X"3D",X"32",X"32",X"C4",X"3A",X"6F",X"ED",X"CB",X"47",X"28",X"20",X"CB",X"4F",X"28",X"1C",
		X"CB",X"A7",X"32",X"6F",X"ED",X"AF",X"32",X"69",X"EF",X"32",X"6B",X"EF",X"32",X"6E",X"EF",X"3E",
		X"20",X"32",X"6F",X"EF",X"21",X"DB",X"C4",X"CD",X"E8",X"9C",X"18",X"1A",X"CB",X"9F",X"32",X"6F",
		X"ED",X"AF",X"32",X"68",X"EF",X"32",X"6A",X"EF",X"32",X"6C",X"EF",X"3E",X"20",X"32",X"6D",X"EF",
		X"21",X"D7",X"C4",X"CD",X"E8",X"9C",X"3A",X"C1",X"C4",X"E6",X"20",X"07",X"07",X"07",X"21",X"28",
		X"9A",X"CD",X"50",X"20",X"7E",X"32",X"71",X"ED",X"21",X"00",X"00",X"22",X"74",X"ED",X"CD",X"5B",
		X"96",X"3E",X"10",X"32",X"D0",X"C4",X"06",X"1E",X"26",X"D0",X"2E",X"0C",X"CB",X"76",X"28",X"FC",
		X"3A",X"C7",X"C4",X"3C",X"32",X"C7",X"C4",X"E5",X"21",X"98",X"7E",X"CD",X"50",X"20",X"7E",X"E1",
		X"32",X"18",X"D0",X"E7",X"10",X"E6",X"E1",X"C9",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",
		X"23",X"36",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"0E",X"0D",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"FF",X"00",X"FF",X"12",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"16",X"15",X"15",X"15",X"15",
		X"15",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"1A",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"1E",X"1D",X"1D",X"1D",
		X"1D",X"1D",X"1D",X"1D",X"1D",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"19",X"00",X"00",X"00",X"19",X"19",X"00",X"00",X"00",
		X"00",X"00",X"19",X"19",X"19",X"19",X"00",X"19",X"19",X"19",X"19",X"00",X"00",X"00",X"00",X"19",
		X"19",X"19",X"19",X"00",X"19",X"19",X"1A",X"19",X"00",X"00",X"00",X"19",X"19",X"1A",X"19",X"03",
		X"03",X"19",X"19",X"19",X"19",X"19",X"00",X"00",X"19",X"19",X"19",X"19",X"03",X"03",X"19",X"19",
		X"19",X"19",X"19",X"00",X"00",X"19",X"19",X"19",X"19",X"19",X"03",X"03",X"1A",X"19",X"1A",X"19",
		X"00",X"00",X"19",X"19",X"1A",X"19",X"19",X"03",X"03",X"19",X"19",X"19",X"1A",X"00",X"00",X"00",
		X"19",X"19",X"19",X"03",X"03",X"19",X"19",X"19",X"19",X"00",X"00",X"00",X"00",X"19",X"19",X"1A",
		X"03",X"03",X"19",X"19",X"19",X"19",X"00",X"00",X"00",X"00",X"00",X"19",X"19",X"19",X"03",X"03",
		X"1A",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"19",X"19",X"03",X"03",X"19",X"19",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"03",X"03",X"19",X"19",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"03",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"D5",X"9E",X"11",X"79",X"EF",X"01",
		X"23",X"00",X"ED",X"B0",X"C9",X"00",X"50",X"00",X"05",X"53",X"53",X"42",X"00",X"45",X"00",X"04",
		X"53",X"4E",X"44",X"00",X"40",X"00",X"03",X"54",X"4F",X"52",X"00",X"35",X"00",X"02",X"4F",X"4E",
		X"4A",X"00",X"30",X"00",X"01",X"41",X"4B",X"52",X"3A",X"66",X"EF",X"A7",X"28",X"14",X"3E",X"10",
		X"32",X"D5",X"C4",X"CD",X"90",X"A4",X"CD",X"9C",X"A4",X"E7",X"3E",X"01",X"32",X"D5",X"C4",X"32",
		X"D0",X"C4",X"3A",X"66",X"EF",X"A7",X"28",X"04",X"06",X"09",X"18",X"02",X"06",X"06",X"FD",X"21",
		X"F2",X"9F",X"CD",X"1D",X"A4",X"3A",X"66",X"EF",X"A7",X"20",X"2D",X"21",X"C2",X"A0",X"11",X"18",
		X"E6",X"0E",X"10",X"CD",X"0D",X"A4",X"21",X"97",X"A0",X"0E",X"08",X"11",X"52",X"E6",X"CD",X"0D",
		X"A4",X"21",X"8D",X"A0",X"11",X"7E",X"E2",X"0E",X"00",X"CD",X"0D",X"A4",X"21",X"72",X"ED",X"7E",
		X"3C",X"FD",X"21",X"FE",X"E0",X"CD",X"2B",X"A5",X"21",X"E8",X"E5",X"11",X"79",X"EF",X"06",X"05",
		X"C5",X"D5",X"E5",X"E5",X"CD",X"39",X"A4",X"E1",X"36",X"00",X"23",X"11",X"80",X"01",X"B7",X"ED",
		X"52",X"36",X"30",X"2B",X"36",X"00",X"E1",X"D1",X"23",X"23",X"23",X"23",X"3E",X"07",X"CD",X"EA",
		X"A3",X"C1",X"10",X"DC",X"06",X"05",X"FD",X"21",X"28",X"E3",X"21",X"7C",X"EF",X"C5",X"E5",X"7E",
		X"FE",X"FF",X"20",X"1C",X"F5",X"C5",X"D5",X"E5",X"FD",X"E5",X"D1",X"1B",X"1B",X"21",X"93",X"A0",
		X"3E",X"42",X"CD",X"EA",X"A3",X"0E",X"10",X"CD",X"0D",X"A4",X"E1",X"D1",X"C1",X"F1",X"18",X"03",
		X"CD",X"2B",X"A5",X"E1",X"3E",X"07",X"CD",X"F2",X"A3",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",
		X"23",X"C1",X"10",X"C9",X"06",X"05",X"21",X"7D",X"EF",X"11",X"28",X"E2",X"C5",X"E5",X"D5",X"06",
		X"03",X"AF",X"12",X"13",X"7E",X"12",X"3E",X"41",X"CD",X"F9",X"A3",X"23",X"10",X"F3",X"D1",X"E1",
		X"C1",X"13",X"13",X"13",X"13",X"3E",X"07",X"CD",X"F2",X"A3",X"10",X"E0",X"3A",X"66",X"EF",X"A7",
		X"C8",X"C9",X"64",X"E5",X"26",X"A0",X"10",X"E8",X"E6",X"37",X"A0",X"00",X"EC",X"E6",X"3B",X"A0",
		X"00",X"F0",X"E6",X"3F",X"A0",X"00",X"F4",X"E6",X"43",X"A0",X"00",X"F8",X"E6",X"47",X"A0",X"00",
		X"D0",X"E5",X"4B",X"A0",X"10",X"14",X"E7",X"5D",X"A0",X"10",X"58",X"E6",X"78",X"A0",X"10",X"06",
		X"42",X"45",X"53",X"54",X"20",X"35",X"10",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"4F",X"55",
		X"4E",X"44",X"20",X"4E",X"41",X"4D",X"45",X"03",X"31",X"53",X"54",X"03",X"32",X"4E",X"44",X"03",
		X"33",X"52",X"44",X"03",X"34",X"54",X"48",X"03",X"35",X"54",X"48",X"11",X"54",X"48",X"45",X"20",
		X"46",X"4F",X"4C",X"4C",X"4F",X"57",X"49",X"4E",X"47",X"20",X"41",X"52",X"45",X"1A",X"54",X"48",
		X"45",X"20",X"52",X"45",X"43",X"4F",X"52",X"44",X"53",X"20",X"4F",X"46",X"20",X"54",X"48",X"45",
		X"20",X"42",X"52",X"41",X"56",X"45",X"53",X"54",X"14",X"46",X"49",X"47",X"48",X"54",X"45",X"52",
		X"53",X"20",X"4F",X"46",X"20",X"41",X"52",X"4B",X"41",X"4E",X"4F",X"49",X"44",X"05",X"52",X"4F",
		X"55",X"4E",X"44",X"03",X"41",X"4C",X"4C",X"15",X"45",X"4E",X"54",X"45",X"52",X"20",X"59",X"4F",
		X"55",X"52",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"21",X"14",X"45",X"4E",
		X"54",X"45",X"52",X"20",X"32",X"55",X"50",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"53",
		X"20",X"21",X"11",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"4F",X"55",X"4E",X"44",X"20",X"20",
		X"4E",X"41",X"4D",X"45",X"21",X"D7",X"C4",X"11",X"9C",X"EF",X"01",X"03",X"00",X"ED",X"B0",X"21",
		X"DB",X"C4",X"11",X"A0",X"EF",X"01",X"03",X"00",X"ED",X"B0",X"21",X"72",X"ED",X"7E",X"47",X"3A",
		X"EF",X"EF",X"FE",X"01",X"20",X"06",X"06",X"FE",X"AF",X"32",X"EF",X"EF",X"78",X"3C",X"32",X"9F",
		X"EF",X"32",X"A3",X"EF",X"3E",X"00",X"32",X"A9",X"EF",X"AF",X"32",X"AA",X"EF",X"32",X"AB",X"EF",
		X"32",X"A7",X"EF",X"32",X"AD",X"EF",X"32",X"AE",X"EF",X"3A",X"C4",X"C4",X"32",X"AF",X"EF",X"3E",
		X"FF",X"32",X"C4",X"C4",X"E7",X"3A",X"7C",X"C4",X"32",X"A4",X"EF",X"CD",X"39",X"A1",X"3A",X"A5",
		X"EF",X"FE",X"05",X"CA",X"96",X"A3",X"C3",X"9D",X"A1",X"3A",X"6F",X"ED",X"21",X"9C",X"EF",X"CB",
		X"4F",X"28",X"03",X"21",X"A0",X"EF",X"06",X"05",X"11",X"95",X"EF",X"CD",X"53",X"A5",X"FE",X"01",
		X"28",X"0C",X"E5",X"EB",X"11",X"07",X"00",X"B7",X"ED",X"52",X"EB",X"E1",X"10",X"ED",X"21",X"A5",
		X"EF",X"70",X"78",X"FE",X"05",X"C8",X"FE",X"04",X"28",X"1D",X"2F",X"E6",X"03",X"3C",X"06",X"07",
		X"CD",X"7A",X"A4",X"E5",X"C1",X"21",X"94",X"EF",X"11",X"9B",X"EF",X"ED",X"B8",X"21",X"03",X"00",
		X"EB",X"B7",X"ED",X"52",X"EB",X"18",X"03",X"11",X"98",X"EF",X"3A",X"6F",X"ED",X"21",X"9F",X"EF",
		X"CB",X"4F",X"28",X"03",X"21",X"A3",X"EF",X"01",X"04",X"00",X"ED",X"B8",X"C9",X"3E",X"0F",X"CD",
		X"AE",X"67",X"3E",X"01",X"32",X"AE",X"EF",X"3A",X"A5",X"EF",X"06",X"07",X"CD",X"7A",X"A4",X"11",
		X"7D",X"EF",X"19",X"01",X"03",X"00",X"3E",X"20",X"CD",X"A8",X"A4",X"3E",X"10",X"32",X"D5",X"C4",
		X"CD",X"90",X"A4",X"CD",X"9C",X"A4",X"E7",X"3E",X"01",X"32",X"D5",X"C4",X"CD",X"F8",X"9E",X"CD",
		X"9D",X"A3",X"3A",X"6F",X"ED",X"11",X"9C",X"EF",X"CB",X"4F",X"28",X"03",X"11",X"A0",X"EF",X"21",
		X"9C",X"E6",X"CD",X"39",X"A4",X"3E",X"30",X"32",X"1D",X"E5",X"3E",X"00",X"32",X"1C",X"E5",X"3A",
		X"6F",X"ED",X"21",X"9F",X"EF",X"CB",X"4F",X"28",X"03",X"21",X"A3",X"EF",X"3A",X"EF",X"EF",X"FE",
		X"01",X"20",X"07",X"3E",X"FF",X"77",X"AF",X"32",X"EF",X"EF",X"7E",X"FD",X"21",X"DC",X"E3",X"FE",
		X"FF",X"20",X"1E",X"F5",X"C5",X"D5",X"E5",X"FD",X"2B",X"FD",X"2B",X"21",X"93",X"A0",X"FD",X"E5",
		X"D1",X"3E",X"42",X"CD",X"EA",X"A3",X"0E",X"10",X"CD",X"0D",X"A4",X"E1",X"D1",X"C1",X"F1",X"18",
		X"03",X"CD",X"2B",X"A5",X"AF",X"32",X"A7",X"EF",X"32",X"A6",X"EF",X"32",X"AC",X"EF",X"01",X"58",
		X"02",X"3E",X"04",X"DF",X"0B",X"79",X"B0",X"CA",X"42",X"A3",X"3A",X"AD",X"EF",X"FE",X"00",X"20",
		X"09",X"21",X"C2",X"01",X"B7",X"ED",X"42",X"CA",X"42",X"A3",X"CD",X"B0",X"A4",X"3A",X"AC",X"EF",
		X"3C",X"32",X"AC",X"EF",X"FE",X"04",X"20",X"1D",X"AF",X"32",X"AC",X"EF",X"21",X"A4",X"EF",X"3E",
		X"FC",X"A6",X"77",X"3A",X"7C",X"C4",X"E6",X"FC",X"96",X"28",X"0A",X"CB",X"7F",X"3A",X"7C",X"C4",
		X"77",X"20",X"31",X"18",X"41",X"21",X"A4",X"EF",X"3A",X"7C",X"C4",X"77",X"3A",X"6F",X"ED",X"21",
		X"10",X"D0",X"CB",X"4F",X"28",X"14",X"3A",X"FF",X"BF",X"FE",X"76",X"20",X"0D",X"3A",X"C1",X"C4",
		X"CB",X"7F",X"28",X"06",X"CB",X"56",X"28",X"30",X"18",X"04",X"CB",X"46",X"28",X"2A",X"AF",X"32",
		X"A8",X"EF",X"18",X"6D",X"3E",X"01",X"32",X"AD",X"EF",X"21",X"A7",X"EF",X"35",X"7E",X"FE",X"FF",
		X"20",X"5F",X"36",X"1C",X"18",X"5B",X"3E",X"01",X"32",X"AD",X"EF",X"21",X"A7",X"EF",X"34",X"7E",
		X"FE",X"1D",X"20",X"4D",X"36",X"00",X"18",X"49",X"3E",X"01",X"32",X"AD",X"EF",X"21",X"A8",X"EF",
		X"CB",X"46",X"C2",X"21",X"A3",X"CB",X"C6",X"3A",X"A6",X"EF",X"CD",X"87",X"A4",X"21",X"9C",X"E2",
		X"B7",X"ED",X"52",X"36",X"10",X"3A",X"A5",X"EF",X"C5",X"06",X"07",X"CD",X"7A",X"A4",X"C1",X"11",
		X"7D",X"EF",X"19",X"3A",X"A6",X"EF",X"CD",X"F2",X"A3",X"3A",X"A7",X"EF",X"11",X"CD",X"A3",X"CD",
		X"EA",X"A3",X"1A",X"77",X"AF",X"32",X"A7",X"EF",X"21",X"A6",X"EF",X"34",X"7E",X"FE",X"03",X"28",
		X"21",X"3A",X"A6",X"EF",X"CD",X"87",X"A4",X"21",X"9C",X"E2",X"23",X"B7",X"ED",X"52",X"3A",X"A7",
		X"EF",X"11",X"CD",X"A3",X"CD",X"EA",X"A3",X"1A",X"77",X"2B",X"3A",X"A9",X"EF",X"77",X"23",X"C3",
		X"41",X"A2",X"E7",X"3A",X"A5",X"EF",X"06",X"07",X"CD",X"7A",X"A4",X"11",X"7D",X"EF",X"19",X"7E",
		X"FE",X"53",X"20",X"14",X"23",X"7E",X"FE",X"45",X"20",X"0E",X"23",X"7E",X"FE",X"58",X"20",X"08",
		X"36",X"21",X"2B",X"36",X"20",X"2B",X"36",X"48",X"CD",X"F8",X"9E",X"01",X"3C",X"00",X"3E",X"02",
		X"DF",X"CD",X"9D",X"A3",X"0B",X"78",X"B1",X"20",X"F5",X"3E",X"0E",X"CD",X"AE",X"67",X"CD",X"9D",
		X"A3",X"AF",X"32",X"A5",X"EF",X"3E",X"78",X"DF",X"3E",X"10",X"32",X"D5",X"C4",X"CD",X"90",X"A4",
		X"E7",X"3E",X"01",X"32",X"D5",X"C4",X"3A",X"AF",X"EF",X"32",X"C4",X"C4",X"C9",X"3A",X"A5",X"EF",
		X"87",X"87",X"21",X"E8",X"E6",X"CD",X"F2",X"A3",X"06",X"18",X"36",X"10",X"3E",X"40",X"CD",X"04",
		X"A4",X"10",X"F7",X"C9",X"3A",X"A5",X"EF",X"87",X"87",X"21",X"E8",X"E6",X"CD",X"F2",X"A3",X"06",
		X"18",X"3A",X"A9",X"EF",X"77",X"3E",X"40",X"CD",X"04",X"A4",X"10",X"F5",X"C9",X"41",X"42",X"43",
		X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",X"4F",X"50",X"51",X"52",X"53",
		X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"2E",X"21",X"20",X"E5",X"26",X"00",X"6F",X"19",X"EB",
		X"E1",X"C9",X"D5",X"16",X"00",X"5F",X"19",X"D1",X"C9",X"E5",X"EB",X"16",X"00",X"5F",X"B7",X"ED",
		X"52",X"EB",X"E1",X"C9",X"D5",X"16",X"00",X"5F",X"B7",X"ED",X"52",X"D1",X"C9",X"46",X"23",X"79",
		X"12",X"13",X"7E",X"12",X"23",X"3E",X"41",X"CD",X"F9",X"A3",X"10",X"F3",X"C9",X"C5",X"FD",X"5E",
		X"00",X"FD",X"56",X"01",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"FD",X"4E",X"04",X"CD",X"0D",X"A4",
		X"C1",X"11",X"05",X"00",X"FD",X"19",X"10",X"E5",X"C9",X"0E",X"30",X"06",X"03",X"E5",X"36",X"00",
		X"23",X"1A",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"81",X"77",X"3E",X"41",X"CD",X"04",
		X"A4",X"36",X"00",X"23",X"1A",X"E6",X"0F",X"81",X"77",X"3E",X"41",X"CD",X"04",X"A4",X"13",X"10",
		X"DD",X"E1",X"23",X"06",X"06",X"7E",X"B9",X"C0",X"1E",X"20",X"79",X"FE",X"30",X"28",X"02",X"1E",
		X"60",X"73",X"3E",X"40",X"CD",X"04",X"A4",X"10",X"EC",X"C9",X"D5",X"26",X"00",X"2E",X"00",X"16",
		X"00",X"5F",X"19",X"10",X"FD",X"D1",X"C9",X"C5",X"06",X"40",X"CD",X"7A",X"A4",X"EB",X"C1",X"C9",
		X"21",X"00",X"E0",X"01",X"FE",X"07",X"3E",X"20",X"CD",X"A8",X"A4",X"C9",X"21",X"00",X"E8",X"01",
		X"3F",X"00",X"3E",X"00",X"CD",X"A8",X"A4",X"C9",X"0B",X"E5",X"D1",X"13",X"77",X"ED",X"B0",X"C9",
		X"F5",X"E5",X"21",X"AA",X"EF",X"34",X"7E",X"FE",X"02",X"20",X"1F",X"AF",X"77",X"21",X"AB",X"EF",
		X"34",X"7E",X"FE",X"01",X"28",X"06",X"FE",X"02",X"28",X"09",X"18",X"0E",X"3E",X"00",X"32",X"A9",
		X"EF",X"18",X"07",X"3E",X"08",X"32",X"A9",X"EF",X"AF",X"77",X"E1",X"F1",X"C9",X"F5",X"E5",X"21",
		X"AA",X"EF",X"34",X"7E",X"FE",X"02",X"20",X"40",X"AF",X"77",X"21",X"AB",X"EF",X"34",X"7E",X"FE",
		X"01",X"28",X"12",X"FE",X"02",X"28",X"15",X"FE",X"03",X"28",X"18",X"FE",X"04",X"28",X"1B",X"FE",
		X"05",X"28",X"1E",X"18",X"23",X"3E",X"00",X"32",X"A9",X"EF",X"18",X"1C",X"3E",X"08",X"32",X"A9",
		X"EF",X"18",X"15",X"3E",X"18",X"32",X"A9",X"EF",X"18",X"0E",X"3E",X"20",X"32",X"A9",X"EF",X"18",
		X"07",X"3E",X"28",X"32",X"A9",X"EF",X"AF",X"77",X"E1",X"F1",X"C9",X"06",X"FF",X"D6",X"0A",X"04",
		X"30",X"FB",X"C6",X"0A",X"4F",X"C5",X"3E",X"30",X"81",X"4F",X"FD",X"71",X"C1",X"FD",X"36",X"C0",
		X"00",X"C1",X"48",X"79",X"FE",X"00",X"C8",X"3E",X"30",X"81",X"4F",X"FD",X"71",X"01",X"FD",X"36",
		X"00",X"00",X"C9",X"C5",X"E5",X"D5",X"06",X"03",X"CD",X"67",X"A5",X"FE",X"02",X"20",X"04",X"13",
		X"23",X"10",X"F5",X"D1",X"E1",X"C1",X"C9",X"1A",X"BE",X"3E",X"00",X"28",X"03",X"30",X"02",X"C9",
		X"3C",X"3C",X"C9",X"79",X"06",X"05",X"3E",X"0A",X"CD",X"AE",X"67",X"3E",X"07",X"F7",X"E7",X"E7",
		X"AF",X"32",X"EF",X"EF",X"CD",X"17",X"21",X"CD",X"D0",X"21",X"3E",X"01",X"32",X"D5",X"C4",X"CD",
		X"D9",X"A5",X"CD",X"35",X"A6",X"CD",X"3F",X"A6",X"CD",X"4B",X"A6",X"3E",X"14",X"DF",X"CD",X"9E",
		X"A7",X"3E",X"07",X"CF",X"E7",X"C9",X"06",X"05",X"3E",X"07",X"F7",X"E7",X"CD",X"D9",X"A5",X"CD",
		X"D0",X"21",X"3E",X"01",X"32",X"EE",X"EF",X"32",X"EF",X"EF",X"CD",X"35",X"A6",X"CD",X"45",X"A6",
		X"CD",X"BE",X"AA",X"CD",X"A8",X"AA",X"CD",X"64",X"A6",X"3E",X"14",X"DF",X"CD",X"9E",X"A7",X"3E",
		X"01",X"32",X"D5",X"C4",X"3E",X"07",X"CF",X"E7",X"C9",X"3A",X"7B",X"C4",X"CB",X"F7",X"CB",X"EF",
		X"32",X"7B",X"C4",X"AF",X"32",X"B3",X"EF",X"32",X"B4",X"EF",X"32",X"B0",X"EF",X"32",X"B1",X"EF",
		X"32",X"B2",X"EF",X"32",X"ED",X"EF",X"32",X"EE",X"EF",X"32",X"B5",X"EF",X"32",X"B6",X"EF",X"32",
		X"B7",X"EF",X"32",X"B8",X"EF",X"32",X"B9",X"EF",X"32",X"BA",X"EF",X"32",X"BB",X"EF",X"32",X"BC",
		X"EF",X"32",X"E4",X"EF",X"32",X"E5",X"EF",X"32",X"E6",X"EF",X"32",X"E7",X"EF",X"32",X"E8",X"EF",
		X"32",X"E9",X"EF",X"32",X"EA",X"EF",X"32",X"EB",X"EF",X"32",X"EC",X"EF",X"32",X"F2",X"EF",X"3E",
		X"45",X"32",X"F1",X"EF",X"C9",X"CD",X"5E",X"A8",X"CD",X"E8",X"A9",X"CD",X"6D",X"A8",X"C9",X"3E",
		X"01",X"32",X"00",X"EC",X"C9",X"3E",X"04",X"32",X"F0",X"EF",X"C9",X"CD",X"A3",X"A6",X"CD",X"E9",
		X"A6",X"CD",X"74",X"A7",X"3A",X"B3",X"EF",X"FE",X"1B",X"C8",X"3A",X"ED",X"EF",X"FE",X"01",X"3E",
		X"01",X"DF",X"18",X"E7",X"3A",X"00",X"EC",X"FE",X"00",X"20",X"1C",X"3A",X"F0",X"EF",X"FE",X"07",
		X"28",X"15",X"21",X"F1",X"EF",X"34",X"3E",X"50",X"BE",X"20",X"0C",X"AF",X"77",X"3A",X"F0",X"EF",
		X"32",X"00",X"EC",X"3C",X"32",X"F0",X"EF",X"CD",X"C5",X"A6",X"CD",X"22",X"A7",X"CD",X"5B",X"A7",
		X"CD",X"74",X"A7",X"3A",X"ED",X"EF",X"FE",X"01",X"3A",X"B3",X"EF",X"FE",X"38",X"C8",X"3E",X"01",
		X"DF",X"18",X"C1",X"3A",X"B0",X"EF",X"47",X"3A",X"B3",X"EF",X"3A",X"B3",X"EF",X"FE",X"03",X"20",
		X"02",X"CB",X"D0",X"3A",X"B3",X"EF",X"FE",X"00",X"20",X"06",X"CB",X"E0",X"AF",X"32",X"E6",X"EF",
		X"78",X"32",X"B0",X"EF",X"C9",X"3A",X"B1",X"EF",X"47",X"3A",X"B3",X"EF",X"FE",X"00",X"20",X"02",
		X"CB",X"F0",X"3A",X"B3",X"EF",X"FE",X"02",X"20",X"02",X"CB",X"D0",X"3A",X"B3",X"EF",X"FE",X"10",
		X"20",X"02",X"CB",X"E8",X"78",X"32",X"B1",X"EF",X"C9",X"3A",X"B0",X"EF",X"CB",X"47",X"C4",X"2A",
		X"AB",X"3A",X"B0",X"EF",X"CB",X"4F",X"C4",X"76",X"AE",X"3A",X"B0",X"EF",X"CB",X"57",X"C4",X"26",
		X"BA",X"3A",X"B0",X"EF",X"CB",X"5F",X"C4",X"D1",X"B3",X"3A",X"B0",X"EF",X"CB",X"67",X"C4",X"B0",
		X"A7",X"3A",X"B0",X"EF",X"CB",X"6F",X"C4",X"BB",X"AF",X"3A",X"B0",X"EF",X"CB",X"77",X"C4",X"FA",
		X"A9",X"C9",X"3A",X"B1",X"EF",X"CB",X"47",X"C4",X"2A",X"AB",X"3A",X"B1",X"EF",X"CB",X"4F",X"C4",
		X"76",X"AE",X"3A",X"B1",X"EF",X"CB",X"57",X"C4",X"26",X"BA",X"3A",X"B1",X"EF",X"CB",X"5F",X"C4",
		X"D1",X"B3",X"3A",X"B1",X"EF",X"CB",X"67",X"C4",X"B0",X"A7",X"3A",X"B1",X"EF",X"CB",X"6F",X"C4",
		X"BB",X"AF",X"3A",X"B1",X"EF",X"CB",X"77",X"C4",X"FA",X"A9",X"C9",X"3A",X"B2",X"EF",X"CB",X"47",
		X"C4",X"B2",X"AB",X"3A",X"B2",X"EF",X"CB",X"4F",X"C4",X"D5",X"AB",X"3A",X"B2",X"EF",X"CB",X"57",
		X"C4",X"76",X"AC",X"C9",X"3A",X"EE",X"EF",X"FE",X"01",X"28",X"0C",X"3A",X"B4",X"EF",X"3C",X"32",
		X"B4",X"EF",X"FE",X"10",X"C0",X"18",X"0A",X"3A",X"B4",X"EF",X"3C",X"32",X"B4",X"EF",X"FE",X"10",
		X"C0",X"3E",X"00",X"32",X"B4",X"EF",X"3A",X"B3",X"EF",X"3C",X"32",X"B3",X"EF",X"C9",X"CD",X"17",
		X"21",X"CD",X"D0",X"21",X"3A",X"7B",X"C4",X"CB",X"B7",X"CB",X"AF",X"32",X"7B",X"C4",X"E7",X"C9",
		X"3A",X"E6",X"EF",X"FE",X"00",X"20",X"09",X"3E",X"04",X"32",X"BB",X"EF",X"21",X"E6",X"EF",X"34",
		X"21",X"BB",X"EF",X"35",X"7E",X"FE",X"02",X"28",X"0D",X"FE",X"00",X"28",X"01",X"C9",X"36",X"04",
		X"DD",X"21",X"30",X"A8",X"18",X"04",X"DD",X"21",X"02",X"A8",X"21",X"E6",X"EF",X"34",X"DD",X"7E",
		X"00",X"FE",X"FF",X"C8",X"11",X"00",X"E0",X"DD",X"66",X"00",X"DD",X"6E",X"01",X"19",X"DD",X"7E",
		X"02",X"07",X"07",X"07",X"47",X"7E",X"E6",X"07",X"B0",X"77",X"DD",X"23",X"DD",X"23",X"DD",X"23",
		X"18",X"DC",X"04",X"34",X"1D",X"04",X"36",X"1D",X"04",X"38",X"1D",X"04",X"6E",X"1D",X"04",X"70",
		X"1D",X"05",X"6E",X"1D",X"05",X"AE",X"1D",X"06",X"F0",X"1D",X"06",X"F2",X"1D",X"06",X"F4",X"1D",
		X"06",X"F6",X"1D",X"07",X"30",X"1D",X"07",X"32",X"1D",X"07",X"34",X"1D",X"07",X"36",X"1D",X"FF",
		X"04",X"34",X"17",X"04",X"36",X"17",X"04",X"38",X"17",X"04",X"6E",X"17",X"04",X"70",X"17",X"05",
		X"6E",X"17",X"05",X"AE",X"17",X"06",X"F0",X"17",X"06",X"F2",X"17",X"06",X"F4",X"17",X"06",X"F6",
		X"17",X"07",X"30",X"17",X"07",X"32",X"17",X"07",X"34",X"17",X"07",X"36",X"17",X"FF",X"21",X"E0",
		X"57",X"CD",X"D1",X"20",X"22",X"C6",X"EF",X"DD",X"21",X"B0",X"A8",X"18",X"0F",X"21",X"E0",X"57",
		X"CD",X"D1",X"20",X"22",X"C6",X"EF",X"DD",X"21",X"DA",X"A8",X"18",X"00",X"DD",X"56",X"04",X"DD",
		X"5E",X"05",X"7A",X"FE",X"FF",X"C8",X"2A",X"C6",X"EF",X"19",X"3E",X"E0",X"DD",X"46",X"02",X"DD",
		X"4E",X"03",X"E5",X"21",X"00",X"E0",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"19",X"EB",X"E1",X"CD",
		X"55",X"22",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",X"CC",
		X"00",X"84",X"0C",X"0C",X"00",X"00",X"03",X"84",X"0C",X"0C",X"00",X"00",X"06",X"84",X"0C",X"04",
		X"00",X"00",X"00",X"9C",X"0C",X"0C",X"00",X"00",X"03",X"9C",X"0C",X"0C",X"00",X"00",X"06",X"9C",
		X"0C",X"04",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"B4",X"06",X"01",X"00",X"00",
		X"00",X"F4",X"06",X"01",X"00",X"0C",X"01",X"34",X"06",X"01",X"00",X"18",X"01",X"72",X"01",X"01",
		X"00",X"2F",X"01",X"74",X"06",X"01",X"00",X"24",X"01",X"B2",X"01",X"01",X"00",X"3B",X"01",X"B4",
		X"06",X"01",X"00",X"30",X"01",X"F4",X"06",X"01",X"00",X"3C",X"02",X"34",X"06",X"01",X"00",X"48",
		X"02",X"76",X"05",X"01",X"00",X"55",X"02",X"B6",X"05",X"01",X"00",X"61",X"02",X"FC",X"02",X"01",
		X"00",X"70",X"03",X"3C",X"02",X"01",X"00",X"7C",X"03",X"7A",X"03",X"01",X"00",X"87",X"03",X"BA",
		X"03",X"01",X"00",X"03",X"03",X"FA",X"03",X"01",X"00",X"0F",X"04",X"3C",X"02",X"01",X"00",X"1C",
		X"04",X"7A",X"03",X"01",X"00",X"27",X"04",X"B6",X"05",X"01",X"00",X"31",X"04",X"F8",X"04",X"01",
		X"00",X"3E",X"05",X"38",X"04",X"01",X"00",X"4A",X"05",X"78",X"04",X"01",X"00",X"56",X"05",X"B6",
		X"05",X"01",X"00",X"61",X"05",X"F6",X"05",X"01",X"00",X"6D",X"06",X"36",X"05",X"01",X"00",X"79",
		X"06",X"76",X"05",X"01",X"00",X"85",X"06",X"B6",X"05",X"01",X"00",X"01",X"06",X"F8",X"04",X"01",
		X"00",X"0E",X"07",X"38",X"04",X"01",X"00",X"1A",X"07",X"74",X"06",X"01",X"00",X"24",X"01",X"66",
		X"01",X"01",X"00",X"29",X"01",X"A6",X"02",X"01",X"00",X"35",X"01",X"E6",X"01",X"01",X"00",X"41",
		X"04",X"E6",X"01",X"01",X"00",X"35",X"04",X"A6",X"01",X"01",X"00",X"41",X"05",X"26",X"01",X"01",
		X"00",X"4D",X"05",X"66",X"01",X"01",X"00",X"59",X"05",X"A6",X"02",X"01",X"00",X"65",X"05",X"E6",
		X"03",X"01",X"00",X"71",X"06",X"26",X"02",X"01",X"00",X"7D",X"06",X"66",X"03",X"01",X"00",X"89",
		X"06",X"A6",X"03",X"01",X"00",X"05",X"06",X"E6",X"04",X"01",X"00",X"11",X"07",X"26",X"05",X"01",
		X"00",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",X"40",X"43",X"CD",X"D1",X"20",X"3E",X"E8",
		X"11",X"66",X"E1",X"01",X"18",X"0B",X"CD",X"55",X"22",X"C9",X"3A",X"E9",X"EF",X"FE",X"00",X"20",
		X"25",X"CD",X"BE",X"AA",X"DD",X"21",X"9F",X"AA",X"DD",X"22",X"D4",X"EF",X"3E",X"1E",X"32",X"BD",
		X"EF",X"3E",X"0C",X"32",X"D8",X"EF",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"05",X"3E",X"04",X"32",
		X"D8",X"EF",X"21",X"E9",X"EF",X"34",X"21",X"BD",X"EF",X"35",X"7E",X"FE",X"00",X"C0",X"3A",X"D8",
		X"EF",X"77",X"21",X"66",X"E1",X"22",X"D6",X"EF",X"01",X"18",X"0B",X"DD",X"2A",X"D4",X"EF",X"DD",
		X"7E",X"00",X"FE",X"FF",X"20",X"2A",X"DD",X"21",X"9F",X"AA",X"3A",X"EE",X"EF",X"FE",X"01",X"28",
		X"0D",X"3A",X"D8",X"EF",X"3D",X"FE",X"06",X"38",X"11",X"32",X"D8",X"EF",X"18",X"12",X"3A",X"D8",
		X"EF",X"3C",X"FE",X"0C",X"D0",X"32",X"D8",X"EF",X"18",X"06",X"3E",X"01",X"32",X"ED",X"EF",X"C9",
		X"C5",X"DD",X"7E",X"00",X"07",X"07",X"07",X"47",X"7E",X"E6",X"07",X"B0",X"77",X"23",X"23",X"C1",
		X"10",X"EE",X"2A",X"D6",X"EF",X"11",X"40",X"00",X"19",X"22",X"D6",X"EF",X"06",X"0B",X"0D",X"20",
		X"DF",X"DD",X"23",X"DD",X"22",X"D4",X"EF",X"C5",X"D5",X"CD",X"6D",X"A8",X"D1",X"C1",X"C9",X"13",
		X"14",X"15",X"16",X"15",X"14",X"13",X"1D",X"FF",X"21",X"80",X"4B",X"CD",X"D1",X"20",X"11",X"A8",
		X"00",X"19",X"11",X"68",X"E3",X"3E",X"E8",X"01",X"06",X"04",X"CD",X"55",X"22",X"C9",X"DD",X"21",
		X"EA",X"AA",X"21",X"60",X"5C",X"CD",X"D1",X"20",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",X"DD",X"56",
		X"02",X"DD",X"5E",X"03",X"19",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"1E",X"1D",X"CD",X"D3",X"BD",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",X"D8",X"04",X"34",X"00",X"01",X"04",X"36",
		X"00",X"02",X"04",X"38",X"00",X"03",X"04",X"6E",X"00",X"05",X"04",X"70",X"00",X"06",X"05",X"6E",
		X"00",X"00",X"05",X"AE",X"00",X"04",X"06",X"F0",X"00",X"08",X"06",X"F2",X"00",X"09",X"06",X"F4",
		X"00",X"0A",X"06",X"F6",X"00",X"0B",X"07",X"30",X"00",X"0C",X"07",X"32",X"00",X"0D",X"07",X"34",
		X"00",X"0E",X"07",X"36",X"00",X"0F",X"FF",X"FF",X"FF",X"FF",X"3A",X"E5",X"EF",X"FE",X"09",X"20",
		X"25",X"3A",X"B0",X"EF",X"CB",X"87",X"CB",X"F7",X"CB",X"A7",X"32",X"B0",X"EF",X"3A",X"EE",X"EF",
		X"FE",X"01",X"C0",X"3A",X"B1",X"EF",X"CB",X"E7",X"CB",X"87",X"CB",X"B7",X"32",X"B1",X"EF",X"CD",
		X"E8",X"A9",X"CD",X"6D",X"A8",X"C9",X"3A",X"E5",X"EF",X"FE",X"00",X"20",X"1D",X"3E",X"03",X"32",
		X"B6",X"EF",X"21",X"80",X"4B",X"CD",X"D1",X"20",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"04",X"11",
		X"A8",X"00",X"19",X"22",X"BE",X"EF",X"21",X"E5",X"EF",X"34",X"3A",X"B6",X"EF",X"3D",X"32",X"B6",
		X"EF",X"FE",X"00",X"C0",X"3E",X"03",X"32",X"B6",X"EF",X"21",X"E5",X"EF",X"34",X"2A",X"BE",X"EF",
		X"11",X"68",X"E3",X"3E",X"E8",X"01",X"06",X"04",X"CD",X"55",X"22",X"EB",X"3A",X"EE",X"EF",X"FE",
		X"01",X"20",X"0B",X"E5",X"CD",X"BE",X"AA",X"E1",X"11",X"30",X"00",X"B7",X"ED",X"52",X"22",X"BE",
		X"EF",X"C9",X"3A",X"EB",X"EF",X"FE",X"00",X"20",X"3D",X"3E",X"05",X"32",X"B7",X"EF",X"21",X"80",
		X"51",X"CD",X"D1",X"20",X"22",X"DA",X"EF",X"21",X"EB",X"EF",X"34",X"DD",X"21",X"55",X"AC",X"DD",
		X"22",X"DC",X"EF",X"18",X"21",X"3A",X"EB",X"EF",X"FE",X"00",X"20",X"1A",X"3E",X"05",X"32",X"B7",
		X"EF",X"21",X"80",X"51",X"CD",X"D1",X"20",X"22",X"DA",X"EF",X"21",X"EB",X"EF",X"34",X"DD",X"21",
		X"64",X"AC",X"DD",X"22",X"DC",X"EF",X"3A",X"B7",X"EF",X"3D",X"32",X"B7",X"EF",X"FE",X"00",X"C0",
		X"DD",X"2A",X"DC",X"EF",X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"0E",X"3A",X"B2",X"EF",X"CB",X"8F",
		X"32",X"B2",X"EF",X"3E",X"01",X"32",X"ED",X"EF",X"C9",X"DD",X"7E",X"00",X"FE",X"EF",X"20",X"0B",
		X"3A",X"B2",X"EF",X"CB",X"87",X"CB",X"D7",X"32",X"B2",X"EF",X"C9",X"DD",X"7E",X"02",X"32",X"B7",
		X"EF",X"21",X"EB",X"EF",X"34",X"2A",X"DA",X"EF",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"19",X"11",
		X"68",X"E3",X"3E",X"E8",X"01",X"06",X"04",X"CD",X"55",X"22",X"DD",X"23",X"DD",X"23",X"DD",X"23",
		X"DD",X"22",X"DC",X"EF",X"C9",X"00",X"18",X"05",X"00",X"30",X"05",X"00",X"48",X"05",X"00",X"60",
		X"0A",X"EF",X"EF",X"FF",X"00",X"60",X"05",X"00",X"48",X"05",X"00",X"30",X"05",X"00",X"18",X"05",
		X"00",X"00",X"78",X"FF",X"FF",X"FF",X"3A",X"EC",X"EF",X"FE",X"00",X"20",X"21",X"3E",X"05",X"32",
		X"B8",X"EF",X"21",X"40",X"60",X"CD",X"BA",X"20",X"22",X"DE",X"EF",X"11",X"36",X"00",X"19",X"22",
		X"E2",X"EF",X"21",X"EC",X"EF",X"34",X"DD",X"21",X"2D",X"AE",X"DD",X"22",X"E0",X"EF",X"3A",X"B8",
		X"EF",X"3D",X"32",X"B8",X"EF",X"FE",X"00",X"C0",X"21",X"EC",X"EF",X"34",X"DD",X"2A",X"E0",X"EF",
		X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"0F",X"3A",X"B2",X"EF",X"CB",X"97",X"CB",X"CF",X"32",X"B2",
		X"EF",X"AF",X"32",X"EB",X"EF",X"C9",X"DD",X"7E",X"03",X"32",X"B8",X"EF",X"DD",X"2A",X"E0",X"EF",
		X"16",X"00",X"DD",X"5E",X"00",X"2A",X"DE",X"EF",X"19",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"1E",
		X"1E",X"3E",X"00",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"DE",X"EF",X"19",X"23",
		X"DD",X"46",X"01",X"DD",X"7E",X"02",X"C6",X"08",X"4F",X"1E",X"1E",X"3E",X"01",X"CD",X"B9",X"BD",
		X"16",X"00",X"DD",X"5E",X"00",X"2A",X"DE",X"EF",X"19",X"23",X"23",X"DD",X"46",X"01",X"DD",X"7E",
		X"02",X"C6",X"10",X"4F",X"1E",X"1E",X"3E",X"02",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",
		X"2A",X"DE",X"EF",X"19",X"23",X"23",X"23",X"DD",X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"4E",X"02",
		X"1E",X"1E",X"3E",X"03",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"DE",X"EF",X"19",
		X"23",X"23",X"23",X"23",X"DD",X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"08",X"4F",
		X"1E",X"1E",X"3E",X"04",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"DE",X"EF",X"19",
		X"23",X"23",X"23",X"23",X"23",X"DD",X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"10",
		X"4F",X"1E",X"1E",X"3E",X"05",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"E2",X"EF",
		X"19",X"DD",X"46",X"01",X"DD",X"4E",X"02",X"1E",X"1E",X"3E",X"0A",X"CD",X"B9",X"BD",X"16",X"00",
		X"DD",X"5E",X"00",X"2A",X"E2",X"EF",X"19",X"23",X"DD",X"46",X"01",X"DD",X"7E",X"02",X"C6",X"08",
		X"4F",X"1E",X"1E",X"3E",X"0B",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"E2",X"EF",
		X"19",X"23",X"23",X"DD",X"46",X"01",X"DD",X"7E",X"02",X"C6",X"10",X"4F",X"1E",X"1E",X"3E",X"0C",
		X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"E2",X"EF",X"19",X"23",X"23",X"23",X"DD",
		X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"4E",X"02",X"1E",X"1E",X"3E",X"0D",X"CD",X"B9",X"BD",X"16",
		X"00",X"DD",X"5E",X"00",X"2A",X"E2",X"EF",X"19",X"23",X"23",X"23",X"23",X"DD",X"7E",X"01",X"C6",
		X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"08",X"4F",X"1E",X"1E",X"3E",X"0E",X"CD",X"B9",X"BD",X"16",
		X"00",X"DD",X"5E",X"00",X"2A",X"E2",X"EF",X"19",X"23",X"23",X"23",X"23",X"23",X"DD",X"7E",X"01",
		X"C6",X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"10",X"4F",X"1E",X"1E",X"3E",X"0F",X"CD",X"B9",X"BD",
		X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"22",X"E0",X"EF",X"C9",X"00",X"80",X"A0",
		X"03",X"06",X"80",X"A0",X"03",X"0C",X"80",X"A0",X"03",X"12",X"80",X"A0",X"03",X"18",X"80",X"A0",
		X"03",X"1E",X"80",X"A0",X"03",X"24",X"80",X"A0",X"03",X"2A",X"80",X"A0",X"03",X"30",X"80",X"A0",
		X"0A",X"2A",X"80",X"A0",X"03",X"24",X"80",X"A0",X"03",X"1E",X"80",X"A0",X"03",X"18",X"80",X"A0",
		X"03",X"12",X"80",X"A0",X"03",X"0C",X"80",X"A0",X"03",X"06",X"80",X"A0",X"03",X"00",X"80",X"A0",
		X"0A",X"00",X"00",X"00",X"01",X"FF",X"3A",X"E7",X"EF",X"FE",X"00",X"20",X"2A",X"3E",X"02",X"32",
		X"00",X"EC",X"3E",X"03",X"32",X"B5",X"EF",X"21",X"E0",X"5C",X"CD",X"BA",X"20",X"22",X"CC",X"EF",
		X"21",X"E7",X"EF",X"34",X"DD",X"21",X"84",X"AF",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"04",X"DD",
		X"21",X"94",X"AF",X"DD",X"22",X"CE",X"EF",X"3A",X"B5",X"EF",X"3D",X"32",X"B5",X"EF",X"FE",X"00",
		X"C0",X"3E",X"03",X"32",X"B5",X"EF",X"21",X"E7",X"EF",X"34",X"DD",X"2A",X"CE",X"EF",X"DD",X"7E",
		X"00",X"FE",X"FF",X"20",X"14",X"3A",X"B0",X"EF",X"CB",X"8F",X"32",X"B0",X"EF",X"3A",X"B1",X"EF",
		X"CB",X"8F",X"32",X"B1",X"EF",X"CD",X"97",X"AF",X"C9",X"DD",X"2A",X"CE",X"EF",X"16",X"00",X"DD",
		X"5E",X"00",X"2A",X"CC",X"EF",X"19",X"3E",X"0B",X"06",X"70",X"0E",X"A4",X"DD",X"5E",X"01",X"CD",
		X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"CC",X"EF",X"19",X"23",X"06",X"70",X"0E",X"AC",
		X"DD",X"5E",X"01",X"3E",X"0C",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"CC",X"EF",
		X"19",X"23",X"23",X"3E",X"0D",X"06",X"70",X"0E",X"B4",X"DD",X"5E",X"01",X"CD",X"B9",X"BD",X"16",
		X"00",X"DD",X"5E",X"00",X"2A",X"CC",X"EF",X"19",X"23",X"23",X"23",X"3E",X"0E",X"06",X"80",X"0E",
		X"A4",X"DD",X"5E",X"01",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"CC",X"EF",X"19",
		X"23",X"23",X"23",X"23",X"3E",X"0F",X"06",X"80",X"0E",X"AC",X"DD",X"5E",X"01",X"CD",X"B9",X"BD",
		X"16",X"00",X"DD",X"5E",X"00",X"2A",X"CC",X"EF",X"19",X"23",X"23",X"23",X"23",X"23",X"3E",X"00",
		X"06",X"80",X"0E",X"B4",X"DD",X"5E",X"01",X"CD",X"B9",X"BD",X"DD",X"23",X"DD",X"23",X"3A",X"EE",
		X"EF",X"FE",X"01",X"20",X"08",X"DD",X"2B",X"DD",X"2B",X"DD",X"2B",X"DD",X"2B",X"DD",X"22",X"CE",
		X"EF",X"C9",X"FF",X"FF",X"00",X"1E",X"06",X"1E",X"0C",X"1E",X"12",X"1E",X"18",X"1E",X"1E",X"1E",
		X"24",X"1E",X"2A",X"1E",X"30",X"1E",X"FF",X"DD",X"21",X"B4",X"AF",X"DD",X"7E",X"00",X"FE",X"FF",
		X"C8",X"11",X"00",X"00",X"21",X"00",X"00",X"DD",X"7E",X"00",X"01",X"00",X"00",X"CD",X"B9",X"BD",
		X"DD",X"23",X"18",X"E7",X"0B",X"0C",X"0D",X"0E",X"0F",X"00",X"FF",X"3A",X"E8",X"EF",X"FE",X"00",
		X"20",X"25",X"3E",X"05",X"32",X"BC",X"EF",X"21",X"C0",X"69",X"CD",X"BA",X"20",X"22",X"D0",X"EF",
		X"21",X"E8",X"EF",X"34",X"DD",X"21",X"D7",X"B0",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"04",X"DD",
		X"21",X"EB",X"B1",X"DD",X"22",X"D2",X"EF",X"3A",X"BC",X"EF",X"3D",X"32",X"BC",X"EF",X"FE",X"00",
		X"C0",X"21",X"E8",X"EF",X"34",X"DD",X"2A",X"D2",X"EF",X"DD",X"7E",X"02",X"FE",X"88",X"20",X"08",
		X"3A",X"B2",X"EF",X"CB",X"C7",X"32",X"B2",X"EF",X"DD",X"2A",X"D2",X"EF",X"3A",X"EE",X"EF",X"FE",
		X"00",X"20",X"1D",X"DD",X"7E",X"01",X"FE",X"60",X"20",X"16",X"3E",X"03",X"32",X"00",X"EC",X"3A",
		X"F2",X"EF",X"FE",X"00",X"20",X"0A",X"3E",X"13",X"CD",X"AE",X"67",X"3E",X"01",X"32",X"F2",X"EF",
		X"DD",X"7E",X"00",X"FE",X"FF",X"20",X"11",X"3A",X"B0",X"EF",X"CB",X"AF",X"32",X"B0",X"EF",X"3A",
		X"B1",X"EF",X"CB",X"AF",X"32",X"B1",X"EF",X"C9",X"DD",X"7E",X"04",X"C6",X"01",X"32",X"BC",X"EF",
		X"DD",X"2A",X"D2",X"EF",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"D0",X"EF",X"19",X"DD",X"46",X"01",
		X"DD",X"4E",X"02",X"DD",X"5E",X"03",X"3E",X"06",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",
		X"2A",X"D0",X"EF",X"19",X"23",X"DD",X"7E",X"01",X"C6",X"00",X"47",X"DD",X"7E",X"02",X"C6",X"08",
		X"4F",X"DD",X"5E",X"03",X"3E",X"07",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"D0",
		X"EF",X"19",X"23",X"23",X"DD",X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"00",X"4F",
		X"DD",X"5E",X"03",X"3E",X"08",X"CD",X"B9",X"BD",X"16",X"00",X"DD",X"5E",X"00",X"2A",X"D0",X"EF",
		X"19",X"23",X"23",X"23",X"DD",X"7E",X"01",X"C6",X"F0",X"47",X"DD",X"7E",X"02",X"C6",X"08",X"4F",
		X"DD",X"5E",X"03",X"3E",X"09",X"CD",X"B9",X"BD",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"DD",X"22",X"D2",X"EF",X"C9",X"00",X"80",X"AC",X"0C",X"01",X"00",X"7F",X"AB",X"0C",
		X"01",X"00",X"7F",X"AB",X"0C",X"01",X"00",X"7E",X"AA",X"0C",X"01",X"00",X"7E",X"A9",X"0C",X"01",
		X"04",X"7D",X"A8",X"0C",X"02",X"04",X"7C",X"A7",X"0C",X"01",X"04",X"7B",X"A6",X"0C",X"01",X"04",
		X"7B",X"A5",X"0C",X"01",X"08",X"7A",X"A4",X"0C",X"01",X"08",X"7A",X"A4",X"0C",X"01",X"08",X"7A",
		X"A3",X"0C",X"01",X"08",X"79",X"A3",X"0C",X"02",X"0C",X"78",X"A2",X"0C",X"02",X"0C",X"78",X"A1",
		X"0C",X"02",X"0C",X"77",X"A0",X"0C",X"01",X"0C",X"77",X"9F",X"0C",X"01",X"10",X"76",X"9E",X"0C",
		X"02",X"10",X"75",X"9D",X"0C",X"02",X"10",X"74",X"9C",X"0C",X"01",X"10",X"74",X"9B",X"0C",X"01",
		X"14",X"73",X"9A",X"0C",X"02",X"14",X"72",X"99",X"0C",X"02",X"14",X"71",X"98",X"0C",X"02",X"14",
		X"71",X"97",X"0C",X"01",X"18",X"70",X"96",X"0C",X"04",X"18",X"6F",X"95",X"0C",X"03",X"1C",X"6E",
		X"94",X"0C",X"02",X"1C",X"6D",X"93",X"0C",X"02",X"1C",X"6C",X"92",X"0C",X"02",X"1C",X"6C",X"91",
		X"0C",X"02",X"20",X"6B",X"8F",X"0C",X"02",X"20",X"6B",X"8E",X"0C",X"03",X"20",X"6A",X"8D",X"0C",
		X"03",X"24",X"69",X"8C",X"0C",X"04",X"24",X"68",X"8B",X"0C",X"04",X"28",X"67",X"8A",X"0C",X"02",
		X"28",X"67",X"89",X"0C",X"03",X"28",X"66",X"88",X"0C",X"03",X"2C",X"65",X"87",X"0C",X"04",X"2C",
		X"65",X"86",X"0C",X"05",X"30",X"64",X"85",X"0C",X"0A",X"34",X"63",X"84",X"0C",X"0B",X"38",X"62",
		X"82",X"0C",X"0C",X"00",X"00",X"00",X"0C",X"20",X"3C",X"60",X"80",X"0C",X"03",X"40",X"60",X"80",
		X"0C",X"03",X"44",X"60",X"80",X"0C",X"03",X"48",X"60",X"80",X"0C",X"03",X"4C",X"60",X"80",X"0C",
		X"06",X"48",X"60",X"80",X"0C",X"03",X"44",X"60",X"80",X"0C",X"03",X"40",X"60",X"80",X"0C",X"03",
		X"3C",X"60",X"80",X"0C",X"03",X"00",X"00",X"00",X"00",X"03",X"FF",X"3C",X"80",X"58",X"0C",X"03",
		X"40",X"80",X"58",X"0C",X"03",X"44",X"80",X"58",X"0C",X"03",X"48",X"80",X"58",X"0C",X"03",X"4C",
		X"80",X"58",X"0C",X"06",X"48",X"80",X"58",X"0C",X"03",X"44",X"80",X"58",X"0C",X"03",X"40",X"80",
		X"58",X"0C",X"03",X"3C",X"80",X"58",X"0C",X"03",X"00",X"00",X"00",X"0C",X"1E",X"50",X"80",X"58",
		X"0C",X"05",X"54",X"80",X"58",X"0C",X"05",X"58",X"80",X"58",X"0C",X"05",X"5C",X"80",X"58",X"0C",
		X"05",X"60",X"80",X"58",X"0C",X"05",X"64",X"80",X"58",X"0C",X"28",X"64",X"80",X"59",X"0C",X"01",
		X"64",X"80",X"5A",X"0C",X"01",X"64",X"80",X"5B",X"0C",X"01",X"64",X"80",X"5C",X"0C",X"01",X"64",
		X"80",X"5D",X"0C",X"01",X"64",X"80",X"5E",X"0C",X"01",X"64",X"80",X"5F",X"0C",X"01",X"64",X"80",
		X"60",X"0C",X"01",X"64",X"80",X"61",X"0C",X"01",X"64",X"80",X"62",X"0C",X"01",X"64",X"80",X"63",
		X"0C",X"01",X"64",X"80",X"64",X"0C",X"01",X"64",X"80",X"65",X"0C",X"01",X"64",X"80",X"66",X"0C",
		X"01",X"64",X"80",X"67",X"0C",X"01",X"64",X"80",X"68",X"0C",X"01",X"64",X"80",X"69",X"0C",X"01",
		X"64",X"80",X"6A",X"0C",X"01",X"64",X"80",X"6B",X"0C",X"01",X"64",X"80",X"6C",X"0C",X"01",X"64",
		X"80",X"6D",X"0C",X"01",X"64",X"80",X"6E",X"0C",X"01",X"64",X"80",X"6F",X"0C",X"01",X"64",X"80",
		X"70",X"0C",X"01",X"64",X"80",X"71",X"0C",X"01",X"64",X"80",X"72",X"0C",X"01",X"64",X"80",X"73",
		X"0C",X"01",X"64",X"80",X"74",X"0C",X"01",X"64",X"80",X"75",X"0C",X"01",X"64",X"80",X"76",X"0C",
		X"01",X"64",X"80",X"77",X"0C",X"01",X"64",X"80",X"78",X"0C",X"01",X"64",X"80",X"79",X"0C",X"01",
		X"64",X"80",X"7A",X"0C",X"01",X"64",X"80",X"7B",X"0C",X"01",X"64",X"80",X"7C",X"0C",X"01",X"64",
		X"80",X"7D",X"0C",X"01",X"64",X"80",X"7E",X"0C",X"01",X"64",X"80",X"7F",X"0C",X"01",X"64",X"80",
		X"80",X"0C",X"01",X"64",X"80",X"81",X"0C",X"01",X"64",X"80",X"82",X"0C",X"01",X"64",X"80",X"83",
		X"0C",X"01",X"64",X"80",X"84",X"0C",X"01",X"64",X"80",X"85",X"0C",X"01",X"64",X"80",X"86",X"0C",
		X"01",X"64",X"80",X"87",X"0C",X"01",X"64",X"80",X"88",X"0C",X"01",X"64",X"80",X"89",X"0C",X"01",
		X"64",X"80",X"8A",X"0C",X"01",X"64",X"80",X"8B",X"0C",X"01",X"64",X"80",X"8C",X"0C",X"01",X"64",
		X"80",X"8D",X"0C",X"01",X"64",X"80",X"8E",X"0C",X"01",X"64",X"80",X"8F",X"0C",X"01",X"64",X"80",
		X"90",X"0C",X"01",X"64",X"80",X"91",X"0C",X"01",X"64",X"80",X"92",X"0C",X"01",X"64",X"80",X"93",
		X"0C",X"01",X"64",X"80",X"94",X"0C",X"01",X"64",X"80",X"95",X"0C",X"01",X"64",X"80",X"96",X"0C",
		X"01",X"64",X"80",X"97",X"0C",X"01",X"64",X"80",X"98",X"0C",X"01",X"64",X"80",X"99",X"0C",X"01",
		X"64",X"80",X"9A",X"0C",X"01",X"64",X"80",X"9B",X"0C",X"01",X"64",X"80",X"9C",X"0C",X"01",X"64",
		X"80",X"9D",X"0C",X"01",X"64",X"80",X"9E",X"0C",X"01",X"64",X"80",X"9F",X"0C",X"01",X"64",X"80",
		X"A0",X"0C",X"01",X"64",X"80",X"A1",X"0C",X"01",X"64",X"80",X"A2",X"0C",X"01",X"64",X"80",X"A3",
		X"0C",X"01",X"64",X"80",X"A4",X"0C",X"01",X"64",X"80",X"A5",X"0C",X"01",X"64",X"80",X"A6",X"0C",
		X"01",X"64",X"80",X"A7",X"0C",X"01",X"64",X"80",X"A8",X"0C",X"01",X"00",X"00",X"00",X"00",X"03",
		X"FF",X"3A",X"E4",X"EF",X"FE",X"06",X"20",X"0A",X"3A",X"B0",X"EF",X"CB",X"C7",X"CB",X"CF",X"32",
		X"B0",X"EF",X"3A",X"E4",X"EF",X"FE",X"00",X"20",X"0E",X"3E",X"01",X"32",X"BA",X"EF",X"21",X"40",
		X"55",X"CD",X"D1",X"20",X"22",X"C8",X"EF",X"21",X"BA",X"EF",X"35",X"C0",X"36",X"01",X"3A",X"EE",
		X"EF",X"FE",X"01",X"28",X"29",X"3A",X"E4",X"EF",X"FE",X"07",X"CC",X"60",X"B9",X"3A",X"E4",X"EF",
		X"FE",X"08",X"CC",X"66",X"B9",X"3A",X"E4",X"EF",X"FE",X"0E",X"20",X"3A",X"CD",X"6C",X"B9",X"3A",
		X"B0",X"EF",X"CB",X"9F",X"CB",X"EF",X"32",X"B0",X"EF",X"AF",X"32",X"E8",X"EF",X"C9",X"3A",X"E4",
		X"EF",X"FE",X"00",X"CC",X"66",X"B9",X"3A",X"E4",X"EF",X"FE",X"07",X"CC",X"60",X"B9",X"3A",X"E4",
		X"EF",X"FE",X"08",X"CC",X"6C",X"B9",X"3A",X"E4",X"EF",X"FE",X"0F",X"20",X"09",X"3A",X"B1",X"EF",
		X"CB",X"9F",X"32",X"B1",X"EF",X"C9",X"3A",X"E4",X"EF",X"87",X"21",X"A8",X"B4",X"5F",X"16",X"00",
		X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"08",X"21",X"C2",X"B4",X"B7",X"ED",X"52",X"18",X"01",X"19",
		X"5E",X"23",X"56",X"D5",X"DD",X"E1",X"21",X"E4",X"EF",X"34",X"DD",X"7E",X"00",X"FE",X"FF",X"C8",
		X"2A",X"C8",X"EF",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"19",X"DD",X"46",X"02",X"DD",X"4E",X"03",
		X"DD",X"5E",X"04",X"DD",X"E5",X"CD",X"D3",X"BD",X"DD",X"E1",X"DD",X"23",X"DD",X"23",X"DD",X"23",
		X"DD",X"23",X"DD",X"23",X"18",X"D4",X"C4",X"B4",X"D4",X"B4",X"F3",X"B4",X"1C",X"B5",X"59",X"B5",
		X"A5",X"B5",X"19",X"B6",X"92",X"B6",X"0B",X"B7",X"84",X"B7",X"FD",X"B7",X"67",X"B8",X"C2",X"B8",
		X"0E",X"B9",X"4B",X"B9",X"00",X"28",X"01",X"98",X"1C",X"00",X"29",X"01",X"58",X"1C",X"00",X"2A",
		X"01",X"18",X"1C",X"FF",X"00",X"00",X"01",X"98",X"0E",X"00",X"01",X"01",X"58",X"0E",X"00",X"02",
		X"01",X"18",X"0E",X"00",X"2B",X"01",X"DA",X"1C",X"00",X"41",X"01",X"9A",X"1C",X"00",X"42",X"01",
		X"5A",X"1C",X"FF",X"00",X"03",X"01",X"98",X"0E",X"00",X"04",X"01",X"58",X"0E",X"00",X"05",X"01",
		X"18",X"0E",X"00",X"06",X"01",X"9A",X"0E",X"00",X"07",X"01",X"5A",X"0E",X"00",X"2B",X"01",X"DA",
		X"1C",X"00",X"44",X"01",X"DC",X"1C",X"00",X"45",X"01",X"9C",X"1C",X"FF",X"00",X"03",X"01",X"98",
		X"0E",X"00",X"04",X"01",X"58",X"0E",X"00",X"05",X"01",X"18",X"0E",X"00",X"08",X"01",X"DA",X"0E",
		X"00",X"09",X"01",X"9A",X"0E",X"00",X"0A",X"01",X"5A",X"0E",X"00",X"0B",X"01",X"DC",X"0E",X"00",
		X"0C",X"01",X"9C",X"0E",X"00",X"43",X"02",X"1C",X"1C",X"00",X"46",X"02",X"5E",X"1C",X"00",X"47",
		X"02",X"1E",X"1C",X"00",X"48",X"01",X"DE",X"1C",X"FF",X"00",X"03",X"01",X"98",X"0E",X"00",X"04",
		X"01",X"58",X"0E",X"00",X"05",X"01",X"18",X"0E",X"00",X"08",X"01",X"DA",X"0E",X"00",X"09",X"01",
		X"9A",X"0E",X"00",X"0A",X"01",X"5A",X"0E",X"00",X"0D",X"02",X"1C",X"0E",X"00",X"0E",X"01",X"DC",
		X"0E",X"00",X"0F",X"01",X"9C",X"0E",X"00",X"10",X"02",X"5E",X"0E",X"00",X"11",X"02",X"1E",X"0E",
		X"00",X"12",X"01",X"DE",X"0E",X"00",X"4A",X"02",X"A0",X"1C",X"00",X"4B",X"02",X"60",X"1C",X"00",
		X"4C",X"02",X"20",X"1C",X"FF",X"00",X"03",X"01",X"98",X"0E",X"00",X"04",X"01",X"58",X"0E",X"00",
		X"05",X"01",X"18",X"0E",X"00",X"08",X"01",X"DA",X"0E",X"00",X"09",X"01",X"9A",X"0E",X"00",X"0A",
		X"01",X"5A",X"0E",X"00",X"0D",X"02",X"1C",X"0E",X"00",X"0E",X"01",X"DC",X"0E",X"00",X"0F",X"01",
		X"9C",X"0E",X"00",X"13",X"02",X"5E",X"0E",X"00",X"14",X"02",X"1E",X"0E",X"00",X"15",X"01",X"DE",
		X"0E",X"00",X"16",X"02",X"A0",X"0E",X"00",X"17",X"02",X"60",X"0E",X"00",X"18",X"02",X"20",X"0E",
		X"00",X"49",X"02",X"E0",X"1C",X"00",X"4D",X"03",X"22",X"1C",X"00",X"4E",X"02",X"E2",X"1C",X"00",
		X"4F",X"02",X"A2",X"1C",X"00",X"50",X"02",X"62",X"1C",X"00",X"52",X"03",X"24",X"1C",X"00",X"53",
		X"02",X"E4",X"1C",X"00",X"53",X"02",X"A4",X"1C",X"FF",X"00",X"03",X"01",X"98",X"0E",X"00",X"04",
		X"01",X"58",X"0E",X"00",X"05",X"01",X"18",X"0E",X"00",X"08",X"01",X"DA",X"0E",X"00",X"09",X"01",
		X"9A",X"0E",X"00",X"0A",X"01",X"5A",X"0E",X"00",X"0D",X"02",X"1C",X"0E",X"00",X"0E",X"01",X"DC",
		X"0E",X"00",X"0F",X"01",X"9C",X"0E",X"00",X"13",X"02",X"5E",X"0E",X"00",X"14",X"02",X"1E",X"0E",
		X"00",X"15",X"01",X"DE",X"0E",X"00",X"19",X"02",X"E0",X"0E",X"00",X"1A",X"02",X"A0",X"0E",X"00",
		X"1B",X"02",X"60",X"0E",X"00",X"1C",X"02",X"20",X"0E",X"00",X"1D",X"03",X"22",X"0E",X"00",X"1E",
		X"02",X"E2",X"0E",X"00",X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",X"62",X"0E",X"00",X"21",X"03",
		X"24",X"0E",X"00",X"22",X"02",X"E4",X"0E",X"00",X"23",X"02",X"A4",X"0E",X"00",X"51",X"03",X"64",
		X"1C",X"FF",X"00",X"03",X"01",X"98",X"0E",X"00",X"04",X"01",X"58",X"0E",X"00",X"05",X"01",X"18",
		X"0E",X"00",X"08",X"01",X"DA",X"0E",X"00",X"09",X"01",X"9A",X"0E",X"00",X"0A",X"01",X"5A",X"0E",
		X"00",X"0D",X"02",X"1C",X"0E",X"00",X"0E",X"01",X"DC",X"0E",X"00",X"0F",X"01",X"9C",X"0E",X"00",
		X"13",X"02",X"5E",X"0E",X"00",X"14",X"02",X"1E",X"0E",X"00",X"15",X"01",X"DE",X"0E",X"00",X"19",
		X"02",X"E0",X"0E",X"00",X"1A",X"02",X"A0",X"0E",X"00",X"1B",X"02",X"60",X"0E",X"00",X"1C",X"02",
		X"20",X"0E",X"00",X"1D",X"03",X"22",X"0E",X"00",X"1E",X"02",X"E2",X"0E",X"00",X"1F",X"02",X"A2",
		X"0E",X"00",X"20",X"02",X"62",X"0E",X"00",X"24",X"03",X"64",X"0E",X"00",X"25",X"03",X"24",X"0E",
		X"00",X"26",X"02",X"E4",X"0E",X"00",X"27",X"02",X"A4",X"0E",X"FF",X"00",X"08",X"01",X"DA",X"0E",
		X"00",X"09",X"01",X"9A",X"0E",X"00",X"0A",X"01",X"5A",X"0E",X"00",X"0D",X"02",X"1C",X"0E",X"00",
		X"0E",X"01",X"DC",X"0E",X"00",X"0F",X"01",X"9C",X"0E",X"00",X"13",X"02",X"5E",X"0E",X"00",X"14",
		X"02",X"1E",X"0E",X"00",X"15",X"01",X"DE",X"0E",X"00",X"19",X"02",X"E0",X"0E",X"00",X"1A",X"02",
		X"A0",X"0E",X"00",X"1B",X"02",X"60",X"0E",X"00",X"1C",X"02",X"20",X"0E",X"00",X"1D",X"03",X"22",
		X"0E",X"00",X"1E",X"02",X"E2",X"0E",X"00",X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",X"62",X"0E",
		X"00",X"24",X"03",X"64",X"0E",X"00",X"25",X"03",X"24",X"0E",X"00",X"26",X"02",X"E4",X"0E",X"00",
		X"27",X"02",X"A4",X"0E",X"00",X"2D",X"01",X"98",X"0E",X"00",X"2E",X"01",X"58",X"0E",X"00",X"2F",
		X"01",X"18",X"0E",X"FF",X"00",X"28",X"01",X"98",X"1C",X"00",X"29",X"01",X"58",X"1C",X"00",X"2A",
		X"01",X"18",X"1C",X"00",X"0D",X"02",X"1C",X"0E",X"00",X"0E",X"01",X"DC",X"0E",X"00",X"0F",X"01",
		X"9C",X"0E",X"00",X"13",X"02",X"5E",X"0E",X"00",X"14",X"02",X"1E",X"0E",X"00",X"15",X"01",X"DE",
		X"0E",X"00",X"19",X"02",X"E0",X"0E",X"00",X"1A",X"02",X"A0",X"0E",X"00",X"1B",X"02",X"60",X"0E",
		X"00",X"1C",X"02",X"20",X"0E",X"00",X"1D",X"03",X"22",X"0E",X"00",X"1E",X"02",X"E2",X"0E",X"00",
		X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",X"62",X"0E",X"00",X"24",X"03",X"64",X"0E",X"00",X"25",
		X"03",X"24",X"0E",X"00",X"26",X"02",X"E4",X"0E",X"00",X"27",X"02",X"A4",X"0E",X"00",X"30",X"01",
		X"DA",X"0E",X"00",X"31",X"01",X"9A",X"0E",X"00",X"32",X"01",X"5A",X"0E",X"FF",X"00",X"2B",X"01",
		X"DA",X"1C",X"00",X"41",X"01",X"9A",X"1C",X"00",X"42",X"01",X"5A",X"1C",X"00",X"33",X"02",X"1C",
		X"0E",X"00",X"34",X"01",X"DC",X"0E",X"00",X"35",X"01",X"9C",X"0E",X"00",X"13",X"02",X"5E",X"0E",
		X"00",X"14",X"02",X"1E",X"0E",X"00",X"15",X"01",X"DE",X"0E",X"00",X"19",X"02",X"E0",X"0E",X"00",
		X"1A",X"02",X"A0",X"0E",X"00",X"1B",X"02",X"60",X"0E",X"00",X"1C",X"02",X"20",X"0E",X"00",X"1D",
		X"03",X"22",X"0E",X"00",X"1E",X"02",X"E2",X"0E",X"00",X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",
		X"62",X"0E",X"00",X"24",X"03",X"64",X"0E",X"00",X"25",X"03",X"24",X"0E",X"00",X"26",X"02",X"E4",
		X"0E",X"00",X"27",X"02",X"A4",X"0E",X"FF",X"00",X"43",X"02",X"1C",X"1C",X"00",X"44",X"01",X"DC",
		X"1C",X"00",X"45",X"01",X"9C",X"1C",X"00",X"36",X"02",X"5E",X"0E",X"00",X"37",X"02",X"1E",X"0E",
		X"00",X"38",X"01",X"DE",X"0E",X"00",X"19",X"02",X"E0",X"0E",X"00",X"1A",X"02",X"A0",X"0E",X"00",
		X"1B",X"02",X"60",X"0E",X"00",X"1C",X"02",X"20",X"0E",X"00",X"1D",X"03",X"22",X"0E",X"00",X"1E",
		X"02",X"E2",X"0E",X"00",X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",X"62",X"0E",X"00",X"24",X"03",
		X"64",X"0E",X"00",X"25",X"03",X"24",X"0E",X"00",X"26",X"02",X"E4",X"0E",X"00",X"27",X"02",X"A4",
		X"0E",X"FF",X"00",X"46",X"02",X"5E",X"1C",X"00",X"47",X"02",X"1E",X"1C",X"00",X"48",X"01",X"DE",
		X"1C",X"00",X"39",X"02",X"E0",X"0E",X"00",X"3A",X"02",X"A0",X"0E",X"00",X"3B",X"02",X"60",X"0E",
		X"00",X"3C",X"02",X"20",X"0E",X"00",X"1D",X"03",X"22",X"0E",X"00",X"1E",X"02",X"E2",X"0E",X"00",
		X"1F",X"02",X"A2",X"0E",X"00",X"20",X"02",X"62",X"0E",X"00",X"24",X"03",X"64",X"0E",X"00",X"25",
		X"03",X"24",X"0E",X"00",X"26",X"02",X"E4",X"0E",X"00",X"27",X"02",X"A4",X"0E",X"FF",X"00",X"49",
		X"02",X"E0",X"1C",X"00",X"4A",X"02",X"A0",X"1C",X"00",X"4B",X"02",X"60",X"1C",X"00",X"4C",X"02",
		X"20",X"1C",X"00",X"4D",X"03",X"22",X"1C",X"00",X"4E",X"02",X"E2",X"1C",X"00",X"4F",X"02",X"A2",
		X"1C",X"00",X"50",X"02",X"62",X"1C",X"00",X"3D",X"03",X"64",X"0E",X"00",X"3E",X"03",X"24",X"0E",
		X"00",X"3F",X"02",X"E4",X"0E",X"00",X"40",X"02",X"A4",X"0E",X"FF",X"00",X"51",X"03",X"64",X"1C",
		X"00",X"52",X"03",X"24",X"1C",X"00",X"53",X"02",X"E4",X"1C",X"00",X"53",X"02",X"A4",X"1C",X"FF",
		X"DD",X"21",X"9F",X"B9",X"18",X"0C",X"DD",X"21",X"CC",X"B9",X"18",X"06",X"DD",X"21",X"F9",X"B9",
		X"18",X"00",X"DD",X"7E",X"02",X"FE",X"FF",X"C8",X"16",X"00",X"DD",X"5E",X"04",X"21",X"00",X"69",
		X"CD",X"BA",X"20",X"19",X"DD",X"7E",X"03",X"DD",X"46",X"00",X"DD",X"4E",X"01",X"DD",X"5E",X"02",
		X"CD",X"B9",X"BD",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"18",X"D3",X"88",
		X"98",X"0D",X"03",X"00",X"98",X"98",X"0D",X"04",X"01",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"0A",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"98",X"0D",X"03",
		X"02",X"98",X"98",X"0D",X"04",X"03",X"78",X"A0",X"0D",X"05",X"04",X"88",X"A0",X"0D",X"06",X"05",
		X"98",X"A0",X"0D",X"07",X"06",X"78",X"A8",X"0D",X"08",X"07",X"88",X"A8",X"0D",X"09",X"08",X"98",
		X"A8",X"0D",X"0A",X"09",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"3A",X"EA",X"EF",X"FE",X"00",X"20",X"28",X"3E",X"01",X"32",
		X"B9",X"EF",X"DD",X"21",X"20",X"BB",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"04",X"DD",X"21",X"2D",
		X"BD",X"DD",X"22",X"C2",X"EF",X"21",X"00",X"67",X"CD",X"BA",X"20",X"22",X"C4",X"EF",X"3A",X"EA",
		X"EF",X"3C",X"32",X"EA",X"EF",X"3A",X"B9",X"EF",X"3D",X"32",X"B9",X"EF",X"FE",X"00",X"C0",X"3E",
		X"01",X"32",X"B9",X"EF",X"DD",X"2A",X"C2",X"EF",X"DD",X"7E",X"02",X"FE",X"FF",X"20",X"11",X"3A",
		X"B0",X"EF",X"CB",X"97",X"32",X"B0",X"EF",X"3A",X"B1",X"EF",X"CB",X"97",X"32",X"B1",X"EF",X"C9",
		X"DD",X"7E",X"03",X"FE",X"04",X"20",X"08",X"3A",X"B1",X"EF",X"CB",X"C7",X"32",X"B1",X"EF",X"DD",
		X"7E",X"03",X"FE",X"03",X"20",X"08",X"3A",X"B1",X"EF",X"CB",X"CF",X"32",X"B1",X"EF",X"DD",X"7E",
		X"03",X"FE",X"02",X"20",X"08",X"3A",X"B1",X"EF",X"CB",X"DF",X"32",X"B1",X"EF",X"DD",X"7E",X"03",
		X"FE",X"01",X"20",X"08",X"3A",X"B0",X"EF",X"CB",X"DF",X"32",X"B0",X"EF",X"16",X"00",X"DD",X"5E",
		X"04",X"2A",X"C4",X"EF",X"19",X"DD",X"7E",X"00",X"C6",X"08",X"47",X"DD",X"4E",X"01",X"DD",X"5E",
		X"02",X"3E",X"01",X"CD",X"B9",X"BD",X"DD",X"2A",X"C2",X"EF",X"16",X"00",X"DD",X"5E",X"04",X"2A",
		X"C4",X"EF",X"19",X"23",X"DD",X"7E",X"00",X"C6",X"08",X"47",X"DD",X"7E",X"01",X"C6",X"08",X"4F",
		X"DD",X"5E",X"02",X"3E",X"02",X"CD",X"B9",X"BD",X"3A",X"EE",X"EF",X"FE",X"01",X"20",X"0D",X"DD",
		X"E5",X"E1",X"11",X"05",X"00",X"B7",X"ED",X"52",X"22",X"C2",X"EF",X"C9",X"11",X"05",X"00",X"DD",
		X"19",X"DD",X"22",X"C2",X"EF",X"C9",X"FF",X"FF",X"FF",X"00",X"20",X"F8",X"40",X"12",X"00",X"00",
		X"98",X"48",X"12",X"00",X"00",X"99",X"48",X"12",X"00",X"00",X"9A",X"48",X"12",X"00",X"00",X"9B",
		X"48",X"12",X"00",X"00",X"9C",X"49",X"12",X"00",X"00",X"9D",X"49",X"12",X"00",X"00",X"9E",X"49",
		X"12",X"00",X"00",X"9F",X"4A",X"12",X"00",X"00",X"A0",X"4A",X"12",X"00",X"00",X"A1",X"4A",X"12",
		X"00",X"00",X"A2",X"4A",X"12",X"00",X"00",X"A3",X"4B",X"12",X"00",X"00",X"A4",X"4B",X"12",X"00",
		X"00",X"A5",X"4C",X"12",X"00",X"00",X"A6",X"4C",X"12",X"00",X"00",X"A7",X"4D",X"12",X"00",X"00",
		X"A8",X"4D",X"12",X"00",X"02",X"A9",X"4D",X"12",X"00",X"02",X"AA",X"4D",X"12",X"00",X"02",X"AB",
		X"4E",X"12",X"00",X"02",X"AC",X"4E",X"12",X"00",X"02",X"AD",X"4E",X"12",X"00",X"02",X"AE",X"4E",
		X"12",X"00",X"02",X"AF",X"4F",X"12",X"00",X"02",X"B0",X"4F",X"12",X"00",X"02",X"B1",X"4F",X"12",
		X"00",X"02",X"B2",X"50",X"12",X"00",X"02",X"B3",X"50",X"12",X"00",X"02",X"B4",X"50",X"12",X"00",
		X"02",X"B5",X"51",X"12",X"00",X"02",X"B6",X"51",X"12",X"00",X"02",X"B7",X"51",X"12",X"00",X"02",
		X"B8",X"51",X"12",X"00",X"04",X"BA",X"52",X"12",X"00",X"04",X"BC",X"52",X"12",X"00",X"04",X"BE",
		X"53",X"12",X"00",X"04",X"C0",X"54",X"12",X"00",X"06",X"C2",X"55",X"12",X"00",X"06",X"C4",X"56",
		X"12",X"00",X"06",X"C6",X"57",X"12",X"00",X"06",X"C8",X"58",X"12",X"00",X"08",X"CA",X"5A",X"12",
		X"01",X"08",X"CC",X"5C",X"12",X"00",X"08",X"CE",X"5E",X"12",X"00",X"08",X"CF",X"60",X"12",X"00",
		X"08",X"D1",X"62",X"12",X"00",X"08",X"D2",X"64",X"12",X"00",X"08",X"D3",X"66",X"12",X"02",X"08",
		X"D3",X"68",X"12",X"00",X"0A",X"D3",X"6A",X"12",X"00",X"0A",X"D3",X"6D",X"12",X"00",X"0A",X"D2",
		X"70",X"12",X"00",X"0C",X"D1",X"73",X"12",X"00",X"0C",X"D0",X"75",X"12",X"00",X"0C",X"CD",X"78",
		X"12",X"00",X"0E",X"CB",X"7A",X"12",X"03",X"0E",X"C8",X"7C",X"12",X"00",X"0E",X"C6",X"7D",X"12",
		X"00",X"0E",X"C3",X"7F",X"12",X"00",X"0E",X"C0",X"80",X"12",X"00",X"10",X"BE",X"81",X"12",X"04",
		X"10",X"BB",X"82",X"12",X"00",X"10",X"B8",X"82",X"12",X"00",X"10",X"B6",X"83",X"12",X"00",X"10",
		X"B3",X"83",X"12",X"00",X"10",X"B0",X"83",X"12",X"00",X"12",X"AC",X"83",X"12",X"00",X"12",X"A8",
		X"83",X"12",X"00",X"12",X"A4",X"83",X"12",X"00",X"12",X"A0",X"83",X"12",X"00",X"14",X"9C",X"82",
		X"12",X"00",X"14",X"98",X"82",X"12",X"00",X"14",X"94",X"81",X"12",X"00",X"14",X"90",X"80",X"12",
		X"00",X"16",X"8C",X"7F",X"12",X"00",X"16",X"88",X"7E",X"12",X"00",X"16",X"84",X"7D",X"12",X"00",
		X"16",X"80",X"7C",X"12",X"00",X"18",X"7C",X"7A",X"12",X"00",X"18",X"78",X"79",X"12",X"00",X"18",
		X"74",X"78",X"12",X"00",X"18",X"70",X"76",X"12",X"00",X"1A",X"6C",X"75",X"12",X"00",X"1A",X"68",
		X"74",X"12",X"00",X"1A",X"64",X"72",X"12",X"00",X"1A",X"60",X"70",X"12",X"00",X"1C",X"5C",X"6E",
		X"12",X"00",X"1C",X"58",X"6C",X"12",X"00",X"1C",X"54",X"6B",X"12",X"00",X"1C",X"50",X"6A",X"12",
		X"00",X"1E",X"4C",X"68",X"12",X"00",X"1E",X"48",X"66",X"12",X"00",X"1E",X"44",X"64",X"12",X"00",
		X"1E",X"40",X"62",X"12",X"00",X"1E",X"3C",X"60",X"12",X"00",X"1E",X"38",X"5D",X"12",X"00",X"1E",
		X"34",X"5A",X"12",X"00",X"1E",X"30",X"58",X"12",X"00",X"1E",X"2C",X"56",X"12",X"00",X"1E",X"28",
		X"54",X"12",X"00",X"1E",X"24",X"52",X"12",X"00",X"1E",X"20",X"50",X"12",X"00",X"1E",X"1C",X"4C",
		X"12",X"00",X"1E",X"10",X"48",X"12",X"00",X"1E",X"0C",X"44",X"12",X"00",X"1E",X"F8",X"40",X"12",
		X"00",X"00",X"FF",X"FF",X"FF",X"00",X"20",X"11",X"75",X"BD",X"21",X"06",X"E7",X"AF",X"CD",X"F1",
		X"21",X"11",X"8E",X"BD",X"21",X"0A",X"E7",X"AF",X"CD",X"F1",X"21",X"11",X"A9",X"BD",X"21",X"0E",
		X"E7",X"AF",X"CD",X"F1",X"21",X"C9",X"11",X"75",X"BD",X"21",X"06",X"E7",X"AF",X"CD",X"F1",X"21",
		X"11",X"8E",X"BD",X"21",X"0A",X"E7",X"AF",X"CD",X"F1",X"21",X"11",X"A9",X"BD",X"21",X"0E",X"E7",
		X"AF",X"CD",X"F1",X"21",X"C9",X"18",X"4D",X"45",X"53",X"53",X"41",X"47",X"45",X"20",X"49",X"4E",
		X"44",X"49",X"43",X"41",X"54",X"49",X"4F",X"4E",X"20",X"41",X"52",X"45",X"41",X"2E",X"1A",X"43",
		X"4F",X"4D",X"49",X"4E",X"47",X"20",X"53",X"4F",X"4F",X"4E",X"21",X"20",X"4E",X"4F",X"57",X"20",
		X"50",X"52",X"49",X"4E",X"54",X"49",X"4E",X"47",X"21",X"0F",X"57",X"41",X"49",X"54",X"20",X"41",
		X"20",X"4D",X"49",X"4E",X"55",X"54",X"45",X"21",X"21",X"E5",X"D5",X"21",X"7D",X"C4",X"07",X"07",
		X"5F",X"16",X"00",X"19",X"71",X"23",X"70",X"23",X"C1",X"79",X"07",X"07",X"07",X"D1",X"B2",X"77",
		X"23",X"73",X"C9",X"E5",X"21",X"00",X"E0",X"09",X"7B",X"07",X"07",X"07",X"C1",X"B0",X"77",X"23",
		X"71",X"C9",X"DD",X"21",X"7D",X"C4",X"DD",X"36",X"00",X"80",X"DD",X"36",X"01",X"80",X"DD",X"36",
		X"04",X"88",X"DD",X"36",X"05",X"80",X"DD",X"36",X"02",X"02",X"DD",X"36",X"03",X"02",X"DD",X"36",
		X"06",X"02",X"DD",X"36",X"07",X"03",X"DD",X"21",X"F3",X"EF",X"DD",X"36",X"02",X"02",X"DD",X"36",
		X"03",X"04",X"DD",X"36",X"04",X"02",X"01",X"00",X"01",X"C5",X"21",X"7D",X"C4",X"DD",X"21",X"F3",
		X"EF",X"CD",X"4A",X"11",X"E7",X"C1",X"78",X"B1",X"20",X"EF",X"25",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0D",X"0E",X"0D",X"0E",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"11",X"11",
		X"12",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"1A",X"19",X"19",X"19",X"1A",
		X"19",X"19",X"1A",X"19",X"19",X"19",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"15",X"15",X"15",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"09",
		X"09",X"09",X"09",X"09",X"09",X"09",X"0A",X"09",X"09",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"09",X"0A",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"12",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",
		X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"16",X"19",X"19",X"19",
		X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"06",X"03",X"7F",X"FF",X"8F",X"7F",X"7F",X"7F",X"06",X"0F",X"7F",X"BF",X"FF",X"0B",X"0B",X"0F",
		X"03",X"07",X"07",X"73",X"33",X"03",X"03",X"07",X"00",X"0C",X"1E",X"0E",X"0F",X"1F",X"07",X"07",
		X"C0",X"C0",X"80",X"80",X"80",X"00",X"00",X"E0",X"FC",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"04",X"0E",X"0E",X"1E",X"1C",X"07",X"0F",X"0F",X"0B",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"70",X"70",X"70",X"38",X"E0",X"F0",X"F0",X"98",X"88",X"00",X"00",X"00",
		X"3C",X"1C",X"1C",X"0E",X"0E",X"07",X"0F",X"1E",X"00",X"1C",X"00",X"0E",X"00",X"07",X"05",X"0A",
		X"38",X"18",X"1C",X"0C",X"0C",X"0C",X"1E",X"3E",X"00",X"18",X"00",X"0C",X"00",X"0C",X"0A",X"16",
		X"03",X"03",X"0E",X"38",X"60",X"00",X"00",X"00",X"00",X"03",X"0E",X"38",X"60",X"00",X"00",X"00",
		X"7F",X"BC",X"BC",X"3C",X"1C",X"08",X"04",X"0F",X"0F",X"67",X"67",X"E7",X"77",X"3F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"80",X"80",X"80",X"80",X"80",X"C0",X"C0",
		X"00",X"00",X"70",X"F8",X"F0",X"70",X"38",X"3C",X"0F",X"3F",X"0F",X"07",X"03",X"70",X"00",X"3C",
		X"00",X"00",X"00",X"00",X"20",X"E0",X"E0",X"E0",X"C0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"1C",X"0E",X"06",X"0E",X"1C",X"00",X"00",X"00",X"00",X"0E",X"02",X"06",X"08",X"00",X"00",X"00",
		X"E0",X"F0",X"F0",X"70",X"38",X"18",X"38",X"78",X"00",X"F0",X"00",X"70",X"00",X"18",X"28",X"30",
		X"01",X"01",X"01",X"03",X"06",X"0C",X"18",X"10",X"00",X"00",X"01",X"03",X"06",X"0C",X"18",X"10",
		X"00",X"00",X"70",X"FC",X"7E",X"7E",X"7F",X"3F",X"0F",X"3F",X"0F",X"03",X"07",X"08",X"12",X"14",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"80",
		X"0F",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"05",X"01",X"00",X"01",X"01",X"00",X"00",X"00",
		X"E0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"A0",X"70",X"20",X"40",X"00",X"00",X"00",X"00",
		X"1C",X"0E",X"7F",X"FF",X"87",X"7F",X"7F",X"7F",X"1C",X"3E",X"7F",X"CF",X"FF",X"07",X"07",X"07",
		X"07",X"07",X"17",X"3F",X"3F",X"06",X"06",X"0F",X"3C",X"7C",X"EC",X"C5",X"47",X"7F",X"0F",X"0F",
		X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"C0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F0",X"E0",X"C0",
		X"03",X"03",X"1F",X"3F",X"7F",X"3F",X"00",X"03",X"04",X"0F",X"00",X"07",X"02",X"00",X"00",X"01",
		X"C0",X"E0",X"F0",X"F8",X"F0",X"E0",X"E0",X"E0",X"30",X"D8",X"28",X"E0",X"00",X"E0",X"E0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"0E",X"0E",X"0E",X"1F",X"1F",X"3F",X"3F",X"1E",X"00",X"00",X"00",
		X"40",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"78",X"80",X"E0",X"00",X"E0",X"00",X"E0",X"E0",X"68",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",X"3E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"0E",X"16",
		X"00",X"00",X"40",X"6C",X"7E",X"7E",X"7C",X"7E",X"7E",X"7F",X"3F",X"13",X"01",X"00",X"00",X"06",
		X"3F",X"3B",X"32",X"70",X"70",X"E0",X"C0",X"00",X"3F",X"01",X"32",X"00",X"70",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"00",X"E0",X"00",X"E0",X"00",X"E0",X"A0",X"F0",
		X"07",X"07",X"0F",X"7F",X"FF",X"07",X"03",X"0F",X"0C",X"3C",X"30",X"00",X"00",X"18",X"1C",X"0F",
		X"90",X"80",X"84",X"8C",X"0C",X"FC",X"F8",X"E0",X"F0",X"F8",X"F8",X"F0",X"F0",X"00",X"00",X"E0",
		X"01",X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"03",X"07",X"07",X"07",X"07",X"3F",X"3F",
		X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"C0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"03",X"03",X"01",X"00",X"00",X"00",X"04",X"03",X"1F",X"1F",X"0F",X"07",X"07",X"07",X"07",X"0F",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"C0",
		X"10",X"18",X"3C",X"7C",X"F0",X"E0",X"F0",X"70",X"0F",X"07",X"03",X"01",X"00",X"E0",X"20",X"50",
		X"38",X"38",X"1C",X"38",X"70",X"00",X"00",X"00",X"20",X"18",X"0C",X"18",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"0F",X"07",X"07",X"07",X"03",X"01",
		X"70",X"30",X"30",X"00",X"00",X"00",X"30",X"C0",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F8",
		X"00",X"00",X"00",X"04",X"0E",X"0F",X"0E",X"0E",X"01",X"03",X"07",X"03",X"01",X"00",X"00",X"00",
		X"00",X"04",X"04",X"0C",X"18",X"38",X"38",X"3C",X"F8",X"F8",X"FC",X"F0",X"F8",X"20",X"30",X"3C",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",X"3E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"0E",X"16",X"00",
		X"07",X"03",X"03",X"03",X"33",X"7B",X"73",X"61",X"04",X"00",X"1C",X"3C",X"0E",X"06",X"06",X"07",
		X"F8",X"F8",X"F8",X"F8",X"C0",X"C6",X"CE",X"FE",X"38",X"28",X"28",X"38",X"7C",X"78",X"70",X"00",
		X"63",X"E0",X"E0",X"1C",X"3F",X"3F",X"1E",X"00",X"03",X"07",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"FC",X"9C",X"1E",X"3E",X"3C",X"70",X"78",X"00",X"00",X"60",X"FC",X"C2",X"38",X"60",X"70",X"00",
		X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",
		X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",
		X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",
		X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",
		X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",
		X"7E",X"60",X"7E",X"03",X"03",X"63",X"3E",X"00",X"7E",X"60",X"7E",X"03",X"03",X"63",X"3E",X"00",
		X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",
		X"7F",X"63",X"06",X"0C",X"18",X"18",X"18",X"00",X"7F",X"63",X"06",X"0C",X"18",X"18",X"18",X"00",
		X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",
		X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",
		X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",
		X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",
		X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",
		X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"3F",X"7F",X"7F",X"7F",X"BF",X"BE",X"00",X"0C",X"3E",X"7E",X"7F",X"7F",X"FF",X"FF",
		X"01",X"01",X"E8",X"FC",X"E2",X"BE",X"7F",X"7F",X"00",X"1E",X"FF",X"3F",X"7F",X"C3",X"80",X"80",
		X"E0",X"F0",X"38",X"1C",X"3E",X"38",X"E3",X"FF",X"00",X"70",X"80",X"DC",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"C3",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"2B",X"2F",
		X"60",X"E0",X"F0",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"10",X"18",X"0C",X"06",X"03",X"01",
		X"81",X"C1",X"E3",X"E2",X"76",X"34",X"1C",X"18",X"01",X"01",X"03",X"02",X"06",X"04",X"04",X"00",
		X"00",X"30",X"38",X"38",X"38",X"38",X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"30",X"18",X"0C",X"06",X"03",X"01",
		X"03",X"07",X"07",X"0E",X"1C",X"38",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"60",X"30",X"18",X"0C",X"04",X"00",X"00",X"C0",X"60",X"30",X"18",X"0C",X"04",X"00",X"00",
		X"80",X"E0",X"38",X"0E",X"03",X"07",X"07",X"03",X"80",X"E0",X"38",X"0E",X"03",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"FC",X"7C",X"1C",X"78",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"03",X"7F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"02",X"03",X"03",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",
		X"07",X"FF",X"06",X"06",X"06",X"06",X"07",X"07",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"78",X"2C",X"26",X"63",X"E1",X"C0",X"00",X"00",X"18",X"0C",X"06",X"03",X"01",X"00",
		X"07",X"FF",X"0E",X"0C",X"1C",X"1C",X"1C",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"3C",X"2E",X"27",X"63",X"40",X"C0",X"80",X"00",X"00",X"20",X"20",X"60",X"40",X"C0",X"80",
		X"00",X"06",X"03",X"7F",X"FF",X"8F",X"7F",X"7F",X"00",X"06",X"0F",X"7F",X"BF",X"FF",X"0B",X"0B",
		X"18",X"1C",X"1E",X"0E",X"1E",X"FC",X"E0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",
		X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"E0",X"F8",X"FE",X"FF",X"FC",X"E0",X"C0",X"E0",X"E0",X"F8",X"FE",X"FF",X"FC",X"F0",X"30",
		X"7F",X"78",X"1C",X"3F",X"7F",X"27",X"03",X"07",X"1C",X"09",X"1F",X"0E",X"6F",X"07",X"07",X"01",
		X"80",X"03",X"0E",X"00",X"80",X"C0",X"C0",X"F0",X"60",X"F3",X"FE",X"F0",X"70",X"B0",X"B0",X"00",
		X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"04",X"05",X"05",
		X"80",X"40",X"40",X"40",X"40",X"00",X"00",X"00",X"70",X"B0",X"B0",X"B0",X"B8",X"F8",X"F8",X"F8",
		X"06",X"07",X"07",X"07",X"07",X"06",X"0C",X"00",X"01",X"06",X"07",X"07",X"07",X"00",X"02",X"3E",
		X"08",X"F8",X"38",X"1C",X"0C",X"0C",X"0C",X"00",X"F0",X"08",X"38",X"1C",X"0C",X"02",X"02",X"1C",
		X"01",X"07",X"1F",X"3F",X"7F",X"7F",X"33",X"3B",X"01",X"07",X"1F",X"3F",X"1F",X"0F",X"13",X"38",
		X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"E0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",
		X"1B",X"1E",X"0F",X"3F",X"77",X"27",X"02",X"07",X"18",X"1D",X"0E",X"0E",X"66",X"00",X"05",X"00",
		X"BE",X"03",X"0E",X"00",X"00",X"00",X"00",X"F0",X"7E",X"F3",X"FE",X"F0",X"F0",X"F0",X"F0",X"00",
		X"03",X"02",X"06",X"14",X"1C",X"1C",X"1C",X"1C",X"04",X"0D",X"09",X"0B",X"13",X"1B",X"1B",X"1B",
		X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"04",X"F0",X"70",X"70",X"78",X"78",X"F8",X"FC",X"F8",
		X"1E",X"19",X"31",X"00",X"00",X"00",X"00",X"00",X"1D",X"00",X"09",X"F8",X"00",X"00",X"00",X"00",
		X"18",X"FC",X"FC",X"E0",X"00",X"00",X"00",X"00",X"E6",X"1A",X"FA",X"E6",X"00",X"00",X"00",X"00",
		X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"07",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"00",
		X"17",X"12",X"11",X"7B",X"F3",X"F4",X"F4",X"7F",X"1C",X"1F",X"1F",X"06",X"4E",X"7F",X"7F",X"90",
		X"E0",X"40",X"80",X"E0",X"FC",X"7E",X"3E",X"FE",X"30",X"F8",X"7C",X"7E",X"72",X"FC",X"FC",X"1C",
		X"16",X"15",X"15",X"15",X"15",X"14",X"15",X"1E",X"79",X"3A",X"1A",X"1A",X"1A",X"1B",X"1A",X"11",
		X"0C",X"00",X"00",X"30",X"70",X"F0",X"70",X"30",X"F2",X"FC",X"F0",X"C0",X"B8",X"78",X"F8",X"F0",
		X"1E",X"1E",X"17",X"17",X"03",X"03",X"06",X"00",X"1F",X"1E",X"17",X"17",X"03",X"00",X"01",X"0F",
		X"30",X"48",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"78",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"33",X"3A",X"3E",X"1E",X"1F",X"06",X"0E",X"1E",X"0C",X"35",X"39",X"1D",X"1C",
		X"80",X"40",X"40",X"40",X"20",X"00",X"02",X"0C",X"78",X"B8",X"BC",X"BC",X"DE",X"FE",X"FC",X"F0",
		X"0F",X"06",X"0E",X"00",X"00",X"00",X"00",X"00",X"0E",X"05",X"01",X"1E",X"00",X"00",X"00",X"00",
		X"FC",X"1E",X"0E",X"0E",X"06",X"06",X"0E",X"00",X"0C",X"1E",X"0E",X"0E",X"06",X"05",X"01",X"1E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"3C",X"38",X"78",X"20",X"C0",X"00",X"1E",X"1E",X"3F",X"18",X"08",X"D0",X"20",X"C0",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"30",X"10",X"10",X"00",X"04",X"0E",X"20",X"20",X"30",X"10",X"10",X"00",X"04",X"0E",
		X"7F",X"78",X"1C",X"0E",X"0F",X"07",X"03",X"07",X"1C",X"09",X"1F",X"0F",X"0F",X"07",X"03",X"01",
		X"80",X"08",X"08",X"08",X"0C",X"84",X"84",X"F6",X"70",X"F8",X"F8",X"F8",X"FC",X"F4",X"F4",X"06",
		X"07",X"0A",X"0A",X"12",X"12",X"1E",X"0E",X"06",X"00",X"05",X"05",X"0D",X"0D",X"11",X"0D",X"05",
		X"02",X"82",X"82",X"80",X"80",X"00",X"08",X"38",X"F2",X"7A",X"7A",X"78",X"78",X"F8",X"F0",X"C8",
		X"03",X"01",X"02",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"07",X"00",X"00",X"00",X"00",
		X"F8",X"B8",X"38",X"38",X"38",X"18",X"10",X"00",X"38",X"B8",X"B8",X"B8",X"00",X"00",X"2C",X"3E",
		X"1B",X"1E",X"0F",X"0F",X"07",X"07",X"02",X"07",X"18",X"1D",X"0E",X"0E",X"06",X"00",X"05",X"00",
		X"08",X"08",X"08",X"0C",X"04",X"04",X"04",X"F6",X"F8",X"F8",X"F8",X"FC",X"F4",X"F4",X"F4",X"06",
		X"1E",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1E",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"10",X"BF",X"C0",X"C0",X"C0",X"9F",X"BF",X"1F",X"00",X"87",X"FC",X"FF",X"FF",X"EF",X"DF",X"EF",
		X"00",X"FF",X"00",X"41",X"63",X"E3",X"FF",X"FF",X"0E",X"FF",X"3F",X"BE",X"9D",X"FD",X"F3",X"F1",
		X"00",X"F8",X"80",X"C0",X"E0",X"F2",X"FE",X"B8",X"00",X"F8",X"00",X"C0",X"E1",X"F1",X"F9",X"BE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"00",X"00",X"01",X"07",X"0F",X"1F",X"3F",X"7F",X"00",
		X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"EC",X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FF",X"00",
		X"03",X"03",X"01",X"02",X"02",X"03",X"1F",X"3F",X"00",X"07",X"0F",X"1F",X"1F",X"3F",X"2F",X"1F",
		X"EE",X"8E",X"0E",X"1E",X"37",X"F7",X"F7",X"7D",X"70",X"F8",X"FE",X"FE",X"DF",X"8F",X"8B",X"E2",
		X"3C",X"24",X"28",X"11",X"01",X"03",X"02",X"06",X"1F",X"1B",X"17",X"07",X"07",X"07",X"07",X"07",
		X"42",X"C0",X"A0",X"A0",X"A0",X"80",X"80",X"8C",X"F8",X"F8",X"DC",X"DC",X"5C",X"7C",X"7C",X"70",
		X"04",X"0F",X"0F",X"07",X"07",X"06",X"0C",X"00",X"07",X"0C",X"0F",X"07",X"07",X"00",X"02",X"3E",
		X"FC",X"9C",X"1C",X"1C",X"0C",X"0C",X"0C",X"00",X"0C",X"1C",X"1C",X"1C",X"0C",X"00",X"02",X"1F",
		X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"3F",
		X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"07",X"07",X"03",
		X"06",X"07",X"03",X"83",X"03",X"03",X"07",X"23",X"C0",X"E0",X"F3",X"73",X"F3",X"F3",X"EF",X"FF",
		X"00",X"00",X"00",X"01",X"01",X"02",X"14",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"41",X"40",X"80",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"1F",X"1E",X"3E",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F8",X"F8",X"7C",X"3C",X"3C",
		X"1C",X"1E",X"0E",X"0E",X"06",X"03",X"07",X"1F",X"1C",X"1E",X"0E",X"0E",X"06",X"03",X"05",X"0B",
		X"1C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0E",X"1F",X"1C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",X"1A",
		X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"18",X"C0",X"E0",X"F0",X"70",X"F0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"31",X"31",X"12",X"04",X"07",X"07",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"3C",X"4C",X"8C",X"0E",X"06",X"00",X"00",X"E0",X"E4",X"FC",X"FE",X"FE",X"FE",X"FE",X"F0",X"E0",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"70",X"F0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"01",X"61",X"62",X"3F",X"3F",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"07",X"0F",
		X"20",X"40",X"80",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"FC",X"7F",X"03",X"07",X"07",X"07",X"07",X"1F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"0F",X"13",X"27",X"27",X"47",X"47",X"42",X"7E",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"7E",
		X"00",X"00",X"60",X"70",X"38",X"3C",X"1C",X"0E",X"3F",X"7F",X"7F",X"7F",X"3F",X"3C",X"1C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"78",X"3C",
		X"06",X"0E",X"3E",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"3E",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"0E",X"0E",X"06",X"07",X"0E",X"18",X"1C",X"1C",X"0E",X"0E",X"06",X"03",X"06",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"3C",X"3F",X"3F",X"7F",X"7E",X"FC",X"F8",X"F8",X"FC",
		X"3E",X"0F",X"07",X"03",X"07",X"0E",X"00",X"00",X"3E",X"0F",X"07",X"03",X"03",X"04",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"03",X"00",X"00",X"03",X"07",X"0F",X"0B",X"08",X"0C",X"07",X"03",
		X"00",X"00",X"00",X"20",X"E8",X"CC",X"0C",X"0C",X"C0",X"E0",X"F0",X"D0",X"10",X"30",X"E0",X"CC",
		X"00",X"00",X"00",X"01",X"12",X"0A",X"0C",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",
		X"2E",X"4E",X"8E",X"06",X"00",X"00",X"00",X"E0",X"FE",X"FE",X"FE",X"FE",X"FC",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",X"0F",X"1F",X"1F",X"3F",X"3E",X"3C",X"3C",X"1C",
		X"1C",X"0E",X"0E",X"06",X"0E",X"1E",X"00",X"00",X"1C",X"0E",X"0E",X"06",X"06",X"1A",X"00",X"00",
		X"0F",X"1F",X"1D",X"38",X"30",X"70",X"F0",X"00",X"0F",X"1F",X"1D",X"38",X"30",X"30",X"50",X"00",
		X"C0",X"E0",X"E0",X"78",X"18",X"38",X"70",X"00",X"C0",X"E0",X"E0",X"78",X"18",X"18",X"30",X"00",
		X"08",X"08",X"24",X"C0",X"03",X"24",X"10",X"10",X"18",X"18",X"3C",X"FF",X"FF",X"3C",X"18",X"18",
		X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",
		X"3F",X"3E",X"60",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"00",X"02",X"04",X"04",X"07",X"FF",X"FF",X"FF",X"0F",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"03",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"00",X"20",X"60",X"40",X"00",
		X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"C0",X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"20",X"60",X"40",X"C0",X"00",X"00",X"00",X"00",X"20",X"60",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"18",X"0C",X"0C",X"06",X"04",X"00",X"00",X"00",X"26",X"73",X"F3",X"F9",X"FB",X"7F",X"3E",
		X"00",X"00",X"F0",X"0C",X"02",X"00",X"01",X"01",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0C",X"1E",X"0F",X"00",X"00",X"F8",X"FC",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"E7",X"FB",
		X"00",X"00",X"00",X"00",X"01",X"63",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"E1",X"FE",X"FF",
		X"00",X"3C",X"FA",X"0F",X"27",X"7B",X"4E",X"00",X"00",X"3C",X"46",X"79",X"3D",X"85",X"7E",X"00",
		X"01",X"07",X"21",X"16",X"08",X"66",X"01",X"27",X"01",X"04",X"3E",X"0B",X"FF",X"19",X"07",X"28",
		X"F8",X"FE",X"FF",X"DF",X"6D",X"7B",X"B6",X"FC",X"F8",X"0E",X"43",X"2D",X"F3",X"85",X"CE",X"7C",
		X"00",X"00",X"08",X"38",X"1C",X"10",X"00",X"00",X"00",X"00",X"08",X"38",X"1C",X"10",X"00",X"00",
		X"00",X"00",X"24",X"18",X"18",X"24",X"00",X"00",X"00",X"00",X"24",X"18",X"18",X"24",X"00",X"00",
		X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"1F",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"1F",
		X"00",X"00",X"80",X"80",X"88",X"90",X"A0",X"C0",X"00",X"00",X"80",X"80",X"88",X"90",X"A0",X"C0",
		X"00",X"00",X"00",X"09",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"09",X"07",X"03",X"00",X"00",
		X"38",X"38",X"78",X"F0",X"E0",X"C0",X"00",X"00",X"38",X"38",X"78",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"18",X"18",X"18",X"00",X"00",X"00",X"20",X"10",X"18",X"18",X"18",
		X"00",X"00",X"38",X"7C",X"7C",X"7C",X"7C",X"38",X"00",X"00",X"08",X"04",X"04",X"04",X"4C",X"38",
		X"07",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"0F",X"06",X"00",X"00",X"00",
		X"E0",X"F8",X"78",X"38",X"10",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"78",X"30",X"00",X"00",X"00",
		X"07",X"0E",X"1F",X"3E",X"3F",X"1F",X"0F",X"77",X"07",X"0E",X"3F",X"7F",X"7F",X"7F",X"3F",X"7F",
		X"78",X"FC",X"FE",X"7C",X"B8",X"DE",X"DF",X"FE",X"78",X"FC",X"FE",X"FE",X"FC",X"FE",X"FF",X"FF",
		X"7F",X"7B",X"77",X"37",X"1B",X"0F",X"06",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1E",X"0C",
		X"FC",X"D8",X"BC",X"FE",X"FE",X"7C",X"38",X"00",X"FF",X"FE",X"FC",X"FE",X"FE",X"FE",X"FC",X"38",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"18",X"99",X"18",X"00",X"00",X"00",X"00",X"00",X"66",X"E7",X"66",X"00",X"00",
		X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"41",X"00",X"3C",X"0C",X"0C",X"3C",X"18",X"3E",X"3E",
		X"38",X"FE",X"4F",X"17",X"6B",X"5F",X"B6",X"3C",X"38",X"06",X"73",X"39",X"95",X"7B",X"4E",X"3C",
		X"18",X"08",X"3C",X"3C",X"7C",X"38",X"10",X"82",X"18",X"18",X"3C",X"34",X"64",X"00",X"6C",X"7C",
		X"00",X"00",X"03",X"03",X"81",X"61",X"18",X"06",X"03",X"07",X"04",X"04",X"86",X"62",X"1B",X"07",
		X"00",X"00",X"00",X"60",X"40",X"10",X"30",X"00",X"00",X"80",X"E0",X"90",X"B8",X"E8",X"C8",X"C0",
		X"80",X"30",X"18",X"00",X"00",X"00",X"00",X"00",X"F8",X"4C",X"64",X"3A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"60",X"18",X"04",X"02",X"39",X"00",X"00",X"80",X"60",X"18",X"04",X"7A",X"C7",
		X"60",X"08",X"12",X"06",X"00",X"00",X"00",X"00",X"9F",X"F7",X"EC",X"78",X"38",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"20",X"00",X"00",X"00",X"C0",X"F0",X"BC",X"9A",X"D1",X"60",X"00",X"00",
		X"00",X"20",X"12",X"04",X"20",X"48",X"04",X"00",X"00",X"62",X"36",X"1C",X"38",X"6C",X"46",X"00",
		X"0F",X"07",X"00",X"00",X"00",X"0C",X"1F",X"3F",X"09",X"0F",X"0F",X"07",X"07",X"0F",X"1F",X"3F",
		X"F8",X"F0",X"30",X"78",X"7C",X"7E",X"3E",X"9C",X"9C",X"FC",X"FC",X"FC",X"FC",X"FE",X"3E",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0B",X"00",X"00",X"00",X"07",X"0F",X"0F",X"09",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"B8",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"9C",X"DC",
		X"0F",X"27",X"30",X"38",X"38",X"3C",X"1E",X"00",X"09",X"2F",X"3F",X"3F",X"3F",X"3F",X"1E",X"00",
		X"F8",X"F0",X"00",X"00",X"00",X"1C",X"3E",X"3F",X"9C",X"FC",X"FC",X"FC",X"FC",X"FC",X"3E",X"3F",
		X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"DF",X"85",
		X"07",X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"00",X"04",X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",
		X"F0",X"F0",X"40",X"40",X"40",X"C0",X"60",X"40",X"70",X"F0",X"F0",X"F8",X"FC",X"3C",X"9C",X"FC",
		X"04",X"00",X"10",X"30",X"21",X"01",X"01",X"01",X"7F",X"7F",X"6F",X"CF",X"DF",X"FF",X"7F",X"1F",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F8",X"FC",X"FE",X"FE",X"FE",X"FC",
		X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"1F",X"1D",X"3D",X"3B",X"7B",X"77",X"EF",
		X"00",X"00",X"80",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"78",X"7C",X"BC",X"BE",X"DE",X"EF",
		X"00",X"00",X"00",X"00",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"07",X"07",
		X"1F",X"1F",X"12",X"12",X"12",X"12",X"12",X"02",X"01",X"13",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"08",X"08",X"08",X"08",X"0C",X"FF",X"FE",X"FC",X"9F",X"1F",X"1F",X"1F",X"1B",
		X"00",X"80",X"00",X"00",X"20",X"20",X"30",X"10",X"F0",X"70",X"F0",X"E0",X"E0",X"E0",X"F0",X"F0",
		X"1C",X"1C",X"3E",X"3E",X"3F",X"3F",X"1F",X"03",X"1B",X"1B",X"3D",X"3D",X"3E",X"3E",X"1F",X"0F",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",
		X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"FF",X"FF",X"FF",X"9F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"60",X"E0",X"60",X"30",X"10",X"F8",X"F8",X"F8",X"98",X"10",X"A0",X"F0",X"F0",
		X"0E",X"0E",X"1E",X"1F",X"1F",X"0F",X"0F",X"07",X"15",X"15",X"0D",X"0E",X"1E",X"0F",X"0F",X"07",
		X"10",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"E0",X"E0",X"F0",X"F0",X"70",X"B8",X"DC",
		X"3C",X"42",X"89",X"85",X"85",X"81",X"42",X"3C",X"00",X"3C",X"76",X"7A",X"7A",X"7E",X"3C",X"00",
		X"3C",X"7E",X"FF",X"FD",X"FD",X"FB",X"76",X"3C",X"00",X"00",X"00",X"02",X"02",X"04",X"08",X"00",
		X"00",X"00",X"00",X"1E",X"03",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"38",X"00",X"00",
		X"00",X"00",X"1C",X"7E",X"27",X"3E",X"00",X"00",X"00",X"00",X"1C",X"02",X"F9",X"4E",X"00",X"00",
		X"00",X"00",X"3C",X"FE",X"2F",X"6B",X"4E",X"00",X"00",X"00",X"3C",X"06",X"31",X"9D",X"76",X"00",
		X"00",X"00",X"F0",X"E0",X"C3",X"07",X"0F",X"0F",X"00",X"00",X"90",X"60",X"03",X"C7",X"EF",X"FF",
		X"00",X"00",X"0F",X"07",X"C3",X"E0",X"F0",X"F0",X"00",X"00",X"09",X"06",X"C0",X"E3",X"F7",X"FF",
		X"0F",X"0F",X"0F",X"07",X"04",X"04",X"04",X"04",X"FD",X"FC",X"F8",X"FC",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"D0",X"40",X"40",X"40",X"40",X"40",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"04",X"00",X"10",X"11",X"11",X"13",X"13",X"FF",X"7F",X"3F",X"1F",X"1F",X"1F",X"1D",X"1D",
		X"40",X"40",X"00",X"08",X"08",X"08",X"88",X"88",X"FF",X"FE",X"FC",X"F8",X"F8",X"F8",X"78",X"78",
		X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",X"1F",X"1D",X"1D",X"3B",X"3B",X"3B",X"77",X"77",X"EF",
		X"80",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",X"F8",X"78",X"78",X"BC",X"BC",X"BC",X"DE",X"DE",X"E7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"FF",
		X"FF",X"41",X"25",X"11",X"09",X"05",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"82",X"A4",X"88",X"90",X"A0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"60",X"30",X"18",X"0C",X"06",X"03",X"00",X"00",X"DF",X"EF",X"F7",X"FB",X"FD",X"FE",
		X"FF",X"00",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"00",X"00",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"FF",X"00",X"06",X"0C",X"18",X"30",X"60",X"C0",X"00",X"00",X"FB",X"F7",X"EF",X"DF",X"BF",X"7F",
		X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"FF",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"DD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"C0",X"C0",X"60",X"60",X"30",X"30",X"00",X"00",X"BF",X"BF",X"DF",X"DF",X"EF",X"EF",
		X"FF",X"00",X"03",X"03",X"06",X"06",X"0C",X"0C",X"00",X"00",X"FD",X"FD",X"FB",X"FB",X"F7",X"F7",
		X"18",X"18",X"0C",X"0C",X"06",X"06",X"03",X"03",X"F7",X"F7",X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",
		X"18",X"18",X"30",X"30",X"60",X"60",X"C0",X"C0",X"EF",X"EF",X"DF",X"DF",X"BF",X"BF",X"7F",X"7F",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"88",X"94",X"94",X"88",X"80",X"80",X"80",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"11",X"29",X"29",X"11",X"01",X"01",X"01",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"BC",X"A6",X"83",X"80",X"80",X"83",X"A6",X"B4",X"83",X"99",X"80",X"99",X"BD",X"BC",X"99",X"88",
		X"FF",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",
		X"FF",X"00",X"82",X"82",X"82",X"82",X"82",X"82",X"00",X"00",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"FF",X"00",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"00",X"00",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",X"D1",X"FF",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"FF",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"FF",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"FF",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"FF",
		X"3C",X"66",X"43",X"00",X"00",X"C3",X"66",X"34",X"C3",X"99",X"80",X"99",X"3D",X"3C",X"99",X"08",
		X"3D",X"65",X"41",X"01",X"01",X"C1",X"65",X"35",X"C1",X"99",X"81",X"99",X"3D",X"3D",X"99",X"09",
		X"80",X"80",X"BC",X"A6",X"83",X"80",X"80",X"FF",X"99",X"93",X"83",X"99",X"BC",X"BF",X"80",X"FF",
		X"00",X"00",X"3C",X"66",X"43",X"00",X"00",X"FF",X"99",X"D3",X"C3",X"99",X"BC",X"FF",X"00",X"FF",
		X"01",X"01",X"3D",X"65",X"41",X"01",X"01",X"FF",X"99",X"D1",X"C1",X"99",X"BD",X"FD",X"01",X"FF",
		X"03",X"1F",X"7B",X"ED",X"75",X"37",X"3E",X"18",X"00",X"01",X"0F",X"3F",X"1F",X"1C",X"00",X"00",
		X"C0",X"F8",X"DE",X"B7",X"AE",X"EC",X"7C",X"18",X"00",X"80",X"F0",X"FC",X"F8",X"38",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"00",X"00",X"40",X"80",X"80",X"40",X"E0",X"E0",X"00",X"00",X"00",X"60",X"60",X"40",X"80",X"9F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"DD",X"DD",X"B9",X"B9",X"76",X"76",
		X"27",X"17",X"97",X"8F",X"CF",X"C7",X"E7",X"E7",X"84",X"84",X"44",X"44",X"A4",X"A4",X"D4",X"D4",
		X"E4",X"E8",X"E9",X"F1",X"F3",X"E3",X"E7",X"E7",X"81",X"81",X"82",X"82",X"85",X"85",X"8B",X"8B",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"BB",X"BB",X"9D",X"9D",X"6E",X"6E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"DF",X"DF",X"9F",X"9F",X"6F",X"6F",
		X"F7",X"F7",X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",X"6C",X"6C",X"B4",X"B4",X"DA",X"DA",X"ED",X"ED",
		X"02",X"44",X"04",X"22",X"87",X"57",X"47",X"2F",X"40",X"23",X"23",X"12",X"14",X"0C",X"0C",X"04",
		X"40",X"82",X"80",X"45",X"E1",X"EA",X"E2",X"F4",X"02",X"64",X"64",X"48",X"88",X"90",X"90",X"80",
		X"EF",X"EF",X"DF",X"DF",X"BF",X"BF",X"7F",X"7F",X"96",X"96",X"AD",X"AD",X"DB",X"DB",X"B7",X"B7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"FB",X"FB",X"F9",X"F9",X"F6",X"F6",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"77",X"77",X"3B",X"3B",X"1D",X"1D",X"0E",X"0E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"EB",X"EB",X"DD",X"DD",X"BE",X"BE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6F",X"6F",X"D7",X"D7",X"BB",X"BB",X"7D",X"7D",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"EE",X"EE",X"DC",X"DC",X"B8",X"B8",X"70",X"70",
		X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",X"07",X"07",X"03",X"03",X"01",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"BF",X"BF",X"DF",X"DF",X"EF",X"EF",
		X"00",X"00",X"02",X"04",X"04",X"02",X"07",X"07",X"00",X"00",X"00",X"03",X"03",X"02",X"04",X"FC",
		X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"02",
		X"FF",X"E4",X"E4",X"E4",X"E4",X"E4",X"E4",X"FF",X"80",X"84",X"84",X"84",X"84",X"84",X"84",X"80",
		X"FF",X"27",X"27",X"27",X"27",X"27",X"27",X"FF",X"04",X"24",X"24",X"24",X"24",X"24",X"24",X"04",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"80",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",
		X"FF",X"01",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"00",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"80",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F6",X"F6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"01",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",
		X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"F9",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",
		X"FF",X"FF",X"FB",X"FB",X"F9",X"F9",X"F9",X"F9",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D6",X"D6",
		X"FF",X"FF",X"FD",X"FD",X"F9",X"F9",X"F9",X"F9",X"EE",X"EE",X"DE",X"DE",X"BE",X"BE",X"76",X"76",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"F7",X"FB",X"FB",X"DD",X"DD",X"DE",X"DE",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"FE",X"FE",X"F1",X"E6",X"C8",X"91",X"22",X"44",X"03",X"0F",X"1F",X"3E",X"78",X"F1",X"E2",X"C4",
		X"88",X"91",X"22",X"44",X"89",X"13",X"A7",X"4F",X"88",X"91",X"22",X"44",X"89",X"13",X"A7",X"4F",
		X"9E",X"3C",X"78",X"F0",X"E0",X"C0",X"80",X"00",X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"9E",X"3E",X"7A",X"F2",X"E2",X"E2",X"E2",X"E2",X"9F",X"3D",X"7F",X"FF",X"FF",X"DF",X"DF",X"DF",
		X"9F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"3F",X"7F",X"FF",X"EF",X"EF",X"AF",X"2F",
		X"7B",X"3E",X"1E",X"0F",X"07",X"03",X"03",X"02",X"FB",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"13",X"8B",X"46",X"22",X"93",X"CA",X"E6",X"F2",X"13",X"8B",X"46",X"22",X"93",X"CA",X"E6",X"F2",
		X"7F",X"7F",X"8F",X"67",X"13",X"8B",X"46",X"22",X"C2",X"F2",X"FA",X"7E",X"1E",X"8F",X"47",X"23",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"02",X"02",X"02",X"02",X"02",X"02",X"82",X"C2",
		X"FB",X"FE",X"FE",X"EF",X"E7",X"E3",X"E3",X"E2",X"FB",X"FE",X"DE",X"DF",X"DF",X"DF",X"DF",X"DF",
		X"FB",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7B",X"3E",X"3E",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"FB",X"3E",X"1E",X"FF",X"07",X"FF",X"FF",X"FF",X"7B",X"FE",X"FE",X"0F",X"FF",X"03",X"FF",X"FF",
		X"9F",X"3E",X"7A",X"FF",X"E2",X"FF",X"FF",X"FF",X"9E",X"3F",X"7F",X"F2",X"FF",X"C2",X"FF",X"FF",
		X"83",X"C3",X"7E",X"02",X"FF",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"FF",X"FF",
		X"FF",X"02",X"02",X"02",X"FF",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"FF",X"FF",
		X"02",X"FF",X"02",X"02",X"FF",X"FF",X"FF",X"FF",X"02",X"FF",X"02",X"02",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"03",X"03",X"03",X"02",X"02",X"02",X"02",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"02",X"02",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"02",X"02",X"FE",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"82",X"82",X"FF",X"82",X"82",X"82",X"82",X"82",
		X"FE",X"82",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"82",X"82",X"FE",X"82",X"82",X"82",X"82",X"82",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"C2",X"0F",X"02",X"02",X"02",X"02",X"02",X"07",X"3F",X"F2",
		X"FF",X"FF",X"FE",X"F2",X"02",X"1B",X"73",X"EF",X"02",X"02",X"03",X"0F",X"FF",X"E6",X"8E",X"12",
		X"DF",X"07",X"03",X"02",X"82",X"A6",X"73",X"FF",X"22",X"FA",X"FE",X"FF",X"7F",X"5B",X"8E",X"02",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"03",X"C2",X"FF",X"02",X"02",X"02",X"82",X"E2",X"FE",X"3F",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7A",X"C7",X"02",X"02",X"02",X"02",X"02",X"03",X"87",X"3A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"FF",X"02",X"02",X"02",X"02",X"02",X"02",X"FA",X"02",
		X"FF",X"F3",X"FB",X"FA",X"FE",X"FE",X"FE",X"FE",X"02",X"0E",X"07",X"07",X"03",X"03",X"03",X"03",
		X"EF",X"27",X"16",X"96",X"AA",X"AA",X"AB",X"A6",X"1A",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"E6",X"C2",X"03",X"03",X"03",X"03",X"03",X"03",X"1B",X"3F",
		X"AB",X"A6",X"AA",X"A2",X"83",X"87",X"1F",X"9F",X"FF",X"FF",X"FF",X"FF",X"FE",X"FA",X"F2",X"F2",
		X"CB",X"E6",X"EA",X"F6",X"F2",X"FA",X"9A",X"8A",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"67",X"77",
		X"23",X"07",X"4F",X"0F",X"2B",X"87",X"2F",X"67",X"FE",X"FE",X"FA",X"F2",X"F6",X"FE",X"FA",X"FA",
		X"CE",X"C6",X"E6",X"E2",X"F2",X"F3",X"3B",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"43",X"4F",X"4F",X"4B",X"4B",X"5E",X"1F",X"1F",X"FE",X"FE",X"FA",X"FE",X"FE",X"FF",X"FB",X"F2",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"C7",X"03",X"3F",X"02",X"02",X"02",X"82",X"C2",X"FA",X"FE",X"FA",
		X"C3",X"03",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"82",X"02",X"02",X"02",X"02",X"02",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"0F",X"87",X"02",X"02",X"02",X"02",X"02",X"82",X"FA",X"FE",
		X"9E",X"CE",X"E3",X"F2",X"FF",X"FE",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"03",X"03",
		X"9F",X"8F",X"66",X"67",X"8B",X"06",X"03",X"F2",X"F2",X"FB",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"87",X"0F",X"1F",X"FF",X"FF",X"07",X"FF",X"1F",X"FE",X"FE",X"FA",X"FA",X"52",X"FA",X"F2",X"E2",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"E3",X"C2",X"FE",X"02",X"02",X"02",X"03",X"03",X"1F",X"3F",X"1F",
		X"F7",X"E6",X"6A",X"2B",X"17",X"07",X"C7",X"27",X"1A",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"CF",X"9F",X"1F",X"3F",X"3F",X"3F",X"7F",X"02",X"72",X"E2",X"E2",X"C2",X"C2",X"C2",X"82",
		X"C3",X"C2",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"03",X"02",X"02",X"02",X"02",X"02",
		X"97",X"67",X"17",X"C7",X"E3",X"FB",X"FA",X"DB",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"0F",X"2F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"67",X"43",X"82",X"82",X"82",X"82",X"82",X"C2",X"DA",X"FE",
		X"C6",X"E2",X"F2",X"F2",X"D6",X"E3",X"F6",X"A6",X"3F",X"3F",X"1F",X"0F",X"2F",X"3F",X"1F",X"5F",
		X"93",X"27",X"57",X"2F",X"4F",X"1F",X"1B",X"13",X"FE",X"FA",X"FA",X"F2",X"F2",X"E2",X"E6",X"EE",
		X"C2",X"F2",X"F2",X"D2",X"92",X"7A",X"FA",X"FA",X"7F",X"3F",X"1F",X"3F",X"7F",X"FF",X"9F",X"0F",
		X"73",X"63",X"67",X"47",X"4F",X"CF",X"9E",X"BA",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F2",X"E3",X"02",X"02",X"02",X"02",X"02",X"03",X"1F",X"3F",
		X"E3",X"F2",X"FA",X"FF",X"FF",X"E2",X"FF",X"FA",X"3F",X"3F",X"1F",X"1F",X"0A",X"1F",X"0F",X"07",
		X"FB",X"F3",X"66",X"E6",X"D3",X"22",X"C2",X"0F",X"0F",X"9F",X"FF",X"DF",X"BF",X"FF",X"FF",X"FF",
		X"3B",X"73",X"C7",X"0F",X"FF",X"7F",X"FF",X"FF",X"FE",X"FE",X"FA",X"F2",X"F2",X"E2",X"C2",X"82",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FB",X"FB",X"F7",X"F7",
		X"E2",X"E6",X"C6",X"E2",X"87",X"D7",X"47",X"2F",X"E2",X"E3",X"E3",X"D2",X"96",X"8E",X"0E",X"06",
		X"47",X"87",X"83",X"47",X"E3",X"EB",X"E2",X"F6",X"07",X"67",X"67",X"4B",X"8B",X"93",X"92",X"82",
		X"FF",X"FF",X"E7",X"C3",X"83",X"83",X"83",X"83",X"02",X"1A",X"3E",X"7E",X"E7",X"DB",X"DB",X"E7",
		X"0A",X"F2",X"EF",X"83",X"02",X"82",X"C2",X"DA",X"F7",X"0F",X"12",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"07",X"02",X"02",X"02",X"02",X"1F",X"3F",X"7B",X"3A",
		X"02",X"03",X"87",X"82",X"E7",X"EE",X"7A",X"73",X"02",X"02",X"7A",X"7F",X"1A",X"13",X"87",X"8E",
		X"FA",X"F2",X"DA",X"1E",X"17",X"03",X"06",X"02",X"02",X"0E",X"27",X"E3",X"EA",X"FE",X"FB",X"FF",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"C2",X"E2",X"F2",X"E2",X"C2",
		X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"3E",
		X"06",X"1F",X"1F",X"3E",X"02",X"BE",X"FF",X"72",X"1B",X"02",X"02",X"03",X"3F",X"43",X"02",X"8F",
		X"FF",X"3F",X"F2",X"13",X"03",X"4F",X"BA",X"FE",X"02",X"C2",X"0F",X"EE",X"FE",X"BE",X"4F",X"33",
		X"02",X"02",X"02",X"FA",X"FB",X"4F",X"03",X"06",X"C2",X"FA",X"FE",X"06",X"06",X"B2",X"FE",X"FA",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"07",X"1F",
		X"7E",X"07",X"03",X"27",X"FF",X"7F",X"F7",X"E2",X"83",X"FA",X"FF",X"DB",X"07",X"8F",X"3F",X"FF",
		X"E2",X"FA",X"FE",X"BF",X"7F",X"8F",X"EE",X"62",X"7F",X"F7",X"C3",X"C7",X"9B",X"FE",X"F3",X"FF",
		X"06",X"02",X"0A",X"FE",X"FA",X"9A",X"3A",X"1F",X"FF",X"FF",X"FF",X"F3",X"07",X"67",X"C7",X"E2",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"F2",X"F2",X"FE",X"FF",X"F2",X"E2",X"FA",X"FE",X"0E",
		X"02",X"A2",X"E3",X"8F",X"FA",X"F2",X"EA",X"FF",X"FF",X"5F",X"1E",X"72",X"1F",X"FF",X"FF",X"FF",
		X"03",X"03",X"CB",X"FF",X"7F",X"3A",X"1E",X"FE",X"FF",X"FF",X"3F",X"FF",X"FE",X"FF",X"E3",X"03",
		X"E2",X"A2",X"E2",X"F2",X"FF",X"7F",X"3F",X"7F",X"FF",X"FF",X"9F",X"0F",X"02",X"82",X"C2",X"82",
		X"1A",X"DF",X"83",X"07",X"83",X"BB",X"FE",X"3E",X"E7",X"22",X"7E",X"FA",X"7E",X"46",X"03",X"C3",
		X"0A",X"F2",X"E6",X"83",X"02",X"02",X"02",X"02",X"F7",X"0F",X"1B",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"7A",X"02",X"22",X"1F",X"06",X"E3",X"63",X"1E",X"86",X"FF",X"DF",X"E2",X"FA",X"1E",X"9E",X"E2",
		X"3F",X"0F",X"9F",X"C7",X"FA",X"F2",X"F2",X"E2",X"F2",X"F2",X"E2",X"FA",X"87",X"0A",X"02",X"02",
		X"E2",X"F2",X"BF",X"1F",X"0A",X"12",X"36",X"02",X"1F",X"0F",X"42",X"E2",X"F7",X"E7",X"02",X"02",
		X"D3",X"82",X"02",X"02",X"02",X"02",X"02",X"02",X"2E",X"7F",X"FF",X"F7",X"E2",X"C2",X"02",X"02",
		X"FE",X"16",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"E2",X"A2",X"02",X"02",X"02",X"02",X"02",
		X"0A",X"0F",X"12",X"02",X"02",X"02",X"02",X"02",X"F7",X"F2",X"6E",X"3E",X"12",X"02",X"02",X"02",
		X"8E",X"FA",X"F2",X"02",X"02",X"02",X"02",X"02",X"72",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"23",X"77",X"3F",X"1F",X"03",X"0F",X"1F",X"3F",X"1E",X"0A",X"42",X"E2",
		X"BF",X"9F",X"0F",X"1F",X"33",X"73",X"E2",X"82",X"4E",X"63",X"F2",X"E2",X"CE",X"8E",X"1F",X"7F",
		X"FA",X"FE",X"FF",X"FB",X"DF",X"8E",X"0E",X"3F",X"07",X"03",X"22",X"36",X"3A",X"7B",X"FB",X"C6",
		X"03",X"03",X"07",X"03",X"E3",X"FF",X"4F",X"03",X"02",X"06",X"1A",X"7E",X"1E",X"02",X"32",X"7E",
		X"83",X"E7",X"FB",X"C2",X"9F",X"FF",X"FF",X"FF",X"7E",X"1A",X"06",X"3F",X"7F",X"F2",X"02",X"02",
		X"3A",X"7E",X"C2",X"E2",X"F3",X"EF",X"9E",X"FE",X"C7",X"83",X"3F",X"1F",X"FF",X"17",X"63",X"03",
		X"3F",X"6E",X"FE",X"1E",X"0F",X"FF",X"FB",X"73",X"C2",X"97",X"07",X"E3",X"F3",X"AB",X"96",X"9F",
		X"0E",X"FF",X"C3",X"0B",X"CF",X"FB",X"F3",X"FF",X"F3",X"02",X"3E",X"F6",X"32",X"86",X"8E",X"C2",
		X"03",X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"3E",X"1E",X"1E",X"06",X"02",X"02",X"02",X"02",
		X"FF",X"F3",X"E2",X"FA",X"FE",X"13",X"3F",X"FE",X"07",X"0F",X"1F",X"07",X"03",X"EE",X"C2",X"03",
		X"FF",X"FF",X"7E",X"1F",X"0F",X"9F",X"BF",X"FF",X"F2",X"FA",X"FF",X"FF",X"FF",X"6F",X"43",X"02",
		X"8F",X"7F",X"06",X"C2",X"FF",X"FF",X"FF",X"FF",X"72",X"82",X"FB",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"02",X"03",X"1E",X"0B",X"07",X"02",X"02",X"02",X"02",X"02",X"03",X"06",X"02",X"02",X"02",X"02",
		X"67",X"C3",X"C2",X"82",X"0E",X"02",X"02",X"02",X"9A",X"3E",X"3F",X"7F",X"F3",X"CF",X"03",X"02",
		X"02",X"C2",X"AA",X"BE",X"EB",X"7F",X"EF",X"63",X"02",X"02",X"43",X"E3",X"16",X"8B",X"52",X"FE",
		X"8A",X"CA",X"CE",X"FA",X"D3",X"4B",X"7B",X"6F",X"02",X"07",X"13",X"07",X"6E",X"B6",X"8E",X"B6",
		X"0A",X"0A",X"EE",X"42",X"6B",X"FB",X"DB",X"9F",X"02",X"17",X"13",X"BF",X"96",X"56",X"B6",X"66",
		X"02",X"03",X"87",X"8B",X"C6",X"CF",X"4E",X"9A",X"02",X"02",X"03",X"06",X"9F",X"BB",X"B7",X"7F",
		X"76",X"1E",X"5F",X"F7",X"F3",X"6A",X"26",X"8E",X"AB",X"E3",X"B7",X"5F",X"EE",X"BF",X"DF",X"FF",
		X"2B",X"9B",X"8E",X"32",X"A7",X"AB",X"4F",X"DE",X"FE",X"FF",X"FB",X"CF",X"7B",X"DF",X"FF",X"FF",
		X"BF",X"DE",X"A6",X"4F",X"BB",X"F3",X"FF",X"F7",X"4E",X"3B",X"DB",X"BB",X"F7",X"FF",X"FF",X"FF",
		X"FE",X"EA",X"4B",X"1B",X"CB",X"A7",X"FF",X"FB",X"B3",X"FF",X"B7",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"62",X"4E",X"D7",X"DE",X"FF",X"EF",X"4B",X"02",X"DF",X"F3",X"BE",X"7F",X"E6",X"3F",X"BE",X"FF",
		X"DE",X"B7",X"BF",X"B7",X"FF",X"DB",X"6A",X"02",X"AB",X"DA",X"63",X"CE",X"AB",X"A6",X"D7",X"FF",
		X"9F",X"B6",X"BB",X"9A",X"DF",X"B7",X"07",X"22",X"F7",X"CB",X"D6",X"67",X"72",X"7A",X"FF",X"FF",
		X"BE",X"D7",X"DF",X"6F",X"FA",X"7F",X"82",X"02",X"67",X"6B",X"6E",X"DA",X"2F",X"9A",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"1F",X"87",X"C3",X"F2",X"02",X"02",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"EB",X"3B",X"33",X"02",X"02",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FA",X"FA",X"9E",X"07",X"02",X"82",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"72",X"73",X"E3",X"E7",X"02",X"02",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"A2",X"F2",X"F3",X"DF",X"8E",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"83",X"0F",X"FF",X"FB",X"33",X"1F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"C7",X"FE",X"CE",X"5F",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"33",X"33",X"67",X"FF",X"D2",X"03",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"DF",X"83",X"07",X"C3",X"FB",X"FF",X"FF",X"E7",X"22",X"7E",X"FA",X"7E",X"4E",X"CF",X"EF",
		X"0A",X"F2",X"EF",X"83",X"02",X"0A",X"8F",X"AF",X"F7",X"0F",X"12",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"E7",X"E7",X"CF",X"DF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"F7",X"A6",X"02",
		X"CF",X"E3",X"7B",X"7F",X"3F",X"BF",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FB",X"77",X"E7",X"62",
		X"C2",X"F2",X"F2",X"FE",X"FF",X"FE",X"EA",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"B7",X"B7",
		X"F7",X"F3",X"37",X"1E",X"0E",X"27",X"FE",X"FE",X"FF",X"FF",X"FF",X"F7",X"F7",X"FB",X"DB",X"97",
		X"C3",X"C3",X"E2",X"72",X"B2",X"FB",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F6",X"E2",
		X"83",X"C7",X"C3",X"FB",X"7E",X"3E",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"F7",X"E7",
		X"F2",X"FA",X"FA",X"FA",X"FB",X"F3",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"86",X"83",X"C3",X"C3",X"87",X"9F",X"9F",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"8A",X"8A",X"8A",X"82",X"82",X"82",X"C2",X"C2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6A",X"62",X"62",X"7E",X"6E",X"6F",X"EF",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"16",X"12",X"02",X"02",X"03",X"03",X"83",X"83",X"EB",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CB",X"AB",X"1B",X"03",X"1B",X"9B",X"9B",X"8B",X"37",X"57",X"E7",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"7F",X"FE",X"7B",X"7E",X"7A",X"F6",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"5B",X"DB",X"FA",X"DE",X"CA",X"AA",X"C2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"82",X"AB",X"AA",X"EA",X"CB",X"CA",X"8A",X"8A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"66",X"66",X"62",X"62",X"6A",X"6A",X"6A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CA",X"63",X"6A",X"4A",X"02",X"22",X"02",X"02",X"B7",X"DE",X"D7",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"43",X"57",X"92",X"0B",X"92",X"87",X"A3",X"53",X"BF",X"AB",X"6F",X"F7",X"6F",X"7B",X"5F",X"AF",
		X"7E",X"FF",X"7B",X"73",X"FF",X"F7",X"7B",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"32",X"96",X"83",X"AB",X"BF",X"7A",X"9A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AE",X"8A",X"9A",X"92",X"D2",X"92",X"92",X"92",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"2F",X"2B",X"23",X"62",X"6A",X"63",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"46",X"23",X"8B",X"23",X"0A",X"12",X"82",X"82",X"BB",X"DE",X"76",X"FE",X"F7",X"EF",X"7F",X"FF",
		X"AB",X"32",X"43",X"E3",X"A7",X"83",X"B7",X"62",X"57",X"CF",X"BF",X"1F",X"5B",X"7F",X"4B",X"9F",
		X"FE",X"F6",X"7F",X"FF",X"FF",X"FF",X"FB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B7",X"6F",X"47",X"D2",X"52",X"7A",X"F3",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"43",X"62",X"EA",X"4A",X"4A",X"0E",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"13",X"13",X"1B",X"57",X"46",X"46",X"47",X"86",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"BE",X"FF",
		X"86",X"02",X"62",X"23",X"07",X"A6",X"EA",X"96",X"FB",X"FF",X"BF",X"DE",X"FA",X"DB",X"97",X"EB",
		X"13",X"83",X"13",X"17",X"43",X"AB",X"63",X"2F",X"EF",X"7F",X"EF",X"EB",X"BF",X"57",X"9F",X"D3",
		X"FA",X"FE",X"FA",X"FF",X"FE",X"F7",X"F7",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"56",X"DA",X"7A",X"D2",X"E2",X"96",X"E6",X"D6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"52",X"12",X"B2",X"6A",X"AA",X"A2",X"A2",X"63",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"12",X"33",X"23",X"2B",X"A3",X"06",X"02",X"02",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"03",X"2B",X"03",X"83",X"82",X"12",X"02",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"EF",X"FF",
		X"83",X"83",X"23",X"83",X"03",X"03",X"83",X"23",X"FF",X"FF",X"DF",X"7F",X"FF",X"FF",X"7F",X"DF",
		X"F7",X"F7",X"F7",X"F7",X"FB",X"FB",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"F7",X"D7",X"97",X"57",X"B6",X"66",X"4E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CB",X"CB",X"CB",X"CB",X"4F",X"4F",X"1E",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CA",X"CA",X"8A",X"8B",X"1A",X"2A",X"2A",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EE",X"6A",X"4E",X"07",X"42",X"4A",X"4B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2B",X"2B",X"2F",X"AB",X"0B",X"03",X"0B",X"4B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"02",X"02",X"02",X"82",X"02",X"82",X"D2",X"02",X"02",X"02",X"02",X"02",X"E2",X"72",X"2A",
		X"1A",X"DF",X"83",X"07",X"83",X"BB",X"FF",X"FF",X"E7",X"22",X"7E",X"FA",X"7E",X"C6",X"C7",X"D7",
		X"0A",X"72",X"EF",X"83",X"42",X"62",X"E2",X"F3",X"F7",X"0F",X"12",X"7E",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"DF",X"83",X"07",X"83",X"BB",X"FF",X"FF",X"E7",X"22",X"7E",X"FA",X"FE",X"C6",X"C3",X"CB",
		X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",X"2F",
		X"E2",X"22",X"02",X"E2",X"02",X"E2",X"E2",X"E2",X"5F",X"DF",X"FF",X"1F",X"FF",X"1F",X"DF",X"DF",
		X"FF",X"FE",X"FA",X"FF",X"FA",X"FF",X"FF",X"FF",X"2E",X"2F",X"2F",X"2A",X"2F",X"2A",X"2F",X"2F",
		X"06",X"03",X"7F",X"FF",X"8F",X"7F",X"7F",X"7F",X"06",X"0F",X"7F",X"BF",X"FF",X"0B",X"0B",X"0F",
		X"03",X"07",X"07",X"73",X"33",X"03",X"03",X"07",X"02",X"0E",X"1E",X"0E",X"0F",X"1F",X"07",X"07",
		X"C2",X"C2",X"82",X"82",X"82",X"02",X"02",X"E2",X"FE",X"FE",X"FE",X"FE",X"FE",X"FA",X"F2",X"E2",
		X"02",X"02",X"02",X"06",X"0E",X"0E",X"1E",X"1E",X"07",X"0F",X"0F",X"0B",X"03",X"02",X"02",X"02",
		X"02",X"02",X"02",X"32",X"72",X"7A",X"7A",X"3A",X"E2",X"F2",X"F2",X"CA",X"8A",X"02",X"02",X"02",
		X"3E",X"1E",X"1E",X"0E",X"0E",X"07",X"0F",X"1E",X"02",X"1E",X"02",X"0E",X"02",X"07",X"07",X"0A",
		X"3A",X"1A",X"1E",X"0E",X"0E",X"0E",X"1E",X"3E",X"02",X"1A",X"02",X"0E",X"02",X"0E",X"0A",X"16",
		X"03",X"03",X"0E",X"3A",X"62",X"02",X"02",X"02",X"02",X"03",X"0E",X"3A",X"62",X"02",X"02",X"02",
		X"7F",X"BE",X"BE",X"3E",X"1E",X"0A",X"06",X"0F",X"0F",X"67",X"67",X"E7",X"77",X"3F",X"0F",X"0F",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"C2",X"02",X"82",X"82",X"82",X"82",X"82",X"C2",X"C2",
		X"02",X"02",X"72",X"FA",X"F2",X"72",X"3A",X"3E",X"0F",X"3F",X"0F",X"07",X"03",X"72",X"02",X"3E",
		X"02",X"02",X"02",X"02",X"22",X"E2",X"E2",X"E2",X"C2",X"E2",X"E2",X"E2",X"C2",X"02",X"02",X"02",
		X"1E",X"0E",X"06",X"0E",X"1E",X"02",X"02",X"02",X"02",X"0E",X"02",X"06",X"0A",X"02",X"02",X"02",
		X"E2",X"F2",X"F2",X"72",X"3A",X"1A",X"3A",X"7A",X"02",X"F2",X"02",X"72",X"02",X"1A",X"2A",X"32",
		X"03",X"03",X"03",X"03",X"06",X"0E",X"1A",X"12",X"02",X"02",X"03",X"03",X"06",X"0E",X"1A",X"12",
		X"02",X"02",X"72",X"FE",X"7E",X"7E",X"7F",X"3F",X"0F",X"3F",X"0F",X"03",X"07",X"0A",X"12",X"16",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"82",X"C2",X"E2",X"E2",X"C2",X"82",X"02",X"02",X"82",
		X"0F",X"03",X"03",X"03",X"03",X"02",X"02",X"02",X"07",X"03",X"02",X"03",X"03",X"02",X"02",X"02",
		X"E2",X"F2",X"E2",X"C2",X"02",X"02",X"02",X"02",X"A2",X"72",X"22",X"42",X"02",X"02",X"02",X"02",
		X"1E",X"0E",X"7F",X"FF",X"87",X"7F",X"7F",X"7F",X"1E",X"3E",X"7F",X"CF",X"FF",X"07",X"07",X"07",
		X"07",X"07",X"17",X"3F",X"3F",X"06",X"06",X"0F",X"3E",X"7E",X"EE",X"C7",X"47",X"7F",X"0F",X"0F",
		X"82",X"82",X"82",X"82",X"02",X"02",X"02",X"C2",X"FA",X"FE",X"FE",X"FE",X"FE",X"F2",X"E2",X"C2",
		X"03",X"03",X"1F",X"3F",X"7F",X"3F",X"02",X"03",X"06",X"0F",X"02",X"07",X"02",X"02",X"02",X"03",
		X"C2",X"E2",X"F2",X"FA",X"F2",X"E2",X"E2",X"E2",X"32",X"DA",X"2A",X"E2",X"02",X"E2",X"E2",X"62",
		X"02",X"02",X"02",X"02",X"02",X"0E",X"0E",X"0E",X"1F",X"1F",X"3F",X"3F",X"1E",X"02",X"02",X"02",
		X"42",X"E2",X"E2",X"E2",X"E2",X"E2",X"F2",X"7A",X"82",X"E2",X"02",X"E2",X"02",X"E2",X"E2",X"6A",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",X"3E",X"02",X"0E",X"02",X"0E",X"02",X"0E",X"0E",X"16",
		X"02",X"02",X"42",X"6E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"3F",X"13",X"03",X"02",X"02",X"06",
		X"3F",X"3B",X"32",X"72",X"72",X"E2",X"C2",X"02",X"3F",X"03",X"32",X"02",X"72",X"22",X"C2",X"02",
		X"02",X"02",X"02",X"02",X"02",X"E2",X"E2",X"E2",X"E2",X"F2",X"F2",X"F2",X"F2",X"02",X"02",X"02",
		X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",X"F2",X"FA",X"02",X"E2",X"02",X"E2",X"02",X"E2",X"A2",X"F2",
		X"07",X"07",X"0F",X"7F",X"FF",X"07",X"03",X"0F",X"0E",X"3E",X"32",X"02",X"02",X"1A",X"1E",X"0F",
		X"92",X"82",X"86",X"8E",X"0E",X"FE",X"FA",X"E2",X"F2",X"FA",X"FA",X"F2",X"F2",X"02",X"02",X"E2",
		X"03",X"03",X"07",X"07",X"07",X"07",X"07",X"03",X"03",X"03",X"07",X"07",X"07",X"07",X"3F",X"3F",
		X"82",X"C2",X"E2",X"E2",X"E2",X"E2",X"E2",X"C2",X"82",X"C2",X"E2",X"E2",X"E2",X"E2",X"E2",X"E2",
		X"03",X"03",X"03",X"02",X"02",X"02",X"06",X"03",X"3F",X"1F",X"1F",X"0F",X"07",X"07",X"07",X"0F",
		X"C2",X"C2",X"82",X"02",X"02",X"02",X"02",X"C2",X"F2",X"FA",X"FA",X"F2",X"E2",X"E2",X"E2",X"C2",
		X"12",X"1A",X"3E",X"7E",X"F2",X"E2",X"F2",X"72",X"0F",X"07",X"03",X"03",X"02",X"E2",X"22",X"52",
		X"3A",X"3A",X"1E",X"3A",X"72",X"02",X"02",X"02",X"22",X"1A",X"0E",X"1A",X"32",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"07",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",
		X"72",X"32",X"32",X"02",X"02",X"02",X"32",X"C2",X"FA",X"FA",X"F2",X"F2",X"F2",X"F2",X"F2",X"FA",
		X"02",X"02",X"02",X"06",X"0E",X"0F",X"0E",X"0E",X"03",X"03",X"07",X"03",X"03",X"02",X"02",X"02",
		X"02",X"06",X"06",X"0E",X"1A",X"3A",X"3A",X"3E",X"FA",X"FA",X"FE",X"F2",X"FA",X"22",X"32",X"3E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"1E",X"3E",X"02",X"0E",X"02",X"0E",X"02",X"0E",X"0E",X"16",X"02",
		X"07",X"03",X"03",X"03",X"33",X"7B",X"73",X"63",X"06",X"02",X"1E",X"3E",X"0E",X"06",X"06",X"07",
		X"FA",X"FA",X"FA",X"FA",X"C2",X"C6",X"CE",X"FE",X"3A",X"2A",X"2A",X"3A",X"7E",X"7A",X"72",X"02",
		X"63",X"E2",X"E2",X"1E",X"3F",X"3F",X"1E",X"02",X"03",X"07",X"0F",X"03",X"02",X"02",X"02",X"02",
		X"FE",X"9E",X"1E",X"3E",X"3E",X"72",X"7A",X"02",X"02",X"62",X"FE",X"C2",X"3A",X"62",X"72",X"02",
		X"1E",X"26",X"63",X"63",X"63",X"32",X"1E",X"02",X"1E",X"26",X"63",X"63",X"63",X"32",X"1E",X"02",
		X"0E",X"1E",X"0E",X"0E",X"0E",X"0E",X"3F",X"02",X"0E",X"1E",X"0E",X"0E",X"0E",X"0E",X"3F",X"02",
		X"3E",X"63",X"07",X"1E",X"3E",X"72",X"7F",X"02",X"3E",X"63",X"07",X"1E",X"3E",X"72",X"7F",X"02",
		X"3F",X"06",X"0E",X"1E",X"03",X"63",X"3E",X"02",X"3F",X"06",X"0E",X"1E",X"03",X"63",X"3E",X"02",
		X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"02",X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"02",
		X"7E",X"62",X"7E",X"03",X"03",X"63",X"3E",X"02",X"7E",X"62",X"7E",X"03",X"03",X"63",X"3E",X"02",
		X"1E",X"32",X"62",X"7E",X"63",X"63",X"3E",X"02",X"1E",X"32",X"62",X"7E",X"63",X"63",X"3E",X"02",
		X"7F",X"63",X"06",X"0E",X"1A",X"1A",X"1A",X"02",X"7F",X"63",X"06",X"0E",X"1A",X"1A",X"1A",X"02",
		X"3E",X"62",X"72",X"3E",X"4F",X"43",X"3E",X"02",X"3E",X"62",X"72",X"3E",X"4F",X"43",X"3E",X"02",
		X"3E",X"63",X"63",X"3F",X"03",X"06",X"3E",X"02",X"3E",X"63",X"63",X"3F",X"03",X"06",X"3E",X"02",
		X"7E",X"63",X"63",X"63",X"7E",X"62",X"62",X"02",X"7E",X"63",X"63",X"63",X"7E",X"62",X"62",X"02",
		X"1E",X"36",X"63",X"63",X"7F",X"63",X"63",X"02",X"1E",X"36",X"63",X"63",X"7F",X"63",X"63",X"02",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"02",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"02",
		X"3E",X"66",X"62",X"3E",X"03",X"63",X"3E",X"02",X"3E",X"66",X"62",X"3E",X"03",X"63",X"3E",X"02",
		X"3F",X"32",X"32",X"3E",X"32",X"32",X"3F",X"02",X"3F",X"32",X"32",X"3E",X"32",X"32",X"3F",X"02",
		X"02",X"46",X"2A",X"12",X"2A",X"46",X"02",X"02",X"02",X"46",X"2A",X"12",X"2A",X"46",X"02",X"02",
		X"02",X"0E",X"3F",X"7F",X"7F",X"7F",X"BF",X"BE",X"02",X"0E",X"3E",X"7E",X"7F",X"7F",X"FF",X"FF",
		X"03",X"03",X"EA",X"FE",X"E2",X"BE",X"7F",X"7F",X"02",X"1E",X"FF",X"3F",X"7F",X"C3",X"82",X"82",
		X"E2",X"F2",X"3A",X"1E",X"3F",X"3F",X"FF",X"FF",X"02",X"72",X"82",X"DE",X"C2",X"C2",X"02",X"02",
		X"02",X"02",X"02",X"02",X"03",X"C3",X"FF",X"FF",X"02",X"02",X"02",X"02",X"03",X"03",X"2B",X"2F",
		X"62",X"E2",X"F2",X"1A",X"0E",X"06",X"03",X"03",X"02",X"02",X"12",X"1A",X"0E",X"06",X"03",X"03",
		X"83",X"C3",X"E3",X"E2",X"76",X"36",X"1E",X"1A",X"03",X"03",X"03",X"02",X"06",X"06",X"06",X"02",
		X"02",X"32",X"3A",X"3A",X"3A",X"3A",X"32",X"72",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"E2",X"E2",X"32",X"1A",X"0E",X"06",X"03",X"03",X"02",X"02",X"32",X"1A",X"0E",X"06",X"03",X"03",
		X"03",X"07",X"07",X"0E",X"1E",X"3A",X"E2",X"C2",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"C2",X"62",X"32",X"1A",X"0E",X"06",X"02",X"02",X"C0",X"60",X"30",X"18",X"0C",X"04",X"00",X"00",
		X"80",X"E0",X"38",X"0E",X"03",X"07",X"07",X"03",X"80",X"E0",X"38",X"0E",X"03",X"00",X"00",X"00",
		X"03",X"03",X"03",X"03",X"03",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"FC",X"7C",X"1C",X"78",X"E0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"03",X"03",X"03",X"7F",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"02",X"02",X"03",X"03",X"00",X"00",X"02",X"02",X"02",X"00",X"00",X"00",
		X"07",X"FF",X"06",X"06",X"06",X"06",X"07",X"07",X"00",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"78",X"2C",X"26",X"63",X"E1",X"C0",X"00",X"00",X"18",X"0C",X"06",X"03",X"01",X"00",
		X"07",X"FF",X"0E",X"0C",X"1C",X"1C",X"1C",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"3C",X"2E",X"27",X"63",X"40",X"C0",X"80",X"00",X"00",X"20",X"20",X"60",X"40",X"C0",X"80",
		X"00",X"06",X"03",X"7F",X"FF",X"8F",X"7F",X"7F",X"00",X"06",X"0F",X"7F",X"BF",X"FF",X"0B",X"0B",
		X"18",X"1C",X"1E",X"0E",X"1E",X"FC",X"E0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"70",X"78",X"78",X"F8",X"F8",X"F8",X"F8",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"F8",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"07",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"FF",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",
		X"10",X"80",X"00",X"44",X"20",X"21",X"70",X"FA",X"10",X"00",X"00",X"44",X"00",X"00",X"40",X"F2",
		X"01",X"40",X"00",X"27",X"4E",X"5C",X"FC",X"FE",X"01",X"00",X"00",X"20",X"02",X"04",X"4C",X"FE",
		X"00",X"10",X"00",X"00",X"00",X"00",X"3C",X"7E",X"10",X"10",X"10",X"10",X"10",X"10",X"3C",X"7E",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"20",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"7D",X"18",X"50",
		X"FC",X"FC",X"7E",X"3E",X"1E",X"02",X"06",X"0C",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"79",X"02",
		X"0F",X"0E",X"1E",X"3C",X"3D",X"7D",X"3D",X"3C",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",
		X"0E",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"0F",X"03",X"07",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"3E",X"1C",X"28",X"70",X"FF",X"FF",X"FF",X"FF",X"3E",X"1C",X"14",X"08",
		X"03",X"06",X"1C",X"19",X"13",X"07",X"0F",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"1F",X"3F",X"7F",
		X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",X"80",
		X"1F",X"3F",X"3E",X"1E",X"0E",X"0C",X"38",X"A0",X"7F",X"FF",X"FE",X"FE",X"7E",X"3C",X"00",X"58",
		X"06",X"0C",X"3C",X"39",X"31",X"13",X"01",X"00",X"1F",X"7F",X"7F",X"7F",X"3F",X"1F",X"0F",X"0F",
		X"30",X"F8",X"FC",X"FC",X"FE",X"FF",X"FE",X"FC",X"F0",X"F8",X"FC",X"FC",X"FF",X"FE",X"FD",X"FA",
		X"00",X"00",X"00",X"F9",X"F1",X"FF",X"7F",X"7F",X"00",X"00",X"00",X"7F",X"1F",X"61",X"80",X"80",
		X"00",X"20",X"78",X"FE",X"00",X"FF",X"FF",X"FF",X"30",X"7C",X"FE",X"FF",X"FF",X"FF",X"1F",X"07",
		X"00",X"00",X"00",X"00",X"01",X"82",X"FD",X"FC",X"00",X"00",X"00",X"80",X"C0",X"F9",X"FE",X"FF",
		X"04",X"0C",X"18",X"30",X"60",X"00",X"00",X"00",X"04",X"0C",X"18",X"30",X"60",X"00",X"00",X"00",
		X"07",X"07",X"0E",X"0E",X"1C",X"1C",X"1C",X"3C",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",
		X"20",X"20",X"20",X"2C",X"0C",X"18",X"38",X"20",X"04",X"04",X"0C",X"10",X"34",X"20",X"18",X"00",
		X"0F",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"07",X"03",X"03",X"43",X"43",X"43",X"C3",X"C3",
		X"46",X"46",X"46",X"46",X"46",X"46",X"46",X"46",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"00",X"00",X"00",X"00",X"3F",X"00",X"1F",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"1F",X"00",
		X"00",X"00",X"00",X"00",X"FC",X"00",X"FE",X"00",X"00",X"00",X"00",X"00",X"FF",X"03",X"FF",X"01",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"06",X"03",X"00",X"00",X"00",X"08",X"08",X"0C",X"06",X"03",
		X"F8",X"F0",X"F0",X"F0",X"F4",X"F0",X"FA",X"F8",X"F8",X"F0",X"00",X"40",X"74",X"10",X"02",X"00",
		X"A0",X"A2",X"67",X"47",X"4F",X"4E",X"1E",X"EC",X"7F",X"7E",X"FF",X"FF",X"FF",X"F2",X"F2",X"EC",
		X"0C",X"1E",X"1E",X"0C",X"00",X"00",X"00",X"00",X"08",X"0E",X"1C",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"18",X"1C",X"1C",X"0E",X"00",X"00",X"00",X"0A",X"17",X"0B",X"17",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"30",X"10",X"98",X"C8",X"00",X"00",X"00",X"20",X"30",X"10",X"98",X"C8",
		X"4C",X"64",X"26",X"32",X"12",X"18",X"08",X"08",X"4C",X"64",X"26",X"33",X"13",X"18",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"18",
		X"08",X"0C",X"04",X"06",X"02",X"03",X"01",X"01",X"08",X"0C",X"04",X"06",X"02",X"03",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"F8",X"F0",X"08",X"18",X"08",X"8C",X"46",X"02",
		X"00",X"03",X"07",X"07",X"03",X"03",X"03",X"01",X"00",X"03",X"07",X"05",X"01",X"00",X"00",X"00",
		X"00",X"1F",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"1F",X"FF",X"FF",X"7F",X"7F",X"3F",X"00",
		X"18",X"18",X"98",X"D8",X"98",X"98",X"30",X"30",X"00",X"20",X"B8",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"18",X"1F",X"0F",X"0F",X"07",X"03",X"03",X"0F",X"0F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",
		X"60",X"40",X"C0",X"E0",X"F0",X"F0",X"FE",X"FF",X"E0",X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",X"F8",
		X"01",X"03",X"07",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"12",X"14",X"01",X"01",X"03",X"03",X"03",X"07",X"0E",X"28",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"01",X"00",X"00",X"00",X"00",X"80",X"40",X"21",X"06",
		X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"7F",X"1F",X"1F",X"0F",X"40",X"80",X"00",X"00",X"30",X"1F",
		X"F8",X"F8",X"F8",X"FC",X"FE",X"FE",X"FC",X"F5",X"80",X"08",X"38",X"C0",X"00",X"01",X"03",X"0A",
		X"00",X"0C",X"3F",X"7F",X"7F",X"7F",X"BF",X"A0",X"00",X"0C",X"3E",X"7E",X"7F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"C1",X"81",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"3F",X"7F",X"FF",X"FF",X"FF",
		X"30",X"7C",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"18",X"64",X"00",X"1C",X"E7",X"E7",
		X"00",X"00",X"00",X"80",X"C1",X"FA",X"FD",X"FC",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"83",
		X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"03",X"07",X"07",X"00",X"00",X"07",X"07",X"03",
		X"06",X"07",X"03",X"83",X"03",X"03",X"07",X"23",X"C0",X"E0",X"F3",X"73",X"F3",X"F3",X"EF",X"FF",
		X"00",X"00",X"00",X"01",X"01",X"02",X"14",X"1F",X"0F",X"1F",X"3F",X"3F",X"3F",X"1F",X"0F",X"07",
		X"41",X"40",X"80",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"1F",X"1F",X"1F",X"1E",X"3E",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F8",X"F8",X"7C",X"3C",X"3C",
		X"1C",X"1E",X"0E",X"0E",X"06",X"03",X"07",X"1F",X"1C",X"1E",X"0E",X"0E",X"06",X"03",X"05",X"0B",
		X"1C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0E",X"1F",X"1C",X"1C",X"1C",X"0C",X"0C",X"0C",X"0C",X"1A",
		X"00",X"00",X"00",X"80",X"00",X"00",X"08",X"18",X"C0",X"E0",X"F0",X"70",X"F0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"31",X"31",X"12",X"04",X"07",X"07",X"0F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"3C",X"4C",X"8C",X"0E",X"06",X"00",X"00",X"E0",X"E4",X"FC",X"FE",X"FE",X"FE",X"FE",X"F0",X"E0",
		X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"70",X"F0",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"01",X"61",X"62",X"3F",X"3F",X"07",X"0F",X"0F",X"1F",X"1F",X"1F",X"07",X"0F",
		X"20",X"40",X"80",X"00",X"00",X"00",X"E0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"01",X"07",X"1F",X"FC",X"7F",X"03",X"07",X"07",X"07",X"07",X"1F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"0F",X"13",X"27",X"27",X"47",X"47",X"42",X"7E",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"7E",
		X"00",X"00",X"60",X"70",X"38",X"3C",X"1C",X"0E",X"3F",X"7F",X"7F",X"7F",X"3F",X"3C",X"1C",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"E0",X"F0",X"F0",X"F0",X"F0",X"F8",X"78",X"3C",
		X"06",X"0E",X"3E",X"00",X"00",X"00",X"00",X"00",X"06",X"0E",X"3E",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"1C",X"0E",X"0E",X"06",X"07",X"0E",X"18",X"1C",X"1C",X"0E",X"0E",X"06",X"03",X"06",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"3C",X"3F",X"3F",X"7F",X"7E",X"FC",X"F8",X"F8",X"FC",
		X"3E",X"0F",X"07",X"03",X"07",X"0E",X"00",X"00",X"3E",X"0F",X"07",X"03",X"03",X"04",X"00",X"00",
		X"00",X"00",X"00",X"04",X"07",X"03",X"00",X"00",X"03",X"07",X"0F",X"0B",X"08",X"0C",X"07",X"03",
		X"00",X"00",X"00",X"20",X"E8",X"CC",X"0C",X"0C",X"C0",X"E0",X"F0",X"D0",X"10",X"30",X"E0",X"CC",
		X"00",X"00",X"00",X"01",X"12",X"0A",X"0C",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",
		X"2E",X"4E",X"8E",X"06",X"00",X"00",X"00",X"E0",X"FE",X"FE",X"FE",X"FE",X"FC",X"F0",X"E0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",X"0F",X"1F",X"1F",X"3F",X"3E",X"3C",X"3C",X"1C",
		X"1C",X"0E",X"0E",X"06",X"0E",X"1E",X"00",X"00",X"1C",X"0E",X"0E",X"06",X"06",X"1A",X"00",X"00",
		X"0F",X"1F",X"1D",X"38",X"30",X"70",X"F0",X"00",X"0F",X"1F",X"1D",X"38",X"30",X"30",X"50",X"00",
		X"C0",X"E0",X"E0",X"78",X"18",X"38",X"70",X"00",X"C0",X"E0",X"E0",X"78",X"18",X"18",X"30",X"00",
		X"08",X"08",X"24",X"C0",X"03",X"24",X"10",X"10",X"18",X"18",X"3C",X"FF",X"FF",X"3C",X"18",X"18",
		X"20",X"40",X"80",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",
		X"3F",X"3E",X"60",X"00",X"00",X"00",X"00",X"00",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"00",X"02",X"04",X"04",X"07",X"FF",X"FF",X"FF",X"0F",X"07",X"07",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",
		X"03",X"06",X"0C",X"00",X"00",X"00",X"00",X"00",X"03",X"06",X"0C",X"00",X"20",X"60",X"40",X"00",
		X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"C0",X"08",X"18",X"10",X"30",X"20",X"60",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"20",X"60",X"40",X"C0",X"00",X"00",X"00",X"00",X"20",X"60",X"40",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"18",X"0C",X"0C",X"06",X"04",X"00",X"00",X"00",X"26",X"73",X"F3",X"F9",X"FB",X"7F",X"3E",
		X"00",X"00",X"F0",X"0C",X"02",X"00",X"01",X"01",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0C",X"1E",X"0F",X"00",X"00",X"F8",X"FC",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"E7",X"FB",
		X"00",X"00",X"00",X"00",X"01",X"63",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"E1",X"FE",X"FF",
		X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",
		X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",
		X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",
		X"00",X"00",X"08",X"38",X"1C",X"10",X"00",X"00",X"00",X"00",X"08",X"38",X"1C",X"10",X"00",X"00",
		X"00",X"00",X"24",X"18",X"18",X"24",X"00",X"00",X"00",X"00",X"24",X"18",X"18",X"24",X"00",X"00",
		X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"1F",X"00",X"00",X"00",X"08",X"04",X"02",X"01",X"1F",
		X"00",X"00",X"80",X"80",X"88",X"90",X"A0",X"C0",X"00",X"00",X"80",X"80",X"88",X"90",X"A0",X"C0",
		X"00",X"00",X"00",X"09",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"09",X"07",X"03",X"00",X"00",
		X"38",X"38",X"78",X"F0",X"E0",X"C0",X"00",X"00",X"38",X"38",X"78",X"F0",X"E0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"20",X"10",X"18",X"18",X"18",X"00",X"00",X"00",X"20",X"10",X"18",X"18",X"18",
		X"00",X"00",X"38",X"7C",X"7C",X"7C",X"7C",X"38",X"00",X"00",X"08",X"04",X"04",X"04",X"4C",X"38",
		X"07",X"0F",X"0F",X"07",X"00",X"00",X"00",X"00",X"07",X"0F",X"1F",X"0F",X"06",X"00",X"00",X"00",
		X"E0",X"F8",X"78",X"38",X"10",X"00",X"00",X"00",X"F0",X"F8",X"F8",X"78",X"30",X"00",X"00",X"00",
		X"07",X"0E",X"1F",X"3E",X"3F",X"1F",X"0F",X"77",X"07",X"0E",X"3F",X"7F",X"7F",X"7F",X"3F",X"7F",
		X"78",X"FC",X"FE",X"7C",X"B8",X"DE",X"DF",X"FE",X"78",X"FC",X"FE",X"FE",X"FC",X"FE",X"FF",X"FF",
		X"7F",X"7B",X"77",X"37",X"1B",X"0F",X"06",X"00",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1E",X"0C",
		X"FC",X"D8",X"BC",X"FE",X"FE",X"7C",X"38",X"00",X"FF",X"FE",X"FC",X"FE",X"FE",X"FE",X"FC",X"38",
		X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",X"1F",
		X"00",X"00",X"00",X"18",X"99",X"18",X"00",X"00",X"00",X"00",X"00",X"66",X"E7",X"66",X"00",X"00",
		X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"01",X"00",X"3C",X"0C",X"0C",X"3C",X"18",X"3E",X"7E",
		X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",
		X"18",X"08",X"3C",X"3C",X"7C",X"38",X"10",X"82",X"18",X"18",X"3C",X"34",X"64",X"00",X"6C",X"7C",
		X"00",X"00",X"03",X"03",X"81",X"61",X"18",X"06",X"03",X"07",X"04",X"04",X"86",X"62",X"1B",X"07",
		X"00",X"00",X"00",X"60",X"40",X"10",X"30",X"00",X"00",X"80",X"E0",X"90",X"B8",X"E8",X"C8",X"C0",
		X"80",X"30",X"18",X"00",X"00",X"00",X"00",X"00",X"F8",X"4C",X"64",X"3A",X"01",X"00",X"00",X"00",
		X"00",X"00",X"80",X"60",X"18",X"04",X"02",X"39",X"00",X"00",X"80",X"60",X"18",X"04",X"7A",X"C7",
		X"60",X"08",X"12",X"06",X"00",X"00",X"00",X"00",X"9F",X"F7",X"EC",X"78",X"38",X"00",X"00",X"00",
		X"00",X"00",X"40",X"60",X"20",X"00",X"00",X"00",X"C0",X"F0",X"BC",X"9A",X"D1",X"60",X"00",X"00",
		X"00",X"20",X"12",X"04",X"20",X"48",X"04",X"00",X"00",X"62",X"36",X"1C",X"38",X"6C",X"46",X"00",
		X"0F",X"07",X"00",X"00",X"00",X"0C",X"1F",X"3F",X"09",X"0F",X"0F",X"07",X"07",X"0F",X"1F",X"3F",
		X"F8",X"F0",X"30",X"78",X"7C",X"7E",X"3E",X"9C",X"9C",X"FC",X"FC",X"FC",X"FC",X"FE",X"3E",X"9C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0B",X"00",X"00",X"00",X"07",X"0F",X"0F",X"09",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"B8",X"00",X"00",X"00",X"F0",X"F8",X"FC",X"9C",X"DC",
		X"0F",X"27",X"30",X"38",X"38",X"3C",X"1E",X"00",X"09",X"2F",X"3F",X"3F",X"3F",X"3F",X"1E",X"00",
		X"F8",X"F0",X"00",X"00",X"00",X"1C",X"3E",X"3F",X"9C",X"FC",X"FC",X"FC",X"FC",X"FC",X"3E",X"3F",
		X"00",X"01",X"03",X"07",X"07",X"07",X"07",X"03",X"07",X"0F",X"1F",X"3E",X"3C",X"1C",X"0C",X"00",
		X"60",X"30",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"FC",X"FF",X"3F",X"3F",X"3E",X"3E",X"3C",
		X"03",X"63",X"F3",X"F2",X"72",X"3A",X"18",X"07",X"3E",X"7E",X"3E",X"3F",X"7F",X"3F",X"1F",X"07",
		X"A0",X"A2",X"67",X"47",X"4F",X"4E",X"1C",X"E0",X"7F",X"7E",X"FC",X"FC",X"FF",X"FE",X"FC",X"E0",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"3F",X"00",X"10",X"12",X"32",X"22",X"22",X"02",X"02",
		X"F0",X"F8",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"10",X"18",X"04",X"02",X"02",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"3F",X"3F",X"3F",X"13",X"28",X"02",X"02",X"02",X"02",X"03",X"01",X"0D",X"14",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"F0",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"8C",X"0E",
		X"06",X"77",X"FB",X"FF",X"7F",X"7E",X"7C",X"39",X"06",X"7F",X"FF",X"BF",X"3F",X"1B",X"1B",X"0F",
		X"00",X"06",X"8E",X"9C",X"3C",X"7C",X"FC",X"F8",X"00",X"20",X"E0",X"D8",X"FC",X"FC",X"FC",X"F8",
		X"1B",X"1B",X"0B",X"09",X"04",X"02",X"01",X"0F",X"0F",X"2F",X"3F",X"3F",X"1F",X"1F",X"0E",X"0E",
		X"F0",X"E0",X"C0",X"80",X"00",X"00",X"FE",X"FF",X"F0",X"E0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"06",X"0C",X"08",X"18",X"88",X"8C",X"46",X"01",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"40",X"60",X"10",X"08",X"04",X"04",X"02",X"02",
		X"FF",X"FF",X"7F",X"7F",X"3E",X"3E",X"08",X"50",X"01",X"00",X"00",X"00",X"00",X"00",X"14",X"2C",
		X"00",X"03",X"07",X"07",X"C3",X"E3",X"FB",X"FD",X"00",X"03",X"07",X"05",X"01",X"60",X"F8",X"FC",
		X"30",X"B8",X"DC",X"FC",X"FC",X"FC",X"F8",X"E0",X"30",X"F9",X"FD",X"FD",X"FF",X"DF",X"DE",X"7E",
		X"FF",X"7F",X"3F",X"0F",X"03",X"02",X"07",X"0F",X"FF",X"7F",X"3F",X"0F",X"03",X"03",X"07",X"03",
		X"00",X"80",X"C0",X"C0",X"C0",X"80",X"0F",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F0",X"F0",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"20",X"A0",X"A0",X"E0",X"C0",X"C0",X"80",
		X"20",X"2C",X"1E",X"1E",X"3E",X"7E",X"FF",X"FF",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"FC",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"F9",X"F1",X"03",X"02",X"00",X"00",X"02",X"03",
		X"1F",X"3F",X"3F",X"3F",X"1F",X"0B",X"20",X"50",X"00",X"00",X"00",X"00",X"00",X"04",X"1C",X"28",
		X"F8",X"F0",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"08",X"18",X"11",X"11",X"11",X"01",X"01",
		X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",X"00",X"08",X"08",X"0C",X"04",X"04",X"02",X"02",
		X"1F",X"0F",X"0F",X"07",X"01",X"02",X"00",X"00",X"01",X"00",X"09",X"03",X"03",X"05",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FC",X"68",X"10",X"80",X"80",X"80",X"80",X"82",X"40",X"50",X"2C",
		X"06",X"77",X"FB",X"FF",X"7F",X"7F",X"7F",X"3C",X"06",X"7F",X"FF",X"BF",X"3F",X"1B",X"1B",X"0F",
		X"60",X"40",X"80",X"80",X"3C",X"7C",X"FC",X"F8",X"00",X"60",X"E0",X"C0",X"FC",X"FC",X"FC",X"F8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"7F",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",
		X"10",X"10",X"10",X"10",X"10",X"10",X"F7",X"00",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"F7",X"00",
		X"1C",X"3F",X"7F",X"7F",X"EF",X"ED",X"A9",X"28",X"63",X"40",X"00",X"00",X"10",X"12",X"56",X"00",
		X"13",X"37",X"FF",X"DF",X"FF",X"FD",X"FF",X"FF",X"6C",X"48",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"8F",X"EF",X"FD",X"FF",X"FF",X"FF",X"FF",X"7A",X"70",X"10",X"00",X"00",X"00",X"00",X"00",
		X"8D",X"DF",X"FD",X"FF",X"DF",X"FF",X"FF",X"FF",X"72",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C3",X"E7",X"FF",X"DF",X"FD",X"FF",X"FF",X"FF",X"3C",X"18",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"70",X"04",X"00",X"50",X"FF",X"FF",X"73",X"20",X"8F",X"FB",X"FF",X"AF",
		X"FF",X"FF",X"FF",X"9F",X"07",X"53",X"80",X"00",X"FF",X"9F",X"0F",X"63",X"F9",X"AC",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"F8",X"E0",X"82",X"2E",X"04",X"FF",X"FD",X"F0",X"C7",X"1F",X"7D",X"D1",X"FB",
		X"FF",X"FF",X"FF",X"E7",X"00",X"0C",X"1C",X"00",X"FF",X"E7",X"42",X"18",X"FF",X"F3",X"E3",X"FF",
		X"30",X"1D",X"06",X"10",X"40",X"E0",X"F9",X"FF",X"CF",X"E2",X"F9",X"EF",X"BF",X"1F",X"06",X"00",
		X"88",X"01",X"00",X"48",X"18",X"BE",X"FE",X"FF",X"77",X"FE",X"FF",X"B7",X"E7",X"41",X"01",X"00",
		X"80",X"90",X"E8",X"20",X"04",X"0C",X"5F",X"FF",X"7F",X"6F",X"17",X"DF",X"FB",X"F3",X"A0",X"00",
		X"60",X"EC",X"70",X"01",X"08",X"DC",X"FF",X"FF",X"9F",X"13",X"8F",X"FE",X"F7",X"23",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"38",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"60",X"C0",X"80",X"82",X"02",X"06",X"3E",X"00",X"83",X"1D",X"3D",X"3C",X"7C",X"78",X"80",X"C1",
		X"00",X"07",X"3D",X"00",X"00",X"00",X"10",X"10",X"FF",X"F8",X"00",X"C2",X"F7",X"F7",X"E7",X"E7",
		X"00",X"00",X"02",X"02",X"06",X"04",X"1C",X"08",X"DB",X"BC",X"7C",X"7C",X"78",X"B9",X"C1",X"E3",
		X"10",X"20",X"C0",X"42",X"03",X"0C",X"00",X"00",X"E7",X"CB",X"1D",X"1C",X"BC",X"C0",X"F3",X"F7",
		X"1E",X"3F",X"7F",X"FF",X"FF",X"ED",X"23",X"01",X"FF",X"FF",X"FF",X"FF",X"F5",X"A1",X"F1",X"F7",
		X"00",X"00",X"02",X"C2",X"F3",X"FF",X"FF",X"FF",X"DB",X"BC",X"7C",X"FC",X"FD",X"FF",X"FF",X"FF",
		X"10",X"20",X"C4",X"76",X"BF",X"EF",X"FD",X"FF",X"E7",X"CB",X"19",X"3A",X"BF",X"EF",X"FF",X"FF",
		X"00",X"00",X"00",X"06",X"CE",X"FB",X"EF",X"FF",X"E3",X"DD",X"BD",X"BC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"07",X"3D",X"0E",X"1F",X"7F",X"EF",X"FF",X"FF",X"F8",X"00",X"CE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"DD",X"00",X"DD",X"00",X"00",X"DD",X"DD",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",
		X"FF",X"80",X"80",X"80",X"FF",X"08",X"08",X"08",X"FF",X"80",X"80",X"80",X"FF",X"08",X"08",X"08",
		X"FF",X"FF",X"FF",X"F7",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"10",X"10",
		X"99",X"FF",X"99",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"99",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"FF",X"00",X"DD",X"00",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",
		X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"5E",X"C3",X"81",X"81",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"7D",X"7C",X"38",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"40",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"30",X"20",X"00",X"00",X"00",X"00",X"00",X"21",X"81",X"81",X"81",X"81",X"85",X"85",X"DD",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"A0",X"B0",X"B8",X"D8",X"E0",X"F8",X"FC",
		X"60",X"FC",X"FD",X"FD",X"FF",X"7F",X"7F",X"70",X"9D",X"1D",X"7D",X"FD",X"FF",X"DF",X"8F",X"8F",
		X"00",X"00",X"00",X"00",X"07",X"18",X"24",X"2E",X"FC",X"FC",X"FE",X"FE",X"F8",X"E7",X"DB",X"D1",
		X"20",X"20",X"20",X"30",X"30",X"30",X"3C",X"3C",X"DF",X"DF",X"DF",X"EF",X"EF",X"EF",X"F3",X"F3",
		X"46",X"4E",X"42",X"40",X"44",X"4C",X"2C",X"2C",X"B9",X"B1",X"BD",X"BE",X"B8",X"B0",X"D0",X"D2",
		X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"30",X"F0",X"F0",X"F0",X"F0",X"B0",X"B0",X"B0",X"B0",
		X"12",X"0D",X"00",X"00",X"C2",X"20",X"02",X"84",X"EC",X"F2",X"FF",X"FF",X"3D",X"DF",X"FC",X"7A",
		X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",X"1C",X"26",X"63",X"63",X"63",X"32",X"1C",X"00",
		X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",X"0C",X"1C",X"0C",X"0C",X"0C",X"0C",X"3F",X"00",
		X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",X"3E",X"63",X"07",X"1E",X"3C",X"70",X"7F",X"00",
		X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",X"3F",X"06",X"0C",X"1E",X"03",X"63",X"3E",X"00",
		X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",X"0E",X"1E",X"36",X"66",X"7F",X"06",X"06",X"00",
		X"7E",X"60",X"7E",X"03",X"03",X"63",X"3E",X"00",X"7E",X"60",X"7E",X"03",X"03",X"63",X"3E",X"00",
		X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",X"1E",X"30",X"60",X"7E",X"63",X"63",X"3E",X"00",
		X"7F",X"63",X"06",X"0C",X"18",X"18",X"18",X"00",X"7F",X"63",X"06",X"0C",X"18",X"18",X"18",X"00",
		X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",X"3C",X"62",X"72",X"3C",X"4F",X"43",X"3E",X"00",
		X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",X"3E",X"63",X"63",X"3F",X"03",X"06",X"3C",X"00",
		X"81",X"81",X"81",X"81",X"81",X"81",X"01",X"01",X"81",X"81",X"81",X"81",X"81",X"81",X"01",X"01",
		X"3F",X"3F",X"3F",X"0F",X"0F",X"07",X"03",X"00",X"C4",X"E2",X"CA",X"F2",X"F4",X"FC",X"FC",X"FF",
		X"00",X"00",X"80",X"80",X"E0",X"E0",X"FD",X"7F",X"00",X"00",X"00",X"00",X"80",X"00",X"3C",X"B9",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"01",X"00",X"00",X"01",X"02",X"06",X"0A",X"0D",X"02",
		X"0D",X"0C",X"10",X"19",X"1B",X"1B",X"3F",X"3F",X"12",X"13",X"0F",X"27",X"27",X"27",X"07",X"07",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",X"1C",X"36",X"63",X"63",X"7F",X"63",X"63",X"00",
		X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",X"7E",X"63",X"63",X"7E",X"63",X"63",X"7E",X"00",
		X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",X"00",X"1E",X"33",X"60",X"60",X"60",X"33",X"1E",X"00",
		X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",X"7C",X"66",X"63",X"63",X"63",X"66",X"7C",X"00",
		X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",X"3F",X"30",X"30",X"3E",X"30",X"30",X"3F",X"00",
		X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",X"7F",X"60",X"60",X"7E",X"60",X"60",X"60",X"00",
		X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",X"00",X"1F",X"30",X"60",X"67",X"63",X"33",X"1F",X"00",
		X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",X"63",X"63",X"63",X"7F",X"63",X"63",X"63",X"00",
		X"1E",X"0C",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",X"1E",X"0C",X"0C",X"0C",X"0C",X"0C",X"1E",X"00",
		X"03",X"03",X"03",X"03",X"03",X"63",X"3E",X"00",X"03",X"03",X"03",X"03",X"03",X"63",X"3E",X"00",
		X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",X"00",X"63",X"66",X"6C",X"78",X"7C",X"6E",X"67",X"00",
		X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"00",X"30",X"30",X"30",X"30",X"30",X"30",X"3F",X"00",
		X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",X"63",X"77",X"7F",X"7F",X"6B",X"63",X"63",X"00",
		X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",X"63",X"73",X"7B",X"7F",X"6F",X"67",X"63",X"00",
		X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"3E",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",
		X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",X"7E",X"63",X"63",X"63",X"7E",X"60",X"60",X"00",
		X"3E",X"63",X"63",X"63",X"6F",X"66",X"3D",X"00",X"3E",X"63",X"63",X"63",X"6F",X"66",X"3D",X"00",
		X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",X"7E",X"63",X"63",X"67",X"7C",X"6E",X"67",X"00",
		X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",X"3C",X"66",X"60",X"3E",X"03",X"63",X"3E",X"00",
		X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"3F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",
		X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",X"63",X"63",X"63",X"63",X"63",X"63",X"3E",X"00",
		X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",X"63",X"63",X"63",X"77",X"3E",X"1C",X"08",X"00",
		X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",X"63",X"63",X"6B",X"7F",X"7F",X"36",X"22",X"00",
		X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",X"63",X"77",X"3E",X"1C",X"3E",X"77",X"63",X"00",
		X"33",X"33",X"12",X"1E",X"0C",X"0C",X"0C",X"00",X"33",X"33",X"12",X"1E",X"0C",X"0C",X"0C",X"00",
		X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",X"7F",X"07",X"0E",X"1C",X"38",X"70",X"7F",X"00",
		X"24",X"24",X"24",X"00",X"00",X"00",X"00",X"00",X"24",X"24",X"24",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",
		X"7F",X"00",X"3E",X"63",X"63",X"63",X"3E",X"00",X"7F",X"00",X"3E",X"63",X"63",X"63",X"3E",X"00",
		X"3C",X"42",X"99",X"A1",X"A1",X"99",X"42",X"3C",X"3C",X"42",X"99",X"A1",X"A1",X"99",X"42",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"63",X"3E",X"30",X"03",X"3F",X"3F",X"30",X"00",X"80",X"C1",X"CF",X"FC",X"C0",X"C0",X"CF",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"3E",X"30",X"8C",X"CE",X"66",X"60",X"C1",X"F9",X"C1",X"CF",X"73",X"31",X"19",X"1F",X"3E",
		X"00",X"C0",X"60",X"30",X"18",X"08",X"18",X"3F",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"E0",X"C8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"78",X"F8",X"D0",X"B0",X"61",X"20",X"C0",X"93",X"B7",X"67",X"4F",X"0F",X"9E",X"DF",X"3F",
		X"C0",X"60",X"23",X"26",X"6C",X"E8",X"69",X"33",X"00",X"80",X"C0",X"C1",X"83",X"27",X"86",X"CC",
		X"7E",X"40",X"60",X"71",X"7F",X"3F",X"1F",X"02",X"01",X"3F",X"1F",X"4E",X"60",X"3E",X"1C",X"01",
		X"0D",X"38",X"D0",X"CD",X"D0",X"42",X"32",X"00",X"F2",X"C7",X"2F",X"B2",X"2F",X"BD",X"CD",X"FF",
		X"02",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"01",X"00",X"02",X"03",X"01",X"00",X"00",X"00",
		X"01",X"73",X"FB",X"FE",X"DC",X"0F",X"07",X"07",X"FE",X"8D",X"24",X"F1",X"DB",X"08",X"07",X"07",
		X"9C",X"F0",X"E0",X"C6",X"1C",X"3C",X"38",X"30",X"63",X"0F",X"5F",X"39",X"E3",X"C3",X"C7",X"CF",
		X"17",X"17",X"72",X"78",X"3C",X"1F",X"1E",X"FC",X"E8",X"E8",X"8D",X"97",X"C3",X"E8",X"E9",X"03",
		X"E1",X"C7",X"8F",X"3F",X"FD",X"FB",X"E6",X"84",X"1E",X"B8",X"73",X"C7",X"1C",X"78",X"E1",X"83",
		X"F9",X"F3",X"E7",X"CF",X"9E",X"3C",X"78",X"F0",X"66",X"CC",X"99",X"33",X"66",X"CC",X"98",X"30",
		X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"30",X"18",X"0C",X"04",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",
		X"05",X"07",X"06",X"0C",X"19",X"3F",X"7F",X"F7",X"F8",X"F8",X"F9",X"F3",X"E6",X"C8",X"9F",X"37",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"07",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",
		X"0C",X"08",X"18",X"10",X"30",X"61",X"41",X"CC",X"03",X"07",X"07",X"0F",X"0F",X"1E",X"3E",X"33",
		X"9C",X"3D",X"79",X"F9",X"E9",X"C9",X"89",X"09",X"63",X"C2",X"96",X"36",X"66",X"C6",X"86",X"06",
		X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"34",X"16",X"17",X"77",X"F3",X"F1",X"C0",X"FF",X"C3",X"E1",X"E4",X"86",X"33",X"F1",X"40",X"00",
		X"38",X"0C",X"06",X"83",X"82",X"C3",X"FF",X"C3",X"C0",X"F0",X"F8",X"7C",X"7D",X"3C",X"81",X"3D",
		X"90",X"80",X"80",X"C1",X"FF",X"FF",X"7E",X"0D",X"6F",X"7F",X"7F",X"3E",X"80",X"FC",X"79",X"02",
		X"02",X"06",X"4E",X"DE",X"8C",X"4C",X"E7",X"83",X"FC",X"F8",X"B2",X"26",X"74",X"B0",X"18",X"7C",
		X"18",X"30",X"20",X"30",X"3F",X"3F",X"1F",X"00",X"07",X"0F",X"1F",X"0F",X"20",X"3F",X"1F",X"00",
		X"13",X"31",X"71",X"FB",X"FF",X"DF",X"8E",X"00",X"EC",X"CE",X"8E",X"24",X"71",X"DF",X"8E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"9C",X"C6",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"38",
		X"00",X"00",X"00",X"07",X"04",X"04",X"FE",X"8C",X"00",X"00",X"00",X"00",X"03",X"03",X"01",X"73",
		X"C3",X"E2",X"60",X"C1",X"03",X"10",X"E1",X"E3",X"BC",X"9D",X"1F",X"3E",X"FC",X"EF",X"1E",X"9C",
		X"C4",X"61",X"E0",X"03",X"9F",X"8F",X"CE",X"C6",X"3B",X"9E",X"1F",X"FC",X"62",X"76",X"37",X"B9",
		X"C7",X"43",X"C6",X"8F",X"98",X"90",X"84",X"1C",X"B9",X"3D",X"38",X"70",X"67",X"6F",X"7B",X"E3",
		X"E0",X"79",X"71",X"F1",X"65",X"05",X"4D",X"CD",X"9F",X"46",X"6E",X"0E",X"9A",X"FA",X"B2",X"32",
		X"19",X"99",X"CB",X"C3",X"E6",X"7F",X"7F",X"3F",X"E6",X"66",X"34",X"BC",X"99",X"40",X"7F",X"3F",
		X"DC",X"9C",X"3C",X"76",X"F7",X"E7",X"C3",X"81",X"23",X"6B",X"CB",X"91",X"34",X"66",X"C3",X"81",
		X"09",X"09",X"09",X"09",X"0D",X"0F",X"0F",X"07",X"06",X"06",X"06",X"06",X"02",X"08",X"0F",X"07",
		X"00",X"00",X"00",X"80",X"E0",X"30",X"10",X"30",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"C0",
		X"F0",X"98",X"08",X"8C",X"04",X"1C",X"3C",X"7C",X"10",X"60",X"F0",X"70",X"F8",X"E0",X"CC",X"80",
		X"F4",X"F4",X"F4",X"A4",X"24",X"24",X"64",X"C4",X"28",X"68",X"C8",X"98",X"18",X"18",X"18",X"38",
		X"C6",X"42",X"03",X"01",X"03",X"FF",X"FF",X"FE",X"38",X"BC",X"FC",X"FE",X"FC",X"01",X"FF",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"F0",X"EF",X"83",X"02",X"80",X"C0",X"DA",X"F7",X"0F",X"10",X"7C",X"FD",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"07",X"00",X"00",X"00",X"00",X"1F",X"3F",X"79",X"38",
		X"00",X"03",X"87",X"80",X"E7",X"EC",X"78",X"71",X"00",X"00",X"78",X"7F",X"18",X"13",X"87",X"8E",
		X"F8",X"F0",X"D8",X"1E",X"17",X"03",X"06",X"02",X"00",X"0C",X"27",X"E1",X"E8",X"FC",X"F9",X"FD",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"3C",
		X"04",X"1F",X"1F",X"3C",X"00",X"BE",X"FF",X"70",X"1B",X"00",X"00",X"03",X"3F",X"41",X"00",X"8F",
		X"FF",X"3F",X"F0",X"13",X"03",X"4F",X"BA",X"FC",X"00",X"C0",X"0F",X"EE",X"FE",X"BC",X"4D",X"33",
		X"00",X"00",X"00",X"F8",X"FB",X"4F",X"01",X"04",X"C0",X"F8",X"FC",X"06",X"04",X"B0",X"FE",X"FA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"07",X"1F",
		X"7C",X"07",X"03",X"27",X"FF",X"7F",X"F5",X"E0",X"83",X"F8",X"FD",X"D9",X"07",X"8F",X"3F",X"FF",
		X"E0",X"F8",X"FE",X"BF",X"7F",X"8F",X"EE",X"60",X"7F",X"F7",X"C1",X"C7",X"99",X"FC",X"F1",X"FF",
		X"06",X"00",X"08",X"FC",X"F8",X"98",X"38",X"1F",X"FF",X"FF",X"FF",X"F3",X"07",X"67",X"C7",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"FE",X"FF",X"F0",X"E0",X"F8",X"FC",X"0C",
		X"00",X"A0",X"E3",X"8F",X"F8",X"F0",X"E8",X"FF",X"FF",X"5F",X"1C",X"70",X"1F",X"FF",X"FF",X"FF",
		X"01",X"01",X"C9",X"FF",X"7D",X"38",X"1C",X"FC",X"FF",X"FF",X"3F",X"FF",X"FE",X"FF",X"E3",X"03",
		X"E0",X"A0",X"E0",X"F0",X"FF",X"7F",X"3F",X"7F",X"FF",X"FF",X"9F",X"0F",X"00",X"80",X"C0",X"80",
		X"1A",X"DF",X"83",X"07",X"81",X"BB",X"FE",X"3E",X"E5",X"20",X"7C",X"F8",X"7E",X"44",X"01",X"C1",
		X"08",X"F0",X"E6",X"83",X"02",X"00",X"00",X"00",X"F7",X"0F",X"19",X"7C",X"FD",X"FF",X"FF",X"FF",
		X"78",X"00",X"20",X"1F",X"06",X"E3",X"63",X"1E",X"86",X"FF",X"DF",X"E0",X"F8",X"1C",X"9C",X"E0",
		X"3F",X"0F",X"9F",X"C5",X"F8",X"F0",X"F0",X"E0",X"F0",X"F0",X"E0",X"FA",X"85",X"08",X"00",X"00",
		X"E2",X"F0",X"BF",X"1F",X"0A",X"10",X"36",X"00",X"1D",X"0F",X"40",X"E0",X"F5",X"E7",X"00",X"00",
		X"D1",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"2E",X"7F",X"FF",X"F7",X"E0",X"C0",X"00",X"00",
		X"FC",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"E0",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"0F",X"12",X"00",X"00",X"00",X"00",X"00",X"F5",X"F0",X"6C",X"3C",X"10",X"00",X"00",X"00",
		X"8C",X"F8",X"F0",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"77",X"3F",X"1F",X"03",X"0F",X"1F",X"3F",X"1E",X"08",X"40",X"E0",
		X"BF",X"9F",X"0D",X"1F",X"31",X"71",X"E0",X"80",X"4C",X"63",X"F2",X"E0",X"CE",X"8E",X"1F",X"7F",
		X"F8",X"FC",X"FF",X"F9",X"DF",X"8E",X"0C",X"3F",X"07",X"03",X"20",X"36",X"38",X"79",X"FB",X"C4",
		X"01",X"01",X"07",X"01",X"E3",X"FF",X"4D",X"01",X"00",X"06",X"18",X"7E",X"1C",X"00",X"32",X"7E",
		X"83",X"E7",X"FB",X"C0",X"9F",X"FF",X"FF",X"FF",X"7C",X"18",X"04",X"3F",X"7F",X"F0",X"00",X"00",
		X"38",X"7C",X"C0",X"E0",X"F3",X"EF",X"9E",X"FC",X"C7",X"83",X"3F",X"1F",X"FF",X"17",X"61",X"03",
		X"3F",X"6E",X"FC",X"1E",X"0F",X"FF",X"F9",X"71",X"C2",X"97",X"07",X"E3",X"F3",X"AB",X"96",X"9F",
		X"0E",X"FF",X"C3",X"09",X"CD",X"F9",X"F3",X"FF",X"F1",X"00",X"3C",X"F6",X"32",X"86",X"8C",X"C0",
		X"01",X"03",X"03",X"01",X"03",X"00",X"00",X"00",X"3E",X"1C",X"1C",X"06",X"00",X"00",X"00",X"00",
		X"FF",X"F1",X"E0",X"F8",X"FE",X"13",X"3F",X"FE",X"07",X"0F",X"1F",X"07",X"01",X"EC",X"C0",X"01",
		X"FF",X"FF",X"7E",X"1F",X"0F",X"9F",X"BF",X"FF",X"F0",X"F8",X"FF",X"FF",X"FF",X"6F",X"43",X"00",
		X"8F",X"7F",X"06",X"C0",X"FF",X"FF",X"FF",X"FF",X"70",X"80",X"F9",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"00",X"03",X"1E",X"09",X"07",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"00",X"00",X"00",X"00",
		X"67",X"C3",X"C2",X"80",X"0C",X"00",X"00",X"00",X"98",X"3C",X"3D",X"7F",X"F3",X"CF",X"03",X"00",
		X"00",X"C2",X"AA",X"BE",X"EB",X"7D",X"ED",X"63",X"00",X"00",X"41",X"E1",X"14",X"8B",X"52",X"FE",
		X"8A",X"CA",X"CE",X"FA",X"D3",X"49",X"79",X"6D",X"02",X"07",X"13",X"07",X"6C",X"B6",X"8E",X"B6",
		X"0A",X"0A",X"EE",X"42",X"6B",X"F9",X"D9",X"9D",X"00",X"15",X"11",X"BD",X"96",X"56",X"B6",X"66",
		X"00",X"03",X"87",X"8B",X"C6",X"CD",X"4E",X"9A",X"00",X"00",X"01",X"04",X"9D",X"BB",X"B5",X"7D",
		X"76",X"1E",X"5D",X"F7",X"F3",X"6A",X"24",X"8E",X"AB",X"E3",X"B7",X"5F",X"EE",X"BF",X"DF",X"FF",
		X"2B",X"9B",X"8E",X"32",X"A5",X"AB",X"4D",X"DC",X"FE",X"FF",X"F9",X"CD",X"7B",X"DF",X"FF",X"FF",
		X"BF",X"DE",X"A6",X"4D",X"BB",X"F1",X"FF",X"F7",X"4C",X"39",X"D9",X"BB",X"F7",X"FF",X"FF",X"FF",
		X"FC",X"EA",X"49",X"19",X"CB",X"A7",X"FF",X"FB",X"B3",X"FD",X"B7",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"62",X"4E",X"D7",X"DE",X"FF",X"ED",X"49",X"00",X"DF",X"F3",X"BE",X"7D",X"E4",X"3F",X"BE",X"FF",
		X"DE",X"B7",X"BD",X"B7",X"FF",X"DB",X"6A",X"02",X"A9",X"DA",X"63",X"CC",X"A9",X"A6",X"D5",X"FF",
		X"9F",X"B6",X"BB",X"9A",X"DF",X"B5",X"05",X"20",X"F5",X"C9",X"D6",X"67",X"72",X"7A",X"FF",X"FF",
		X"BE",X"D7",X"DD",X"6F",X"FA",X"7F",X"82",X"00",X"65",X"69",X"6E",X"DA",X"2F",X"98",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"1F",X"87",X"C1",X"F0",X"00",X"00",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CF",X"EB",X"3B",X"33",X"00",X"00",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"F8",X"9E",X"07",X"00",X"82",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"70",X"71",X"E1",X"E5",X"00",X"02",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F3",X"A0",X"F0",X"F3",X"DF",X"8E",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"81",X"0F",X"FF",X"F9",X"31",X"1F",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"83",X"C7",X"FE",X"CC",X"5F",X"FF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"33",X"67",X"FD",X"D0",X"03",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1A",X"DF",X"83",X"07",X"C1",X"FB",X"FF",X"FF",X"E5",X"20",X"7C",X"F8",X"7E",X"4C",X"CD",X"ED",
		X"08",X"F0",X"EF",X"83",X"02",X"08",X"8D",X"AF",X"F7",X"0F",X"10",X"7C",X"FD",X"FF",X"FF",X"FF",
		X"E7",X"E7",X"CF",X"DF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FB",X"F7",X"A4",X"00",
		X"CF",X"E3",X"79",X"7D",X"3F",X"BF",X"9F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FB",X"77",X"E7",X"62",
		X"C0",X"F0",X"F0",X"FE",X"FF",X"FC",X"E8",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"B7",X"B7",
		X"F7",X"F3",X"35",X"1C",X"0C",X"25",X"FE",X"FE",X"FF",X"FF",X"FF",X"F7",X"F7",X"FB",X"D9",X"95",
		X"C3",X"C1",X"E0",X"70",X"B0",X"F9",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F6",X"E2",
		X"83",X"C7",X"C3",X"F9",X"7C",X"3C",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"F7",X"E5",
		X"F2",X"F8",X"F8",X"F8",X"F9",X"F1",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"84",X"81",X"C1",X"C3",X"87",X"9F",X"9F",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"88",X"88",X"88",X"80",X"80",X"80",X"C0",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"68",X"60",X"60",X"7C",X"6E",X"6F",X"EF",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"14",X"10",X"00",X"00",X"01",X"01",X"83",X"83",X"EB",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CB",X"AB",X"1B",X"03",X"1B",X"99",X"99",X"8B",X"37",X"57",X"E7",X"FF",X"F7",X"FF",X"FF",X"FF",
		X"F7",X"7D",X"FE",X"79",X"7E",X"7A",X"F6",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"59",X"DB",X"FA",X"DE",X"CA",X"A8",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"82",X"A9",X"AA",X"EA",X"C9",X"C8",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"64",X"64",X"62",X"62",X"68",X"68",X"68",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C8",X"61",X"68",X"48",X"00",X"20",X"00",X"00",X"B7",X"DE",X"D7",X"F7",X"FF",X"FF",X"FF",X"FF",
		X"41",X"55",X"90",X"09",X"90",X"85",X"A3",X"53",X"BF",X"AB",X"6F",X"F7",X"6F",X"7B",X"5F",X"AF",
		X"7E",X"FF",X"7B",X"73",X"FF",X"F5",X"7B",X"7D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AA",X"32",X"96",X"83",X"AB",X"BF",X"7A",X"9A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AC",X"8A",X"9A",X"92",X"D2",X"92",X"92",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"2D",X"29",X"21",X"60",X"6A",X"63",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"21",X"89",X"21",X"08",X"12",X"82",X"80",X"BB",X"DE",X"76",X"FE",X"F7",X"ED",X"7D",X"FF",
		X"A9",X"30",X"41",X"E1",X"A5",X"81",X"B5",X"60",X"57",X"CF",X"BF",X"1F",X"5B",X"7F",X"4B",X"9F",
		X"FE",X"F6",X"7F",X"FF",X"FF",X"FF",X"FB",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B5",X"6D",X"45",X"D0",X"52",X"7A",X"F3",X"62",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"43",X"62",X"E8",X"4A",X"48",X"0C",X"28",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"11",X"19",X"55",X"44",X"44",X"45",X"84",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"BE",X"FF",
		X"84",X"00",X"60",X"21",X"05",X"A4",X"E8",X"94",X"FB",X"FF",X"BF",X"DE",X"FA",X"DB",X"97",X"EB",
		X"13",X"83",X"11",X"15",X"43",X"A9",X"61",X"2D",X"EF",X"7F",X"EF",X"EB",X"BF",X"57",X"9F",X"D3",
		X"F8",X"FE",X"FA",X"FF",X"FC",X"F7",X"F5",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"56",X"DA",X"7A",X"D0",X"E2",X"94",X"E6",X"D4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"50",X"10",X"B2",X"68",X"A8",X"A0",X"A0",X"61",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"12",X"33",X"23",X"29",X"A1",X"04",X"00",X"02",X"FF",X"FE",X"FF",X"F7",X"FF",X"FF",X"FF",X"FD",
		X"49",X"01",X"29",X"01",X"81",X"80",X"10",X"00",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"EF",X"FF",
		X"83",X"83",X"23",X"83",X"03",X"03",X"83",X"23",X"FF",X"FF",X"DF",X"7F",X"FF",X"FF",X"7F",X"DF",
		X"F5",X"F5",X"F5",X"F5",X"FB",X"FB",X"FD",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"F5",X"D5",X"95",X"55",X"B4",X"64",X"4C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CB",X"CB",X"C9",X"C9",X"4D",X"4D",X"1C",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CA",X"C8",X"8A",X"89",X"1A",X"2A",X"2A",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EE",X"6A",X"4C",X"05",X"40",X"48",X"49",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"2B",X"2B",X"2F",X"AB",X"0B",X"03",X"0B",X"4B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"D0",X"00",X"00",X"00",X"00",X"00",X"E0",X"70",X"28",
		X"18",X"DF",X"81",X"07",X"81",X"BB",X"FF",X"FF",X"E7",X"20",X"7E",X"F8",X"7E",X"C4",X"C5",X"D5",
		X"08",X"70",X"EF",X"83",X"42",X"60",X"E0",X"F1",X"F7",X"0F",X"10",X"7C",X"FD",X"FF",X"FF",X"FF",
		X"18",X"DF",X"83",X"07",X"81",X"BB",X"FF",X"FF",X"E7",X"20",X"7C",X"F8",X"FE",X"C4",X"C1",X"CB",
		X"00",X"03",X"03",X"07",X"07",X"0F",X"3F",X"3F",X"1F",X"1C",X"1C",X"18",X"18",X"71",X"43",X"C3",
		X"00",X"00",X"00",X"04",X"00",X"01",X"04",X"10",X"03",X"03",X"07",X"0B",X"0F",X"1E",X"1B",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
