library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity eprom_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of eprom_3 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"00",X"C0",X"E0",X"00",X"00",X"28",X"FE",X"FE",X"28",X"FE",X"FE",X"28",X"00",
		X"08",X"5C",X"54",X"FE",X"54",X"74",X"20",X"00",X"84",X"4A",X"24",X"10",X"48",X"A4",X"42",X"00",
		X"0A",X"04",X"6E",X"9A",X"B2",X"72",X"0C",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",
		X"00",X"00",X"82",X"C6",X"7C",X"38",X"00",X"00",X"00",X"38",X"7C",X"C6",X"82",X"00",X"00",X"00",
		X"00",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"10",X"10",X"7C",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"02",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"10",X"10",X"54",X"10",X"10",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"6C",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"6E",X"02",X"00",X"00",
		X"00",X"82",X"C6",X"6C",X"38",X"10",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"00",X"10",X"38",X"6C",X"C6",X"82",X"00",X"00",X"60",X"F0",X"DA",X"CA",X"CA",X"E0",X"60",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"82",X"82",X"FE",X"FE",X"00",X"00",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"0F",X"07",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"C0",X"60",X"70",X"58",X"5C",X"56",X"53",X"51",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"FF",X"60",X"30",X"18",X"0C",X"06",X"03",X"01",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"FF",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"5C",X"57",X"51",X"50",X"50",X"50",
		X"FF",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FE",X"FD",X"F4",X"FF",X"E4",X"D5",X"50",X"D0",X"70",X"58",X"4C",X"FE",X"46",X"57",
		X"10",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"C4",X"FF",X"C4",X"D5",X"C4",X"FF",X"C4",X"D5",X"45",X"FF",X"45",X"55",X"44",X"FF",X"44",X"55",
		X"02",X"03",X"81",X"81",X"81",X"81",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",
		X"C4",X"FF",X"E4",X"F5",X"F4",X"FF",X"FC",X"FF",X"45",X"FF",X"45",X"57",X"46",X"FE",X"4C",X"58",
		X"81",X"03",X"02",X"02",X"02",X"06",X"04",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"07",X"03",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"F0",X"D0",X"50",X"50",X"50",X"50",X"51",X"57",
		X"08",X"18",X"10",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5C",X"F0",X"FF",X"50",X"50",X"50",X"50",X"50",
		X"00",X"00",X"F0",X"18",X"0C",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"01",X"03",X"07",X"0F",X"50",X"50",X"F0",X"D0",X"D0",X"50",X"50",X"51",
		X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"53",X"56",X"5C",X"58",X"70",X"7F",X"50",X"50",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"50",X"50",X"50",X"FF",X"50",X"50",
		X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"50",X"50",X"50",X"50",X"50",X"7F",X"70",X"58",
		X"01",X"01",X"01",X"01",X"01",X"FD",X"18",X"30",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"00",X"5C",X"56",X"53",X"51",X"50",X"50",X"D0",X"50",
		X"60",X"C0",X"80",X"00",X"00",X"01",X"03",X"06",X"30",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"00",X"00",X"20",X"70",X"F8",X"FC",X"FE",X"FF",X"30",X"10",X"08",X"04",X"02",X"01",X"03",X"06",
		X"0C",X"18",X"30",X"70",X"D8",X"8C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"8C",X"D8",X"70",X"70",X"50",X"50",X"50",X"50",
		X"01",X"03",X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"51",X"50",X"50",X"50",X"50",X"50",X"50",X"50",
		X"80",X"C0",X"60",X"30",X"18",X"0C",X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"01",X"03",X"07",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"50",X"FF",X"01",X"03",X"06",X"8C",X"D8",X"70",
		X"01",X"FF",X"8C",X"06",X"03",X"01",X"03",X"06",X"80",X"C0",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"FF",X"7F",X"3F",X"1F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"DF",X"CF",X"87",X"FF",X"FF",X"70",X"50",X"50",X"50",X"50",X"51",X"50",X"50",
		X"0C",X"18",X"30",X"60",X"C0",X"80",X"C0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"50",X"50",X"50",X"50",X"FF",X"50",
		X"30",X"18",X"0C",X"06",X"03",X"01",X"FF",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"50",X"50",X"50",X"50",X"50",X"50",X"7F",X"70",
		X"01",X"01",X"01",X"01",X"01",X"01",X"FD",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",X"00",X"58",X"5C",X"56",X"53",X"51",X"50",X"50",X"D0",
		X"30",X"60",X"C0",X"80",X"00",X"00",X"01",X"03",X"60",X"30",X"18",X"30",X"60",X"C0",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"30",X"10",X"08",X"04",X"02",X"01",X"00",
		X"06",X"0C",X"18",X"30",X"60",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"80",X"80",X"FF",X"80",X"FF",X"00",
		X"FE",X"01",X"00",X"00",X"FF",X"FF",X"01",X"FE",X"AA",X"00",X"55",X"55",X"AA",X"AA",X"00",X"AA",
		X"3F",X"C0",X"80",X"80",X"FF",X"BF",X"C0",X"3F",X"52",X"53",X"50",X"58",X"5F",X"60",X"3F",X"00",
		X"B1",X"B1",X"52",X"7E",X"52",X"52",X"52",X"52",X"0C",X"B1",X"0C",X"B1",X"B1",X"B1",X"B1",X"B1",
		X"B1",X"B1",X"B1",X"B1",X"0C",X"B1",X"0C",X"B1",X"52",X"52",X"52",X"7E",X"72",X"B1",X"B1",X"B1",
		X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"52",X"00",X"3F",X"68",X"50",X"53",X"53",X"53",X"52",
		X"00",X"FF",X"80",X"80",X"FF",X"80",X"FF",X"00",X"FE",X"01",X"00",X"00",X"FF",X"FF",X"01",X"FE",
		X"AA",X"55",X"55",X"55",X"FF",X"FF",X"55",X"AA",X"3F",X"C0",X"80",X"80",X"FF",X"BF",X"C0",X"3F",
		X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"80",X"7F",X"20",X"20",X"FF",X"E0",X"7F",X"80",
		X"BF",X"00",X"40",X"40",X"BF",X"BF",X"00",X"BF",X"80",X"00",X"41",X"41",X"80",X"80",X"00",X"80",
		X"FE",X"00",X"01",X"01",X"FE",X"FE",X"00",X"FE",X"00",X"FF",X"02",X"02",X"FF",X"02",X"FF",X"00",
		X"E0",X"1F",X"08",X"08",X"FF",X"F8",X"1F",X"E0",X"2F",X"00",X"50",X"50",X"2F",X"2F",X"00",X"2F",
		X"FA",X"00",X"05",X"05",X"FA",X"FA",X"00",X"FA",X"03",X"FC",X"08",X"08",X"FF",X"0B",X"FC",X"03",
		X"F8",X"07",X"02",X"02",X"FF",X"FE",X"07",X"F8",X"0B",X"00",X"14",X"14",X"0B",X"0B",X"00",X"0B",
		X"E8",X"00",X"14",X"14",X"E8",X"E8",X"00",X"E8",X"0F",X"F0",X"20",X"20",X"FF",X"2F",X"F0",X"0F",
		X"FC",X"03",X"01",X"01",X"FF",X"FF",X"03",X"FC",X"1F",X"E0",X"40",X"40",X"FF",X"5F",X"E0",X"1F",
		X"05",X"00",X"CA",X"0A",X"15",X"05",X"00",X"05",X"00",X"00",X"C0",X"01",X"12",X"0C",X"00",X"00",
		X"D0",X"00",X"28",X"29",X"D2",X"D4",X"00",X"D0",X"05",X"00",X"1A",X"4A",X"85",X"05",X"00",X"05",
		X"00",X"00",X"10",X"48",X"84",X"01",X"00",X"00",X"D0",X"00",X"28",X"28",X"D4",X"D1",X"00",X"D0",
		X"05",X"00",X"0A",X"1A",X"25",X"C5",X"00",X"05",X"00",X"00",X"0C",X"10",X"21",X"C0",X"00",X"00",
		X"D0",X"00",X"2C",X"28",X"D1",X"D0",X"00",X"D0",X"05",X"00",X"0A",X"8A",X"45",X"15",X"00",X"05",
		X"00",X"00",X"01",X"84",X"48",X"10",X"00",X"00",X"D0",X"00",X"29",X"2C",X"D0",X"D0",X"00",X"D0",
		X"B9",X"B9",X"5A",X"7E",X"52",X"52",X"52",X"52",X"1C",X"B9",X"1C",X"B9",X"B9",X"B9",X"B9",X"B9",
		X"B9",X"B9",X"B9",X"B9",X"1C",X"B9",X"1C",X"B9",X"52",X"52",X"52",X"7E",X"7A",X"B9",X"B9",X"B9",
		X"BD",X"BD",X"5A",X"7E",X"52",X"52",X"52",X"52",X"3C",X"BD",X"3C",X"BD",X"BD",X"BD",X"BD",X"BD",
		X"BD",X"BD",X"BD",X"BD",X"3C",X"BD",X"3C",X"BD",X"52",X"52",X"52",X"7E",X"7A",X"BD",X"BD",X"BD",
		X"FF",X"FF",X"7E",X"7E",X"52",X"52",X"52",X"52",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"52",X"52",X"52",X"7E",X"7E",X"FF",X"FF",X"FF",
		X"7E",X"7E",X"3C",X"7E",X"52",X"52",X"52",X"52",X"FF",X"7E",X"FF",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"FF",X"7E",X"FF",X"7E",X"52",X"52",X"52",X"7E",X"3C",X"7E",X"7E",X"7E",
		X"FF",X"FF",X"7E",X"7E",X"52",X"52",X"52",X"52",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"52",X"52",X"52",X"7E",X"7E",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"FF",X"FF",X"FF",X"83",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"FF",X"FF",X"C1",X"81",X"81",X"81",X"81",X"83",X"83",
		X"81",X"81",X"81",X"83",X"83",X"83",X"83",X"FF",X"FF",X"01",X"81",X"81",X"81",X"81",X"81",X"81",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"01",X"FF",X"FF",X"83",X"83",X"83",X"83",X"03",X"03",
		X"83",X"83",X"83",X"03",X"03",X"03",X"03",X"0F",X"FF",X"FF",X"83",X"83",X"83",X"83",X"83",X"83",
		X"18",X"2C",X"00",X"5C",X"5C",X"5C",X"5C",X"7E",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"7E",X"5C",X"5C",X"5C",X"5C",X"6E",X"2C",X"18",
		X"FF",X"DF",X"FF",X"BF",X"BF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"BF",X"BF",X"BF",X"DF",
		X"0E",X"5F",X"FF",X"BF",X"BE",X"7F",X"0F",X"0F",X"0F",X"0F",X"0E",X"7F",X"BF",X"BF",X"BE",X"50",
		X"FF",X"DF",X"FF",X"BF",X"BF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"BF",X"BF",X"BF",X"DF",
		X"3C",X"1C",X"08",X"00",X"07",X"0F",X"1F",X"3F",X"03",X"07",X"0F",X"1F",X"FF",X"EF",X"C7",X"C3",
		X"3C",X"1C",X"08",X"00",X"07",X"0F",X"1F",X"3F",X"03",X"07",X"0F",X"1F",X"FF",X"EF",X"C7",X"C3",
		X"7F",X"1F",X"07",X"01",X"03",X"07",X"0F",X"1F",X"81",X"87",X"1E",X"7E",X"3C",X"1C",X"08",X"00",
		X"7F",X"1F",X"07",X"01",X"03",X"07",X"0F",X"1F",X"81",X"87",X"1E",X"7E",X"3C",X"1C",X"08",X"00",
		X"FF",X"EF",X"C7",X"C3",X"81",X"87",X"1E",X"7E",X"07",X"0F",X"1F",X"3F",X"7F",X"1F",X"07",X"01",
		X"FF",X"EF",X"C7",X"C3",X"81",X"87",X"1E",X"7E",X"07",X"0F",X"1F",X"3F",X"7F",X"1F",X"07",X"01",
		X"28",X"24",X"E1",X"31",X"13",X"D6",X"16",X"16",X"66",X"DE",X"90",X"20",X"2F",X"48",X"48",X"52",
		X"0C",X"08",X"46",X"66",X"24",X"04",X"64",X"E4",X"80",X"98",X"19",X"10",X"9C",X"9B",X"90",X"84",
		X"32",X"E2",X"41",X"49",X"88",X"92",X"83",X"00",X"52",X"63",X"38",X"80",X"C6",X"39",X"00",X"06",
		X"06",X"02",X"33",X"B1",X"81",X"CC",X"06",X"33",X"46",X"67",X"30",X"98",X"CC",X"60",X"20",X"02",
		X"1C",X"36",X"33",X"A1",X"E1",X"26",X"1C",X"00",X"26",X"21",X"23",X"3E",X"E0",X"60",X"64",X"C4",
		X"70",X"E0",X"86",X"06",X"60",X"70",X"C0",X"93",X"73",X"30",X"0C",X"CE",X"E3",X"00",X"7C",X"1E",
		X"C0",X"18",X"1C",X"CC",X"03",X"33",X"36",X"30",X"9E",X"92",X"C2",X"40",X"1F",X"71",X"60",X"60",
		X"93",X"49",X"40",X"12",X"13",X"71",X"6C",X"5C",X"8F",X"E0",X"70",X"37",X"8F",X"06",X"F2",X"C2",
		X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"AF",X"FF",X"01",X"7F",X"7F",X"FF",X"60",X"6F",X"6F",
		X"FB",X"39",X"FF",X"FF",X"FF",X"00",X"FF",X"F1",X"D7",X"52",X"FF",X"FF",X"FF",X"13",X"D7",X"D7",
		X"AF",X"AF",X"EF",X"EF",X"EF",X"E4",X"BF",X"84",X"FF",X"EF",X"EF",X"EF",X"EF",X"EF",X"EF",X"AF",
		X"FF",X"DF",X"FF",X"DF",X"EF",X"F5",X"FF",X"FF",X"F7",X"56",X"57",X"57",X"DF",X"DF",X"D0",X"77",
		X"FF",X"80",X"FF",X"BF",X"FF",X"BF",X"86",X"B7",X"AF",X"AF",X"AF",X"AF",X"A8",X"AB",X"AB",X"BD",
		X"FF",X"FF",X"FF",X"FF",X"4D",X"5F",X"59",X"FF",X"D7",X"7F",X"D7",X"D7",X"57",X"F7",X"57",X"D7",
		X"B7",X"FA",X"FF",X"FF",X"FE",X"AF",X"AF",X"FF",X"AF",X"A5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DB",X"3F",X"FB",X"FB",X"3B",X"FB",X"FB",X"FB",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"00",X"DD",X"EA",X"EE",X"E8",X"EB",X"08",X"FF",X"3F",X"BE",
		X"FF",X"FF",X"20",X"AE",X"20",X"FF",X"E0",X"3B",X"EF",X"EF",X"AF",X"AF",X"A0",X"FF",X"00",X"FF",
		X"DD",X"DD",X"DD",X"DD",X"1D",X"FF",X"BF",X"BF",X"BE",X"BE",X"BF",X"BF",X"BE",X"FB",X"FF",X"F7",
		X"CC",X"77",X"9B",X"ED",X"75",X"D6",X"FA",X"EA",X"0F",X"EF",X"0F",X"BF",X"8F",X"EF",X"88",X"BA",
		X"BF",X"BF",X"03",X"FA",X"FB",X"FA",X"FB",X"FA",X"F7",X"F7",X"FF",X"3B",X"7E",X"3F",X"FF",X"BE",
		X"E8",X"EF",X"FA",X"D6",X"75",X"ED",X"9B",X"77",X"82",X"FA",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"3E",X"FA",X"0A",X"EE",X"EA",X"EA",X"EE",X"EA",
		X"CF",X"DF",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FA",X"0A",X"EA",X"E8",X"EF",X"EF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"24",X"12",X"01",X"01",X"19",X"A1",X"00",X"73",X"21",X"01",X"82",X"80",X"00",X"02",X"00",
		X"00",X"63",X"21",X"25",X"C4",X"00",X"01",X"03",X"00",X"80",X"80",X"A0",X"A4",X"78",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"05",X"1F",X"A1",X"00",X"7F",X"25",X"25",X"A2",X"80",X"00",X"23",X"21",
		X"25",X"67",X"25",X"25",X"FC",X"24",X"21",X"03",X"00",X"A0",X"A7",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"24",X"7E",X"A5",X"A5",X"7F",X"A5",X"00",X"FF",X"A5",X"25",X"FF",X"81",X"81",X"FB",X"A1",
		X"25",X"F7",X"25",X"A5",X"FD",X"A4",X"21",X"67",X"00",X"A5",X"EF",X"A5",X"A5",X"7A",X"24",X"18",
		X"18",X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"18",
		X"00",X"08",X"00",X"58",X"58",X"00",X"58",X"7E",X"00",X"58",X"58",X"00",X"58",X"58",X"00",X"58",
		X"58",X"00",X"58",X"58",X"00",X"58",X"58",X"00",X"7E",X"58",X"00",X"58",X"58",X"00",X"08",X"00",
		X"18",X"2C",X"00",X"5C",X"5C",X"5C",X"5C",X"7E",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"7E",X"5C",X"5C",X"5C",X"5C",X"6E",X"2C",X"18",
		X"00",X"00",X"00",X"18",X"2C",X"00",X"5C",X"5C",X"58",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"5C",X"5C",X"6E",X"2C",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"18",X"2C",X"00",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"6E",X"2C",X"18",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",
		X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"59",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"7E",X"59",X"59",X"59",X"59",X"5F",X"59",X"59",X"59",
		X"59",X"59",X"59",X"5F",X"59",X"59",X"59",X"59",X"30",X"30",X"10",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"7E",X"51",X"51",X"51",X"51",X"50",X"59",X"59",X"59",
		X"59",X"59",X"59",X"50",X"51",X"51",X"51",X"51",X"30",X"30",X"30",X"30",X"10",X"08",X"00",X"00",
		X"00",X"18",X"30",X"30",X"30",X"30",X"30",X"7E",X"59",X"59",X"59",X"59",X"5F",X"59",X"59",X"59",
		X"59",X"59",X"59",X"5F",X"59",X"59",X"59",X"59",X"30",X"30",X"30",X"30",X"30",X"10",X"08",X"00",
		X"00",X"08",X"3E",X"78",X"38",X"38",X"38",X"7E",X"59",X"59",X"59",X"59",X"5F",X"59",X"59",X"59",
		X"59",X"59",X"59",X"5F",X"59",X"59",X"59",X"59",X"7E",X"38",X"38",X"38",X"78",X"3E",X"08",X"04",
		X"00",X"00",X"1C",X"38",X"70",X"34",X"34",X"7E",X"59",X"59",X"59",X"59",X"5E",X"59",X"59",X"59",
		X"59",X"59",X"59",X"5E",X"59",X"59",X"59",X"59",X"7E",X"34",X"34",X"70",X"78",X"2C",X"14",X"08",
		X"00",X"00",X"1E",X"3E",X"7C",X"3C",X"3C",X"7E",X"59",X"59",X"59",X"59",X"5E",X"59",X"59",X"59",
		X"59",X"59",X"59",X"5E",X"59",X"59",X"59",X"59",X"7E",X"3C",X"3C",X"7C",X"7E",X"2E",X"14",X"08",
		X"18",X"2C",X"20",X"7C",X"5E",X"5D",X"5C",X"7E",X"79",X"59",X"59",X"59",X"5D",X"5F",X"59",X"59",
		X"59",X"59",X"79",X"D9",X"79",X"59",X"5B",X"5D",X"7E",X"5C",X"5C",X"7E",X"5C",X"6E",X"2C",X"18",
		X"18",X"2C",X"24",X"7C",X"5E",X"5D",X"5C",X"7E",X"79",X"59",X"59",X"79",X"5D",X"DF",X"59",X"59",
		X"59",X"59",X"7F",X"D9",X"79",X"59",X"5B",X"5D",X"7E",X"5C",X"7C",X"7E",X"5D",X"7E",X"2C",X"18",
		X"00",X"40",X"60",X"30",X"10",X"80",X"40",X"00",X"80",X"80",X"00",X"40",X"C0",X"80",X"00",X"00",
		X"83",X"08",X"0C",X"04",X"61",X"F0",X"50",X"00",X"01",X"00",X"06",X"66",X"B0",X"C0",X"E2",X"42",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"40",X"E0",X"F0",X"A0",X"C0",X"C0",X"80",X"00",X"00",X"40",X"20",X"00",X"80",X"C0",X"40",X"00",
		X"71",X"AF",X"15",X"21",X"03",X"01",X"20",X"60",X"C0",X"84",X"02",X"02",X"05",X"80",X"80",X"86",
		X"00",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"02",
		X"80",X"00",X"00",X"00",X"40",X"E0",X"40",X"80",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"02",X"04",X"20",X"30",X"10",X"00",X"81",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"03",X"19",X"0C",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"18",X"0C",X"00",X"00",X"00",
		X"3C",X"81",X"00",X"0C",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"04",X"0E",X"04",X"00",X"00",
		X"06",X"0D",X"0B",X"00",X"00",X"00",X"06",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"20",X"70",X"30",X"80",X"40",X"A0",X"C0",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"0C",X"0C",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"1C",X"0B",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"40",X"00",X"20",X"30",X"10",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"02",X"04",X"08",X"00",X"00",X"00",X"30",X"00",X"01",X"70",X"E0",X"00",X"00",X"00",X"00",
		X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"20",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"30",X"18",X"08",X"00",
		X"0C",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"41",X"40",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"08",X"00",X"20",X"30",X"10",X"20",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"10",X"20",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"20",X"70",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",
		X"00",X"00",X"01",X"02",X"1C",X"3F",X"47",X"03",X"23",X"32",X"00",X"05",X"01",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"38",X"18",X"18",X"98",X"F0",X"F0",X"38",X"18",X"18",X"98",X"10",X"20",X"00",
		X"00",X"00",X"01",X"0F",X"1F",X"23",X"01",X"11",X"19",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E0",X"70",X"B0",X"F0",X"F8",X"1C",X"0C",X"8C",X"CC",X"08",X"10",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"1F",X"23",X"01",X"11",X"19",X"00",X"02",X"04",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"F8",X"1C",X"0C",X"8C",X"CC",X"08",X"10",X"80",X"00",
		X"00",X"07",X"0F",X"11",X"00",X"08",X"0C",X"00",X"09",X"11",X"00",X"08",X"0C",X"00",X"01",X"00",
		X"00",X"00",X"80",X"C0",X"F8",X"FC",X"8E",X"06",X"46",X"66",X"84",X"C8",X"C0",X"80",X"00",X"00",
		X"00",X"07",X"0F",X"11",X"00",X"08",X"0C",X"07",X"0F",X"11",X"00",X"08",X"0C",X"00",X"01",X"00",
		X"00",X"00",X"80",X"C0",X"F8",X"FC",X"8E",X"06",X"C6",X"E6",X"C4",X"C8",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"03",X"07",X"08",X"01",X"0E",X"1F",X"23",X"01",X"11",X"19",X"01",X"02",X"00",X"00",
		X"00",X"00",X"80",X"F0",X"F8",X"1C",X"0C",X"8C",X"CC",X"88",X"90",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"0E",X"1F",X"23",X"01",X"11",X"19",X"01",X"02",X"00",X"00",
		X"00",X"00",X"00",X"70",X"F8",X"1C",X"0C",X"8C",X"CC",X"88",X"90",X"F0",X"30",X"20",X"40",X"00",
		X"00",X"00",X"01",X"02",X"1C",X"3F",X"47",X"03",X"23",X"33",X"02",X"05",X"01",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"38",X"18",X"18",X"98",X"10",X"30",X"38",X"18",X"18",X"98",X"10",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"04",X"00",X"02",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"40",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"04",X"00",X"00",X"10",X"00",X"00",X"04",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"08",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"08",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"00",X"01",X"00",X"10",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"10",X"00",X"01",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"07",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"00",
		X"01",X"07",X"0F",X"1E",X"3C",X"78",X"F0",X"F0",X"78",X"78",X"3C",X"3C",X"1E",X"1E",X"0F",X"00",
		X"F0",X"B0",X"38",X"18",X"1C",X"0C",X"0E",X"06",X"07",X"02",X"04",X"08",X"10",X"20",X"00",X"00",
		X"02",X"07",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7C",X"3C",X"1C",X"0C",X"04",X"00",
		X"80",X"C0",X"E0",X"F0",X"F8",X"EC",X"CC",X"8C",X"0C",X"0C",X"0C",X"18",X"30",X"60",X"C0",X"80",
		X"01",X"07",X"07",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"C0",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",X"07",X"02",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",
		X"03",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"7F",X"3F",X"1E",X"0E",X"04",X"00",
		X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"FF",X"C2",X"86",X"84",X"0C",X"08",X"18",X"10",X"00",X"00",
		X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1E",X"0E",X"00",X"00",
		X"E0",X"F0",X"F8",X"FC",X"FC",X"7E",X"BE",X"86",X"84",X"8C",X"0C",X"08",X"10",X"20",X"00",X"00",
		X"00",X"03",X"0F",X"03",X"1D",X"3E",X"3E",X"7F",X"7F",X"7F",X"3E",X"3E",X"1C",X"00",X"00",X"00",
		X"00",X"E0",X"F0",X"F8",X"F8",X"F8",X"7C",X"3C",X"3C",X"18",X"18",X"18",X"10",X"20",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"07",X"19",X"3C",X"7E",X"7F",X"7F",X"73",X"33",X"3F",X"1F",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"7C",X"7C",X"BC",X"B8",X"B8",X"B0",X"40",X"00",X"00",
		X"00",X"01",X"07",X"1F",X"23",X"00",X"18",X"3C",X"3E",X"3F",X"33",X"13",X"1F",X"06",X"00",X"00",
		X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"7C",X"7C",X"3C",X"3C",X"38",X"38",X"70",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"3C",X"F8",X"3E",X"0F",X"03",X"00",X"00",X"00",X"00",
		X"70",X"70",X"F0",X"F0",X"F8",X"E8",X"F8",X"F8",X"7C",X"7C",X"BC",X"FC",X"FC",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"0F",X"3B",X"6D",X"37",X"1B",X"0D",X"07",X"03",X"01",X"00",
		X"00",X"60",X"78",X"1C",X"3C",X"FC",X"78",X"68",X"78",X"70",X"50",X"F0",X"E0",X"E0",X"A0",X"80",
		X"00",X"03",X"03",X"00",X"0E",X"0F",X"3F",X"3F",X"15",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"02",
		X"00",X"00",X"C0",X"70",X"1C",X"8E",X"FE",X"1C",X"38",X"B8",X"F0",X"E0",X"E0",X"C0",X"80",X"00",
		X"00",X"01",X"07",X"1F",X"3F",X"2F",X"37",X"17",X"15",X"1F",X"0F",X"0F",X"0D",X"07",X"07",X"04",
		X"00",X"80",X"C0",X"60",X"B0",X"F8",X"FC",X"FE",X"3C",X"38",X"70",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"03",X"07",X"07",X"07",X"0F",X"0F",X"0C",X"1C",X"1E",X"1E",X"3C",X"3F",X"3E",X"00",X"00",
		X"F0",X"F0",X"F8",X"E8",X"E8",X"FC",X"F4",X"54",X"7C",X"3E",X"1E",X"FE",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"07",X"1C",X"3F",X"FD",X"37",X"1D",X"06",X"03",X"00",X"00",X"00",
		X"00",X"18",X"78",X"E8",X"A8",X"38",X"78",X"F8",X"F8",X"78",X"E8",X"E8",X"B8",X"F8",X"60",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0E",X"38",X"FF",X"3D",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"3C",X"FC",X"BC",X"3C",X"7C",X"78",X"F8",X"E8",X"F8",X"F0",X"F0",X"F0",X"70",X"40",
		X"00",X"01",X"03",X"07",X"0F",X"1F",X"3D",X"7B",X"3D",X"0F",X"03",X"01",X"00",X"00",X"00",X"00",
		X"A0",X"E0",X"E0",X"F0",X"50",X"50",X"78",X"68",X"68",X"FC",X"FC",X"BC",X"18",X"60",X"00",X"00",
		X"02",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"14",X"3C",X"3F",X"0E",X"0E",X"00",X"03",X"00",X"00",
		X"80",X"C0",X"E0",X"A0",X"F0",X"F8",X"28",X"3C",X"1E",X"FE",X"0C",X"30",X"C0",X"00",X"00",X"00",
		X"05",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"17",X"15",X"3F",X"2F",X"3F",X"1F",X"07",X"00",X"00",
		X"00",X"80",X"C0",X"E0",X"F0",X"78",X"3C",X"3E",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"3E",X"3F",X"3C",X"1E",X"1E",X"1F",X"0D",X"0F",X"0F",X"07",X"07",X"07",X"03",X"00",
		X"00",X"00",X"00",X"E0",X"FE",X"1E",X"3E",X"7C",X"54",X"F4",X"FC",X"E8",X"E8",X"F8",X"F0",X"F0",
		X"00",X"00",X"00",X"03",X"0F",X"3E",X"78",X"40",X"1F",X"63",X"1C",X"06",X"00",X"00",X"00",X"00",
		X"0C",X"3E",X"7E",X"FF",X"33",X"01",X"01",X"01",X"1F",X"1F",X"1E",X"0E",X"30",X"7C",X"18",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"19",X"30",X"67",X"5F",X"71",X"8E",X"00",X"00",X"00",X"00",X"00",
		X"18",X"3C",X"7C",X"66",X"C6",X"02",X"03",X"0F",X"1F",X"1F",X"0F",X"0F",X"00",X"0E",X"1C",X"00",
		X"00",X"00",X"04",X"06",X"0E",X"1B",X"13",X"23",X"2F",X"5D",X"33",X"4C",X"A0",X"00",X"00",X"00",
		X"10",X"30",X"78",X"78",X"C8",X"8C",X"0C",X"84",X"86",X"1E",X"3E",X"3F",X"3F",X"02",X"1E",X"00",
		X"00",X"00",X"00",X"07",X"0F",X"19",X"31",X"60",X"5C",X"70",X"8E",X"00",X"00",X"00",X"00",X"00",
		X"18",X"3C",X"6C",X"46",X"C6",X"82",X"03",X"03",X"01",X"21",X"E1",X"E1",X"F0",X"00",X"38",X"00",
		X"00",X"00",X"00",X"03",X"0F",X"3D",X"78",X"40",X"19",X"61",X"18",X"05",X"00",X"00",X"00",X"00",
		X"0C",X"3E",X"66",X"C3",X"83",X"01",X"01",X"01",X"81",X"81",X"80",X"00",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"0F",X"A1",X"4D",X"31",X"18",X"08",X"00",X"00",X"00",X"00",
		X"1E",X"3F",X"7B",X"71",X"01",X"01",X"01",X"00",X"C0",X"C2",X"C0",X"40",X"80",X"40",X"20",X"00",
		X"00",X"00",X"70",X"7E",X"7F",X"9F",X"23",X"50",X"2C",X"36",X"18",X"0C",X"08",X"00",X"00",X"00",
		X"0F",X"0F",X"1E",X"1E",X"82",X"80",X"00",X"64",X"78",X"78",X"78",X"B0",X"D0",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"7F",X"7F",X"0F",X"A0",X"4C",X"37",X"18",X"0E",X"00",X"00",X"00",X"00",
		X"1E",X"3F",X"5F",X"0F",X"01",X"01",X"01",X"00",X"10",X"1E",X"3C",X"5C",X"E8",X"70",X"30",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"7E",X"7E",X"7E",X"7E",X"7E",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"FC",X"FC",X"7C",X"7C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"BC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"7E",X"7E",X"7E",X"7C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3C",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"7C",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"BC",X"BC",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"7E",X"7C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"7C",X"7C",X"7C",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"7C",X"7C",X"7C",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"BC",X"FC",X"FC",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3E",X"3E",X"3E",X"3C",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"FC",X"FC",X"FC",X"7C",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"FC",X"FC",X"FC",X"BC",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"7E",X"7E",X"7E",X"7E",X"7C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3E",X"3E",X"3E",X"3E",X"3E",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"BC",X"FC",X"FC",X"FC",X"FC",X"FC",X"BC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"00",X"18",X"3C",X"3C",X"7C",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"3C",X"3C",X"3C",X"18",X"00",
		X"7C",X"E6",X"82",X"82",X"9A",X"BE",X"FE",X"CE",X"CE",X"FE",X"FE",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"86",X"8E",X"9E",X"9A",X"9E",X"9E",X"9E",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"82",X"82",X"86",X"86",X"86",X"86",X"86",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"82",X"82",X"82",X"82",X"C2",X"C2",X"82",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"82",X"C2",X"C2",X"C2",X"E2",X"E2",X"C2",X"82",X"82",X"82",X"A6",X"5C",
		X"7C",X"E6",X"82",X"82",X"E2",X"F2",X"F2",X"B2",X"FA",X"FA",X"F2",X"82",X"82",X"82",X"A6",X"5C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",X"06",X"60",X"60",X"60",X"00",
		X"00",X"03",X"07",X"07",X"0F",X"2D",X"2D",X"4C",X"00",X"ED",X"ED",X"00",X"4C",X"2D",X"2D",X"0C",
		X"C0",X"F0",X"F8",X"F8",X"FC",X"FC",X"7C",X"FC",X"38",X"F8",X"F0",X"00",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"08",X"01",X"14",X"04",X"08",X"18",X"1D",X"00",X"0D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"40",X"00",X"90",X"30",X"B0",X"20",X"00",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"05",X"07",X"0C",X"0B",X"01",X"07",X"02",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"80",X"40",X"20",X"E0",X"30",X"B0",X"20",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"1B",X"0C",X"0D",X"0E",X"1E",X"08",X"0A",X"0C",X"0F",X"09",X"10",X"00",X"00",
		X"00",X"00",X"08",X"90",X"F0",X"B0",X"D0",X"90",X"58",X"B0",X"90",X"F0",X"D8",X"80",X"00",X"00",
		X"00",X"00",X"00",X"26",X"4C",X"40",X"00",X"00",X"03",X"01",X"08",X"0C",X"04",X"10",X"08",X"00",
		X"00",X"00",X"20",X"18",X"08",X"40",X"E0",X"60",X"40",X"08",X"08",X"10",X"10",X"00",X"60",X"C0",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"80",X"A0",X"40",X"80",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",
		X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"82",X"BA",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"BA",X"82",X"FE",X"A2",X"EA",X"EA",X"A2",X"FE",X"D7",X"D7",X"D7",X"D7",X"FF",X"C3",X"FF",X"DB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"22",X"AA",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"9E",X"1F",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5E",X"5E",X"DF",X"59",X"58",X"D9",X"F8",X"F9",
		X"DD",X"DD",X"F9",X"2F",X"08",X"2E",X"0E",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"F9",X"D9",X"59",X"59",X"D9",X"59",X"59",X"F9",
		X"2F",X"2F",X"28",X"2F",X"28",X"2E",X"2E",X"28",X"FF",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FB",
		X"DF",X"DF",X"DF",X"DF",X"68",X"6A",X"68",X"6C",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"9F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"34",X"B6",X"B7",X"B7",X"B7",X"FF",X"FF",X"FF",X"47",X"B7",X"43",X"8B",X"A1",X"C5",X"D1",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"5F",X"DF",X"F0",X"FA",
		X"D2",X"92",X"AC",X"14",X"41",X"1A",X"A0",X"8A",X"87",X"1C",X"65",X"D9",X"23",X"27",X"8F",X"1F",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"F0",X"DA",X"5A",X"50",X"DF",X"59",X"56",X"F9",
		X"28",X"A1",X"0F",X"E8",X"6E",X"0E",X"DE",X"14",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F6",X"F8",X"F1",X"F7",X"FF",X"FF",X"FB",
		X"37",X"74",X"F5",X"B5",X"B5",X"B4",X"B7",X"B4",X"FF",X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",
		X"B6",X"B4",X"37",X"6C",X"6E",X"68",X"6F",X"D9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7E",X"FE",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FE",X"F9",X"F5",X"EC",X"FD",X"FC",X"F1",X"C5",X"14",X"41",X"0A",X"B0",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"BF",X"69",X"13",X"97",X"27",X"2E",X"49",X"FD",X"FE",X"F7",X"E7",X"DB",X"A4",X"44",X"59",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"4F",X"E3",X"68",X"CA",X"92",X"C4",
		X"45",X"34",X"52",X"0A",X"68",X"83",X"1F",X"7F",X"23",X"A7",X"8F",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"80",X"55",X"FD",X"FE",X"F7",X"E7",X"89",X"10",X"A1",X"13",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"4F",X"E3",X"68",X"CA",X"92",X"C4",
		X"00",X"55",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"46",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"ED",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"80",X"55",X"FD",X"FE",X"F7",X"E7",X"89",X"10",X"A1",X"13",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DD",X"B1",X"7F",X"CA",X"6A",X"EF",X"E8",X"EA",
		X"00",X"55",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"46",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F4",X"D4",X"B7",X"74",X"94",X"77",X"FF",X"FF",X"5F",X"5F",X"DF",X"5F",X"7F",X"C3",X"FF",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"77",X"94",X"74",X"B7",X"D4",X"F4",X"FF",X"D7",X"D7",X"57",X"57",X"FF",X"43",X"7F",X"FB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"FF",X"E2",X"E8",X"E2",X"E8",X"E2",X"E8",X"FD",X"FE",X"AB",X"A3",X"8B",X"A3",X"8B",X"A3",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"E2",X"E8",X"E2",X"E8",X"E2",X"F4",X"F1",X"F4",X"8B",X"A3",X"8B",X"A1",X"45",X"53",X"47",X"53",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F1",X"F4",X"F1",X"F4",X"FA",X"F8",X"FA",X"F8",X"47",X"53",X"4B",X"23",X"FF",X"43",X"FF",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FA",X"F8",X"FD",X"FC",X"FD",X"FC",X"FD",X"FE",X"D7",X"57",X"57",X"57",X"7F",X"43",X"7F",X"3B",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"8D",X"36",X"87",X"53",X"42",X"1A",X"A2",X"89",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FF",X"FC",X"F8",X"F8",X"FC",X"A1",X"8D",X"D1",X"C4",X"50",X"47",X"53",X"6B",
		X"A4",X"A4",X"A4",X"FF",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"23",X"2B",X"23",X"EB",X"FF",X"43",X"7F",X"57",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"FF",X"88",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"F5",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"57",X"57",X"57",X"7F",X"C3",X"FF",X"BB",
		X"88",X"88",X"88",X"88",X"FF",X"80",X"FF",X"F7",X"F5",X"F5",X"F5",X"F5",X"FF",X"E1",X"FF",X"EF",
		X"FF",X"FF",X"FD",X"FD",X"FD",X"FD",X"FF",X"FF",X"BD",X"F6",X"77",X"71",X"75",X"71",X"EA",X"E3",
		X"F7",X"F7",X"77",X"FF",X"A4",X"FF",X"A4",X"A4",X"DF",X"BF",X"7F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E8",X"E2",X"E8",X"D6",X"C2",X"FF",X"FF",X"FF",
		X"A4",X"A4",X"A4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",X"07",X"3F",X"F1",X"FF",X"FC",X"FC",X"FE",X"8F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"1F",X"1F",X"FF",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"FE",X"FC",X"FC",X"FC",X"FF",X"FC",X"FC",X"FC",X"7E",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",
		X"FC",X"FC",X"FC",X"FF",X"FC",X"FC",X"FC",X"FE",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",X"FB",X"E1",X"E1",X"E1",X"E3",X"FF",X"1F",X"1F",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"8F",X"FE",X"FC",X"FC",X"FF",X"F1",X"3F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"1F",X"1F",X"3F",
		X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"C0",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"07",X"0F",X"1E",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"1F",X"1F",X"1E",X"0F",X"07",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"3F",X"1F",X"1F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",
		X"80",X"C0",X"C0",X"E0",X"F0",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"07",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E4",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"10",X"10",X"11",X"FE",X"1E",X"1F",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"C6",X"8C",X"9C",X"BC",X"7C",X"3C",X"1C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"3C",X"7C",X"BC",X"9C",X"8C",X"C6",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1E",X"FE",X"11",X"10",X"10",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E4",X"E4",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"D6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E9",X"FC",X"F6",X"F5",X"F2",X"9E",X"8F",X"8F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",X"E5",X"82",X"02",X"03",
		X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"03",X"03",X"03",X"07",X"07",X"07",X"06",X"04",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"04",X"06",X"07",X"07",X"07",X"03",X"03",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"02",X"82",X"E5",X"F9",X"F9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"8F",X"9E",X"F2",X"F5",X"F6",X"FC",X"E9",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"D6",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E4",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EF",X"F5",X"AD",X"AF",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"4F",X"56",X"D3",X"D2",X"D2",X"5A",X"5F",X"5F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"5F",X"5A",X"D2",X"D2",X"D3",X"56",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",X"AF",X"AD",X"F5",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"E4",X"DF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FC",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"C8",X"7F",X"FF",X"FF",X"C4",X"22",X"2F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"8F",X"87",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"87",X"8F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FC",X"FF",
		X"FF",X"2F",X"22",X"C4",X"FF",X"FF",X"7F",X"C8",X"FF",X"FF",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F8",X"FF",X"FF",X"FF",X"FC",X"FE",X"FF",X"FF",X"79",X"FB",X"FF",X"C7",X"03",X"0E",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"FF",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"FC",X"FC",X"FF",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FF",X"FF",X"FF",X"F8",
		X"FE",X"FE",X"0E",X"03",X"C7",X"FF",X"FB",X"79",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7F",X"00",X"00",X"00",X"00",X"00",X"0F",X"FD",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6B",X"F4",X"7C",X"B3",X"F7",X"F9",X"E9",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"DF",X"D7",X"CF",X"CE",X"EE",X"FE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"EE",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EF",X"EE",X"FE",X"EE",X"EE",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"FE",X"EE",X"CE",X"CF",X"D7",X"DF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FB",X"E9",X"F9",X"F7",X"B3",X"7C",X"F4",X"6B",X"7F",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FD",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"F4",X"FC",X"F3",X"F7",X"F9",X"F9",X"FB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F9",X"F9",X"F7",X"F3",X"FC",X"F4",X"EB",
		X"FF",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",X"00",X"00",X"07",X"18",X"73",X"9F",X"3F",X"FF",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F2",X"C1",X"E3",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"FC",X"FC",X"FF",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FD",X"FE",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FE",X"FD",X"FC",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FF",X"FC",X"FC",X"F8",X"F8",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"E3",X"C1",X"F2",X"FE",
		X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",X"FF",X"3F",X"9F",X"73",X"18",X"07",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"C7",X"00",X"00",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"C7",X"83",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"07",X"00",X"00",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"78",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"0C",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"3E",X"7F",X"3E",X"1C",X"08",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"08",X"04",X"04",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"04",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"10",X"10",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"10",X"08",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"1C",X"3E",X"7F",X"3E",X"1C",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"18",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FC",X"FB",X"D6",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",
		X"00",X"00",X"07",X"18",X"73",X"9F",X"3F",X"FF",X"00",X"C0",X"40",X"60",X"E0",X"F0",X"F0",X"88",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"D1",X"3F",X"FC",X"7C",X"FE",X"8F",
		X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",X"FC",X"37",X"2F",X"5F",X"7F",X"7B",X"73",X"57",
		X"FF",X"A4",X"24",X"3F",X"FF",X"FF",X"FF",X"FF",X"E9",X"FC",X"F6",X"F5",X"F2",X"9E",X"8F",X"8F",
		X"5F",X"E4",X"7F",X"FF",X"7F",X"3E",X"BE",X"FF",X"C8",X"7F",X"FF",X"FF",X"C4",X"22",X"2F",X"FF",
		X"79",X"FB",X"FF",X"C7",X"03",X"0E",X"FE",X"FE",X"6B",X"F4",X"7C",X"B3",X"F7",X"F9",X"E9",X"FB",
		X"FE",X"F2",X"C1",X"E3",X"FF",X"FF",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"F2",
		X"5F",X"7F",X"5F",X"7F",X"7B",X"F3",X"A7",X"A7",X"1F",X"1F",X"FF",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"A7",X"BD",X"F9",X"F9",X"F9",X"FF",X"F9",X"F9",
		X"F0",X"10",X"10",X"11",X"FE",X"1E",X"1F",X"1F",X"FF",X"FF",X"F9",X"F9",X"65",X"82",X"02",X"03",
		X"FF",X"FF",X"FF",X"6F",X"75",X"AD",X"AF",X"2F",X"0F",X"8F",X"87",X"FE",X"3E",X"1F",X"9F",X"9F",
		X"FF",X"FF",X"FF",X"3F",X"1F",X"1F",X"3F",X"C9",X"F7",X"DF",X"D7",X"CF",X"CE",X"EE",X"FE",X"EE",
		X"8F",X"B8",X"F8",X"FC",X"7C",X"7F",X"7C",X"FC",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"EE",X"FC",X"FC",X"FC",X"BF",X"BC",X"FC",X"BC",X"7E",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"07",X"0F",X"1E",X"1F",X"1F",X"F9",X"FF",X"F7",X"78",X"88",X"9F",X"F1",X"91",
		X"EE",X"46",X"8C",X"9C",X"BC",X"7C",X"3C",X"1C",X"03",X"03",X"03",X"07",X"07",X"07",X"06",X"04",
		X"4F",X"56",X"D3",X"D2",X"D2",X"5A",X"5F",X"5F",X"6F",X"4F",X"47",X"A7",X"7F",X"E7",X"E7",X"E7",
		X"88",X"88",X"88",X"9F",X"E4",X"C4",X"C4",X"C4",X"EF",X"EE",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",
		X"7C",X"7C",X"7C",X"7D",X"7E",X"FC",X"7C",X"7C",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"BC",X"FC",X"BC",X"BF",X"FC",X"FC",X"FC",X"EE",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"1F",X"1F",X"1E",X"0F",X"07",X"00",X"00",X"00",X"91",X"F1",X"9F",X"88",X"78",X"F7",X"FF",X"F9",
		X"1C",X"3C",X"7C",X"BC",X"9C",X"8C",X"46",X"EE",X"04",X"06",X"07",X"07",X"07",X"03",X"03",X"03",
		X"5F",X"5F",X"5A",X"D2",X"D2",X"D3",X"56",X"4F",X"E7",X"E7",X"E7",X"7F",X"A7",X"47",X"4F",X"6F",
		X"C4",X"C4",X"C4",X"E4",X"9F",X"88",X"88",X"88",X"EE",X"EE",X"EF",X"EE",X"FE",X"EE",X"EE",X"EF",
		X"7C",X"7C",X"FC",X"7E",X"7D",X"7C",X"7C",X"7C",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"A7",X"A7",X"F3",X"7B",X"7F",X"5F",X"7F",X"5F",X"FB",X"E1",X"E1",X"E1",X"E3",X"FF",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"F9",X"F9",X"FF",X"F9",X"F9",X"F9",X"BD",X"A7",
		X"1F",X"1F",X"1E",X"FE",X"11",X"10",X"10",X"F0",X"03",X"02",X"82",X"65",X"F9",X"F9",X"FF",X"FF",
		X"2F",X"AF",X"AD",X"75",X"6F",X"FF",X"FF",X"FF",X"9F",X"9F",X"1F",X"3E",X"FE",X"87",X"8F",X"0F",
		X"C9",X"3F",X"1F",X"1F",X"3F",X"FF",X"FF",X"FF",X"EE",X"FE",X"EE",X"CE",X"CF",X"D7",X"DF",X"F7",
		X"FC",X"7C",X"7F",X"7C",X"FC",X"F8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"8F",X"FE",X"7C",X"FC",X"3F",X"D1",X"3F",X"07",
		X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",X"57",X"73",X"7B",X"7F",X"5F",X"2F",X"37",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"24",X"A4",X"FF",X"8F",X"8F",X"9E",X"F2",X"F5",X"F6",X"FC",X"E9",
		X"FF",X"BE",X"3E",X"7F",X"FF",X"7F",X"E4",X"5F",X"FF",X"2F",X"22",X"C4",X"FF",X"FF",X"7F",X"C8",
		X"FE",X"FE",X"0E",X"03",X"C7",X"FF",X"FB",X"79",X"FB",X"E9",X"F9",X"F7",X"B3",X"7C",X"F4",X"6B",
		X"1F",X"9F",X"FF",X"FF",X"E3",X"C1",X"F2",X"FE",X"F2",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"D6",X"FB",X"FC",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"9F",X"73",X"18",X"07",X"00",X"00",X"88",X"F0",X"F0",X"E0",X"60",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"BF",X"DF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FE",X"F7",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",
		X"00",X"00",X"07",X"18",X"73",X"9F",X"3F",X"FF",X"00",X"C0",X"40",X"60",X"E0",X"F0",X"F0",X"88",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"D1",X"3F",X"FC",X"7C",X"FE",X"8F",
		X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",X"FC",X"37",X"2F",X"5F",X"7F",X"7B",X"73",X"57",
		X"FF",X"A8",X"28",X"7F",X"FF",X"FF",X"FF",X"FF",X"F9",X"BC",X"9F",X"FC",X"FE",X"FF",X"F9",X"F9",
		X"5F",X"E4",X"7F",X"FF",X"7F",X"3E",X"BF",X"FF",X"C8",X"7F",X"FF",X"FF",X"C4",X"22",X"2F",X"FF",
		X"79",X"FB",X"FF",X"C7",X"03",X"0E",X"FE",X"FE",X"6B",X"F4",X"7C",X"B3",X"F7",X"F9",X"E9",X"FB",
		X"FE",X"F2",X"C1",X"E3",X"FF",X"FF",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"F2",
		X"5F",X"7F",X"5F",X"7F",X"7B",X"F3",X"A7",X"A7",X"1F",X"1F",X"FF",X"E3",X"E1",X"E1",X"E1",X"FB",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"A7",X"BD",X"F9",X"F9",X"FB",X"FD",X"F9",X"F9",
		X"90",X"10",X"10",X"11",X"FE",X"1E",X"1F",X"1E",X"7C",X"7F",X"7D",X"FC",X"64",X"83",X"03",X"03",
		X"FF",X"FF",X"FF",X"BF",X"FF",X"AF",X"2B",X"45",X"8F",X"8F",X"C7",X"FE",X"1E",X"0F",X"8F",X"5F",
		X"FF",X"FF",X"FF",X"3F",X"1F",X"1F",X"3F",X"C9",X"F7",X"DF",X"D7",X"CF",X"CE",X"EE",X"FE",X"EE",
		X"8F",X"B8",X"F8",X"FC",X"7C",X"7F",X"7C",X"FC",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"EE",X"FC",X"FC",X"FC",X"BF",X"BC",X"FC",X"BC",X"7E",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",
		X"00",X"00",X"00",X"07",X"0F",X"1E",X"1F",X"1F",X"F9",X"FF",X"F7",X"78",X"88",X"9F",X"F1",X"91",
		X"EE",X"44",X"8C",X"98",X"B8",X"78",X"38",X"38",X"03",X"03",X"03",X"07",X"07",X"07",X"06",X"04",
		X"47",X"C5",X"C4",X"C6",X"C6",X"47",X"47",X"47",X"6F",X"27",X"E3",X"B3",X"BF",X"F3",X"F3",X"F3",
		X"88",X"88",X"88",X"9F",X"E4",X"C4",X"C4",X"C4",X"EF",X"EE",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",
		X"7C",X"7C",X"7C",X"7D",X"7E",X"FC",X"7C",X"7C",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"BC",X"FC",X"BC",X"BF",X"FC",X"FC",X"FC",X"EE",X"7E",X"7E",X"7E",X"FE",X"7E",X"7E",X"7E",X"7E",
		X"1F",X"1F",X"1E",X"0F",X"07",X"00",X"00",X"00",X"91",X"F1",X"9F",X"88",X"78",X"F7",X"FF",X"F9",
		X"38",X"38",X"78",X"B8",X"98",X"8C",X"44",X"EE",X"04",X"06",X"07",X"07",X"07",X"03",X"03",X"03",
		X"47",X"47",X"47",X"C6",X"C6",X"C4",X"C5",X"47",X"F3",X"F3",X"F3",X"BF",X"B3",X"E3",X"27",X"6F",
		X"C4",X"C4",X"C4",X"E4",X"9F",X"88",X"88",X"88",X"EE",X"EE",X"EF",X"EE",X"FE",X"EE",X"EE",X"EF",
		X"7C",X"7C",X"FC",X"7E",X"7D",X"7C",X"7C",X"7C",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"A7",X"A7",X"F3",X"7B",X"7F",X"5F",X"7F",X"5F",X"FB",X"E1",X"E1",X"E1",X"E3",X"FF",X"1F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"F9",X"F9",X"FD",X"FB",X"F9",X"F9",X"BD",X"A7",
		X"1E",X"1F",X"1E",X"FE",X"11",X"10",X"10",X"90",X"03",X"03",X"83",X"64",X"FC",X"7D",X"7F",X"7C",
		X"45",X"2B",X"AF",X"FF",X"BF",X"FF",X"FF",X"FF",X"5F",X"8F",X"0F",X"1E",X"FE",X"C7",X"8F",X"8F",
		X"C9",X"3F",X"1F",X"1F",X"3F",X"FF",X"FF",X"FF",X"EE",X"FE",X"EE",X"CE",X"CF",X"D7",X"DF",X"F7",
		X"FC",X"7C",X"7F",X"7C",X"FC",X"F8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"8F",X"FE",X"7C",X"FC",X"3F",X"D1",X"3F",X"07",
		X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",X"57",X"73",X"7B",X"7F",X"5F",X"2F",X"37",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"28",X"A8",X"FF",X"F9",X"F9",X"FF",X"FE",X"FC",X"9F",X"BC",X"F9",
		X"FF",X"BF",X"3E",X"7F",X"FF",X"7F",X"E4",X"5F",X"FF",X"2F",X"22",X"C4",X"FF",X"FF",X"7F",X"C8",
		X"FE",X"FE",X"0E",X"03",X"C7",X"FF",X"FB",X"79",X"FB",X"E9",X"F9",X"F7",X"B3",X"7C",X"F4",X"6B",
		X"1F",X"9F",X"FF",X"FF",X"E3",X"C1",X"F2",X"FE",X"F2",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"06",X"01",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"BF",X"FF",X"00",X"00",X"00",X"00",X"00",X"F7",X"FE",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"9F",X"73",X"18",X"07",X"00",X"00",X"88",X"F0",X"F0",X"E0",X"60",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"BF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",
		X"00",X"00",X"07",X"18",X"73",X"9F",X"3F",X"FF",X"00",X"C0",X"40",X"60",X"E0",X"F0",X"F0",X"88",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"D1",X"3F",X"FC",X"78",X"FE",X"9F",
		X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",X"FB",X"27",X"3F",X"7F",X"73",X"57",X"A7",X"AF",
		X"FF",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"FF",X"7D",X"F3",X"FE",X"EF",X"EF",X"FF",X"3D",
		X"5F",X"E4",X"FF",X"FF",X"7F",X"FE",X"FF",X"FF",X"C8",X"7F",X"FF",X"FF",X"C2",X"21",X"1F",X"FF",
		X"79",X"FB",X"FF",X"C7",X"03",X"0E",X"FE",X"FE",X"6B",X"F4",X"7C",X"B3",X"F7",X"F9",X"E9",X"FB",
		X"FE",X"F2",X"C1",X"E3",X"FF",X"FF",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"F2",
		X"5F",X"7E",X"5F",X"7F",X"7F",X"F7",X"AF",X"AF",X"1F",X"3F",X"FF",X"E3",X"C1",X"C2",X"C2",X"FA",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"B9",X"F9",X"7A",X"72",X"73",X"7E",X"F2",X"72",
		X"10",X"10",X"10",X"17",X"FE",X"3F",X"5E",X"4C",X"3C",X"3C",X"3E",X"FE",X"C7",X"02",X"03",X"02",
		X"FF",X"BF",X"BF",X"BF",X"FF",X"BC",X"36",X"4B",X"8F",X"87",X"C7",X"FE",X"BF",X"1F",X"0F",X"3F",
		X"FF",X"FF",X"FF",X"1F",X"0F",X"0F",X"BF",X"C9",X"F7",X"DF",X"D7",X"CF",X"CE",X"EE",X"FE",X"EE",
		X"8F",X"B8",X"F8",X"FC",X"7C",X"7F",X"7C",X"FC",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"EE",X"F8",X"F8",X"F8",X"BF",X"B8",X"F8",X"B8",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"07",X"0F",X"1E",X"1F",X"1F",X"F2",X"7F",X"F7",X"79",X"92",X"FE",X"A2",X"22",
		X"84",X"8C",X"18",X"B8",X"F8",X"F8",X"78",X"38",X"03",X"03",X"03",X"07",X"07",X"06",X"04",X"04",
		X"45",X"C4",X"C2",X"C3",X"82",X"81",X"81",X"81",X"C7",X"C3",X"A3",X"53",X"DF",X"F9",X"F9",X"F9",
		X"C4",X"C4",X"E4",X"FF",X"E2",X"E2",X"E2",X"E2",X"EF",X"EE",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",
		X"7C",X"7C",X"7C",X"7D",X"7E",X"FC",X"7C",X"7C",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"B8",X"F8",X"B8",X"BF",X"F8",X"F8",X"F8",X"EE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"1F",X"1F",X"1E",X"0F",X"07",X"00",X"00",X"00",X"22",X"A2",X"FE",X"92",X"79",X"F7",X"7F",X"F2",
		X"38",X"78",X"F8",X"F8",X"B8",X"18",X"8C",X"84",X"04",X"04",X"06",X"07",X"07",X"03",X"03",X"03",
		X"81",X"81",X"81",X"82",X"C3",X"C2",X"C4",X"45",X"F9",X"F9",X"F9",X"DF",X"53",X"A3",X"C3",X"C7",
		X"E2",X"E2",X"E2",X"E2",X"FF",X"E4",X"C4",X"C4",X"EE",X"EE",X"EF",X"EE",X"FE",X"EE",X"EE",X"EF",
		X"7C",X"7C",X"FC",X"7E",X"7D",X"7C",X"7C",X"7C",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"AF",X"AF",X"F7",X"7F",X"7F",X"5F",X"7E",X"5F",X"FA",X"C2",X"C2",X"C1",X"E3",X"FF",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"72",X"F2",X"7E",X"73",X"72",X"7A",X"F9",X"B9",
		X"4C",X"5E",X"3F",X"FE",X"17",X"10",X"10",X"10",X"02",X"03",X"02",X"C7",X"FE",X"3E",X"3C",X"3C",
		X"4B",X"36",X"BC",X"FF",X"BF",X"BF",X"BF",X"FF",X"3F",X"0F",X"1F",X"BF",X"FE",X"C7",X"87",X"8F",
		X"C9",X"BF",X"0F",X"0F",X"1F",X"FF",X"FF",X"FF",X"EE",X"FE",X"EE",X"CE",X"CF",X"D7",X"DF",X"F7",
		X"FC",X"7C",X"7F",X"7C",X"FC",X"F8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"9F",X"FE",X"78",X"FC",X"3F",X"D1",X"3F",X"07",
		X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",X"AF",X"A7",X"57",X"73",X"7F",X"3F",X"27",X"FB",
		X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"FF",X"3D",X"FF",X"EF",X"EF",X"FE",X"F3",X"7D",X"FF",
		X"FF",X"FF",X"FE",X"7F",X"FF",X"FF",X"E4",X"5F",X"FF",X"1F",X"21",X"C2",X"FF",X"FF",X"7F",X"C8",
		X"FE",X"FE",X"0E",X"03",X"C7",X"FF",X"FB",X"79",X"FB",X"E9",X"F9",X"F7",X"B3",X"7C",X"F4",X"6B",
		X"1F",X"9F",X"FF",X"FF",X"E3",X"C1",X"F2",X"FE",X"F2",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"9F",X"73",X"18",X"07",X"00",X"00",X"88",X"F0",X"F0",X"E0",X"60",X"40",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"BF",X"00",X"00",X"00",X"00",X"00",X"F8",X"FC",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"7E",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F5",X"16",X"00",X"00",X"00",X"00",X"00",X"01",X"82",X"C6",
		X"00",X"00",X"07",X"18",X"73",X"9F",X"3F",X"FF",X"00",X"C0",X"40",X"60",X"E0",X"F0",X"F0",X"88",
		X"00",X"00",X"01",X"07",X"0B",X"14",X"14",X"2B",X"07",X"3F",X"D1",X"3F",X"FC",X"78",X"FE",X"9F",
		X"FF",X"CB",X"2C",X"10",X"A0",X"40",X"40",X"80",X"FB",X"27",X"3F",X"7F",X"73",X"57",X"A7",X"AF",
		X"FF",X"24",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"FF",X"7D",X"F3",X"FE",X"EF",X"EF",X"FF",X"3D",
		X"5F",X"E4",X"FF",X"FF",X"7F",X"FE",X"FF",X"FF",X"C8",X"7F",X"FF",X"FF",X"C2",X"21",X"1F",X"FF",
		X"79",X"FB",X"FF",X"C7",X"03",X"0E",X"FE",X"FE",X"6B",X"F4",X"7C",X"B3",X"F7",X"F9",X"E9",X"FB",
		X"FE",X"F2",X"C1",X"E3",X"FF",X"FF",X"9F",X"1F",X"08",X"08",X"78",X"FC",X"FC",X"FC",X"FE",X"F2",
		X"5F",X"7E",X"5F",X"7F",X"7F",X"F7",X"AF",X"AF",X"1F",X"3F",X"FF",X"E3",X"C1",X"C2",X"C2",X"FA",
		X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"B9",X"F9",X"7A",X"72",X"73",X"7E",X"F2",X"72",
		X"10",X"10",X"10",X"17",X"FE",X"3F",X"5E",X"4C",X"3C",X"3C",X"3E",X"FE",X"C7",X"02",X"03",X"02",
		X"FF",X"BF",X"BF",X"BF",X"FF",X"BF",X"27",X"41",X"8F",X"87",X"C7",X"FF",X"9F",X"EF",X"DF",X"EF",
		X"FF",X"FF",X"FF",X"1F",X"0F",X"8F",X"BF",X"C9",X"F7",X"DF",X"D7",X"CF",X"CE",X"EE",X"FE",X"EE",
		X"8F",X"B8",X"F8",X"FC",X"7C",X"7F",X"7C",X"FC",X"82",X"82",X"42",X"42",X"7F",X"C1",X"41",X"21",
		X"EE",X"F8",X"F8",X"F8",X"BF",X"B8",X"F8",X"B8",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"00",X"07",X"0F",X"1E",X"1F",X"1F",X"F2",X"7F",X"F7",X"79",X"92",X"FE",X"A2",X"22",
		X"84",X"8C",X"18",X"B8",X"F8",X"F8",X"78",X"38",X"03",X"03",X"03",X"07",X"07",X"06",X"04",X"04",
		X"40",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"D7",X"4B",X"65",X"35",X"2A",X"16",X"12",X"12",
		X"C4",X"E4",X"E4",X"FF",X"E2",X"F2",X"F2",X"F2",X"EF",X"EE",X"EE",X"FE",X"EE",X"EF",X"EE",X"EE",
		X"7C",X"7C",X"7C",X"7D",X"7E",X"FC",X"7C",X"7C",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",X"21",
		X"B8",X"F8",X"B8",X"BF",X"F8",X"F8",X"F8",X"EE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FE",
		X"1F",X"1F",X"1E",X"0F",X"07",X"00",X"00",X"00",X"22",X"A2",X"FE",X"92",X"79",X"F7",X"7F",X"F2",
		X"38",X"78",X"F8",X"F8",X"B8",X"18",X"8C",X"84",X"04",X"04",X"06",X"07",X"07",X"03",X"03",X"03",
		X"80",X"80",X"80",X"80",X"C0",X"C0",X"C0",X"40",X"12",X"12",X"16",X"2A",X"35",X"65",X"4B",X"D7",
		X"F2",X"F2",X"F2",X"E2",X"FF",X"E4",X"E4",X"C4",X"EE",X"EE",X"EF",X"EE",X"FE",X"EE",X"EE",X"EF",
		X"7C",X"7C",X"FC",X"7E",X"7D",X"7C",X"7C",X"7C",X"21",X"21",X"21",X"21",X"FF",X"21",X"21",X"21",
		X"AF",X"AF",X"F7",X"7F",X"7F",X"5F",X"7E",X"5F",X"FA",X"C2",X"C2",X"C1",X"E3",X"FF",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"72",X"F2",X"7E",X"73",X"72",X"7A",X"F9",X"B9",
		X"4C",X"5E",X"3F",X"FE",X"17",X"10",X"10",X"10",X"02",X"03",X"02",X"C7",X"FE",X"3E",X"3C",X"3C",
		X"41",X"27",X"BF",X"FF",X"BF",X"BF",X"BF",X"FF",X"EF",X"DF",X"EF",X"9F",X"FF",X"C7",X"87",X"8F",
		X"C9",X"BF",X"8F",X"0F",X"1F",X"FF",X"FF",X"FF",X"EE",X"FE",X"EE",X"CE",X"CF",X"D7",X"DF",X"F7",
		X"FC",X"7C",X"7F",X"7C",X"FC",X"F8",X"B8",X"8F",X"21",X"41",X"C1",X"7F",X"42",X"42",X"82",X"82",
		X"2B",X"14",X"14",X"0B",X"07",X"01",X"00",X"00",X"9F",X"FE",X"78",X"FC",X"3F",X"D1",X"3F",X"07",
		X"80",X"40",X"40",X"A0",X"10",X"2C",X"CB",X"FF",X"AF",X"A7",X"57",X"73",X"7F",X"3F",X"27",X"FB",
		X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"24",X"FF",X"3D",X"FF",X"EF",X"EF",X"FE",X"F3",X"7D",X"FF",
		X"FF",X"FF",X"FE",X"7F",X"FF",X"FF",X"E4",X"5F",X"FF",X"1F",X"21",X"C2",X"FF",X"FF",X"7F",X"C8",
		X"FE",X"FE",X"0E",X"03",X"C7",X"FF",X"FB",X"79",X"FB",X"E9",X"F9",X"F7",X"B3",X"7C",X"F4",X"6B",
		X"1F",X"9F",X"FF",X"FF",X"E3",X"C1",X"F2",X"FE",X"F2",X"FE",X"FC",X"FC",X"FC",X"78",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"07",X"01",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FC",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"F5",X"0F",X"00",X"00",X"00",X"00",X"00",X"C6",X"82",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"3F",X"9F",X"73",X"18",X"07",X"00",X"00",X"88",X"F0",X"F0",X"E0",X"60",X"40",X"C0",X"00",
		X"00",X"20",X"00",X"40",X"40",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"40",X"40",X"40",X"20",
		X"01",X"03",X"07",X"3F",X"7F",X"1F",X"07",X"01",X"01",X"81",X"00",X"7E",X"20",X"00",X"08",X"00",
		X"03",X"01",X"01",X"1F",X"C1",X"81",X"07",X"43",X"05",X"01",X"01",X"3F",X"01",X"01",X"07",X"01",
		X"81",X"87",X"1E",X"7E",X"3C",X"0C",X"08",X"00",X"01",X"01",X"03",X"1F",X"FF",X"EF",X"C7",X"C3",
		X"03",X"07",X"0F",X"3F",X"03",X"01",X"05",X"01",X"01",X"01",X"00",X"7E",X"0C",X"04",X"00",X"00",
		X"03",X"01",X"01",X"1F",X"7D",X"6D",X"45",X"41",X"07",X"0F",X"1F",X"3F",X"0D",X"09",X"01",X"01",
		X"00",X"03",X"00",X"98",X"CC",X"60",X"20",X"02",X"00",X"80",X"01",X"10",X"00",X"01",X"00",X"04",
		X"8F",X"00",X"00",X"37",X"81",X"00",X"32",X"42",X"61",X"00",X"00",X"CE",X"01",X"00",X"0C",X"06",
		X"46",X"67",X"30",X"98",X"4C",X"60",X"20",X"00",X"00",X"00",X"01",X"10",X"9C",X"9B",X"90",X"84",
		X"83",X"00",X"00",X"37",X"83",X"00",X"70",X"40",X"61",X"00",X"00",X"CE",X"03",X"00",X"60",X"10",
		X"46",X"01",X"00",X"98",X"4C",X"60",X"20",X"00",X"80",X"98",X"19",X"10",X"8C",X"09",X"00",X"00",
		X"31",X"02",X"47",X"57",X"DF",X"DF",X"D0",X"77",X"17",X"00",X"C1",X"FF",X"61",X"01",X"45",X"55",
		X"87",X"01",X"01",X"D7",X"C1",X"81",X"17",X"57",X"45",X"01",X"01",X"D7",X"01",X"01",X"07",X"C7",
		X"F7",X"56",X"57",X"57",X"5D",X"4D",X"40",X"65",X"55",X"00",X"83",X"FF",X"FF",X"13",X"D7",X"D7",
		X"C3",X"07",X"07",X"D7",X"83",X"01",X"55",X"55",X"45",X"01",X"01",X"D7",X"07",X"07",X"43",X"D1",
		X"77",X"00",X"01",X"57",X"5D",X"4D",X"40",X"65",X"D7",X"52",X"FF",X"FF",X"8D",X"01",X"41",X"53",
		X"09",X"83",X"07",X"BF",X"8F",X"EF",X"88",X"BA",X"27",X"81",X"81",X"AF",X"20",X"61",X"00",X"7D",
		X"88",X"00",X"00",X"EA",X"C0",X"81",X"27",X"67",X"00",X"00",X"00",X"FF",X"01",X"01",X"8F",X"C7",
		X"0F",X"EF",X"0F",X"BF",X"0D",X"6D",X"08",X"28",X"6D",X"01",X"83",X"AF",X"A0",X"FF",X"00",X"FF",
		X"E0",X"02",X"0A",X"EA",X"80",X"01",X"6D",X"6D",X"00",X"00",X"00",X"FF",X"0F",X"07",X"E3",X"F1",
		X"07",X"01",X"01",X"BF",X"0D",X"6D",X"08",X"28",X"EF",X"EF",X"AF",X"AF",X"80",X"09",X"00",X"73",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"EA",X"6E",X"10",X"8A",X"01",X"FC",X"E7",X"00",X"C4",X"80",X"01",X"62",X"45",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FD",
		X"F9",X"E3",X"80",X"3F",X"FF",X"FF",X"BF",X"FF",X"80",X"DF",X"7F",X"1F",X"C0",X"0D",X"E9",X"DD",
		X"08",X"28",X"8F",X"18",X"07",X"8F",X"87",X"C0",X"0B",X"1F",X"DF",X"7F",X"FF",X"FF",X"BF",X"27",
		X"FF",X"FF",X"FF",X"FE",X"FD",X"FA",X"F8",X"F8",X"FF",X"E7",X"B0",X"C0",X"00",X"00",X"01",X"00",
		X"FF",X"BF",X"27",X"05",X"1A",X"21",X"FA",X"DB",X"FC",X"FF",X"F9",X"FB",X"BE",X"B1",X"8A",X"D1",
		X"F7",X"4F",X"BB",X"CF",X"3F",X"7F",X"7F",X"7F",X"C0",X"DD",X"E3",X"FF",X"FF",X"FF",X"F7",X"FF",
		X"16",X"E1",X"FD",X"F0",X"FC",X"FD",X"FF",X"FF",X"F9",X"B9",X"DE",X"E7",X"FA",X"39",X"F0",X"FC",
		X"F0",X"F0",X"F0",X"F0",X"F8",X"F0",X"FC",X"FC",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"A3",X"7E",X"1B",X"00",X"78",X"7D",X"0A",X"4B",X"E5",X"63",X"10",X"3A",X"51",X"A2",X"E5",X"C5",
		X"8F",X"DE",X"55",X"55",X"7F",X"7F",X"7D",X"4B",X"FF",X"6F",X"CB",X"E7",X"39",X"DF",X"07",X"21",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"77",X"FB",X"FF",X"FF",X"FF",X"FF",X"DF",X"AF",X"F7",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"C0",X"BD",X"F0",X"FF",X"FF",X"FF",
		X"08",X"21",X"47",X"9F",X"FF",X"FF",X"FF",X"FF",X"0D",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B7",X"89",X"F7",X"ED",X"E7",X"DC",X"97",X"28",X"D1",X"E4",X"BB",X"05",X"F1",X"47",X"18",X"3C",
		X"FF",X"FF",X"FF",X"7F",X"E3",X"8F",X"FE",X"FF",X"BE",X"FC",X"FD",X"FB",X"F4",X"C7",X"15",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"FF",X"EF",X"FE",X"FF",X"FF",X"FF",X"E0",X"E3",X"FE",X"FE",X"20",X"80",X"FF",X"FF",
		X"BF",X"3F",X"4F",X"EE",X"FB",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"F7",X"E7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"C1",X"DB",X"FE",X"FF",X"FF",X"FF",X"E3",X"FB",X"FD",X"FE",X"3E",X"C4",X"E1",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"F8",X"C6",X"30",X"EF",X"FF",X"FF",X"FF",X"7B",X"FC",X"20",X"20",X"E8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"FF",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"F3",X"F7",X"EF",X"EF",X"DF",X"DF",X"BF",
		X"FD",X"FF",X"FE",X"FF",X"FF",X"FD",X"F9",X"FA",X"E3",X"F9",X"7E",X"E3",X"FB",X"87",X"BF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FF",X"FC",X"DF",X"B4",X"6E",X"FF",X"FF",X"EE",X"FE",
		X"07",X"D2",X"13",X"02",X"D4",X"BD",X"25",X"28",X"7F",X"FD",X"0B",X"70",X"26",X"1E",X"DF",X"50",
		X"FF",X"FF",X"7F",X"1E",X"EE",X"89",X"2E",X"E4",X"3F",X"33",X"7B",X"53",X"FF",X"DF",X"69",X"37",
		X"F8",X"F8",X"7D",X"51",X"59",X"4D",X"D1",X"3C",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FF",X"FF",X"DC",X"FF",X"F6",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"6F",X"08",X"3E",X"13",X"12",X"E7",X"04",X"83",X"02",X"2D",X"00",X"8B",X"A1",X"F1",X"60",X"41",
		X"81",X"08",X"9B",X"B4",X"6C",X"80",X"D1",X"21",X"64",X"10",X"33",X"50",X"46",X"AB",X"20",X"3F",
		X"65",X"84",X"82",X"30",X"00",X"84",X"19",X"00",X"0F",X"61",X"C6",X"4C",X"23",X"09",X"20",X"6E",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"C0",X"F0",X"E9",X"FF",X"FA",X"FF",
		X"44",X"00",X"00",X"07",X"BD",X"EF",X"3F",X"FF",X"E8",X"F6",X"4B",X"9F",X"7F",X"FF",X"FF",X"FF",
		X"86",X"F1",X"F7",X"FA",X"FE",X"FF",X"FF",X"FF",X"7F",X"BF",X"FF",X"DF",X"FF",X"FF",X"CF",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F2",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7D",X"F8",X"DC",X"E0",X"E8",X"F0",X"F0",X"F8",
		X"FF",X"7B",X"7F",X"00",X"A8",X"40",X"1F",X"07",X"FF",X"FF",X"7F",X"17",X"BF",X"7F",X"FF",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"44",X"DB",X"E0",X"FC",X"FF",X"FF",X"FF",X"FF",X"5F",X"E0",X"00",X"00",X"F0",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"67",X"80",X"20",X"FF",X"FF",X"FF",X"FC",X"01",X"F7",X"C7",X"24",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EB",X"B9",X"4D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"E0",X"E0",X"CA",X"80",X"E0",X"07",X"80",
		X"41",X"30",X"03",X"00",X"08",X"00",X"00",X"00",X"FF",X"3F",X"C3",X"7C",X"08",X"8E",X"0F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"F7",X"EF",X"FF",X"F5",X"EF",X"1F",X"70",X"C1",X"8E",X"3F",X"21",
		X"DF",X"FF",X"FA",X"10",X"23",X"A0",X"17",X"0B",X"FF",X"FF",X"3F",X"3F",X"13",X"8F",X"94",X"66",
		X"FF",X"FE",X"FE",X"F7",X"E4",X"03",X"7E",X"40",X"00",X"11",X"28",X"9C",X"08",X"04",X"0A",X"34",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"DE",X"FE",X"D6",X"DF",X"FF",X"FF",X"FF",X"FF",X"41",X"4D",X"4B",X"AF",X"C0",X"E2",X"1F",X"CC",
		X"01",X"18",X"C2",X"00",X"87",X"8F",X"8F",X"4B",X"F7",X"BA",X"02",X"02",X"B0",X"30",X"11",X"AC",
		X"26",X"B1",X"41",X"FF",X"C1",X"F3",X"6F",X"9C",X"32",X"F1",X"FE",X"F0",X"E6",X"F8",X"E0",X"41",
		X"80",X"40",X"80",X"58",X"00",X"20",X"18",X"C0",X"20",X"04",X"08",X"00",X"02",X"3F",X"14",X"08",
		X"F4",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"03",X"E5",X"00",X"B3",X"BF",X"DD",X"FF",X"FF",
		X"60",X"C3",X"F8",X"F4",X"5F",X"FF",X"FF",X"FF",X"14",X"FF",X"BF",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"E8",X"E1",X"F4",X"F8",X"FC",X"FC",X"FE",X"9F",X"3F",X"FF",X"16",X"A0",X"3F",X"FF",X"70",
		X"A8",X"D8",X"E0",X"0F",X"00",X"80",X"20",X"01",X"00",X"00",X"20",X"38",X"00",X"01",X"1C",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"02",X"1C",X"1B",X"A7",X"9C",X"C0",X"CE",X"E1",
		X"00",X"00",X"C0",X"A0",X"00",X"00",X"00",X"59",X"02",X"01",X"00",X"00",X"C0",X"63",X"21",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"BF",X"70",X"FC",X"FF",X"FF",X"FF",X"FF",X"07",X"C0",X"00",X"7E",X"F8",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"C0",X"E0",X"00",X"C0",X"E0",X"00",X"00",X"28",X"FE",X"FE",X"28",X"FE",X"FE",X"28",X"00",
		X"08",X"5C",X"54",X"FE",X"54",X"74",X"20",X"00",X"84",X"4A",X"24",X"10",X"48",X"A4",X"42",X"00",
		X"0A",X"04",X"6E",X"9A",X"B2",X"72",X"0C",X"00",X"00",X"00",X"00",X"00",X"E0",X"D0",X"00",X"00",
		X"00",X"00",X"82",X"C6",X"7C",X"38",X"00",X"00",X"00",X"38",X"7C",X"C6",X"82",X"00",X"00",X"00",
		X"00",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"10",X"10",X"7C",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0E",X"02",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"10",X"10",X"54",X"10",X"10",X"00",X"00",
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"6C",X"6C",X"00",X"00",X"00",X"00",X"00",X"00",X"6C",X"6E",X"02",X"00",X"00",
		X"00",X"82",X"C6",X"6C",X"38",X"10",X"00",X"00",X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"00",
		X"00",X"10",X"38",X"6C",X"C6",X"82",X"00",X"00",X"60",X"F0",X"DA",X"CA",X"CA",X"E0",X"60",X"00",
		X"3C",X"42",X"81",X"A5",X"A5",X"99",X"42",X"3C",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"92",X"FE",X"FE",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"FE",X"FE",X"1C",X"38",X"1C",X"FE",X"FE",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"E0",X"F0",X"1E",X"1E",X"F0",X"E0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"82",X"82",X"FE",X"FE",X"00",X"00",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"78",X"FC",X"7E",X"3F",X"7F",X"BF",X"1F",X"1F",X"00",X"01",X"00",X"00",X"80",X"C1",X"E2",X"E0",
		X"F0",X"F8",X"FC",X"7E",X"FF",X"7F",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"2F",X"27",X"47",X"43",X"43",X"01",X"01",
		X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"3F",X"5F",X"4F",X"8F",X"87",X"87",X"00",X"00",
		X"E0",X"E0",X"F0",X"F0",X"D8",X"18",X"1C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"3F",X"32",X"64",X"64",X"E8",X"E8",X"F0",X"F1",X"FF",X"00",X"00",X"00",X"00",X"C0",X"C0",X"E0",
		X"C0",X"04",X"03",X"00",X"01",X"0F",X"3F",X"FF",X"4F",X"40",X"98",X"78",X"FC",X"FC",X"FE",X"FE",
		X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0F",X"1E",
		X"01",X"03",X"03",X"E3",X"F7",X"FF",X"8F",X"0F",X"E0",X"E3",X"C3",X"C7",X"E7",X"DF",X"DF",X"EF",
		X"E0",X"70",X"3F",X"9F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F8",X"F8",X"FC",X"FC",
		X"00",X"00",X"FF",X"E0",X"10",X"10",X"08",X"08",X"08",X"04",X"FC",X"0C",X"34",X"04",X"1A",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"34",X"27",X"2B",X"5B",X"7B",X"77",X"77",X"0F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"EF",X"EF",X"BD",X"BD",X"DE",X"DE",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"FE",X"FE",X"BF",X"DF",X"DF",X"EF",X"AF",X"B7",X"04",X"05",X"02",X"22",X"A1",X"91",X"DF",X"C8",
		X"01",X"FF",X"00",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"80",X"80",X"40",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"6F",X"6F",X"6F",X"3F",X"3F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"ED",X"EE",X"F6",X"D6",X"F7",X"FB",X"FB",X"FD",X"FD",X"FE",X"FE",
		X"BF",X"DF",X"DF",X"D7",X"D7",X"FB",X"FB",X"FB",X"D7",X"DB",X"EB",X"ED",X"DD",X"DA",X"BA",X"BD",
		X"E8",X"E4",X"B7",X"70",X"D8",X"B7",X"E7",X"68",X"40",X"40",X"E0",X"20",X"1F",X"FF",X"E0",X"30",
		X"10",X"10",X"08",X"08",X"F4",X"FC",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"0F",X"07",X"03",X"03",X"03",X"03",X"D7",X"DF",X"EF",X"EF",X"FF",X"BE",X"BE",X"D6",
		X"7E",X"7E",X"7E",X"7E",X"7D",X"FD",X"ED",X"ED",X"FA",X"F6",X"B6",X"B6",X"DE",X"DE",X"EC",X"6C",
		X"FD",X"FB",X"7B",X"7F",X"3D",X"3D",X"1C",X"1C",X"5C",X"BC",X"FE",X"FE",X"BF",X"7F",X"FF",X"FF",
		X"10",X"18",X"08",X"0C",X"04",X"06",X"82",X"83",X"08",X"08",X"04",X"04",X"02",X"82",X"F9",X"41",
		X"80",X"80",X"40",X"40",X"20",X"20",X"10",X"10",X"00",X"00",X"00",X"00",X"40",X"40",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"D6",X"DB",X"DB",X"DD",X"BD",X"BD",X"BD",X"BD",X"F7",X"F7",X"FB",X"FB",X"FB",X"FB",X"FB",X"FB",
		X"6C",X"AC",X"AC",X"DC",X"D8",X"D8",X"C8",X"88",X"8C",X"8C",X"44",X"44",X"24",X"26",X"14",X"14",
		X"7F",X"7F",X"3E",X"3C",X"51",X"52",X"28",X"29",X"C1",X"C1",X"E0",X"E0",X"70",X"70",X"BF",X"3F",
		X"7C",X"A0",X"BE",X"C0",X"7F",X"00",X"FF",X"FF",X"88",X"88",X"87",X"44",X"C2",X"02",X"FF",X"FF",
		X"30",X"C0",X"03",X"0C",X"33",X"CF",X"FF",X"FF",X"00",X"E0",X"20",X"F0",X"F0",X"E0",X"C0",X"80",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",
		X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",
		X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",X"14",X"14",X"13",X"13",X"A7",X"A7",X"63",X"63",
		X"7F",X"FF",X"FF",X"FF",X"DF",X"DF",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"BF",X"BF",X"DF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FB",X"FB",X"FD",X"FD",X"FF",X"FE",X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"A3",X"A3",X"97",X"97",X"AF",X"2F",X"17",X"17",X"C6",X"C7",X"A3",X"A3",X"91",X"91",X"88",X"88",
		X"FF",X"FF",X"B7",X"B7",X"DB",X"DB",X"FF",X"FF",X"EF",X"FF",X"FB",X"FB",X"FD",X"FD",X"FF",X"FF",
		X"F0",X"F0",X"70",X"70",X"B8",X"B8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"07",X"0F",X"07",X"03",X"07",X"0B",X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",
		X"85",X"C4",X"84",X"88",X"88",X"88",X"88",X"88",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",
		X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",X"0B",X"0B",X"49",X"29",X"31",X"19",X"1F",X"0F",
		X"C4",X"C4",X"E2",X"E2",X"F1",X"F1",X"F9",X"F9",X"FF",X"E3",X"D1",X"B7",X"A7",X"A7",X"E3",X"E3",
		X"FF",X"FE",X"FD",X"FB",X"FA",X"FA",X"FE",X"FE",X"FC",X"3C",X"1C",X"7C",X"7C",X"7C",X"3C",X"3E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"12",X"02",X"02",X"02",X"02",X"06",X"04",X"05",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"88",X"90",X"50",X"50",X"70",X"50",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"0F",X"07",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"F1",X"F8",X"F8",X"F0",X"F0",X"E0",
		X"3E",X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"3E",X"00",X"00",X"00",X"80",X"80",X"00",X"00",X"00",
		X"05",X"05",X"05",X"03",X"03",X"00",X"01",X"01",X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",
		X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",
		X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",X"FF",X"FF",X"7F",X"BF",X"DF",X"DF",X"DF",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"BF",X"73",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"FF",X"FF",X"3F",X"03",X"30",X"60",X"00",X"00",
		X"FE",X"FE",X"FE",X"FE",X"3E",X"1C",X"08",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BF",X"7F",X"7F",X"3F",X"03",X"03",X"01",X"01",
		X"74",X"32",X"E2",X"E1",X"E1",X"E1",X"F1",X"F2",X"51",X"11",X"10",X"04",X"44",X"42",X"22",X"21",
		X"7F",X"3F",X"BF",X"BF",X"FF",X"FF",X"FF",X"7F",X"E0",X"E8",X"E8",X"E4",X"C4",X"C2",X"C2",X"C2",
		X"00",X"20",X"00",X"07",X"78",X"7F",X"78",X"7F",X"24",X"24",X"42",X"82",X"01",X"81",X"78",X"87",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"FA",X"FA",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"11",X"11",X"09",X"29",X"24",X"14",X"12",X"0A",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C2",X"C2",X"84",X"84",X"84",X"84",X"80",X"90",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8B",X"8B",X"53",X"55",X"25",X"25",X"15",X"15",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"77",X"91",X"89",X"C9",X"C9",X"E1",X"E1",X"F3",X"F3",
		X"FF",X"FF",X"C3",X"C0",X"C0",X"C0",X"8F",X"8F",X"FF",X"FF",X"FF",X"3F",X"1F",X"1E",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"1F",X"07",X"01",X"00",X"00",X"00",X"00",
		X"08",X"08",X"04",X"04",X"82",X"86",X"4F",X"5F",X"FB",X"FB",X"FB",X"FB",X"77",X"07",X"07",X"07",
		X"FB",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"88",X"8B",X"D7",X"D7",X"DF",X"FF",X"FF",X"FF",
		X"7E",X"FE",X"FE",X"FC",X"FC",X"FC",X"BC",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"7F",X"EF",X"DF",X"BF",X"BF",X"9F",X"9F",
		X"87",X"87",X"CF",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"0F",X"0F",X"14",X"14",X"0A",X"0A",X"85",X"85",X"B1",X"30",X"58",X"98",X"2F",X"4F",X"1F",X"3F",
		X"FF",X"1F",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",X"1E",X"FF",X"FF",X"FF",X"FF",
		X"80",X"40",X"40",X"20",X"E0",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"44",X"29",X"29",X"18",X"18",X"08",X"08",
		X"FF",X"FF",X"F7",X"F7",X"F3",X"F3",X"F1",X"F1",X"FF",X"FF",X"EF",X"EF",X"F7",X"F7",X"BF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FB",X"FF",X"F8",X"FC",X"FC",X"FE",X"7E",X"7E",X"FE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"03",X"03",X"01",X"01",X"00",X"00",X"E8",X"E8",X"E4",X"E4",X"E2",X"E2",X"F1",X"F1",
		X"ED",X"ED",X"76",X"76",X"3F",X"3F",X"3F",X"38",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"DE",X"DC",X"6E",X"6E",X"FF",X"FF",X"FF",X"8F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"78",X"78",X"3C",X"3C",X"00",X"00",X"00",X"00",X"B4",X"AD",X"69",X"69",X"78",X"78",X"78",X"7D",
		X"7F",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"47",X"DF",X"9F",X"9F",X"8F",X"8F",X"8F",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"FC",X"FC",X"F8",X"70",X"00",
		X"5F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"00",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"FA",X"79",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"B9",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"CC",X"B4",X"A8",X"98",X"88",X"88",X"88",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"88",X"94",X"50",X"50",X"72",X"51",X"70",X"E0",
		X"7B",X"7B",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"EF",X"E9",X"DC",X"DC",X"DE",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"FA",X"79",X"79",X"C6",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"B9",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"CE",X"B5",X"A8",X"98",X"98",X"A8",X"C9",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"8A",X"94",X"5A",X"52",X"72",X"51",X"71",X"E1",
		X"7B",X"7B",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E1",X"F2",X"FD",X"EF",X"E9",X"DC",X"DC",X"DE",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"C1",X"D0",X"F8",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E0",X"EE",X"47",X"43",X"82",X"84",X"CC",X"FC",
		X"12",X"72",X"89",X"D9",X"5D",X"3D",X"3E",X"1E",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"FE",X"9F",X"03",X"01",X"00",X"90",X"D0",X"D0",
		X"0E",X"0F",X"07",X"85",X"C1",X"F5",X"E3",X"F5",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"81",X"87",X"0F",X"1A",X"11",X"51",X"60",X"E0",
		X"F9",X"8B",X"0B",X"07",X"07",X"07",X"87",X"CF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"C0",X"C1",X"E2",X"EE",X"E8",X"DC",X"DC",X"DE",
		X"F7",X"37",X"1F",X"0F",X"0E",X"06",X"1E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DE",X"FC",X"FC",X"F8",X"F9",X"FD",X"DC",X"20",X"2C",X"6E",X"DF",X"DF",X"DC",X"DC",X"BE",
		X"12",X"72",X"89",X"59",X"5D",X"BD",X"3E",X"3F",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DD",X"EF",X"EE",X"F6",X"B7",X"B7",X"D5",X"D1",X"BF",X"BF",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",
		X"17",X"87",X"CF",X"F1",X"F9",X"F9",X"F9",X"F1",X"95",X"A4",X"22",X"22",X"22",X"02",X"82",X"84",
		X"E8",X"E0",X"E1",X"E9",X"FF",X"FF",X"FF",X"FE",X"0F",X"CF",X"BF",X"BF",X"3F",X"3F",X"1F",X"9F",
		X"F1",X"F3",X"EF",X"E3",X"E1",X"C1",X"C1",X"E3",X"84",X"84",X"84",X"D0",X"F7",X"EF",X"EF",X"AF",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"03",X"17",X"17",X"29",X"E8",X"DC",X"DC",X"D0",
		X"E7",X"E7",X"F7",X"EF",X"1E",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D8",X"F8",X"F9",X"F8",X"F0",X"B0",X"90",X"D4",
		X"08",X"30",X"F0",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"E7",X"E3",X"C3",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"E7",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E0",X"EC",X"6E",X"5F",X"DF",X"DF",X"DF",X"BF",
		X"72",X"12",X"1B",X"1B",X"0D",X"8D",X"86",X"86",X"80",X"80",X"20",X"20",X"10",X"91",X"91",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"BF",X"BF",X"BF",X"BF",X"7F",X"7F",X"BF",X"DF",
		X"C6",X"E7",X"EF",X"F1",X"F9",X"F9",X"F9",X"F1",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"CE",X"8E",X"8F",X"8F",X"9F",X"FF",X"FF",X"FE",X"EF",X"CF",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"F1",X"F3",X"E3",X"E7",X"E7",X"E7",X"EB",X"F3",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"AF",
		X"FE",X"FE",X"FC",X"FD",X"D8",X"E8",X"E1",X"F1",X"E3",X"F7",X"F7",X"E9",X"E8",X"FC",X"DC",X"DE",
		X"E3",X"E3",X"E3",X"E3",X"06",X"EE",X"7E",X"1C",X"2F",X"2F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EB",X"DB",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"FA",X"E7",X"C3",X"E1",X"B2",X"90",X"D4",
		X"88",X"70",X"10",X"90",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EE",X"EC",X"E8",X"ED",X"F6",X"F7",X"F7",X"B7",X"BF",X"5F",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E0",X"EC",X"6E",X"5F",X"DF",X"DF",X"DF",X"BF",
		X"15",X"74",X"8A",X"5A",X"5D",X"BD",X"BE",X"BE",X"80",X"80",X"60",X"60",X"30",X"31",X"D1",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"BF",X"BF",X"BF",X"BF",X"7F",X"7F",X"BF",X"DF",
		X"D6",X"E7",X"EF",X"F1",X"F9",X"F9",X"F9",X"F1",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"E6",X"E3",X"E3",X"F7",X"FF",X"FF",X"FE",X"EF",X"CF",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"F1",X"F3",X"E3",X"E7",X"E7",X"E7",X"E7",X"E7",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FE",X"DC",X"EE",X"EF",X"F7",X"E3",X"F7",X"F7",X"E9",X"68",X"3C",X"1C",X"9E",
		X"E7",X"E7",X"F7",X"EF",X"1F",X"FF",X"7F",X"1C",X"0F",X"0F",X"5C",X"9B",X"B7",X"B7",X"A7",X"A7",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B3",X"96",X"D6",
		X"88",X"70",X"10",X"10",X"88",X"88",X"CA",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"58",X"D8",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E0",X"EC",X"6E",X"5F",X"DF",X"DF",X"DF",X"BF",
		X"12",X"72",X"89",X"59",X"5D",X"BD",X"BE",X"BE",X"E0",X"F0",X"60",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"BF",X"BF",X"BF",X"BF",X"7F",X"7F",X"BF",X"DF",
		X"D6",X"E7",X"EF",X"F1",X"F9",X"F9",X"F9",X"F1",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"EF",X"CF",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"F1",X"F3",X"E3",X"E7",X"E7",X"E7",X"E7",X"E7",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E3",X"F7",X"F7",X"E9",X"E8",X"DC",X"DC",X"BE",
		X"E7",X"E7",X"F7",X"EF",X"1E",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"37",X"57",X"57",X"57",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"19",X"B8",X"F8",X"F8",X"F0",X"B0",X"91",X"D7",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E0",X"EC",X"6E",X"5F",X"DF",X"DF",X"DF",X"BF",
		X"12",X"72",X"89",X"59",X"5D",X"BD",X"BE",X"BE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"BF",X"BF",X"BF",X"BF",X"7F",X"7F",X"BF",X"DF",
		X"D6",X"E7",X"EF",X"F1",X"F9",X"F9",X"F9",X"F1",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"EF",X"CF",X"3F",X"3F",X"3F",X"3F",X"5F",X"DF",
		X"F1",X"F3",X"E3",X"E7",X"E7",X"E7",X"E7",X"E7",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E3",X"F7",X"F7",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"E7",X"E7",X"F7",X"EF",X"1E",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"C4",X"84",X"88",X"88",X"88",X"88",X"88",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"88",X"90",X"50",X"50",X"70",X"50",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"C4",X"84",X"88",X"88",X"80",X"80",X"80",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"88",X"90",X"50",X"50",X"70",X"50",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"C4",X"84",X"80",X"84",X"84",X"84",X"84",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"84",X"84",X"50",X"50",X"70",X"50",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"CF",X"87",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"85",X"C0",X"80",X"80",X"80",X"82",X"80",X"80",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"80",X"90",X"50",X"50",X"70",X"50",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"FB",X"BB",X"5B",X"DB",X"EF",X"EF",X"EF",X"EF",X"F6",X"F7",X"F7",X"B7",X"BF",X"DF",X"DE",X"FC",
		X"08",X"88",X"D0",X"F0",X"D1",X"11",X"10",X"10",X"12",X"12",X"15",X"25",X"22",X"22",X"A1",X"81",
		X"EF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FC",X"F8",X"78",X"61",X"C2",X"C5",X"C7",X"83",
		X"12",X"72",X"89",X"39",X"FD",X"FD",X"FE",X"FE",X"80",X"80",X"20",X"20",X"10",X"11",X"11",X"11",
		X"DF",X"EF",X"EF",X"F7",X"B7",X"B7",X"D5",X"D5",X"81",X"C0",X"80",X"80",X"80",X"80",X"80",X"80",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"5B",X"15",X"24",X"22",X"22",X"22",X"02",X"82",X"84",
		X"EE",X"EE",X"EF",X"EF",X"FF",X"FF",X"FF",X"FE",X"80",X"80",X"40",X"40",X"60",X"40",X"70",X"E0",
		X"5B",X"43",X"7F",X"7F",X"7F",X"7F",X"3F",X"DF",X"84",X"84",X"84",X"90",X"97",X"8F",X"8F",X"8F",
		X"FE",X"FE",X"FE",X"FF",X"DF",X"EF",X"EF",X"F7",X"E0",X"F0",X"F9",X"E9",X"E8",X"DC",X"DC",X"DE",
		X"EF",X"FF",X"FF",X"FF",X"FE",X"FE",X"7E",X"1C",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"EF",X"DF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"D9",X"F8",X"F8",X"F8",X"F0",X"B0",X"90",X"D4",
		X"88",X"70",X"10",X"10",X"88",X"88",X"4A",X"52",X"3B",X"3C",X"3F",X"3F",X"3F",X"5F",X"7F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"12",X"08",X"04",X"02",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"12",X"08",X"04",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"C8",X"60",X"20",X"30",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"98",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"62",X"23",X"31",X"18",X"08",X"00",X"02",
		X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"98",X"00",X"80",X"80",X"C0",X"60",X"30",X"10",X"00",
		X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"04",X"87",X"83",X"C0",X"60",X"30",X"10",X"04",X"00",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"60",X"30",X"10",
		X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",
		X"02",X"03",X"81",X"80",X"C0",X"60",X"30",X"10",X"00",X"00",X"80",X"C0",X"60",X"30",X"10",X"00",
		X"30",X"18",X"0C",X"0C",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",
		X"00",X"00",X"80",X"C0",X"60",X"30",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"18",X"0C",X"0C",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"80",X"C0",X"C0",X"60",
		X"00",X"00",X"80",X"C0",X"60",X"30",X"18",X"0C",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"60",X"30",X"18",X"1C",X"0E",X"06",X"03",X"07",X"03",X"01",X"00",X"00",X"00",X"80",X"C0",
		X"00",X"80",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",
		X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"10",X"10",X"18",X"1C",X"0E",
		X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"10",X"1C",X"1E",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"04",X"07",X"03",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"02",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"03",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"18",X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"1C",X"1E",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"8F",X"77",X"E3",X"F7",X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"F1",X"F8",X"F8",X"F0",X"F0",X"E0",X"3E",X"7F",X"7F",X"FF",X"FF",X"7F",X"7F",X"3E",
		X"FB",X"FB",X"FB",X"FB",X"77",X"07",X"07",X"07",X"0F",X"0F",X"1C",X"1B",X"17",X"17",X"47",X"47",
		X"FF",X"FF",X"7F",X"BF",X"DF",X"DF",X"DF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B4",X"AD",X"69",X"69",X"78",X"78",X"78",X"7D",X"7F",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"47",X"DF",X"9F",X"9F",X"8F",X"8F",X"8F",X"DF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"05",X"03",X"03",X"01",X"01",X"00",X"00",X"00",X"FC",X"FE",X"FE",X"FC",X"FC",X"F8",X"70",X"00",
		X"5F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"00",X"C0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",
		X"00",X"01",X"06",X"18",X"01",X"02",X"04",X"08",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"74",X"BA",X"59",X"54",X"94",X"92",X"12",X"11",X"11",X"10",X"00",X"00",X"00",X"00",
		X"F8",X"00",X"E0",X"18",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"18",X"07",X"00",X"1F",
		X"00",X"00",X"00",X"00",X"08",X"88",X"88",X"48",X"49",X"29",X"2A",X"9A",X"5D",X"2E",X"FD",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"10",X"20",X"40",X"80",X"18",X"60",X"80",X"00",
		X"00",X"01",X"06",X"18",X"61",X"02",X"04",X"08",X"11",X"21",X"02",X"02",X"04",X"04",X"00",X"00",
		X"7F",X"BF",X"74",X"BA",X"59",X"54",X"94",X"92",X"12",X"11",X"11",X"10",X"10",X"10",X"10",X"10",
		X"FF",X"00",X"E0",X"1C",X"02",X"80",X"40",X"20",X"10",X"08",X"00",X"80",X"80",X"40",X"00",X"00",
		X"00",X"00",X"02",X"01",X"01",X"00",X"10",X"08",X"04",X"02",X"01",X"40",X"38",X"07",X"00",X"FF",
		X"08",X"08",X"08",X"08",X"08",X"88",X"88",X"48",X"49",X"29",X"2A",X"9A",X"5D",X"2E",X"FD",X"FE",
		X"00",X"00",X"00",X"20",X"40",X"40",X"80",X"88",X"10",X"20",X"40",X"86",X"18",X"60",X"80",X"00",
		X"00",X"01",X"06",X"18",X"01",X"02",X"04",X"08",X"01",X"01",X"02",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"BF",X"74",X"BA",X"59",X"54",X"94",X"92",X"12",X"11",X"11",X"10",X"00",X"00",X"00",X"00",
		X"FC",X"00",X"E0",X"18",X"00",X"80",X"40",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"02",X"01",X"00",X"18",X"07",X"00",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"48",X"49",X"29",X"2A",X"9A",X"5D",X"2E",X"FD",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"10",X"20",X"40",X"80",X"18",X"60",X"80",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"C0",X"40",X"40",X"60",X"20",X"30",X"10",X"18",X"0C",X"06",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"81",X"FF",X"1C",
		X"01",X"01",X"01",X"03",X"02",X"02",X"06",X"04",X"0C",X"08",X"18",X"30",X"60",X"C0",X"00",X"00",
		X"00",X"00",X"03",X"06",X"0C",X"18",X"10",X"30",X"20",X"60",X"40",X"40",X"C0",X"80",X"80",X"80",
		X"1C",X"FF",X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"60",X"30",X"18",X"08",X"0C",X"04",X"06",X"02",X"02",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"24",X"24",X"22",X"42",X"42",X"41",X"41",X"41",X"41",X"41",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"20",X"20",X"20",X"20",X"10",X"11",X"11",X"09",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"04",X"04",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"06",X"00",X"00",X"00",X"00",X"00",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"C0",X"C0",X"C0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"60",X"E0",X"E0",X"E0",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"60",X"70",X"F0",X"F0",X"F0",X"30",X"00",X"C0",X"00",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"60",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"18",X"E0",X"10",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"01",X"06",X"03",X"02",X"01",X"00",X"00",X"00",X"30",X"18",X"0C",X"00",
		X"14",X"3A",X"7D",X"FC",X"FC",X"F8",X"78",X"30",X"B0",X"A8",X"40",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"07",X"0B",X"04",X"02",X"02",X"01",X"60",X"60",X"30",X"30",X"10",X"00",
		X"0A",X"3A",X"FD",X"FD",X"FC",X"FC",X"F8",X"78",X"30",X"A0",X"80",X"00",X"40",X"20",X"00",X"00",
		X"00",X"00",X"13",X"0F",X"07",X"03",X"05",X"05",X"04",X"20",X"23",X"23",X"11",X"11",X"10",X"00",
		X"00",X"1A",X"FA",X"FA",X"FD",X"FD",X"F8",X"F0",X"E0",X"C0",X"40",X"00",X"80",X"00",X"80",X"00",
		X"00",X"39",X"1F",X"0F",X"07",X"07",X"05",X"25",X"20",X"22",X"12",X"11",X"01",X"00",X"00",X"00",
		X"00",X"80",X"0C",X"0C",X"0C",X"06",X"06",X"80",X"80",X"80",X"80",X"00",X"40",X"C0",X"80",X"00",
		X"30",X"3D",X"1F",X"0F",X"07",X"03",X"03",X"01",X"01",X"11",X"02",X"02",X"02",X"02",X"00",X"00",
		X"00",X"80",X"00",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"06",X"07",X"03",X"03",X"03",X"03",X"01",X"05",X"07",X"07",X"07",X"07",X"0E",X"0C",X"00",
		X"00",X"00",X"40",X"E0",X"E0",X"F0",X"E8",X"E8",X"D0",X"D0",X"D0",X"A0",X"A0",X"00",X"00",X"00",
		X"02",X"03",X"03",X"03",X"03",X"03",X"07",X"03",X"03",X"07",X"07",X"07",X"02",X"00",X"00",X"00",
		X"00",X"00",X"80",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"03",X"00",X"00",X"00",X"01",X"03",X"07",X"0E",X"18",X"00",X"00",
		X"80",X"80",X"80",X"F0",X"EC",X"BC",X"FC",X"78",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"70",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"C0",X"E0",X"70",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"C0",X"E0",X"F0",X"38",X"18",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"3C",X"1C",X"0E",X"07",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"F0",X"78",X"3C",X"1E",X"0F",X"07",
		X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"78",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"01",X"03",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",
		X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"80",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"03",X"03",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"A0",X"A0",X"C0",X"C0",X"60",X"60",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"06",X"02",X"03",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",X"40",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A0",X"F0",X"C0",X"20",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1A",X"1D",X"0E",X"17",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E0",X"F0",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"0F",X"06",X"0F",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"A0",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"F0",X"60",X"70",X"18",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0E",X"06",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D0",X"60",X"20",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"0C",X"0E",X"03",X"06",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"A0",X"20",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"03",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"40",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"80",X"40",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"40",X"40",X"40",
		X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"E0",X"C0",X"60",X"40",X"40",
		X"00",X"00",X"06",X"03",X"07",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"C0",X"80",X"C0",X"80",
		X"05",X"03",X"0E",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"40",
		X"00",X"05",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",
		X"01",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"00",X"00",X"02",X"00",X"00",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"00",X"02",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"80",X"00",X"00",
		X"01",X"00",X"04",X"02",X"00",X"04",X"01",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"05",X"00",X"04",X"02",X"01",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"80",X"00",X"80",X"40",X"80",
		X"01",X"02",X"04",X"03",X"00",X"04",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"80",X"40",X"80",X"00",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"05",X"02",X"05",X"02",X"01",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"40",X"80",X"40",X"80",X"40",X"80",
		X"05",X"06",X"05",X"03",X"02",X"04",X"05",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"C0",X"80",X"40",X"80",X"80",X"40",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"01",X"01",X"03",X"01",X"01",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"80",X"40",X"40",X"40",X"40",
		X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"40",X"40",X"40",X"40",X"80",X"00",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FE",X"E0",X"CE",X"7F",X"00",X"FF",X"FF",X"F9",X"38",X"78",X"FF",X"00",X"20",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"F0",X"E3",X"C0",X"E0",X"C3",X"58",X"00",X"00",
		X"E0",X"FF",X"00",X"04",X"82",X"FB",X"58",X"3F",X"07",X"F9",X"20",X"01",X"7D",X"0B",X"F5",X"DB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FB",X"FF",X"FF",X"FF",X"FD",X"FB",X"58",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"1F",X"FD",X"FF",X"4C",X"FF",X"FF",X"FF",X"7F",X"FF",X"37",X"8F",X"B9",
		X"FF",X"F0",X"F0",X"F0",X"E0",X"B8",X"BF",X"FC",X"BC",X"00",X"00",X"20",X"00",X"00",X"00",X"00",
		X"07",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"CD",X"0C",X"F0",X"1A",X"03",X"10",X"02",X"00",
		X"EF",X"F2",X"F8",X"FF",X"BF",X"BF",X"BF",X"BF",X"FF",X"7F",X"1F",X"9E",X"80",X"C3",X"E2",X"C6",
		X"F4",X"3D",X"00",X"3F",X"BF",X"FF",X"7F",X"BF",X"12",X"5F",X"03",X"F9",X"FE",X"FA",X"FF",X"FF",
		X"52",X"F1",X"FA",X"FD",X"3E",X"BE",X"FE",X"F3",X"00",X"88",X"C0",X"C0",X"00",X"A0",X"6D",X"33",
		X"00",X"00",X"03",X"00",X"00",X"07",X"81",X"81",X"0C",X"02",X"80",X"00",X"3F",X"00",X"FF",X"83",
		X"FF",X"DF",X"FD",X"F8",X"EC",X"FC",X"FE",X"FF",X"C6",X"CE",X"16",X"27",X"BD",X"C6",X"31",X"F9",
		X"3F",X"F3",X"63",X"7C",X"18",X"A0",X"FF",X"08",X"7F",X"5E",X"AE",X"A4",X"E0",X"03",X"1F",X"FF",
		X"83",X"8D",X"B5",X"FF",X"99",X"40",X"40",X"80",X"20",X"03",X"1E",X"80",X"46",X"DC",X"03",X"39",
		X"01",X"00",X"00",X"00",X"00",X"00",X"FB",X"F0",X"80",X"04",X"01",X"7F",X"22",X"0F",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"91",X"C4",X"E0",X"E6",X"E0",X"E8",X"F0",X"FC",X"CF",X"3C",X"17",X"03",X"60",X"38",X"F8",X"00",
		X"F8",X"03",X"FF",X"FE",X"7F",X"00",X"10",X"02",X"3B",X"B3",X"00",X"00",X"80",X"38",X"7F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"79",X"07",X"BF",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"80",X"11",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FE",X"F8",
		X"FF",X"FF",X"FB",X"CE",X"C0",X"00",X"04",X"04",X"FF",X"FC",X"FF",X"00",X"00",X"00",X"80",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"A8",X"C1",X"80",X"97",X"81",X"8F",X"17",
		X"00",X"76",X"57",X"D8",X"FF",X"D0",X"FB",X"FF",X"80",X"02",X"60",X"88",X"74",X"08",X"E8",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"D8",X"7C",X"CF",X"C6",X"E2",X"FC",X"F6",
		X"3F",X"41",X"3F",X"30",X"49",X"70",X"8F",X"AF",X"FF",X"FF",X"BF",X"3F",X"EB",X"0B",X"DA",X"89",
		X"FF",X"FE",X"FE",X"EB",X"EB",X"0E",X"41",X"4B",X"1B",X"5F",X"5F",X"FF",X"DF",X"76",X"FF",X"FF",
		X"FE",X"F7",X"FF",X"FF",X"FF",X"FD",X"FF",X"FF",X"00",X"FC",X"E0",X"F0",X"E0",X"E0",X"7A",X"FC",
		X"F7",X"FF",X"FF",X"FF",X"F7",X"FF",X"FF",X"FF",X"CA",X"C5",X"F5",X"F9",X"D3",X"E2",X"8F",X"4C",
		X"EC",X"2F",X"B9",X"9F",X"1F",X"94",X"DD",X"4F",X"00",X"88",X"13",X"1B",X"98",X"10",X"88",X"F8",
		X"A7",X"E3",X"7F",X"7F",X"43",X"C7",X"DF",X"83",X"17",X"EF",X"C7",X"DB",X"C7",X"DF",X"6F",X"D7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"F7",X"C0",X"FE",X"F0",X"F0",X"E4",X"E0",X"FC",X"D0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"B8",X"8E",X"83",X"E1",X"F9",X"FF",X"FF",
		X"AD",X"C4",X"4E",X"EF",X"C4",X"FF",X"FF",X"FF",X"74",X"33",X"37",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"D5",X"E7",X"FB",X"FD",X"FD",X"FF",X"FF",X"FF",X"8C",X"6F",X"17",X"89",X"01",X"80",X"80",X"85",
		X"FC",X"FF",X"7D",X"FB",X"5D",X"00",X"92",X"10",X"A0",X"40",X"00",X"80",X"40",X"00",X"00",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"40",X"E0",X"E0",X"F0",X"F8",X"FC",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"1B",X"19",X"34",X"4C",X"5D",X"38",X"53",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"FC",X"EF",X"FE",X"FF",X"FF",X"FF",X"2F",X"4A",X"15",X"92",X"D0",X"BE",X"F3",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7F",X"EE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E2",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"1E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"79",
		X"FF",X"DD",X"FF",X"BF",X"BF",X"DF",X"EF",X"DF",X"7F",X"E1",X"F2",X"F2",X"F0",X"22",X"B3",X"EA",
		X"AB",X"CA",X"01",X"70",X"26",X"69",X"EA",X"9B",X"FF",X"7F",X"3E",X"7A",X"34",X"25",X"80",X"36",
		X"80",X"00",X"00",X"20",X"5C",X"07",X"82",X"1D",X"00",X"00",X"00",X"02",X"BF",X"F5",X"00",X"C4",
		X"01",X"00",X"00",X"E0",X"FF",X"FF",X"3F",X"07",X"F8",X"2C",X"00",X"00",X"F8",X"7F",X"CB",X"E7",
		X"FF",X"BF",X"FF",X"DF",X"FF",X"FF",X"FD",X"FF",X"FF",X"F4",X"FD",X"DD",X"F8",X"FF",X"3F",X"BD",
		X"F6",X"18",X"02",X"93",X"9B",X"CF",X"BF",X"FF",X"79",X"83",X"33",X"F2",X"F8",X"F0",X"FC",X"F9",
		X"A2",X"AE",X"5C",X"7B",X"67",X"CE",X"9A",X"77",X"01",X"F2",X"FF",X"E8",X"8F",X"7D",X"E2",X"C7",
		X"00",X"22",X"FD",X"BA",X"E7",X"45",X"8F",X"BF",X"17",X"6F",X"6F",X"2E",X"6F",X"DD",X"F8",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"BF",X"7F",X"FF",X"7F",X"3E",X"9F",X"E7",X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"00",X"FC",X"FF",X"FF",X"7F",X"DF",X"EB",X"E7",X"CF",X"1C",X"80",X"D8",X"B3",X"77",X"70",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F9",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B7",X"5F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"FE",X"F1",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"C0",X"FD",X"1F",X"03",X"E1",X"7C",X"13",X"0F",X"1D",X"21",X"98",X"04",X"00",X"FF",X"FE",
		X"FF",X"FF",X"FF",X"FD",X"FF",X"F4",X"F1",X"E0",X"FF",X"FF",X"BE",X"FF",X"00",X"78",X"C7",X"33",
		X"FF",X"FF",X"FF",X"D3",X"05",X"A6",X"ED",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"5F",X"9E",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"D0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"1F",X"07",X"03",X"00",X"00",X"00",X"18",
		X"E8",X"F1",X"E0",X"C2",X"82",X"A2",X"82",X"81",X"C7",X"04",X"38",X"3C",X"3F",X"7B",X"BF",X"FC",
		X"B7",X"7C",X"30",X"1A",X"89",X"FD",X"88",X"38",X"E5",X"3D",X"9B",X"DF",X"25",X"9D",X"1D",X"B8",
		X"00",X"80",X"C2",X"E2",X"6E",X"F7",X"F0",X"8E",X"00",X"03",X"73",X"40",X"3F",X"8F",X"10",X"03",
		X"07",X"E6",X"03",X"FF",X"FF",X"FF",X"00",X"B3",X"C9",X"07",X"FE",X"FF",X"FE",X"FC",X"00",X"F8",
		X"E1",X"F0",X"F8",X"F8",X"F4",X"F9",X"FF",X"FF",X"3E",X"AA",X"63",X"11",X"0D",X"00",X"FF",X"DD",
		X"36",X"BF",X"5F",X"19",X"EC",X"3B",X"EF",X"FF",X"FB",X"5B",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"0D",X"1D",X"00",X"00",X"00",X"00",X"00",X"01",X"83",X"17",X"18",X"01",X"01",X"00",X"77",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"F3",X"EF",X"DE",X"9E",X"FF",X"FD",X"21",X"00",X"F1",X"07",X"3F",X"6F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FD",X"FA",X"FD",X"F7",X"FF",X"FE",
		X"67",X"FE",X"49",X"1F",X"FF",X"18",X"80",X"1F",X"BF",X"F0",X"F8",X"1F",X"FE",X"0F",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FE",X"FC",X"D8",X"A0",X"C0",X"B9",X"01",X"84",X"71",X"07",
		X"E0",X"01",X"00",X"31",X"2C",X"30",X"49",X"57",X"1D",X"C3",X"38",X"C7",X"06",X"FE",X"FE",X"FF",
		X"FF",X"7F",X"E7",X"3F",X"00",X"F8",X"60",X"30",X"DF",X"B9",X"4F",X"76",X"FB",X"14",X"FC",X"FF",
		X"E0",X"98",X"60",X"E7",X"87",X"40",X"01",X"C7",X"FF",X"E7",X"07",X"03",X"C8",X"E0",X"F9",X"1F",
		X"FE",X"FD",X"F0",X"F8",X"F0",X"F0",X"F0",X"FC",X"08",X"08",X"0C",X"12",X"11",X"00",X"19",X"01",
		X"83",X"47",X"C8",X"F2",X"25",X"1C",X"6F",X"FF",X"49",X"8B",X"03",X"51",X"07",X"0F",X"C3",X"FF",
		X"B9",X"98",X"CF",X"CF",X"8F",X"0D",X"81",X"73",X"FD",X"F6",X"FF",X"FE",X"FC",X"EA",X"FC",X"F3",
		X"C2",X"46",X"08",X"4A",X"E1",X"03",X"60",X"C0",X"E7",X"7E",X"00",X"06",X"F0",X"F0",X"3C",X"0F",
		X"FC",X"F8",X"FE",X"FD",X"FE",X"FF",X"FF",X"FF",X"11",X"0A",X"06",X"00",X"C0",X"FF",X"FB",X"FF",
		X"11",X"B3",X"F9",X"00",X"00",X"80",X"FF",X"F7",X"FE",X"F9",X"C4",X"17",X"16",X"BB",X"EF",X"FF",
		X"EF",X"C1",X"19",X"DE",X"7F",X"FF",X"FF",X"FF",X"FB",X"D3",X"EA",X"78",X"BF",X"FF",X"F6",X"FF",
		X"00",X"0D",X"FE",X"FF",X"80",X"78",X"7C",X"97",X"23",X"FD",X"01",X"FB",X"0F",X"61",X"00",X"81",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D0",X"E0",X"F9",X"F7",X"F8",X"FE",X"FC",X"FF",
		X"FF",X"7F",X"00",X"87",X"2B",X"FC",X"F0",X"00",X"F8",X"CF",X"1F",X"8F",X"F8",X"47",X"17",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E3",X"3E",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"1F",X"7E",X"03",X"87",X"D8",X"F8",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"E3",X"8C",
		X"FF",X"FF",X"FF",X"F1",X"4C",X"7C",X"7F",X"78",X"FF",X"FF",X"4D",X"53",X"67",X"00",X"FF",X"2D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FE",X"FF",X"FF",X"FF",X"F4",X"03",X"FF",X"DA",X"AF",X"77",X"81",X"FB",
		X"46",X"96",X"2C",X"7F",X"BF",X"BF",X"FE",X"04",X"38",X"70",X"E2",X"B9",X"FF",X"BF",X"3B",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"F6",X"ED",X"FF",X"FF",X"F0",X"FF",X"60",X"9F",X"7C",X"80",
		X"FF",X"FF",X"FF",X"E7",X"FA",X"03",X"17",X"39",X"FF",X"FF",X"FF",X"FF",X"7F",X"BF",X"CF",X"05",
		X"FC",X"FD",X"F4",X"F7",X"FE",X"EB",X"E7",X"43",X"04",X"FF",X"F9",X"F9",X"00",X"F7",X"E0",X"A4",
		X"FE",X"F1",X"9F",X"E9",X"10",X"C0",X"E2",X"63",X"27",X"42",X"F2",X"64",X"40",X"A7",X"B8",X"CC",
		X"F7",X"F4",X"AB",X"AD",X"BA",X"FF",X"FC",X"F6",X"41",X"40",X"8A",X"16",X"A6",X"98",X"20",X"02",
		X"83",X"C7",X"00",X"87",X"C9",X"81",X"CF",X"C8",X"83",X"11",X"A8",X"DC",X"28",X"A8",X"90",X"18",
		X"59",X"93",X"4F",X"13",X"27",X"27",X"03",X"57",X"1E",X"81",X"7F",X"18",X"6F",X"80",X"70",X"80",
		X"AD",X"20",X"FF",X"23",X"FF",X"00",X"0F",X"00",X"99",X"17",X"FE",X"16",X"7F",X"02",X"20",X"00",
		X"F7",X"E8",X"FA",X"C0",X"F6",X"E3",X"FC",X"FF",X"3F",X"1D",X"1F",X"00",X"1F",X"FF",X"F0",X"FF",
		X"BF",X"37",X"70",X"B7",X"73",X"29",X"FF",X"FF",X"80",X"87",X"2F",X"FF",X"7F",X"FF",X"FF",X"FF",
		X"9D",X"27",X"D8",X"C7",X"F7",X"FD",X"FC",X"FF",X"F9",X"B4",X"5C",X"0E",X"90",X"C8",X"7F",X"1F",
		X"BF",X"FD",X"7D",X"ED",X"10",X"20",X"FF",X"FE",X"EB",X"E1",X"65",X"2A",X"02",X"0F",X"C0",X"BC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FE",X"FD",X"FF",X"FF",X"FE",X"FF",X"C0",X"EF",X"08",X"A8",X"FB",X"EE",X"12",X"36",
		X"03",X"EF",X"FF",X"00",X"0B",X"3E",X"A8",X"50",X"20",X"1F",X"C0",X"C0",X"7C",X"72",X"27",X"DF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"40",X"F7",X"9D",X"F5",X"F6",X"FF",X"FF",X"FF",
		X"98",X"FC",X"F7",X"82",X"7F",X"9F",X"F8",X"FF",X"0B",X"FD",X"59",X"FD",X"87",X"E1",X"04",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FF",X"FC",X"F3",X"E0",X"F8",X"FE",X"C1",X"3F",X"1F",X"FF",X"7F",X"0F",X"5F",
		X"00",X"C0",X"FC",X"1F",X"FF",X"FF",X"7F",X"03",X"0F",X"01",X"00",X"81",X"FF",X"FF",X"BE",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FE",X"FD",X"FF",X"FF",X"FB",X"DE",X"E0",X"83",X"18",X"C1",
		X"FF",X"FF",X"FD",X"06",X"81",X"03",X"86",X"1C",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"3D",X"47",
		X"C0",X"80",X"86",X"00",X"00",X"00",X"80",X"E0",X"10",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"7F",X"07",X"03",X"06",X"82",X"03",X"14",
		X"F8",X"FC",X"F3",X"F0",X"E4",X"E0",X"E0",X"E0",X"16",X"1B",X"78",X"01",X"00",X"00",X"00",X"00",
		X"0B",X"C3",X"96",X"76",X"5D",X"62",X"1E",X"5B",X"34",X"42",X"71",X"9E",X"9E",X"A0",X"83",X"0C",
		X"30",X"D8",X"30",X"08",X"9C",X"29",X"E0",X"18",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"04",X"00",X"02",X"00",X"00",X"00",X"FC",X"07",X"02",X"00",X"06",X"7F",
		X"E0",X"F4",X"FA",X"FD",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"80",X"70",X"DF",X"FF",
		X"87",X"39",X"0B",X"16",X"0D",X"77",X"FF",X"FF",X"A4",X"5F",X"7D",X"FF",X"FE",X"FF",X"FF",X"FF",
		X"00",X"C4",X"00",X"18",X"81",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"1F",X"03",X"03",X"02",X"02",X"02",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F0",X"E8",X"F4",X"FF",X"FC",X"FF",X"FF",X"03",X"01",X"13",X"08",X"00",X"90",X"7F",X"FF",
		X"F0",X"C1",X"7F",X"7F",X"FF",X"FB",X"FF",X"F8",X"7F",X"FF",X"FF",X"FF",X"FF",X"FD",X"E3",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F5",
		X"FF",X"FF",X"FF",X"FE",X"FD",X"F5",X"97",X"2E",X"EF",X"D2",X"E9",X"DB",X"87",X"F1",X"39",X"47",
		X"18",X"7F",X"FE",X"E7",X"71",X"AE",X"FF",X"DE",X"3C",X"9E",X"7C",X"B8",X"A0",X"41",X"82",X"84",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C9",X"C0",X"0C",X"50",X"93",X"A8",X"8C",X"DF",
		X"5C",X"3C",X"F6",X"EA",X"9B",X"E5",X"87",X"F7",X"9A",X"7E",X"7F",X"FD",X"FF",X"FD",X"C9",X"FB",
		X"72",X"0C",X"EF",X"FF",X"FF",X"11",X"CF",X"AF",X"C5",X"EF",X"80",X"FF",X"FF",X"FF",X"3F",X"2C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"FA",X"EF",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"F9",X"DE",X"EC",X"FD",X"FE",X"FF",X"FF",X"FF",X"D9",X"3F",X"63",X"79",X"BF",X"43",X"5E",X"B0",
		X"0E",X"1F",X"0D",X"0F",X"83",X"86",X"2F",X"4F",X"FA",X"FE",X"5F",X"FF",X"7F",X"FF",X"8E",X"E3",
		X"BC",X"9F",X"FF",X"C2",X"B1",X"AE",X"8A",X"F6",X"F9",X"FF",X"FC",X"05",X"80",X"BC",X"A5",X"88",
		X"FB",X"FF",X"FF",X"EF",X"EF",X"FF",X"F7",X"F7",X"FF",X"DF",X"EF",X"FF",X"FE",X"FE",X"FE",X"FF",
		X"F2",X"F5",X"C8",X"F3",X"52",X"DB",X"F9",X"FE",X"04",X"E0",X"D8",X"00",X"FA",X"8F",X"83",X"E3",
		X"17",X"09",X"15",X"4D",X"0A",X"86",X"85",X"C8",X"C7",X"47",X"EF",X"DF",X"FF",X"BF",X"7F",X"FF",
		X"FA",X"F9",X"F7",X"F6",X"FA",X"FD",X"F7",X"FF",X"A2",X"7E",X"CB",X"44",X"65",X"F7",X"5F",X"1F",
		X"FF",X"FF",X"FF",X"FB",X"FD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3E",X"ED",
		X"F8",X"F7",X"F6",X"EF",X"01",X"88",X"00",X"3F",X"DF",X"BF",X"63",X"04",X"C6",X"2F",X"B7",X"6F",
		X"D5",X"8D",X"4B",X"B0",X"F0",X"F0",X"F9",X"FE",X"FF",X"FF",X"3F",X"7F",X"5F",X"FF",X"8F",X"AF",
		X"FF",X"FF",X"F3",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",X"14",X"80",X"FE",X"FC",X"F8",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"3F",X"DB",X"C4",X"FE",X"FF",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"EB",X"3C",X"26",X"07",X"88",X"FF",X"FF",X"FF",X"F2",X"7B",X"1C",X"20",X"08",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"63",X"00",X"81",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
