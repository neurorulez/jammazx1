-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "051117A0704D8044A14D22900410110F864E82D12E050080A76135DFDEA3F339";
    attribute INIT_01 of inst : label is "67D8F7E7918CFFEF2CDFF801541802AA9AAAAAA7C6A27D2F83FA42EF8F01523D";
    attribute INIT_02 of inst : label is "8E38D0DE43C9754B9ADC09E9013813D202790540D70B019B5DECC3AAA7B314D6";
    attribute INIT_03 of inst : label is "53E823E803E823E803E823E803E823E803D343D22397D9446ED9CA21BBE34D9B";
    attribute INIT_04 of inst : label is "A60509A154C050C230983C4FE954B51C8724E5107A2019A4C9B210130DF15553";
    attribute INIT_05 of inst : label is "A8C5463A39D1E8DBB27257DC2D0FB0BB2167D45A7F69785A2A0AA4012E35588A";
    attribute INIT_06 of inst : label is "A6A80A6C7308B6AB0C3E90244B28892FC4090F336492C90C9030EDD893242218";
    attribute INIT_07 of inst : label is "1C6AB170141D94A4749B5D62903152801B1EC229AA252E66116C0B5445067308";
    attribute INIT_08 of inst : label is "1C0444055B7372818812B379ACD3EE82410126C6300283180141085450B62304";
    attribute INIT_09 of inst : label is "4CD0F3A9CCEEA7333A9CCEB92CCAECBFCE4FE051444025FC4788888888888A09";
    attribute INIT_0A of inst : label is "222292427AC040AA0A00220002BB4ACACACA69869AA8AAAEEBAE8ABAA69AF8BA";
    attribute INIT_0B of inst : label is "2978C5806132BA08228B00B8D949951450245F4B37DE7F844587E1A2811259AE";
    attribute INIT_0C of inst : label is "AAAAAAAA8080C4EFAD9A00011244C4088C4D140902E90FC92596D9F624801011";
    attribute INIT_0D of inst : label is "2B4F59BF6B75D0FBA15A7AE511C4B2478C106D9B27B24998CC4018B980C086AA";
    attribute INIT_0E of inst : label is "0E86BA8CA3A8C3042BD3B58A881D10AD3D66BDACD541EA8569EBB4ED62A20744";
    attribute INIT_0F of inst : label is "BB90008814D6C496184DA8EDEC777B211212D29092C389251DBEC4C64405E480";
    attribute INIT_10 of inst : label is "EB624B089B51DBF036C476EAD8EEF6422216948496104928EDCC01A4C76E2863";
    attribute INIT_11 of inst : label is "AC8214361B7B0924B9FCF000F70879E0781E0780031BBB7C9D3D999599944005";
    attribute INIT_12 of inst : label is "A3124A3B7A99968F368E8D0A8D880D3BB18F31C62EFBEA1605A44382F5DB0BD2";
    attribute INIT_13 of inst : label is "26D476F7331FD264B46348476F5124A3B7A9997CDBA3136A3B7B998E9534DE93";
    attribute INIT_14 of inst : label is "84F4677555755556AA9D4E9D14470BAA081295150E9C223B79B76B4636D8EDEE";
    attribute INIT_15 of inst : label is "D93B4C93B4C88E35BA534FB22EE4EEE15E06FAD2FAD2BA92BA92B9373DC38144";
    attribute INIT_16 of inst : label is "F8DBF1B7E1951477EF8FDF1FBE3F7C6EF8DDF2038A3B9DC67B13FDDC505A9924";
    attribute INIT_17 of inst : label is "AC39D9718EEB0E765C60DB6D00514D78627AC14000151A7AC9CFBF1F7E3EFC7D";
    attribute INIT_18 of inst : label is "8C6231FAC73991C88A528C8D1052956DB492222000000590C420204081022DBB";
    attribute INIT_19 of inst : label is "922EA9AE8C7ACC7AEC7ACC7AEF0BFE40125D0C3F640082F82C0000BCBA398CC5";
    attribute INIT_1A of inst : label is "0121AF24975102A32635464C59A5EA285CDC4CB337132ECDC4CB337132EB0632";
    attribute INIT_1B of inst : label is "8CF91763BB9264A2945B6406E8A516D9301FBA45AC63141C048592A76416C507";
    attribute INIT_1C of inst : label is "77C8EBB807BD50F87136891BBF0C30C21E602C0A0F692BCE6610596227F38708";
    attribute INIT_1D of inst : label is "0CDDDC924776E362DF14D5AF004000C0A1FD83FA5D3D24F4DA610103A889C149";
    attribute INIT_1E of inst : label is "9F3F4FF9BED93388E98C75D452495249524AA482A9DDDD111190393A69A69A5B";
    attribute INIT_1F of inst : label is "B924924230F3A243A468985DD0AF08DA1D903F5B433815AB4875B3E5F9855548";
    attribute INIT_20 of inst : label is "4A02942528493FE340555351F5F36FB94999939924C9132250540CA082201187";
    attribute INIT_21 of inst : label is "25920B3E9A29683104929A4CC000CE6575AA0AA098CE19679797979797934929";
    attribute INIT_22 of inst : label is "3A36ECE2E9192F06123CDCE7A24065939C324027620023FBFE8AC42D82B80229";
    attribute INIT_23 of inst : label is "91C9643A121A1D1E8F47A1848430C30C229D07486EEEE888889E4358B7DDD6FB";
    attribute INIT_24 of inst : label is "F242CA2388A2D79D1EC5E992B871BA8B26592490F0A10E848024F2592C964723";
    attribute INIT_25 of inst : label is "BF9F7929B286F74BA7CFE96E9427B259F325B250327BEA311888B0B6B0DCACB6";
    attribute INIT_26 of inst : label is "97433B2592592C85674BA43A5D08EC964964B2159D2EF81937FD29F282F64B26";
    attribute INIT_27 of inst : label is "FDAE39F377F01C718F6F3E35CF8FFD480735EE7F3C4C964D7DEC965C9DD2E90E";
    attribute INIT_28 of inst : label is "F7B6AADACD85B84798AFF1E76F50306842074F33ED5893E5416C8909F4EE7A07";
    attribute INIT_29 of inst : label is "FC0C8D0BA9D8051188126C008880220A200094A8A39AE9B0D94D34D3BE5C16F7";
    attribute INIT_2A of inst : label is "B67E7CD4D7D3F86577268AE2E2B7C5618D320909E79EAAD1007C073287DB5FFD";
    attribute INIT_2B of inst : label is "3B0A98A6E6433329999A235CE811A66508D33A2A00A4D310D9C49B7BB6B8EE84";
    attribute INIT_2C of inst : label is "E7AE99D87515151514D3F18285FD467572527B7702DB500000000D715D487593";
    attribute INIT_2D of inst : label is "7D2C2BA888889DFBFC7FDDF852E9B17CD6E971DFB43716CF3246B63DFACB8D3F";
    attribute INIT_2E of inst : label is "9CB31109C23D772213C672CC442708F5CD99FAEA7EBA9BAEA7EBA9F5A9FFE428";
    attribute INIT_2F of inst : label is "19001D35B430C8FD4F7CAD370FF53DF2B70E74FA1F08816213413E9A7BC884F1";
    attribute INIT_30 of inst : label is "A855805621045C538EE8202027003FE7741002A40890B385B9953B3988180040";
    attribute INIT_31 of inst : label is "1FC78F13C21E4CA739DF2C8F13B8A03943A222C042CB1DFB0AF0F40110220440";
    attribute INIT_32 of inst : label is "EA0007C622E25051E1E8BEACCCCCCCC067A9050041041020F500C86080260800";
    attribute INIT_33 of inst : label is "9CE739CE739CE7154119FCABC5507E7F7FF445198B98B1110067E2FC540308B9";
    attribute INIT_34 of inst : label is "DD9EF8BB2F97FC05FF807BF08ABDF7C2BF6DDFD7EE6BCDDEA58D63420090A6CD";
    attribute INIT_35 of inst : label is "DEB004FD30D4DF90139D0663C926CE004042300E51373222AAAD73BEBD241EE1";
    attribute INIT_36 of inst : label is "1017081704170217011700970057FFC7ABEBABEEEE98C0008119842604FAABAE";
    attribute INIT_37 of inst : label is "CD42EE0445DC0ABA4E2BA42997D8753C7C70E9C1F18B85570057801740172017";
    attribute INIT_38 of inst : label is "CAAB9395476780A7CBE751D4501D8176EF8B1F5FFB070E5CBAA5E907A4168047";
    attribute INIT_39 of inst : label is "FBFB182A80003BAAABFFFFE3D3BF111F6E07333929DF4ED4F46A701864F541D9";
    attribute INIT_3A of inst : label is "09090003800042C042C0D310400000022A00E8AD62147BEAFBDFFFD9FF89F8F3";
    attribute INIT_3B of inst : label is "1117404052ED961119BBB0556837E007C17F0FC7EFDB7A89D61740C059900C01";
    attribute INIT_3C of inst : label is "39903870005CB83FE007A0105A56819FF0487B5AB105E854F6A4826F411C4441";
    attribute INIT_3D of inst : label is "5DC06464655101C0262E803983A72E0B8017057928AB556529DFD7F5C3970E1C";
    attribute INIT_3E of inst : label is "6464655180D69B019191955555555571029001ED5B4C6DBA48665D6597597597";
    attribute INIT_3F of inst : label is "F78100000000000000000004E8EC4EA283B13A8A0EC4EA283BAAAAD6D31501C0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "D60FAD542CD83676770085BB20A48347E2061F49F2162C04B5289E7E7E66232B";
    attribute INIT_01 of inst : label is "496F101050C0082008E20801995000CCD333333A485098C9664044444C71E808";
    attribute INIT_02 of inst : label is "815160979AF1543A87D40A63012814C6025E04203E44410562B71006C29C4961";
    attribute INIT_03 of inst : label is "62DC1ADC1ADC3ADC3ADC1ADC1ADC3ADC3ABAFAA11A8D8BAC4A951D612CC04892";
    attribute INIT_04 of inst : label is "486FAA37FE87FECAEF500589A154172851B86DB6274AABF5E2363AD7C050199A";
    attribute INIT_05 of inst : label is "111889C446222D432865E807F7D882639F5FF727216785AFD6A7539F3B61A5FB";
    attribute INIT_06 of inst : label is "7691C97EFF2C669FAE7370306FF33A4993D9F8846C92592B5BFD326C2CD949E3";
    attribute INIT_07 of inst : label is "F3B272D8CBF1D75AD4BB49CEC943D24F9FBFCB19A4648FF658EDFA48A4AF7F2C";
    attribute INIT_08 of inst : label is "967E92FF308637698CBFB24DAD9648D56AB4EDBD29FCCA94DE647D367DB7530B";
    attribute INIT_09 of inst : label is "18A2285221D148874D231F466F15919FD0CE1E4BC44406A82288080808008821";
    attribute INIT_0A of inst : label is "594829BF9F000000AA88938458201141414015F75DF5DF79369B6DA69F7DE787";
    attribute INIT_0B of inst : label is "D6822EE901ACEB6FB45DA9609653E9F69A9BA4B6880D1230F9F3E6B5F51649A5";
    attribute INIT_0C of inst : label is "55555555B3ED90E92CB20002400D3ADA0AF5AFA8A24DDF6B3496CB25576DF22A";
    attribute INIT_0D of inst : label is "64D592C5AC9E392C7366ACB6C9FECF2AEBAA8002552494665BCFB24CEDAD9155";
    attribute INIT_0E of inst : label is "E4C82E7B1667906FD0AB52ED5CD2B993565B76B3FBE7B7CD9AB26BD4BF5F3CBE";
    attribute INIT_0F of inst : label is "046E31252B293960CAB277132B8804C62FB525276439524E60659194ADAE22EA";
    attribute INIT_10 of inst : label is "35BCB0616DEE261E5B7B890F67101BCE594B6B7B21C296F3030BCA5B9810F64C";
    attribute INIT_11 of inst : label is "DAB134E4E44666DA2431864F206CBCF4BD2F4BD3D8B24C82AA42377656296550";
    attribute INIT_12 of inst : label is "5E2494C0C028329B3B8ACECACE4ACE4CCCC098130B4D93BA7A3E644F09653C0F";
    attribute INIT_13 of inst : label is "5B6B898250E72DDB4B44B79810225B4C0C1282B926CE2C95C4C02869C6C90326";
    attribute INIT_14 of inst : label is "200AA0CC502AAAA8AA92E1365B27D03B6CB28BF66939001CF6DDB5945B771204";
    attribute INIT_15 of inst : label is "766CBB265B964FA0ECEC922C89114197B1B1A5858DADA5858DADA780532D22FC";
    attribute INIT_16 of inst : label is "B2AD6F4EC87B2FD4B5793A52D5E4E95B57B3A75097DACCB2258527662FA7C259";
    attribute INIT_17 of inst : label is "CBAF364D699269CC974AB2CB958699D6CCD45B5555423CA39B28D6F0ECA35BC3";
    attribute INIT_18 of inst : label is "718DC25585FA5F526C2ED716E7617792CBE44C4C8C8C8E4F08B24599166A0926";
    attribute INIT_19 of inst : label is "C081B34922A491AC91A4B1ACB26C009DAC82E10106664DBC5993916F64CE330B";
    attribute INIT_1A of inst : label is "5A5ADF386ABEF81CC8F03991F65E0CC4912311A449C4E912311AC49C4EB055A5";
    attribute INIT_1B of inst : label is "C454BACC00268BA734E6C8B029CD39F3D2C0459FFEF734D1696D276F49EDCF34";
    attribute INIT_1C of inst : label is "8C2D1EE9F0632934F8C8B1609155D55C811264A6609F8295E099525A490C2225";
    attribute INIT_1D of inst : label is "B2600125B888E8B72DB938786CE6DE99B2032E072DA3968E434CF674044D3CB7";
    attribute INIT_1E of inst : label is "A1FF5FCC452A4625925B58BFD597D59FD59DAB3D7C26262626F90264B6592DAC";
    attribute INIT_1F of inst : label is "F8F78F303448D0EADA3DF7967B51F97FD67B472FFAC778ADDF4B7F000025555A";
    attribute INIT_20 of inst : label is "DF5FBE9F7D00802600199A63EA97A1F36C0081080840568872780EE502B281A2";
    attribute INIT_21 of inst : label is "1B4B600123E4F47D91242C999B6D99DA40145145111C8095ADE5ADE5ADE0024F";
    attribute INIT_22 of inst : label is "07848339E38803E2BFC408552C9D61C149A49D602529340200F9F6740F96D942";
    attribute INIT_23 of inst : label is "2C322F05CB258651699C5C22C90C10C10EA208ACB5353313130126A585B430B6";
    attribute INIT_24 of inst : label is "F70BD5F7F1E49F970097F53D41BC15D450A6592C0C32C7E93B5BC4ABE320B4CA";
    attribute INIT_25 of inst : label is "A824C6E04EE9C8984C121311374E45C24C5C45DDADE554D66B8773EA59BD5D63";
    attribute INIT_26 of inst : label is "31996CDC6FE6E372D8984FC4C2679170BE8B85CF266323E800066646EDC9B8DE";
    attribute INIT_27 of inst : label is "A6CAD3008012C396549071D93FD54694B2CA10F583B170BD51117093B66633D3";
    attribute INIT_28 of inst : label is "FCB25B48A06AB1FB8450FBFFC60D7AE5396B00FA026127008C9011926910EFD2";
    attribute INIT_29 of inst : label is "713338DB04E374AA25AEFC00A0A000888820465BB668A696723DE3CF0CD498AA";
    attribute INIT_2A of inst : label is "32F0003E415FF96FBCCFEEE56403CAE647DD5CD0040BFF1BF2F8FCFCF8D35039";
    attribute INIT_2B of inst : label is "315BA5F191B8C8D444673732371B991A8DC88CF367514536104AE048ADCC28E4";
    attribute INIT_2C of inst : label is "0F9AE18AD66226626754DA653B6664B491EC5DF467217800003BAE5327B3075C";
    attribute INIT_2D of inst : label is "B1B24CDF5F5F6A1DBD1780F8E79693AB2CB2A2A90AE5E29702A05277F592F01C";
    attribute INIT_2E of inst : label is "E1A4C5F7BDC7589BE7398EB117DE730D2D2E693D8A4F6293D9A4F66F7600164C";
    attribute INIT_2F of inst : label is "8112846BAD750AFA5AB5CF5E23E96AD73E2355FB4B71A9D3FD8814316066F9DE";
    attribute INIT_30 of inst : label is "12A79B9E66ACC9715548202025924BEB82335466C51A642DED818792C01CA052";
    attribute INIT_31 of inst : label is "208B32245EB0518059F33D11C1A9B4EACE485FCFFD96F6DECFF3AE6A2544A995";
    attribute INIT_32 of inst : label is "140000209D1991141E07414848484841288827A4C1441515E59309854A689CC9";
    attribute INIT_33 of inst : label is "B5AD6B5AD6B5AF940A861355E502818480785082746754147A981D0510408746";
    attribute INIT_34 of inst : label is "5B1761ED6DBD571355CC2B747DEE7A4BFBA5B2B47792A8ED4ED39CA7395B4A35";
    attribute INIT_35 of inst : label is "0127CDFE4C2DCBFC882232971A83116E7CAE0AC2441F67E1FFE3662802420AC2";
    attribute INIT_36 of inst : label is "00250025002500250025002500250025892D144050540111D545444454FAAF80";
    attribute INIT_37 of inst : label is "8BE2F00D85E059B8D01BE24925875B075C825A09C06B80D50025002500250025";
    attribute INIT_38 of inst : label is "C18DB3830B272067C625A169501ED158B311D41FF9A74A953CC9F027C0DF00E9";
    attribute INIT_39 of inst : label is "6684672AAAAA011557FFFFDEF87F3BE52E3729B84DE64EBEEE5F70001CF0D2C9";
    attribute INIT_3A of inst : label is "51110003D519139391111B586A00002A2225AD48B50904178402181710FC11B0";
    attribute INIT_3B of inst : label is "54162A256C011BBBB8000433197C3F007F408020103FF4A1D3F2418092534F49";
    attribute INIT_3C of inst : label is "A9E1AB500355B821E035C000301C33092DA8026B259D865804C155AB83CC5150";
    attribute INIT_3D of inst : label is "7955775D623F1E4EA0B008C7CBA76E1A80370DD224075EE94495374DDAA56ADD";
    attribute INIT_3E of inst : label is "775D623F9FDDD555DD7588FFFFFFFEF23CD23F8CC46CD1234CDE7DF79F7DE79F";
    attribute INIT_3F of inst : label is "100100000000000000000025AD887AEBA6216BAEB887AE9A62EEBBF3BAFF9B55";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "21DAFAE8C11C44FE3844C1BC90341147F206090252F48950240C2A2E2E774932";
    attribute INIT_01 of inst : label is "B88C9142D02462A52EAFF0FE1E60FCF0E43C3C238802B4E468C008C4514F3518";
    attribute INIT_02 of inst : label is "8D32A01662CC5602AB140ECD80281D9B0059860158C140125E56501AC9594BC0";
    attribute INIT_03 of inst : label is "83B823B803B823B823B823B823B803B802F9C2E8A39C71A42E044D20AD07170A";
    attribute INIT_04 of inst : label is "18E7864F7C5F7C42AE75C44BAFFF5F0F7FBE69B92D802FFFF48522A5F32E9E1C";
    attribute INIT_05 of inst : label is "998CCC7663B37CFE96D363D8C8C514A31D77F7E5A04678BBDAF44618AE5539CB";
    attribute INIT_06 of inst : label is "24C44C6A5A1B24CAFB2ED5753FC609CE326DC48C6D96596B1EEC4CD1D13563C1";
    attribute INIT_07 of inst : label is "9A5B2E788B89B73394B7C933A44893071A9686CD31260B443648E36226255A1B";
    attribute INIT_08 of inst : label is "28AF334997CC33B1263493EF64F24AED72DBB875283A62943D306C1C64A11283";
    attribute INIT_09 of inst : label is "A208079B45FE6D17F1B55D906DC6499FDACEB94DCCCE8EAAEDBB3BB33BB336DA";
    attribute INIT_0A of inst : label is "9B1CA9247710000000E4CB40DC8852D2D2D2B12492C92CB2CB2CB24B28A20A28";
    attribute INIT_0B of inst : label is "C65737B783BB93ACB16F7131DDCF65861DC626CDFC9FDB7930F84004C7325B65";
    attribute INIT_0C of inst : label is "AAAAAAAAE736B84B64B25042EA04AB6F1B20263D86FCCF793DB249251126998C";
    attribute INIT_0D of inst : label is "2ECE5870E6C38C87193672E89D486DA72EB8C4CB9292DCCFA21E673EF6B6FAAA";
    attribute INIT_0E of inst : label is "BC60BACEB38EE96713B973E1C6438C9B3967CFBF1E323C65D9CB1F3DDCF999F3";
    attribute INIT_0F of inst : label is "D99BBDC10C8E8CC369C999E464F33377B33191D1D84DB9A33C8EC6E7252CDA72";
    attribute INIT_10 of inst : label is "47474133DA3BE8A2768EFA298DF766AD724C8E8C8361ED1DF44443B4EFAA9837";
    attribute INIT_11 of inst : label is "6CC1963716E38B6CBAE6AB0E86A634D5B56D5B579CDB92099B6EB8971C8C315E";
    attribute INIT_12 of inst : label is "26334679571A86B46E805B891B891B939B0B616C2C5F69CC759932CCB6BA32DC";
    attribute INIT_13 of inst : label is "768EFAAE35B89A74764768EFA2E3B477D571ADC4D336334679571A9D636DEED3";
    attribute INIT_14 of inst : label is "7436633555755557D53CB4D9A635160C462049972C3E8EF609A7474C769DF55C";
    attribute INIT_15 of inst : label is "99BA4E93B6EC6A471336DEB9DFB8C669C1BA0E2E262626060E0E0ECE3CD13265";
    attribute INIT_16 of inst : label is "DDD3B1A364FB266ECE8D8D1B9B7776ECE8D8D35993170BC2F303DCCC37656936";
    attribute INIT_17 of inst : label is "8CBB9C65DCE32E671D72FF68C3C840C00642624000003672EDDD3B1A36366EED";
    attribute INIT_18 of inst : label is "5AE5779EFE7B09984772C1BB323B9729B7BB3BB8D9C8DF1E33191336688A6DB3";
    attribute INIT_19 of inst : label is "63E6B3CEC970EA70EA78EA78E9EC1F463B09345E1230E44CE4193B13D06B95DC";
    attribute INIT_1A of inst : label is "1D1990187299B633A20E46665C8FA4662A381C3A8E070EA3C1E3A8F078E9F739";
    attribute INIT_1B of inst : label is "FBA37D679D98760F81F164BF43E07C18A2F9D76D6A5200547460D28434408215";
    attribute INIT_1C of inst : label is "0FEED537DAFD8C94DBDFC9853E18E387CEE26FFC666ECECD8A0C1C626F679DDB";
    attribute INIT_1D of inst : label is "3DBCECDB4F3ACBCF937CDE5088B3678C9981F3E589F2C7CB53F39978B30FC646";
    attribute INIT_1E of inst : label is "BDEADAACF5BB6E64C66C63A627652764276A4EC8563773BFFB4C993B49249B33";
    attribute INIT_1F of inst : label is "A4C30D717469937BB24FDD988B2349D3188B243A6311748F4C61CF9080322A9B";
    attribute INIT_20 of inst : label is "1B86372C6E40DFC3409E1C802997C7034B85C55A0AC2469CA15CDEA336A18BA3";
    attribute INIT_21 of inst : label is "BFF32FADB32566B0C508A926649265712DE79E79EE5F48CFF7B7BFFFF7B9548B";
    attribute INIT_22 of inst : label is "9D97E78963DA89A3FFD956B32CDDC3629526DD800108302964C9D30BB7FF6B3F";
    attribute INIT_23 of inst : label is "986C261241924D36CA6D268A645965145AF73FC61DFB9D9BB9CE4AD917FCE2FF";
    attribute INIT_24 of inst : label is "F69DD8C7F460DF9F14D7F1BC546494C5176DA490101916CE8C741A0D26C34522";
    attribute INIT_25 of inst : label is "ECD32D38B876A34FB06969EEC3A51B7D31B7BA0E3A501528948471388CBD9D39";
    attribute INIT_26 of inst : label is "DF4DB9A7DA2D3EDB734FB45A7DB6E6DF48B6FA6DCDBE9918332DBAF076A34FB2";
    attribute INIT_27 of inst : label is "59B73C5333F2CCFB9DABB664E978A8D8BF76AAF89CE6DF45DEC6DF6CDCDBE936";
    attribute INIT_28 of inst : label is "F029482223D8893033C07AF39A0C42830846027C38523704C0DC991B4DAAF37E";
    attribute INIT_29 of inst : label is "5DB84CC82D0A758F76CC8000AA00880A0880664B306454565B30C35C8694D811";
    attribute INIT_2A of inst : label is "10B3366F091FF16F184F443CFCA4793C975A70C511855503E4F8E6A6F0B6D629";
    attribute INIT_2B of inst : label is "085EB4CBBAB59D52EEA43AF7665D73BA2EBDDD3B96454830628CE1693AD14CE4";
    attribute INIT_2C of inst : label is "AFA63042D333377735D7A747BFD66FE7E3FEF5F545BA7955557EAF93FBFCF0C6";
    attribute INIT_2D of inst : label is "3DBB8EFFF55FFF76FEDFDCF8B7FFA2EDBFFFDB77FEDFF8DC32CEF65FF7FFF901";
    attribute INIT_2E of inst : label is "16B911C9E629623393CC52C4673798A599BB3FDFCFF7F7FDFCFF7F7BFF0017A7";
    attribute INIT_2F of inst : label is "8A51C46A8C532A0DCEB4FB0C00373AD3EC0311FA7D1D8D57378018217A88E6F3";
    attribute INIT_30 of inst : label is "93378CDE02644F1B514D7465769017EB8210AA058B033F4834AB9308E5BC76D1";
    attribute INIT_31 of inst : label is "05DD9B35D7BF0D90A0E007008BA0A43EC354D5C08493DBC345F0FA33266CDC99";
    attribute INIT_32 of inst : label is "EA00001362E6311001F8BEA848484844063009205B45B7011180E0635206AC48";
    attribute INIT_33 of inst : label is "8B4AD2B4AD2B4FE5B45BEEABF96D7EFBFFFF5A4D8BBAA3D68567E2FF188C58B9";
    attribute INIT_34 of inst : label is "5A80315C6C2AA65900D83B264C0EEA4EF3BD874F76C75EEDF79DEE718E736F7B";
    attribute INIT_35 of inst : label is "20498BD7100CA3E4CB66B3E768AA15B2603504C2CE3D3B2155636815B3630EC0";
    attribute INIT_36 of inst : label is "0015001500150015001500150017FFD5E05EEFBD40811414540FAD6FBBEEAAE1";
    attribute INIT_37 of inst : label is "4722C924059208B9C90BFC90952857347E49F925C9A38B050015001500150015";
    attribute INIT_38 of inst : label is "D60503AC0A07811743D5C570701F515AB40A565403050A54AF05F947E05F806A";
    attribute INIT_39 of inst : label is "020480FFFFFFFAEAA800003553C0004F0E07A2B995E92E70FE38700468EB0281";
    attribute INIT_3A of inst : label is "D0504093C14B8101010112123F00003BBB88CB418718001580220428101A172A";
    attribute INIT_3B of inst : label is "55462A649EA89DAAADAAA80F048015002A800000000001FC240EC30112395443";
    attribute INIT_3C of inst : label is "A898295000543821E007E020B58C580618082C74C28A5F9C58E3CFD024005545";
    attribute INIT_3D of inst : label is "715FB9318F59D9220C3422D5E3970E0B8007057722945C4DC21C5715CA972A54";
    attribute INIT_3E of inst : label is "B9318F59599CF17EE4C63D555555556B3298330CF54CC1EA78CD71C71D75D75C";
    attribute INIT_3F of inst : label is "07800000000000000000000CC900CCBFFC03B2FFD00ECBDF40AFFAFF9E49CD5F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "4C555141100144CCDB46019C90103107D3860C9A44EB8955060448C8C9D69822";
    attribute INIT_01 of inst : label is "0DEED3F7A88452BF272C50001F8000FF003FC01E26F9401537C604C2C0B5CAB4";
    attribute INIT_02 of inst : label is "8518305602C1550AAB540AC500B8158A017805015B0300084AF6C3066BDB0D02";
    attribute INIT_03 of inst : label is "0298029822980298029802980298029802B8C398428E21042A284820BD800203";
    attribute INIT_04 of inst : label is "ECB4EB2A4A9A4A8A1FB9CF84C40011A1382A829F01CA941A3603A06741041FE0";
    attribute INIT_05 of inst : label is "88C446223111950D48A3BD94D6D150370F6BF56F814682E0DC37EB0D8AE421F5";
    attribute INIT_06 of inst : label is "275C4C1DAD332754014ED569D05A11BF524EFE042CB249517145C8919125BCB8";
    attribute INIT_07 of inst : label is "FDE543E753FDFF6284BEC9F32478D337C76BCCCDD7263DBE666AF2AE261BED33";
    attribute INIT_08 of inst : label is "BED2D249DA940726C6FCB65B64B24EE773DB29F2D6BE6D6B5F37F5EBBCBD19CB";
    attribute INIT_09 of inst : label is "00001B0BE49E2FD278BE49DE21C7E0841E41BE38CCC8EDF8EF3B3BBBB333BCD3";
    attribute INIT_0A of inst : label is "3368ADB53B8010504472E780CA8D52929292A208200200000000000000000000";
    attribute INIT_0B of inst : label is "E7DA63A9101DF16556C76BD80ECD3EAACA8E36DDFD9E49D0BCD3260750064967";
    attribute INIT_0C of inst : label is "FFFFFFFF2B76D0092492EBBB46008F6A06303A83A0DADBDB3C92492711A49DF9";
    attribute INIT_0D of inst : label is "768BEE3856E1EDC3DBB45F5DAADCFFA5D59CC6C97292CEED272FA21E36F693FF";
    attribute INIT_0E of inst : label is "ED6EDCF735CD7933695CAF72F6E5EDFA2FB8C15B06B60D6ED17DC70ADC3DB87B";
    attribute INIT_0F of inst : label is "99DEB7A92D8ECC836CDD99E574F33BF7F73DB1D9D06D9BB33CAE5452D1284068";
    attribute INIT_10 of inst : label is "C7666131BB33CAE26ECCF2A1B9E677EFEA6D8ECCC360DD99E5444376CF221A27";
    attribute INIT_11 of inst : label is "7F55AAF2DB6D5925948CDB6F45B6CB6ACAB6ACABCDD57209917C98AB4B8DB474";
    attribute INIT_12 of inst : label is "363766791B10A400470511E011E151FBBBAF75EEB7FB49AD7BFA34FD2CB6B4ED";
    attribute INIT_13 of inst : label is "6ECCF236214ADA766646ECCF2B63766791B10AD6D3363766791B10A6E124ECD3";
    attribute INIT_14 of inst : label is "2C624A2800222220002B749D72E34A1656C6AFA165958AA2ADA7664C6ED9E46C";
    attribute INIT_15 of inst : label is "DC9F07C9E27186E3BC925CD68D10945D85982C2C2C2C2C0C040405D428BB2BAC";
    attribute INIT_16 of inst : label is "5A54B4A96C8E3A8ADAB5F5EB6A96952D2A5A54F95D7D6A5A9602B8B80FEFE9A6";
    attribute INIT_17 of inst : label is "E71C8F38E479C723CA3B4932DB4DAC8DE6843BB5555F428450B56B6BD7D5AD2A";
    attribute INIT_18 of inst : label is "EF57AABA7AFD6CBB6A5D78F91F52EAED24DAA2222E3B3DE5F3DB9E2C58ADF7D1";
    attribute INIT_19 of inst : label is "EA24D99495567756775677567F3E1746330D36018BB5D75F57D975DF1EBD5EA8";
    attribute INIT_1A of inst : label is "9BDB982E3AFBBB2777E66FEFAB7FB556E79B4D1DE6D34779B4D1DE6D347D1A97";
    attribute INIT_1B of inst : label is "3BBFA7EFDD9FB5D4FA9FEC1F753EA7BB907D927FF6B730AE6F6ED273B45CCE2B";
    attribute INIT_1C of inst : label is "C7553B65FBFCACF871DD4EB324796597CEFA5AFD6FEDC0CE03EDABA82F75CCFD";
    attribute INIT_1D of inst : label is "9FBEECFACF3256E4FAA7EEEC88B765CD5A439217896BC5AF12DB1F363BCB47C6";
    attribute INIT_1E of inst : label is "92BFCFF5F8B976A75A752DBAE264E265E269C4CBFE5111D9996D99B24936D23B";
    attribute INIT_1F of inst : label is "E1D71C7158231B896371CBAB8F7749F54B8F743FA971FE87F52D5FE1C8955541";
    attribute INIT_20 of inst : label is "9DD73B8E7740CA02801FE00249314059358D81D80EC054689114562014800AC1";
    attribute INIT_21 of inst : label is "6495492C99702218D508A937679EECA924C71C71DDCACCDA7A7A72323239548B";
    attribute INIT_22 of inst : label is "133B4419C1D805BE3B8006A74EF840489416F842A121D42B6E5C636D5AE7634B";
    attribute INIT_23 of inst : label is "9068345A65BA6934CA6D36C16E11451409DDF566EA888EA888CE034B3368866D";
    attribute INIT_24 of inst : label is "FE8CFA67B00677CC064DF49518449CC71A3924D0705B06CE8C761B0DA4C26532";
    attribute INIT_25 of inst : label is "67FFFD183C6A6F47FFFFE8DFE3437B3FFFB37F8D953403BFDF8C23284D130B00";
    attribute INIT_26 of inst : label is "8FDC5FA1FF3D1FF8BF43FE7A3FF17EC7FCF67FE2FD1FFA50B3BD1E34686F47FC";
    attribute INIT_27 of inst : label is "5D65AB5B32A85CEFC9A33674E03CBE5E1DFEE24C7CEE8FD8CFFE8FFD2BD0FB9E";
    attribute INIT_28 of inst : label is "FA487C0A35DF33987FDF8A986F2DC39DEF740755EFDCE6DC705B8F0BE5E25D54";
    attribute INIT_29 of inst : label is "01D196D7F9FB3AA226CA6802000022000200CA759541D41A7875C71CDAAAB4FF";
    attribute INIT_2A of inst : label is "50F71C4C3242FCC4C784570FC7F41F87C28DF6D990091141707E7E60FC2C9105";
    attribute INIT_2B of inst : label is "B16D3CEB3BA59DD2EEEEDDE754AEF3A2577DD1B3FA7549B54587FB331D52C7F8";
    attribute INIT_2C of inst : label is "C4463D8B71111555198739539EB5DB792197AC0D5BFAC955557FF48A4A5EA887";
    attribute INIT_2D of inst : label is "EF397FF5555FDFCE7E4FCD7E334FA5D6FA4B75DCADBB384F55EAB4ADEF5D9940";
    attribute INIT_2E of inst : label is "C4D7B8D96789AF61B2CF135EC3759E26B09BD252F494B9252E494B98CBFFE972";
    attribute INIT_2F of inst : label is "01404C29C47101FC460CB92D13E1983AE11258F82D5C8C323340192495DC6CB3";
    attribute INIT_30 of inst : label is "47299CA26264441A40082021346207E5402222D2C74B700571B3111CC8AC0290";
    attribute INIT_31 of inst : label is "144489154D32CC943C6383024A80B8F40F9440CA9687BC87A4F3C072CE51CA3B";
    attribute INIT_32 of inst : label is "1400000C1519434A0005414848484850679C09840A40A405A190C160506720A1";
    attribute INIT_33 of inst : label is "AB4A56B4A56B4FDAA02DFD55F6A8037F7FFDA03074CD416800181D00B7302546";
    attribute INIT_34 of inst : label is "32C2624D1D617CC4FFE816355FAE0A68DFB396D2F486C5E91E7694AD6B5B2F46";
    attribute INIT_35 of inst : label is "201C9BFDF04D72AA2CEC1E4748AA45B32E3484E0F40525700060E53C996A0588";
    attribute INIT_36 of inst : label is "1017081704170217011700970055FFD5D3C6BBEEBAFAEBAEF80BBEAF5A040030";
    attribute INIT_37 of inst : label is "03024504048A08ABC50AE00217C05110582958A5E80B84170057801740172017";
    attribute INIT_38 of inst : label is "C8070B900E178007CB47F1FC501F917AF6005417FB152A142FF5F817E01F804B";
    attribute INIT_39 of inst : label is "0404848000005015555555414400001D2E1750B885EC2E32EE19701402E40385";
    attribute INIT_3A of inst : label is "83435002120242424242511A1500001416169481871804158422100010001504";
    attribute INIT_3B of inst : label is "455280038112604442444D80FC402A0055408020102491F74D54860200359213";
    attribute INIT_3C of inst : label is "B98029500054A8202015E000BA046E6005F580870E7311E301123810320C0015";
    attribute INIT_3D of inst : label is "51FFBB192FAA1BA28EBE2A76BB972A0A8017054221087E494057D5F54A952E54";
    attribute INIT_3E of inst : label is "BB192FAA9A94B7FEEC64BE8000000092B48F356A7E685DF37C54514515555555";
    attribute INIT_3F of inst : label is "04010000000000000000001694C36956130DA5504C36954130BAAE5C968979FF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "1101141041010066D191D51802828A204020DD8EC3E200A15A53C02C2D440D33";
    attribute INIT_01 of inst : label is "E07617FF8904429F6C2050FFE000FF0007C000123AAD81D116342626C9557054";
    attribute INIT_02 of inst : label is "006B0000E81D00A80440000000800000010380A022069E45243BA78008EE8221";
    attribute INIT_03 of inst : label is "F861E860E860E860E860E860E860E860E8030801C8000A8A208114508010D080";
    attribute INIT_04 of inst : label is "504924049224922F79260BE08D55E85011AF80C2AD000C1628642D5460A8E000";
    attribute INIT_05 of inst : label is "998CCD776BBB23480100892290915B5052983180B404AEE406C118B3D26AA990";
    attribute INIT_06 of inst : label is "C033432848AEC03440D3602404140883209028C8082400004441332526CE0521";
    attribute INIT_07 of inst : label is "5080CA56025126DB0024804CDB4680D48A102BB00CC189015D829119A18508AE";
    attribute INIT_08 of inst : label is "8028A092614834D8058B25A2416000341E66D08A10A45908522D13460B04D22A";
    attribute INIT_09 of inst : label is "00000089D59A2756689C59AA61B631801EC03022C44604AC2280800000000A00";
    attribute INIT_0A of inst : label is "52510602401515005039F944CD06840404048800000000000000000000000000";
    attribute INIT_0B of inst : label is "90840ACE330D28C10D15CA5186840831C701A9324B45B6218921155133348048";
    attribute INIT_0C of inst : label is "000000006ED920700901FBA88004019418AA899926909412480090005A592762";
    attribute INIT_0D of inst : label is "C7F00260C68B0B16163F8012A8386C380134C8884AB6DA88801C542019196000";
    attribute INIT_0E of inst : label is "B0598581605A110263346355A5AB4B1FC009A31AAD2D5A58FE004C18D16162C2";
    attribute INIT_0F of inst : label is "11252B31C92928400492510650822484652925254800124A20C81B309D3AC04A";
    attribute INIT_10 of inst : label is "1494208124A20C8A492883312104494ACE492928400C92510671724908339384";
    attribute INIT_11 of inst : label is "1A3161E0CCD874D3076312E95125A28BB2ECBA2A402049032378B00242212D58";
    attribute INIT_12 of inst : label is "802494419421082B010F8053805380464648C919216DA1214A572D6B4804ED2B";
    attribute INIT_13 of inst : label is "4928832842142489508C928832824944194210A12480249441942101036D8924";
    attribute INIT_14 of inst : label is "E00A8C0082FD7D7DD50283224AA0D50945ED0260C3B10441C2489520C9210650";
    attribute INIT_15 of inst : label is "2384E1304E1541860236D8850AA91803C7AA3E1E3E1E3E3E1E3E1C484006A099";
    attribute INIT_16 of inst : label is "C3C7878F08A209EE3E7C3C7878F0F1E1E3C3C51104D85D174504644424A40649";
    attribute INIT_17 of inst : label is "410582082C1041608208DB6CB38290E685EC482AAABF41A41C3CF8F8F0F1E1E3";
    attribute INIT_18 of inst : label is "18D46A96F6406D93666E15DBBB33709B6FB7777BABAFA8690C9664C993219330";
    attribute INIT_19 of inst : label is "24511B013688168816881688161551B5A104800BE22F54E55175D539056351AA";
    attribute INIT_1A of inst : label is "7312DCEB2826CC4000488000C2EEA445E7B2D985ECB6617B2D985ECB66110085";
    attribute INIT_1B of inst : label is "311E279C156F10C438879899610C21E7826510296350BA8DCC4E4D3593642CA3";
    attribute INIT_1C of inst : label is "AD0341552B66CC4A431C3864C99E79E78BBFEDC4E13E47024C0B06186D5408B1";
    attribute INIT_1D of inst : label is "1720AB6828A290C43221CA0268AD974B16A94CACA4D6535109AF57AD4EE6D5D5";
    attribute INIT_1E of inst : label is "34AA8AA440B1685415610AA1C03640364034806C40BBBBBBBB8B164DB6C924A1";
    attribute INIT_1F of inst : label is "61C34D31A208DDB8DBB7C6022ED1B178C22ED66E1845CAC5C3089F2420088003";
    attribute INIT_20 of inst : label is "846919D611970AB56AE000FA26614B0B220400400A0050503BAB4B54D2DA0D10";
    attribute INIT_21 of inst : label is "5A0852526042B358B85506181201800FEDBEF965B0D88CB63636363636319115";
    attribute INIT_22 of inst : label is "13FEC4D980C01DB86B5004333EC9C320C756C9C17515052E981072C25C0D9242";
    attribute INIT_23 of inst : label is "082400C9296924821100800058830C1009334CC599999999998BB427FED89FDB";
    attribute INIT_24 of inst : label is "098C2412C014C05814E00DC35298211451E000080816A12B6B40000020402412";
    attribute INIT_25 of inst : label is "564C0211C2480884422610B112504522C052C4498D05402010830AA00B02C2E8";
    attribute INIT_26 of inst : label is "08A2044221A211050884434422081148868A4414221164610AA215CA4A088441";
    attribute INIT_27 of inst : label is "5649C05022A2408AD0B233192534A648985AF2D4262309A2A8230992422114D1";
    attribute INIT_28 of inst : label is "0808150C0872D38383B062CA42891A2318E80855300B120266584CCB44F2CD58";
    attribute INIT_29 of inst : label is "D948209C5602A22553282688000011200805001C8C1091001070D34C048A0388";
    attribute INIT_2A of inst : label is "54BF5C6E3068028040C1DD0D05489AC440EB6C959A11051C17011420C9BEDC6D";
    attribute INIT_2B of inst : label is "E1423334AB1A518D0AE3841453860AA9C1011073211822278D8C6F6F3956CC68";
    attribute INIT_2C of inst : label is "804E370A033333333186014985E056636B927C0B019644000011104EDA4A7986";
    attribute INIT_2D of inst : label is "9C18566AAAA00806C2D85E0130CB60CCB6CB10458E9734CA38E66C1806DB9A1E";
    attribute INIT_2E of inst : label is "630C689110C618D122218C31A2544318699336D24DB4936D24DB4939C9000850";
    attribute INIT_2F of inst : label is "0D1A092102A9D7F505082429ABD4942895AAE085A0D85EA9A26C02AA6A344888";
    attribute INIT_30 of inst : label is "0DA0568174CA91A961420202068B401451AA679CB9F32037200884C55E969A5A";
    attribute INIT_31 of inst : label is "A4CD9B3D2C23F23F3EEBD75A794D42A02A0CE4298F9A11A2040A815A1BC3686D";
    attribute INIT_32 of inst : label is "EA000040CAE4FC820012BEA84848485FB8B0A356E94694178D5B2594457802D5";
    attribute INIT_33 of inst : label is "38C6B1AD6358C7888B1612ABE2228584807A29038B76BC8A02E7E2FF6AA112B9";
    attribute INIT_34 of inst : label is "E8CDB35670EA80BA00687D643148EB24E696373CC2973985673DCF7BDCF7244C";
    attribute INIT_35 of inst : label is "00039B50480E921A0C20191512C080CA0E5C92A5A81058420043A855B92A1F59";
    attribute INIT_36 of inst : label is "00000000000000000000000000000000021EEAFBBBABEEBAA80EBAFEFFBFBB80";
    attribute INIT_37 of inst : label is "6C2034A94069520214A01CD9C8C50A0106A40290244808900000000000000000";
    attribute INIT_38 of inst : label is "11282022404020000C080601A060020002572003FC8000000004BB52ED43B880";
    attribute INIT_39 of inst : label is "440010BBBBBBBEEFB844446156C0045801C08E00100180C00060001210189010";
    attribute INIT_3A of inst : label is "40C0C04040004040404041507F00002A9DF527A38E38002A0020040800100004";
    attribute INIT_3B of inst : label is "9AAA7DF87AEDFFBBBFBBB07FFEAA2A0055408020102491FFE998CC040027C041";
    attribute INIT_3C of inst : label is "01388000010080800012EE20040F901FF8007FF8F1FCEC00FFE5FFEFC55F2AAA";
    attribute INIT_3D of inst : label is "005FFFF747C3331A8CBCAAF41800000000000005870502841602008000100000";
    attribute INIT_3E of inst : label is "FFF747C3B201A57FFFDD1F7FFFFFFF3E250624040C0110401110000001041041";
    attribute INIT_3F of inst : label is "90800000000000000000003725A172551E85C9547A172551E8FFFF003486365F";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "AF8FAAABFFAD95EEF3C2E51924C0E208440C95194A0C2BE5140035D151664B03";
    attribute INIT_01 of inst : label is "01071850BA08CDA14DE0E800000000000000002AAAABBAB17EEC3EE771AA8FAA";
    attribute INIT_02 of inst : label is "800000540281500A8054000000A8000001500000020E1E0000838780020E0000";
    attribute INIT_03 of inst : label is "0281E280E280E280E280E280E280E280E2800280028000002A000000A800000A";
    attribute INIT_04 of inst : label is "D61A65A1A621A6084B15DEEAA955501DBDFF8B8272754C1E3996760EE0790000";
    attribute INIT_05 of inst : label is "998889666A222B420840C8049493227546C82B9072D4CAA26E5B39871868A132";
    attribute INIT_06 of inst : label is "EDB35B01082EEDB14AC370301294880A249B70992492490A51691225244C0821";
    attribute INIT_07 of inst : label is "E106D29022E096CB2D92498EDB46B6C580400BBB6CED91085DDAB6D9AD91882E";
    attribute INIT_08 of inst : label is "8A24A4937D291249159993F9249249B4DA26731C202D5A1016ACBB56DBA0D64A";
    attribute INIT_09 of inst : label is "00000C5B4C136D704DB5C10101349C001000D2E3E66466042200888888880A20";
    attribute INIT_0A of inst : label is "5653A44BC2551555003E54048184C6C6C6C60000000000000000000000000000";
    attribute INIT_0B of inst : label is "94848ECE416CCE796D1DCA50B6400F3DF330A0324000122488A5451931124924";
    attribute INIT_0C of inst : label is "00000000AA5BA449249315509C4401BC88A8C98B224A96C92492492452593762";
    attribute INIT_0D of inst : label is "D4ECF64894A24B4496A767B28A194CD67B34C192D726439490CCCCE10989E400";
    attribute INIT_0E of inst : label is "B2592D2B4AD0B20643244A5125A24B53B3D92252892D125A9D9EC91294496892";
    attribute INIT_0F of inst : label is "366E33214B6B6B24F196D20E8106CDE764216D6D249EB2DA41D2B1159D6B4D4A";
    attribute INIT_10 of inst : label is "35B5927B2DA41D1A4B690741620D9BCEC84B6B6B24F596D20E93525B90749688";
    attribute INIT_11 of inst : label is "C9BD7DA58042D2002D4192D94925A69BA6E9AB6E6676CD939801032256292D59";
    attribute INIT_12 of inst : label is "CF25B483A59A33C42BA14AE94AE80ACECED9DB3B6B209139CC52AF29D268A729";
    attribute INIT_13 of inst : label is "4B69074B34606DDB59E4B69074B25B483A59A3836ECF25B483A59A393249336E";
    attribute INIT_14 of inst : label is "789A68CD552A802AAA969976CA28748955BD32647903201486DDB59ECB720E96";
    attribute INIT_15 of inst : label is "36ADAB6AD8B450966424932D3264D19381AC2C2C0C0C2C2C2C0C0E6B3326AC99";
    attribute INIT_16 of inst : label is "9285250A490049A49429285250A4A1494292840224C2D5B46C93132254953259";
    attribute INIT_17 of inst : label is "DB6D06DB6836DB41B6DC9244B113B28D958D89FFFFE835D8B1685250A4A14942";
    attribute INIT_18 of inst : label is "52954A04B4024D0264CC9512A326649248A4444028282A410C9664C993234120";
    attribute INIT_19 of inst : label is "384BB06B706DB06DB06DB06DB52989B5AC9679676AAE94A941ADA52A054A552A";
    attribute INIT_1A of inst : label is "9292D4AAAD264C8E4C891C99568E75558082C16C20B05B082C16C20B05B205AC";
    attribute INIT_1B of inst : label is "62282D18326C0B0520A51E208148290608876190210820BA4A482F400B6A082E";
    attribute INIT_1C of inst : label is "B899C0992D020C424A2ABB6E8314514493B2F4A5699C6280008B73CA499A3101";
    attribute INIT_1D of inst : label is "92019365906C58A5282959036BAC94AB57A60F28DBB46ED0876E16A54EDDA5A4";
    attribute INIT_1E of inst : label is "D52AEAAD04386948B4AB5A54A1B6A1B6A1BD436D53222222228B226DB6DB6DA5";
    attribute INIT_1F of inst : label is "AAEBAEBB70A4D19ADA3356566A589B22566A5A254ACD4B0489598C0120222A8D";
    attribute INIT_20 of inst : label is "AECB4C9299C03D27400000066D94D790A81611602B086AD2B336FA64BE921B85";
    attribute INIT_21 of inst : label is "4006501A6654B65EBC2784D55B6D575A4934D34D2B01B694242424242426C225";
    attribute INIT_22 of inst : label is "2184984988E020B02321EB616C40443D6D428045650964DCD1956AE6DDC5B652";
    attribute INIT_23 of inst : label is "649249ECF56CF67B3D9ECF2559A7965973222895911115555513262D84931092";
    attribute INIT_24 of inst : label is "0BAD2EB0DE45885209A20D4B64611194D0A249248496492B6B5B2D926B2596CB";
    attribute INIT_25 of inst : label is "652A26E4454E09B8CD9537132A704CC6A4CC4CA96F0414E673A362D5AB32DADD";
    attribute INIT_26 of inst : label is "719D2CDC64A6E33A59B8C94DC676B33192998CED66E35398C6C6E6454E09B8CE";
    attribute INIT_27 of inst : label is "A64733BC65D8D11AD2F47B58BD774692225B9416C6B3719CC8B37189D66E3253";
    attribute INIT_28 of inst : label is "036C11860672A5046DBFB36F75C9C3918C4640EEC28485103056070A49140F59";
    attribute INIT_29 of inst : label is "7504109BD4E6AE14C928182000003300000014906D819800E0BAEBAF6CB82A44";
    attribute INIT_2A of inst : label is "79B12092955207A2C4E056EF67535E2608CE649756AFAA9CB703B841DAF7C2B8";
    attribute INIT_2B of inst : label is "A706A19C6DCE36E71951AD8DA9B2C65CD9632E772D9C10A4D849E848AFEC29F8";
    attribute INIT_2C of inst : label is "204BA538133332222575B055293AB42257A44A8A1504AC00002BEBBE96945934";
    attribute INIT_2D of inst : label is "9492445555555FF4C2D85D03A6824A8824820C012985AC96A69449520492D701";
    attribute INIT_2E of inst : label is "EBACE59635D759CB2C6BAEB39648D75D792A24B4892D224B4892D22D52001264";
    attribute INIT_2F of inst : label is "1BD2110BC6F961F8ED0E75BB27F3B439D726B801FD9DDCF732483AEADA72CB1A";
    attribute INIT_30 of inst : label is "5CAE92BA64CC943F4802020200D2441CCB22E7DEBD7BCA374800001065F497D2";
    attribute INIT_31 of inst : label is "2A891226C63D5A239DFBBF145F99C4C48C9DE509DDC4A4349503125EBB576AED";
    attribute INIT_32 of inst : label is "14000033251A0A201FE941484848485FACFD2A24DF45F4399793B9C4126C2CE9";
    attribute INIT_33 of inst : label is "3AD631AD6B18C7A834D9EF55EA0D7E7BFFF8A2CC75994828FD181D020882C946";
    attribute INIT_34 of inst : label is "A50748A55315D23BAA0634D5B1F10DC4D4DA458C98E59931F7B9CF73DCF7488D";
    attribute INIT_35 of inst : label is "0003A8D2448AA0482C315834B2E0064AC81F06C169107251FFDA982922408D20";
    attribute INIT_36 of inst : label is "00050005000500050005000500050005000ABABBEBFAAFEABC0FEBAFBBBABE90";
    attribute INIT_37 of inst : label is "00024021448042A8002A80001500500050004001400A80150005000500050005";
    attribute INIT_38 of inst : label is "40202280404500050005054150541150A2005457F8050A142FF143150C543800";
    attribute INIT_39 of inst : label is "0000003EBEBEEAFEBD0505250780004D2BC5002801400A00A000500000A01011";
    attribute INIT_3A of inst : label is "0080804240400000000001C0C0000015402E89C5861800000020000000000000";
    attribute INIT_3B of inst : label is "300A00000003FF00000002BEFCAA00000000781C00000155CE1F18080065C001";
    attribute INIT_3C of inst : label is "A80029500054282020050E0000047FFDFBFCFFFFFFFFFCFFFFEAFBF7E55F7C00";
    attribute INIT_3D of inst : label is "C755555547D2131A8C942AD75A852A0A8015054000005000001415054A952A54";
    attribute INIT_3E of inst : label is "555547D21209655555551F2AAAAAAB42E7F7A41EE5DA932ECA91C71C70C30C30";
    attribute INIT_3F of inst : label is "BA810000000000000000002C898EE8B5963B22D658EE8B5963BBEEB92C82B355";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "14041111455C4854594650D49B333DB7922366D84E0190B0C9642BEDEDE27919";
    attribute INIT_01 of inst : label is "FC81F97288E67FE56C2FF800000000000000002BEAABBEF54356426224110501";
    attribute INIT_02 of inst : label is "7FFFFF43E07D0FE07F43FFFFFE87FFFFFD0FFFFFFB2301FFFE40C07FF9031FFF";
    attribute INIT_03 of inst : label is "007E007F007F007F007F007F007F007F007FE07FE07FFFFFA1FFFFFE87FFFFE8";
    attribute INIT_04 of inst : label is "AD72CB372C972CE50E983AABA400005C57181C993DC518142C820682C1040000";
    attribute INIT_05 of inst : label is "CCE666333199B66F6DEF25B2C2CDD9121D34236F3E46788CDB36EB5D416605ED";
    attribute INIT_06 of inst : label is "846E0E9DEF9984645B9EC00402CA1B2CD240C6442492491B112CE89191A4259C";
    attribute INIT_07 of inst : label is "98C19B60038C9FB084924939B63C1397277BE6611B876DE73308E237075E6F99";
    attribute INIT_08 of inst : label is "082E5248C69433208734124924924CC261D9887108B870845C38666D36738333";
    attribute INIT_09 of inst : label is "0000171B549C6D1271B4499025C6C0849A42B838666640A80008000000000A00";
    attribute INIT_0A of inst : label is "0128892631051555559500001289438383823000000000000000000000000000";
    attribute INIT_0B of inst : label is "463A61A1031891061AC325298C5960C3088612DB2C924990E490F1C4E3324927";
    attribute INIT_0C of inst : label is "00000000832450C924935551460D86421E0E27188648C2492492492709348CD8";
    attribute INIT_0D of inst : label is "821B082C42316E62DC10D84801E4270D841246CD32B6DCC8CE2E221C36761000";
    attribute INIT_0E of inst : label is "0D75D1B46D1B491B0912210897112E086C20B108C5B98B70436104884225C44B";
    attribute INIT_0F of inst : label is "9991AF856C84848207C908E45C733214F0AD90909040F9211C8B4C4A74043861";
    attribute INIT_10 of inst : label is "C24241079211C8E16484722D98E6646BE16C84848207C908E45C1B24472258E3";
    attribute INIT_11 of inst : label is "2C61C33A132D0925D0BE5BAC65B77BE9FA3E9FA72981320C736C9CCBA9CEB886";
    attribute INIT_12 of inst : label is "20B242391A728E852CA14B280B294B31310620C414B64D846118398C6592318C";
    attribute INIT_13 of inst : label is "64847234E519922424164847234B242391A728CC9120B242391A7286C924CC91";
    attribute INIT_14 of inst : label is "0C61CB35D7AAAA80AA99E68920078B1C070F89D18614823719224241E488E469";
    attribute INIT_15 of inst : label is "C8D2348D23400F4B99925CD28D138668141080808080A0A0A0A0A394ECD34274";
    attribute INIT_16 of inst : label is "C8D191A32481A71666CC8D191A32346468C8D009D3A5374DD20EB8980A4ACDA6";
    attribute INIT_17 of inst : label is "041188208C4104620820DB62E0E89894C614643FFFE03651428D999A32346468";
    attribute INIT_18 of inst : label is "8C462262C6032D8D623348D11B119A5B6C16666008080B2CE25D1224489524B1";
    attribute INIT_19 of inst : label is "C2B4519493D043D043D043D04B03EE431209045F623A26F05C8981BC72311889";
    attribute INIT_1A of inst : label is "58590208329D2377B336EF662915066733180C10C603043180C10C6030490A53";
    attribute INIT_1B of inst : label is "644CADA39991A4758EB0A1EE5D63AC2857B99243BDEF8F096163901EE401E1C2";
    attribute INIT_1C of inst : label is "76C4EE4D919869B3299B60DB264924924E6B46BE6E4B865C622E0C342E638225";
    attribute INIT_1D of inst : label is "585CCC92473246358DAC2CEFD03B608E1DFD99FF093F84FE1278DC3339899716";
    attribute INIT_1E of inst : label is "BF55D575BCB974A34A14A50A3240324032406480BC111111116E9D924924921A";
    attribute INIT_1F of inst : label is "31C71C7922630A55214A292985264585298523B1A530A47634A46CC1F615554B";
    attribute INIT_20 of inst : label is "19B4336866469FF17B0000036F50D70130CCC0C8D66096E8F88E4918934C4913";
    attribute INIT_21 of inst : label is "2D910B2491066530E4688D2EE492ECA36DC71C71DC4A48E6363636363639449A";
    attribute INIT_22 of inst : label is "D096E465F448C23E128746260CC031C8C406C033702E13FB2441C3992D3A411B";
    attribute INIT_23 of inst : label is "9048361201D209048241208874D345144D1104470888888888CE919896DC92DB";
    attribute INIT_24 of inst : label is "0E0938E5B372E85B36DA19AE99C48C430A592498785D96C48624120DA4824522";
    attribute INIT_25 of inst : label is "6497790A7063F643244BC85C830FB2197321720C11F817BDCEBE4DA84EA393A1";
    attribute INIT_26 of inst : label is "8640532393190C81A647263219014C8E4C643206990CB8723339087061F64326";
    attribute INIT_27 of inst : label is "59BDEDF3BBE7DE6D0D23B467C758B8D9ECA4A258B8CC864CCDCC865C2991C98C";
    attribute INIT_28 of inst : label is "0618430223C982103260E0CA5EAC64C5295DB76C3D6313ACECDD9C9BADA25086";
    attribute INIT_29 of inst : label is "5EB04EC87408224A26C7DA88000099800004CA401B40F4121871C71CD5080E11";
    attribute INIT_2A of inst : label is "58F3366C024503CB64450629A1D05320A14352CC738D55E2E881E630F79247E8";
    attribute INIT_2B of inst : label is "91093C4332A19910CC8CDAE7548D73AA46B9D1218344683248A4797939744C60";
    attribute INIT_2C of inst : label is "A44C3C8861111111198649058DC2365363B6708B05B6340000140B06DAD92587";
    attribute INIT_2D of inst : label is "5ADB076000000AB6C2D85C81B2CB62ECB6CB32EDECB7B2CA10E22C5A16DBDD03";
    attribute INIT_2E of inst : label is "045332C9C608A665938C114CCB2718228593B6D6EDB5BB6D6EDB5BB9DBFFF326";
    attribute INIT_2F of inst : label is "490C4E2B63EFCB0216896ACDDC18DA2DADDE0C84E6582E30B770069A3B9964E3";
    attribute INIT_30 of inst : label is "1603680D32236D8927FB13131399AE1EE2D9B2018307B38CB1FFFFC80C93126C";
    attribute INIT_31 of inst : label is "DEE58B9BDACF4CD6448C94EE294C363AB3205526A48B199B0508EB202C0580B0";
    attribute INIT_32 of inst : label is "EA00000C1AE18A220006BEA8484848406790CDBB49849885B5CCE4781BA6374E";
    attribute INIT_33 of inst : label is "8E739CC6318C67A08027FDFFE82001FF7FFA2831DE67E08A0067F7F8222C26B9";
    attribute INIT_34 of inst : label is "F205F959392B3A3655C42E686C7EE7C1EF2F0642E66645CCCEF79DEF7BCF6E46";
    attribute INIT_35 of inst : label is "0018082B3841CF600EEE1E42482201B02024090274330D200061C315B3600B80";
    attribute INIT_36 of inst : label is "FFC0FFC0FFC0FFC0FFC0FFC0FFC0FFC0FFD41011545110005401141440401570";
    attribute INIT_37 of inst : label is "FF803FDE007FBC07FFC07FFFD0FD0FFC0FFC3FF03FE07FC0FFC0FFC0FFC0FFC0";
    attribute INIT_38 of inst : label is "3FDFC07FBF80FFC0FFC000000F00000E1DFF400007D0A14280043C90F243C7FF";
    attribute INIT_39 of inst : label is "00000000154015001550054404001510A000FE07F03F81F81FFC0FFFF81FEFE0";
    attribute INIT_3A of inst : label is "408080420000404040404140400000000023905830C200000000000000000000";
    attribute INIT_3B of inst : label is "555600000003FC0000000E3EFCAA000000400800100000A2B01FD01000250041";
    attribute INIT_3C of inst : label is "87FE050FFC0287801FD0F1FFFFE47BFDFB1FFFFFF3FFFC1FFFE2FBF7E557D555";
    attribute INIT_3D of inst : label is "4980222222B858F0828A08AB7040A1E07FD0F03FFFFD0FFFFF43C0F02840A142";
    attribute INIT_3E of inst : label is "222222B8586C520088888A80000000CA30CD30CC9248C93248C2492492492492";
    attribute INIT_3F of inst : label is "E78000000000000000000021925A393CB168E4F2C5A193CB160550A58A18E880";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "51454144004D2844E5C2009249111507C20527D80E055008812221C7C6913819";
    attribute INIT_01 of inst : label is "0180F95290047FE5248DF80000000000000000141504400825D244C004542140";
    attribute INIT_02 of inst : label is "000000280D01A005002800000050000000A000000101000000C0400003010000";
    attribute INIT_03 of inst : label is "05000D000D000D000D000D000D000D000D000D000D0000001400000050000005";
    attribute INIT_04 of inst : label is "214208342094208418DC35444D55555D06109904981053E1C282268680020000";
    attribute INIT_05 of inst : label is "88C446223111B86D6DAD45B6868550211090022E9E4478C50180805009440506";
    attribute INIT_06 of inst : label is "24880895A50024805A1A50145688092DC00906002492490A1428A10202800518";
    attribute INIT_07 of inst : label is "18C21B60020C9E10049249220030121425694009222464A200488244045A2500";
    attribute INIT_08 of inst : label is "802C4001161012008400924924924CA25148A04319A0418CD020083040D20102";
    attribute INIT_09 of inst : label is "00001289544A2551289544B218A2487B4A3CA050222022060008888888888000";
    attribute INIT_0A of inst : label is "0021800072150505114000000385C6C6C6C60000000000000000000000000000";
    attribute INIT_0B of inst : label is "04184080012892082281060894484104100C167B64925B814480A188011249A6";
    attribute INIT_0C of inst : label is "000000008212C04924935551020485280C0C4008024882492492492600001010";
    attribute INIT_0D of inst : label is "060D142C46316862D03068A000AC66868A16C28EB29248884C28003812D28000";
    attribute INIT_0E of inst : label is "8544E8BA2E8BA11A09162318B43168183450911844A08940C1A28488C225044A";
    attribute INIT_0F of inst : label is "1101ED052A400000068000C55862203DA1AD48000000500018A9AA2D4020A041";
    attribute INIT_10 of inst : label is "A000000500018AD1C00062AD50C4407B436A400000028000C54A0E00862A5443";
    attribute INIT_11 of inst : label is "A481041D172E9B6CE9BAEA38AEB45D70DC771DC62552A904D92A845AB54AA0C2";
    attribute INIT_12 of inst : label is "00E00031595C1D452A040A940A954AA8A88510A21A925D14C5102388F6DA2388";
    attribute INIT_13 of inst : label is "C00062B2B8294940001C00062B2E00031595C14A4A00E00031595C1FAB6DAA4A";
    attribute INIT_14 of inst : label is "0451611228000000AA95D25480028908040790088A0A0015149400014010C565";
    attribute INIT_15 of inst : label is "54E93A4E93A0050C89B6CAEA0402D220100880808080A0A0A0A0A352B440C401";
    attribute INIT_16 of inst : label is "6060C0C18080C0132346060C0C18183030606001602EB3ACE90B54540C2FA492";
    attribute INIT_17 of inst : label is "0A28F05147828A3C14504926842108B84438844AAAA03441A7468C8C18183030";
    attribute INIT_18 of inst : label is "8C462362430228C5422188D11A110C492412222008080A28C450204081166C9E";
    attribute INIT_19 of inst : label is "A612E05A4160A360A360A360A123E4000000009E622206706889819CA231188D";
    attribute INIT_1A of inst : label is "D0D082410100804200308400753C844433B05828EC160A3B05828EC160A10D6B";
    attribute INIT_1B of inst : label is "444CA983110180750EA181EC5D43A860C7B1100694A504134343029AC0114104";
    attribute INIT_1C of inst : label is "7A48FEDD09B568A02911811DF7DF7DF60A2FC2B4442B42C8F828145625430225";
    attribute INIT_1D of inst : label is "5458880006224E350DA870FF0021208811FD83FE893F44FD5260502320099414";
    attribute INIT_1E of inst : label is "2E551558B9933083A83AD49C10011001100A2002FA11111111E814A924924909";
    attribute INIT_1F of inst : label is "90820821102A8D3691A6743546150D4E354611A8C6A8C23518D568C0F0055542";
    attribute INIT_20 of inst : label is "0A8215042AC05FE3550000014DC2B6007A8C81CC064002A05016402890040881";
    attribute INIT_21 of inst : label is "65920936F20424108C018404400045D124820820884508A2121212121211C001";
    attribute INIT_22 of inst : label is "109254E5504C0E26121446260840A388C40240A3602823FFB481420B2DA1200B";
    attribute INIT_23 of inst : label is "000012000100000000000018404008208611044408888888888A030892489249";
    attribute INIT_24 of inst : label is "00090284834A680A065A00A81B601882891000086850B24000000004A0000402";
    attribute INIT_25 of inst : label is "98023018A0435406040180E8021AA0302203A00828A9423118C8402008201021";
    attribute INIT_26 of inst : label is "0C006A0101101801D40202203003A804044060035018105822301AA041540605";
    attribute INIT_27 of inst : label is "5085B1F223E7886E042A30408240B049EDC0AA2090880C0B30880C0835008088";
    attribute INIT_28 of inst : label is "0228010611418308370088108E28204D6B568508052100A6464CC8C9A4AA21C2";
    attribute INIT_29 of inst : label is "0C8006887408240002474000000000000000AD08A120D2115820820850100E11";
    attribute INIT_2A of inst : label is "187334440AC6030A24010619D1D033108001428C718C00C280818630C70007C0";
    attribute INIT_2B of inst : label is "92839AA6AA935549AAAA68D562146AB90A355821040C0022C884593911B44444";
    attribute INIT_2C of inst : label is "A0049C94311111111C92DB0484C222D1231230810492200000000B06484B2C93";
    attribute INIT_2D of inst : label is "4ACA832000000AB240480C00905922459259B2CCA43296581242244A02494F03";
    attribute INIT_2E of inst : label is "12EA02810425D40502084BA80A0410974CB19242649099242649099089FFF2A5";
    attribute INIT_2F of inst : label is "09040A0A61C5E20638F342F24C0863C50A4E4C00C2502850A49006BA5B014082";
    attribute INIT_30 of inst : label is "19020418200525180002020203949418A30000848912B349B00000180C811204";
    attribute INIT_31 of inst : label is "5E64C993909E4456C40480AE0888B53283105510000B190B0504CA90320640C8";
    attribute INIT_32 of inst : label is "00000040E00E0000001800084848484063A044A148048005358468280A221448";
    attribute INIT_33 of inst : label is "0C6318C6318C67A88B1A12ABEA228684807AA3032BBAAAA882884A800A011802";
    attribute INIT_34 of inst : label is "4000F81121037A37550008188038A4C3EA0C0AC7426ACE848E739CEF7BCE2443";
    attribute INIT_35 of inst : label is "00100C2A28414E400AAA16202060089044110440501626215501031491200200";
    attribute INIT_36 of inst : label is "001A001A001A001A001A001A001A001A003501000011155540011404F5554010";
    attribute INIT_37 of inst : label is "00288000510000D0000D00001A00A001A00180068015002A001A001A001A001A";
    attribute INIT_38 of inst : label is "80000500000A000A000AFABEA0ABE2A140002BA8001A3468D002800A00280000";
    attribute INIT_39 of inst : label is "000000001555EABFE955502412801542140A0050028014014000A00001400002";
    attribute INIT_3A of inst : label is "0101000100000000000003001500001555615848100000000000000000000000";
    attribute INIT_3B of inst : label is "0003FFFFFFFC03FFFFFFF1C102AA000000000000000000A8BFE0002000250003";
    attribute INIT_3C of inst : label is "5000D0A001A85040000A0000000F840204E000000C0003E0001D040815560000";
    attribute INIT_3D of inst : label is "5980222222F150C1FBEBFF29450A1405000A02800000A00000280A02850A1428";
    attribute INIT_3E of inst : label is "222222F150E8420088888BD5555555EA209021CCDA4889324886596596596596";
    attribute INIT_3F of inst : label is "FF8100000000000000000023580215982008566080215982004001B508308180";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
