-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0008000000000016080000000000640000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0A98008101800639C780D2002440E60008780000090102B4964000000040E800";
    attribute INIT_02 of inst : label is "6FFF606009FF3FFFFFE20909FD60FFF8903302BF1E00C8338FA6FE8000B4CC33";
    attribute INIT_03 of inst : label is "0EAA020002007FFCA200000000C02FF5003F000B050F0038FC00E000F0502C00";
    attribute INIT_04 of inst : label is "00000FFFAFC000000000FFF000000000000500FF55000000FF50FFFF00000000";
    attribute INIT_05 of inst : label is "9E000007500099C0EAAB2BE83FAA000005FF0000FC0000005000000003FA0000";
    attribute INIT_06 of inst : label is "03C0F57CF03C15E0F028157C7D543F80F0287D5005F8B5780F000F8070B42D60";
    attribute INIT_07 of inst : label is "0005039901E000B02AA800000B400E00000003C0014000007800B578F50C2578";
    attribute INIT_08 of inst : label is "F0B455E0003C557C00F055F0783C2D7CA0B4B5E0F03CB57CF57C2DE0D743B55E";
    attribute INIT_09 of inst : label is "F03CB578FD3CF0BCF13CF8BC00F000F02F7C783CF828F0000F005F50F03CF03C";
    attribute INIT_0A of inst : label is "7DF4F03C1FD0F03CF03CF03C0F005F50F0282D782F7CB57C0099D000157CB57C";
    attribute INIT_0B of inst : label is "15540000B50099B00C000A8009000008003002A001F8FD540F00F0F0BDF8F8BC";
    attribute INIT_0C of inst : label is "1E003000000C000C000000010000EAAA00B4000C0000AAAB0000400030003000";
    attribute INIT_0D of inst : label is "00000000000C000D00000000300002AA00000000000CAA800000000030007000";
    attribute INIT_0E of inst : label is "00B4000C000CAA871E0030003000D2AA0000AAAA00000000000C000C30003000";
    attribute INIT_0F of inst : label is "000000000000AAAF000000000000FAAA000C000C000C000F300030003000F000";
    attribute INIT_10 of inst : label is "002F000C000CAAFFF80030003000FFAA000000000000D0000000000000000007";
    attribute INIT_11 of inst : label is "002F00000000AAFFF80000000000FFAA002F000C000C00FFF80030003000FF00";
    attribute INIT_12 of inst : label is "003F000C000DAAFFFFFC3000FF50FFFFF80000000000FF00002F0000000000FF";
    attribute INIT_13 of inst : label is "000500FF003F0000003F00000005AAFFFFFC0000FF50FFFF003F000C000D00FF";
    attribute INIT_14 of inst : label is "03FF000C005F0FFFFFC03000F500FFF003FF000C005FAFFFFFC03000F500FFFA";
    attribute INIT_15 of inst : label is "005F0FFFF500FFF003FF0000FFC0000003FF0000005FAFFFFFC00000F500FFFA";
    attribute INIT_16 of inst : label is "FC0000005000FFAAFC0030007000FF003FFF000C05FFFFFFFC0030007000FFAA";
    attribute INIT_17 of inst : label is "03FF0000005F0FFFFFC00000F500FFF05000FF00FC0000003FFF000005FFFFFF";
    attribute INIT_18 of inst : label is "002B000000002FFFC00000000000C0003FFF00BF050F3FFCFFFEAFA02140EDBE";
    attribute INIT_19 of inst : label is "0C33000001400C330CD0000050400CC02D99D02A07B9399999B8A8079BD0999C";
    attribute INIT_1A of inst : label is "03FF0000005F0FFFFFC00000F500FFF0003F0000000500FFFFFC0000FF50FFFF";
    attribute INIT_1B of inst : label is "0000000000000007000000000000D0003FFF000005FFFFFFFC0000005000FF00";
    attribute INIT_1C of inst : label is "BD0002BF07F83F550FC0E000001557FCFFE00000005F07FF0FF8FFFFFFFF03FE";
    attribute INIT_1D of inst : label is "30C000000600000018000000000C00C00030000000240040000200000006200C";
    attribute INIT_1E of inst : label is "0000000003D9D000005F0F9999C000071FE8002BFF4002BF003FFE802FC0D7F4";
    attribute INIT_1F of inst : label is "FFFF0000FFFC0000FFF00000FFC00000FF000000FC000000F0000000C0000000";
    attribute INIT_20 of inst : label is "57FA00010000FE08AFD50000000000BF00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "07FA00030000FE08AFD00000000000BF000000AAF40000000000AA00001F0000";
    attribute INIT_22 of inst : label is "01F0293CBFD4FCC00000400000000000000028AAF40000000000AA28001F0000";
    attribute INIT_23 of inst : label is "01F0293CBFD4FC000000540000000000000000000000000034003000078003FA";
    attribute INIT_24 of inst : label is "00FC003CAB40FA800000000000000000000000000000000034003000278023FA";
    attribute INIT_25 of inst : label is "000002A0340000000000A8080278000000000000000000003C00F0001FFA00AA";
    attribute INIT_26 of inst : label is "0007003FFFF00000C000FFA00000000007A000000000300002F4000000000030";
    attribute INIT_27 of inst : label is "0007003FFD7400008000FFFF0000000000030AFF00000000D000FC0C0FFF0000";
    attribute INIT_28 of inst : label is "000202D700000000F000FE0403F000000002FFFF00000000D000FC061D7F0000";
    attribute INIT_29 of inst : label is "030B0BD700000000FC00FF8001E0F0000E00005700000000AFF4FC043000A4FC";
    attribute INIT_2A of inst : label is "FFFFFFFFFFD4A8008000F000000000000E00021F00030002AFE0FC00F00090F0";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFEAFF00FFC0F40000000002000F00000000FFFFFFFF07FF002A";
    attribute INIT_2C of inst : label is "000002FF2FFF00000000FF80FFF8000000FF03FF001F0000FFFFFFFFFFFFABFF";
    attribute INIT_2D of inst : label is "02FF3FFFFFFF0000FF80FFFCFFFF000007FF001F00003FFFFFD0F4000000FFFC";
    attribute INIT_2E of inst : label is "00C200B7000500008300FE00500000007FFF0FFF0005FFFFFFFDFFF05000FFFF";
    attribute INIT_2F of inst : label is "006B03F30000002AE900FFC00000A8000B580F1C00000000BE0ED6C300000000";
    attribute INIT_30 of inst : label is "3C333C7300000000FC0E5B0350000000001503F9A28000BF5400FFC0028AFE00";
    attribute INIT_31 of inst : label is "03D0015400050000C000BFC054B40000B58BF1CD00000000FE1F6F0F50140030";
    attribute INIT_32 of inst : label is "3737333315150000370F330C1515000000030F0F005F0000FD8485C040000280";
    attribute INIT_33 of inst : label is "00001207000000000000F6550000000000007F65000000000000500000000000";
    attribute INIT_34 of inst : label is "727D7472686E2F8A373FBFE00B6FFFE000004087000000000000F95500000000";
    attribute INIT_35 of inst : label is "003F0038050F000BFC002C00F050E000003F0038000F280BFC002C00F000E028";
    attribute INIT_36 of inst : label is "0EAA7FFC20002000A2002FF50C0000001FFF207A00000A8080000FC057F82000";
    attribute INIT_37 of inst : label is "F2DE3E507EB72FF85EBD29FFA2F82BF80EAA7FFC02000200A2002FF500C00000";
    attribute INIT_38 of inst : label is "000900030000000B900000000000E000F4BF3D9838660BFA39F097DF81BC2BE0";
    attribute INIT_39 of inst : label is "0004000F000300010000F000C00000000000000F000300024000F000C0000000";
    attribute INIT_3A of inst : label is "FFFE002F3FF80000FD60D5A007FFBE8002C70794FC1EBE00FD940780543E00A0";
    attribute INIT_3B of inst : label is "0010009F000000000000C0000000000000000000020002800034000003F80000";
    attribute INIT_3C of inst : label is "0B0F1BF8001D0000FEA09FF475000000009C00F20000000072004D0000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000008000000200002200210000008800008";
    attribute INIT_3E of inst : label is "0000000400000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "3D1D707F5AFF000007420387541F2FF88074D0B5D47E2FE0A07C203DAAFE0000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "001E000000000024900000000000420000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "049A014B0001088BF4300860050025E0001300800000029F9D0000800000DF00";
    attribute INIT_02 of inst : label is "3FFF06FF90909FFFFFF4FE900606FFD1C0332D00017F67F3CC330078FD40C7D9";
    attribute INIT_03 of inst : label is "BFFC010001000D551FFA00C0000051000035287F0003002F5C00FD28C000F800";
    attribute INIT_04 of inst : label is "00010015FFF000008000500000EA000A0002003F00ABFFA04000FFFC00000000";
    attribute INIT_05 of inst : label is "99C0A000000B99001EB4D55715FF000000013EAA540000008000FC000FFF0000";
    attribute INIT_06 of inst : label is "01401E0015502ABC1550B55414003C7815502F8055547E8055500F000540F03C";
    attribute INIT_07 of inst : label is "E000007900100B4000002AA8040001E000000060000002800550FAB415501AF4";
    attribute INIT_08 of inst : label is "5540A83C00142ABC55502AF00554F03C1540003C15547ABC5014F03C7AADEB83";
    attribute INIT_09 of inst : label is "1550F03C5014FBFC5014FFFC555000F0541407BC1550F00055500F005014FABC";
    attribute INIT_0A of inst : label is "1010FBBC0100F8BC1550F03C05000F0015502AB45414F83C0399000A0014F03C";
    attribute INIT_0B of inst : label is "00002AA8000B9BC00E800C001000009002B0003055541F8005003AC050141FD0";
    attribute INIT_0C of inst : label is "01553000000E000C00000000000000005540000C0000000000000000B0003000";
    attribute INIT_0D of inst : label is "00020000000C000CD555000030002D0055570000000C00788000000030003000";
    attribute INIT_0E of inst : label is "554B000C000C0078E155300030002D000000000055550000000C000C30003000";
    attribute INIT_0F of inst : label is "555F000000000000F555000000000000000F000C000C000CF000300030003000";
    attribute INIT_10 of inst : label is "55FF000C000C001FFF5530003000F400E000000000000000000B000000000000";
    attribute INIT_11 of inst : label is "55FF00000000001FFF5500000000F40000FF000C000C001FFF0030003000F400";
    attribute INIT_12 of inst : label is "55FF000E000C003FFFFFFFA03000FFFCFF0000000000F40000FF00000000001F";
    attribute INIT_13 of inst : label is "0000003F00FF000A55FF000A0000003FFFFFFFA00000FFFC00FF000E000C003F";
    attribute INIT_14 of inst : label is "0FFF00AF000C03FFFFF0FA003000FFC05FFF00AF000C03FFFFF5FA003000FFC0";
    attribute INIT_15 of inst : label is "000003FF0000FFC00FFF00AFFFF0FA005FFF00AF000003FFFFF5FA000000FFC0";
    attribute INIT_16 of inst : label is "FF15A0000000FC00FF00B0003000FC00FFFF0AFF000C3FFFFF55B0003000FC00";
    attribute INIT_17 of inst : label is "0FFF00AF000003FFFFF0FA000000FFC00000FC00FF00A000FFFF0AFF00003FFF";
    attribute INIT_18 of inst : label is "02FF000000005555C0002000000040001FFF0FFF00B71FFFFFFFFFF8FE80C7FD";
    attribute INIT_19 of inst : label is "0C33028000000C330CC0A08000000CC039990BD9E0151D99999C9DE0540B99B4";
    attribute INIT_1A of inst : label is "0FFF00AF000003FFFFF0FA000000FFC000FF000A0000003FFFFFFFA00000FFFC";
    attribute INIT_1B of inst : label is "000B000000000000E000000000000000FFFF0AFF00003FFFFF00A0000000FC00";
    attribute INIT_1C of inst : label is "FEAA2FD000540F80ABF07E000000007E1FFCFFC0000101FF0FFCFFF5FFFFE3FF";
    attribute INIT_1D of inst : label is "1A40202A005A000003008000AA900043009000090A9000020809000000A9400C";
    attribute INIT_1E of inst : label is "000000000D9900ADE000039999F0FA0000550BF50000BFF4EBFC05FE15000BD0";
    attribute INIT_1F of inst : label is "0000FFFF0000FFFC0000FFF00000FFC00000FF000000FC000000F0000000C000";
    attribute INIT_20 of inst : label is "0105000000005F8650400000000002F500000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0105000100005F8650400000000002F50000AB4030000000000001EA000C0000";
    attribute INIT_22 of inst : label is "003C02F0FCC07FE800000000000000000000AB4030000000000001EA000C0000";
    attribute INIT_23 of inst : label is "003C02F0FC007FE8000000000000000000000000000000003000380003F50B40";
    attribute INIT_24 of inst : label is "003018B4540401F8000000000000000000000000000000003000380013F51B40";
    attribute INIT_25 of inst : label is "00002FF5F000000000005780043C000000000000000000003000380001500B50";
    attribute INIT_26 of inst : label is "000B0AFD50410078E8005000400000000055000000003C00F5400000000000FC";
    attribute INIT_27 of inst : label is "000B02FF0000007EFEA0550000002A00002B000500010000E0007FA141052D00";
    attribute INIT_28 of inst : label is "00AB0D0000000000FC085FF800FC30000ABF0055000000A8E008FF800000BD00";
    attribute INIT_29 of inst : label is "012F0D0000000003FC005FD000F0F00001EB000100000000FD08F000000003F0";
    attribute INIT_2A of inst : label is "FFFFFFFF5400FFE8F00040000000000007EB030700000000FF40FC00F00002D0";
    attribute INIT_2B of inst : label is "FFFFFFFFFFD5FFFFFFC0FF000000F800000F000100000000FFFFFFFF00152BFF";
    attribute INIT_2C of inst : label is "002F0BFF3FFF0000F800FFE0FFFC0000037F00FF0000002FFFFFFFFF57FFFFFF";
    attribute INIT_2D of inst : label is "0FFFBFFFFFFF000AFFF0FFFEFFFFA00001FF000000001FFFFF4000000000FFF4";
    attribute INIT_2E of inst : label is "00150079007A00BF5400FD00AD00FE003FFF01FF0000FFFFFFFCFF400000FFFF";
    attribute INIT_2F of inst : label is "00AA005E007A00D5AA00F500AD0057000F2C07A400000000FFC37D0D00000000";
    attribute INIT_30 of inst : label is "3CB31E9300000000FF03FC0D0000A00000B7007F01FF00C2FE00FD00FF408300";
    attribute INIT_31 of inst : label is "0F0F0003000000AF4AC0E74801408000F2CF7A4700000000FF0FFD2F0030A028";
    attribute INIT_32 of inst : label is "33333B3B00002A2A330C3B0C00002A0802A803E00000000A7BC0C0000000A878";
    attribute INIT_33 of inst : label is "048B000000000000F6A0000000000000BF6A0000000000000000000000000000";
    attribute INIT_34 of inst : label is "D45DB22407F4BD7706F4DBDE5AF4EFFC080B000000000000F9A0000000000000";
    attribute INIT_35 of inst : label is "0035002F0003287F5C00F800C000FD280035142F0003007F5C00F814C000FD00";
    attribute INIT_36 of inst : label is "BFFC0D55100010001FFA510000000C0007FD000500103FFE3804FFE000140000";
    attribute INIT_37 of inst : label is "1E1281C901402D7D4978CB747F54F1FFBFFC0D55010001001FFA5100000000C0";
    attribute INIT_38 of inst : label is "000300000000000FC00000000000F0001E4DF21705FA3F1B46FC376FFD40FFFC";
    attribute INIT_39 of inst : label is "000B000600030000E000600000004000000B000900030008E000900000001000";
    attribute INIT_3A of inst : label is "1F5F0AF507F42FE0F87C0BFE00547FF00BD6286F0500792B13D02E400015E3FE";
    attribute INIT_3B of inst : label is "000D000000000000E4000000000000000000000007D00F4000000080005000F8";
    attribute INIT_3C of inst : label is "2FF9057F000500AE1FDCF0D00000B80002DB000700000002A780D00000008000";
    attribute INIT_3D of inst : label is "00010000000000005000000000000000000008D0000021800000002C000000C4";
    attribute INIT_3E of inst : label is "000C000000000000000000000000000000090000000000000000000000000000";
    attribute INIT_3F of inst : label is "F082F03F01500BF8830F0BFA0000FFF4F030ABF0000557EF703FF03807FDABE0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "000800000000001B008000000000F40000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0A98008101900633A700D2006040E600087800000901022F1E40000000407000";
    attribute INIT_02 of inst : label is "6232606009FF33333A220909FD6033782FFF000001FF3FFFFFF80000FF40FFFC";
    attribute INIT_03 of inst : label is "0400BF80BF800A0F07400A803FF0D0001400BE001F400A07001400BE01F4D0A0";
    attribute INIT_04 of inst : label is "005F0000FFC00000F5000000003F0000000000FFAAFC00000000FFFF00000000";
    attribute INIT_05 of inst : label is "9900000F506099002BE800000055000005FFFFFF000000005000FF0003FF0000";
    attribute INIT_06 of inst : label is "03C0F57CF03C15E0F028157C7D543F80F0287D5005F8B5780F000F8070B42D60";
    attribute INIT_07 of inst : label is "0905009901E000B02AA800000B400E00000003C0014000007800B578F50C2578";
    attribute INIT_08 of inst : label is "F0B455E0003C557C00F055F0783C2D7CA0B4B5E0F03CB57CF57C2DE0D743B55E";
    attribute INIT_09 of inst : label is "F03CB578FD3CF0BCF13CF8BC00F000F02F7C783CF828F0000F005F50F03CF03C";
    attribute INIT_0A of inst : label is "7DF4F03C1FD0F03CF03CF03C0F005F50F0282D782F7CB57C0049F000157CB57C";
    attribute INIT_0B of inst : label is "15540000006099000C000A8009000008003002A001F8FD540F00F0F0BDF8F8BC";
    attribute INIT_0C of inst : label is "E000C000000300030000000000001555000B00030000555400000000C000C000";
    attribute INIT_0D of inst : label is "000000000003000200000000C000FD55000000000003557F00000000C0008000";
    attribute INIT_0E of inst : label is "000B00030003557FE000C000C000FD55000055550000000000030003C000C000";
    attribute INIT_0F of inst : label is "0000000000005557000000000000D5550003000300030007C000C000C000D000";
    attribute INIT_10 of inst : label is "002F0003000355FBF800C000C000FF55000000000000D0000000000000000007";
    attribute INIT_11 of inst : label is "002F0000000055FBF80000000000FF55002F0003000300FBF800C000C000FF00";
    attribute INIT_12 of inst : label is "003F0003000755F9FFFCC000FF50FFFFF80000000000FF00002F0000000000FB";
    attribute INIT_13 of inst : label is "000500F9003F0000003F0000000555F9FFFC0000FF50FFFF003F0003000700F9";
    attribute INIT_14 of inst : label is "03FF0003005F0F9FFFC0C000F500FFF003FF0003005F5F9FFFC0C000F500FFF5";
    attribute INIT_15 of inst : label is "005F0F9FF500FFF003FF0000FFC0000003FF0000005F5F9FFFC00000F500FFF1";
    attribute INIT_16 of inst : label is "FC0000005000FF55FC00C000D000FF003FFF000305FFF9FFFC00C000D000FF55";
    attribute INIT_17 of inst : label is "03FF0000005F0F9FFFC00000F500FFF05000FF00FC0000003FFF000005FFF9FF";
    attribute INIT_18 of inst : label is "002B000000002FFFF00000003000F0003FDD00BF05003FD37FFEAFA0DD4047FE";
    attribute INIT_19 of inst : label is "0C33000001400C330CD0000050400CC00199F000081909999980000F91209990";
    attribute INIT_1A of inst : label is "03FF0000005F0FFFFFC00000F500FFF0003E0000000500FEA07C0000FF50A03F";
    attribute INIT_1B of inst : label is "000000000000000800000000000020003EA0000005FFFEA07C00000050003F00";
    attribute INIT_1C of inst : label is "024000001800C0AA30000000006AA8000000000001A018007000000000000400";
    attribute INIT_1D of inst : label is "0F0002FF01FE000007F8E800AFF0003F3FC002BEFFD0FFAF3FFD00280FF8D3F0";
    attribute INIT_1E of inst : label is "000000000099F000090101999800000F20100000009000000040000000302809";
    attribute INIT_1F of inst : label is "FFFF0000FFFC0000FFF00000FFC00000FF000000FC000000F0000000C0000000";
    attribute INIT_20 of inst : label is "F800000A00000008002F80000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "F800000000010008002F0000000000000000BF00003D0000000000FE7C000000";
    attribute INIT_22 of inst : label is "00002900002A03FE00003400000000000000BF00003D0000000000FE7C000000";
    attribute INIT_23 of inst : label is "00002900002A03FE0000034000000000000000000000000000A000E0F800BC00";
    attribute INIT_24 of inst : label is "00020003000800000000000000000000000000000000000000A000E0F800BC00";
    attribute INIT_25 of inst : label is "0000001F0000000000005007020000000000000000000000002F000000000005";
    attribute INIT_26 of inst : label is "14000000000F00023C000000F000A000000000000000C0F0000000000000000F";
    attribute INIT_27 of inst : label is "00000000000000007FC00000FF000000003C0000000F000A0014000CF0008000";
    attribute INIT_28 of inst : label is "0AA01D0002800000000001FD0000000003FD000000FF00000000000600000000";
    attribute INIT_29 of inst : label is "0FF400000A00000002FE00000000000000003FA800000380000001FD0000A400";
    attribute INIT_2A of inst : label is "FFFEFFFFFFD4A8008000F0000000000000000BE001540E02000002FE00009000";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFEAFF00FFC0F40000000002000F00000000FFFFFFFF17FF002A";
    attribute INIT_2C of inst : label is "000002FF2FFF00000000FF80FFF8000000FF033F001F0000FFFFFFFFFFFFABFF";
    attribute INIT_2D of inst : label is "02FF3FFFFFFF0000FF80FFFCFFFF000007FF001F00003FFFFFD0F4000000FFFC";
    attribute INIT_2E of inst : label is "0B0201400000000080E00140000000007FFF0FFF0005FFFFFFFDFDF05000FFFF";
    attribute INIT_2F of inst : label is "2FAB000000000000EAF8000000000000000F001F007F00004000000040000000";
    attribute INIT_30 of inst : label is "003C007C01FF002800000000000000002FFF000000000000FFF8000000000000";
    attribute INIT_31 of inst : label is "00000EFF00000000FF00400000000000007C007C01FF00280000000000000000";
    attribute INIT_32 of inst : label is "3737333315150000370F330C151500000BFC000F000000000000FA00BD000000";
    attribute INIT_33 of inst : label is "000A800700000000A000F95000000000AA007F95000000000000000000000000";
    attribute INIT_34 of inst : label is "0D828B8D17910000C8C04000F4900000000A210700000000A000F65000000000";
    attribute INIT_35 of inst : label is "14000A071F40BE000014D0A001F400BE14000A071F40BE000014D0A001F400BE";
    attribute INIT_36 of inst : label is "04000A0FBF80BF800740D0003FF00A800600FF0500BF000B00B8F055C000F800";
    attribute INIT_37 of inst : label is "0D2101AF01400000A140D6005D00000004000A0FBF80BF800740D0003FF00A80";
    attribute INIT_38 of inst : label is "000600000000003B600000000000EC000B40026707990000C60068207E400000";
    attribute INIT_39 of inst : label is "0000003F000300080000FC00C00010000000003F000300040000FC00C0004000";
    attribute INIT_3A of inst : label is "00000000000000000000000000000000003B006F000000009240FC0000000000";
    attribute INIT_3B of inst : label is "027B06EC09060000BB00BD6000C0200000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "6BF47F87097F201A1FE962FDFD60A40801FF09FF09110008FF40BF6060600000";
    attribute INIT_3D of inst : label is "0002000F00000000A000FC000000000020000040C60124062000000002190244";
    attribute INIT_3E of inst : label is "000A001F00000000A000F40000000000000A001F000000008000FC0000000000";
    attribute INIT_3F of inst : label is "3FFF7FFF7FFF0000FFFFFFFF541F2FF8FFFFFFFFD47F2FE0FFFCFFFDFFFE0000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0095008000000024900000000000460000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "041301CB00010849F6302860050023F0001E0080000002099D00008000009B00";
    attribute INIT_02 of inst : label is "333306FF909091313534FE90060631113FFF02FF00001FFFFFFCFF800000FFF4";
    attribute INIT_03 of inst : label is "050F7F407F400800E0003FF005400B80000FFF4C00003FE0F00031FF00000BFC";
    attribute INIT_04 of inst : label is "000003EAF540FA000000AFC000FF000000000001FFFF00000000550000000000";
    attribute INIT_05 of inst : label is "9900A090000F92001FF40000EA000AFF00003FFFAB00A0000000FC00015F00AF";
    attribute INIT_06 of inst : label is "01401E0015502ABC1550B55414003C7815502F8055547E8055500F000540F03C";
    attribute INIT_07 of inst : label is "F000009900100B4000002AA8040001E000000060000002800550FAB415501AF4";
    attribute INIT_08 of inst : label is "5540A83C00142ABC55502AF00554F03C1540003C15547ABC5014F03C7AADEB83";
    attribute INIT_09 of inst : label is "1550F03C5014FBFC5014FFFC555000F0541407BC1550F00055500F005014FABC";
    attribute INIT_0A of inst : label is "1010FBBC0100F8BC1550F03C05000F0015502AB45414F83C009906000014F03C";
    attribute INIT_0B of inst : label is "00002AA8000F99000E800C001000009002B0003055541F8005003AC050141FD0";
    attribute INIT_0C of inst : label is "FEAAC000000100030000000000000000AABF000300000000000000004000C000";
    attribute INIT_0D of inst : label is "00000000000300032AAA0000C000D000AAA800000003000700000000C000C000";
    attribute INIT_0E of inst : label is "AABF000300030007FEAAC000C000D00000000000AAAA000000030003C000C000";
    attribute INIT_0F of inst : label is "AAAB000000000000EAAA000000000000000B000300030003E000C000C000C000";
    attribute INIT_10 of inst : label is "AAF700030003001FFFAAC000C000F400E000000000000000000B000000000000";
    attribute INIT_11 of inst : label is "AAF700000000001FFFAA00000000F40000F700030003001FFF00C000C000F400";
    attribute INIT_12 of inst : label is "AAF3000B0003003EFFFFFFA0C000FFFCFF0000000000F40000F700000000001F";
    attribute INIT_13 of inst : label is "0002003E00F3000AAAF3000A0002003EFFFFFFA04000FFFC00F3000B0003003E";
    attribute INIT_14 of inst : label is "0F3F00AF000303EFFFF0FA00C000FFC0AF3F00AF000303EFFFFAFA00C000FFC0";
    attribute INIT_15 of inst : label is "000103EF8000FFC00F3F00AFFFF0FA008F3F00AF000103EFFFFAFA008000FFC0";
    attribute INIT_16 of inst : label is "FFAAA0008000FC00FF00E000C000FC00F3FF0AFF00033EFFFFAAE000C000FC00";
    attribute INIT_17 of inst : label is "0F3F00AF000103EFFFF0FA008000FFC08000FC00FF00A000F3FF0AFF00013EFF";
    attribute INIT_18 of inst : label is "02FF000000005555F0000000000070001FE00FFF00001FC00FFFFFF801003BFD";
    attribute INIT_19 of inst : label is "0C33028000000C330CC0A08000000CC009990489F000019999909810000F9980";
    attribute INIT_1A of inst : label is "0FFF00AF000103FFFFF0FA008000FFC000FD000A0002003D503FFFA0400050BC";
    attribute INIT_1B of inst : label is "00000000000000010000000000004000FD500AFF00013D503F00A0008000BC00";
    attribute INIT_1C of inst : label is "0100002501A83000040080000000018060000000000606003000000A00000000";
    attribute INIT_1D of inst : label is "05000FD500050BE000FE7F80554002BCFF420FF41540FFFDF7F40BFF01540BF0";
    attribute INIT_1E of inst : label is "0000000000990600F0000019998080900580000A5500000900035A002AC04024";
    attribute INIT_1F of inst : label is "0000FFFF0000FFFC0000FFF00000FFC00000FF000000FC000000F0000000C000";
    attribute INIT_20 of inst : label is "7C0000010000A006003D00000000000A00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "7C00000A0000A006003D80000000000A00005400000000000000001500000000";
    attribute INIT_22 of inst : label is "0000000003FD0015200000000000000000005400000000000000001500000000";
    attribute INIT_23 of inst : label is "0000000003FD00150200000000000000000000000000000000D000507C00F400";
    attribute INIT_24 of inst : label is "000F1800A00B00000000000000000000000000000000000000D000507C00F400";
    attribute INIT_25 of inst : label is "000000000000000000000000040300000000000000000000C0F00000002F0000";
    attribute INIT_26 of inst : label is "000000020007A80710008000D000FC00000A00000000001F0000000000000001";
    attribute INIT_27 of inst : label is "0000000000007C0003402800FD00BF80000400020007003F00008001D000D02A";
    attribute INIT_28 of inst : label is "3F5400000340000002FE00000000000001C00028007D02FE000800000000003D";
    attribute INIT_29 of inst : label is "07D000000D0002A801FD0000000000002E0005500000014002FE000000000000";
    attribute INIT_2A of inst : label is "FFFFFFFF5400FFE8F00040000000000000000FF800000500000001FD00000000";
    attribute INIT_2B of inst : label is "FFFFFFFFFFD5FFFFFFC0FF000000F800000F000100000000FFFFFFFF00152BFF";
    attribute INIT_2C of inst : label is "002F0BFF3FFF0000F800FFE0FFFC0000037F00E70000002FFFFFFFFF57FFFFFF";
    attribute INIT_2D of inst : label is "0FFFBFFFFFFF000AFFF0FFFEFFFFA00001FF000000001FFFFF4000000000FFF4";
    attribute INIT_2E of inst : label is "0FFF000000000000FFF00000000000003FFF01FD0000FFFFFFFC5B400000FFFF";
    attribute INIT_2F of inst : label is "1F5500000000020055F4000000000080002F000F000000BF0000800000008000";
    attribute INIT_30 of inst : label is "00BC003C001402FF00000000000000001F4000000000020201F4000000008080";
    attribute INIT_31 of inst : label is "000F07FC00000000F500000000007E0000BC00BC001402FF0000000000000000";
    attribute INIT_32 of inst : label is "33333B3B00002A2A330C3B0C00002A080DFF0000000000008000FF0000000000";
    attribute INIT_33 of inst : label is "820B000500000000F9A0500000000000BF9A5500000000000000000000000000";
    attribute INIT_34 of inst : label is "2BA24DDB00000288F900242005001000410B000500000000F6A0500000000000";
    attribute INIT_35 of inst : label is "000F3FE00000FF4CF0000BFC000031FF000F3FE00000FF4CF0000BFC000031FF";
    attribute INIT_36 of inst : label is "050F08007F407F40E0000B8005403FF0BA0F1408001F0063C1FF0000C000F400";
    attribute INIT_37 of inst : label is "01ED2E3600000282B680348000000E00050F08007F407F40E0000B8005403FF0";
    attribute INIT_38 of inst : label is "000300000000003FC00000000000FC0001B20DE8000500E4B900C89000000000";
    attribute INIT_39 of inst : label is "003B000900000002EC00900000008000003B000600000000EC00600000008000";
    attribute INIT_3A of inst : label is "00000000000000000000000000000000002F024600000600EE00D90000000000";
    attribute INIT_3B of inst : label is "06F600B7000006847F4067000000909000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "BF4697F8102506BFE1FE2FD65804FE901BF402FF0000068B5FE0F7800000E290";
    attribute INIT_3D of inst : label is "000F000100000000FC0050000000000000001000110096090038088101940013";
    attribute INIT_3E of inst : label is "003F000000000000FC00000000000000003F000100000000F800500000000000";
    attribute INIT_3F of inst : label is "FFFFFFFF01500BF8FFFFFFFF0000FFFEFFFFFFFF0005FFEFFFFFFFF807FDABE0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
